

module top
(
  i,
  o
);

  input [6399:0] i;
  output [6399:0] o;

  bsg_flatten_2D_array
  wrapper
  (
    .i(i),
    .o(o)
  );


endmodule



module bsg_flatten_2D_array
(
  i,
  o
);

  input [6399:0] i;
  output [6399:0] o;
  wire [6399:0] o;
  assign o[6399] = i[6399];
  assign o[6398] = i[6398];
  assign o[6397] = i[6397];
  assign o[6396] = i[6396];
  assign o[6395] = i[6395];
  assign o[6394] = i[6394];
  assign o[6393] = i[6393];
  assign o[6392] = i[6392];
  assign o[6391] = i[6391];
  assign o[6390] = i[6390];
  assign o[6389] = i[6389];
  assign o[6388] = i[6388];
  assign o[6387] = i[6387];
  assign o[6386] = i[6386];
  assign o[6385] = i[6385];
  assign o[6384] = i[6384];
  assign o[6383] = i[6383];
  assign o[6382] = i[6382];
  assign o[6381] = i[6381];
  assign o[6380] = i[6380];
  assign o[6379] = i[6379];
  assign o[6378] = i[6378];
  assign o[6377] = i[6377];
  assign o[6376] = i[6376];
  assign o[6375] = i[6375];
  assign o[6374] = i[6374];
  assign o[6373] = i[6373];
  assign o[6372] = i[6372];
  assign o[6371] = i[6371];
  assign o[6370] = i[6370];
  assign o[6369] = i[6369];
  assign o[6368] = i[6368];
  assign o[6367] = i[6367];
  assign o[6366] = i[6366];
  assign o[6365] = i[6365];
  assign o[6364] = i[6364];
  assign o[6363] = i[6363];
  assign o[6362] = i[6362];
  assign o[6361] = i[6361];
  assign o[6360] = i[6360];
  assign o[6359] = i[6359];
  assign o[6358] = i[6358];
  assign o[6357] = i[6357];
  assign o[6356] = i[6356];
  assign o[6355] = i[6355];
  assign o[6354] = i[6354];
  assign o[6353] = i[6353];
  assign o[6352] = i[6352];
  assign o[6351] = i[6351];
  assign o[6350] = i[6350];
  assign o[6349] = i[6349];
  assign o[6348] = i[6348];
  assign o[6347] = i[6347];
  assign o[6346] = i[6346];
  assign o[6345] = i[6345];
  assign o[6344] = i[6344];
  assign o[6343] = i[6343];
  assign o[6342] = i[6342];
  assign o[6341] = i[6341];
  assign o[6340] = i[6340];
  assign o[6339] = i[6339];
  assign o[6338] = i[6338];
  assign o[6337] = i[6337];
  assign o[6336] = i[6336];
  assign o[6335] = i[6335];
  assign o[6334] = i[6334];
  assign o[6333] = i[6333];
  assign o[6332] = i[6332];
  assign o[6331] = i[6331];
  assign o[6330] = i[6330];
  assign o[6329] = i[6329];
  assign o[6328] = i[6328];
  assign o[6327] = i[6327];
  assign o[6326] = i[6326];
  assign o[6325] = i[6325];
  assign o[6324] = i[6324];
  assign o[6323] = i[6323];
  assign o[6322] = i[6322];
  assign o[6321] = i[6321];
  assign o[6320] = i[6320];
  assign o[6319] = i[6319];
  assign o[6318] = i[6318];
  assign o[6317] = i[6317];
  assign o[6316] = i[6316];
  assign o[6315] = i[6315];
  assign o[6314] = i[6314];
  assign o[6313] = i[6313];
  assign o[6312] = i[6312];
  assign o[6311] = i[6311];
  assign o[6310] = i[6310];
  assign o[6309] = i[6309];
  assign o[6308] = i[6308];
  assign o[6307] = i[6307];
  assign o[6306] = i[6306];
  assign o[6305] = i[6305];
  assign o[6304] = i[6304];
  assign o[6303] = i[6303];
  assign o[6302] = i[6302];
  assign o[6301] = i[6301];
  assign o[6300] = i[6300];
  assign o[6299] = i[6299];
  assign o[6298] = i[6298];
  assign o[6297] = i[6297];
  assign o[6296] = i[6296];
  assign o[6295] = i[6295];
  assign o[6294] = i[6294];
  assign o[6293] = i[6293];
  assign o[6292] = i[6292];
  assign o[6291] = i[6291];
  assign o[6290] = i[6290];
  assign o[6289] = i[6289];
  assign o[6288] = i[6288];
  assign o[6287] = i[6287];
  assign o[6286] = i[6286];
  assign o[6285] = i[6285];
  assign o[6284] = i[6284];
  assign o[6283] = i[6283];
  assign o[6282] = i[6282];
  assign o[6281] = i[6281];
  assign o[6280] = i[6280];
  assign o[6279] = i[6279];
  assign o[6278] = i[6278];
  assign o[6277] = i[6277];
  assign o[6276] = i[6276];
  assign o[6275] = i[6275];
  assign o[6274] = i[6274];
  assign o[6273] = i[6273];
  assign o[6272] = i[6272];
  assign o[6271] = i[6271];
  assign o[6270] = i[6270];
  assign o[6269] = i[6269];
  assign o[6268] = i[6268];
  assign o[6267] = i[6267];
  assign o[6266] = i[6266];
  assign o[6265] = i[6265];
  assign o[6264] = i[6264];
  assign o[6263] = i[6263];
  assign o[6262] = i[6262];
  assign o[6261] = i[6261];
  assign o[6260] = i[6260];
  assign o[6259] = i[6259];
  assign o[6258] = i[6258];
  assign o[6257] = i[6257];
  assign o[6256] = i[6256];
  assign o[6255] = i[6255];
  assign o[6254] = i[6254];
  assign o[6253] = i[6253];
  assign o[6252] = i[6252];
  assign o[6251] = i[6251];
  assign o[6250] = i[6250];
  assign o[6249] = i[6249];
  assign o[6248] = i[6248];
  assign o[6247] = i[6247];
  assign o[6246] = i[6246];
  assign o[6245] = i[6245];
  assign o[6244] = i[6244];
  assign o[6243] = i[6243];
  assign o[6242] = i[6242];
  assign o[6241] = i[6241];
  assign o[6240] = i[6240];
  assign o[6239] = i[6239];
  assign o[6238] = i[6238];
  assign o[6237] = i[6237];
  assign o[6236] = i[6236];
  assign o[6235] = i[6235];
  assign o[6234] = i[6234];
  assign o[6233] = i[6233];
  assign o[6232] = i[6232];
  assign o[6231] = i[6231];
  assign o[6230] = i[6230];
  assign o[6229] = i[6229];
  assign o[6228] = i[6228];
  assign o[6227] = i[6227];
  assign o[6226] = i[6226];
  assign o[6225] = i[6225];
  assign o[6224] = i[6224];
  assign o[6223] = i[6223];
  assign o[6222] = i[6222];
  assign o[6221] = i[6221];
  assign o[6220] = i[6220];
  assign o[6219] = i[6219];
  assign o[6218] = i[6218];
  assign o[6217] = i[6217];
  assign o[6216] = i[6216];
  assign o[6215] = i[6215];
  assign o[6214] = i[6214];
  assign o[6213] = i[6213];
  assign o[6212] = i[6212];
  assign o[6211] = i[6211];
  assign o[6210] = i[6210];
  assign o[6209] = i[6209];
  assign o[6208] = i[6208];
  assign o[6207] = i[6207];
  assign o[6206] = i[6206];
  assign o[6205] = i[6205];
  assign o[6204] = i[6204];
  assign o[6203] = i[6203];
  assign o[6202] = i[6202];
  assign o[6201] = i[6201];
  assign o[6200] = i[6200];
  assign o[6199] = i[6199];
  assign o[6198] = i[6198];
  assign o[6197] = i[6197];
  assign o[6196] = i[6196];
  assign o[6195] = i[6195];
  assign o[6194] = i[6194];
  assign o[6193] = i[6193];
  assign o[6192] = i[6192];
  assign o[6191] = i[6191];
  assign o[6190] = i[6190];
  assign o[6189] = i[6189];
  assign o[6188] = i[6188];
  assign o[6187] = i[6187];
  assign o[6186] = i[6186];
  assign o[6185] = i[6185];
  assign o[6184] = i[6184];
  assign o[6183] = i[6183];
  assign o[6182] = i[6182];
  assign o[6181] = i[6181];
  assign o[6180] = i[6180];
  assign o[6179] = i[6179];
  assign o[6178] = i[6178];
  assign o[6177] = i[6177];
  assign o[6176] = i[6176];
  assign o[6175] = i[6175];
  assign o[6174] = i[6174];
  assign o[6173] = i[6173];
  assign o[6172] = i[6172];
  assign o[6171] = i[6171];
  assign o[6170] = i[6170];
  assign o[6169] = i[6169];
  assign o[6168] = i[6168];
  assign o[6167] = i[6167];
  assign o[6166] = i[6166];
  assign o[6165] = i[6165];
  assign o[6164] = i[6164];
  assign o[6163] = i[6163];
  assign o[6162] = i[6162];
  assign o[6161] = i[6161];
  assign o[6160] = i[6160];
  assign o[6159] = i[6159];
  assign o[6158] = i[6158];
  assign o[6157] = i[6157];
  assign o[6156] = i[6156];
  assign o[6155] = i[6155];
  assign o[6154] = i[6154];
  assign o[6153] = i[6153];
  assign o[6152] = i[6152];
  assign o[6151] = i[6151];
  assign o[6150] = i[6150];
  assign o[6149] = i[6149];
  assign o[6148] = i[6148];
  assign o[6147] = i[6147];
  assign o[6146] = i[6146];
  assign o[6145] = i[6145];
  assign o[6144] = i[6144];
  assign o[6143] = i[6143];
  assign o[6142] = i[6142];
  assign o[6141] = i[6141];
  assign o[6140] = i[6140];
  assign o[6139] = i[6139];
  assign o[6138] = i[6138];
  assign o[6137] = i[6137];
  assign o[6136] = i[6136];
  assign o[6135] = i[6135];
  assign o[6134] = i[6134];
  assign o[6133] = i[6133];
  assign o[6132] = i[6132];
  assign o[6131] = i[6131];
  assign o[6130] = i[6130];
  assign o[6129] = i[6129];
  assign o[6128] = i[6128];
  assign o[6127] = i[6127];
  assign o[6126] = i[6126];
  assign o[6125] = i[6125];
  assign o[6124] = i[6124];
  assign o[6123] = i[6123];
  assign o[6122] = i[6122];
  assign o[6121] = i[6121];
  assign o[6120] = i[6120];
  assign o[6119] = i[6119];
  assign o[6118] = i[6118];
  assign o[6117] = i[6117];
  assign o[6116] = i[6116];
  assign o[6115] = i[6115];
  assign o[6114] = i[6114];
  assign o[6113] = i[6113];
  assign o[6112] = i[6112];
  assign o[6111] = i[6111];
  assign o[6110] = i[6110];
  assign o[6109] = i[6109];
  assign o[6108] = i[6108];
  assign o[6107] = i[6107];
  assign o[6106] = i[6106];
  assign o[6105] = i[6105];
  assign o[6104] = i[6104];
  assign o[6103] = i[6103];
  assign o[6102] = i[6102];
  assign o[6101] = i[6101];
  assign o[6100] = i[6100];
  assign o[6099] = i[6099];
  assign o[6098] = i[6098];
  assign o[6097] = i[6097];
  assign o[6096] = i[6096];
  assign o[6095] = i[6095];
  assign o[6094] = i[6094];
  assign o[6093] = i[6093];
  assign o[6092] = i[6092];
  assign o[6091] = i[6091];
  assign o[6090] = i[6090];
  assign o[6089] = i[6089];
  assign o[6088] = i[6088];
  assign o[6087] = i[6087];
  assign o[6086] = i[6086];
  assign o[6085] = i[6085];
  assign o[6084] = i[6084];
  assign o[6083] = i[6083];
  assign o[6082] = i[6082];
  assign o[6081] = i[6081];
  assign o[6080] = i[6080];
  assign o[6079] = i[6079];
  assign o[6078] = i[6078];
  assign o[6077] = i[6077];
  assign o[6076] = i[6076];
  assign o[6075] = i[6075];
  assign o[6074] = i[6074];
  assign o[6073] = i[6073];
  assign o[6072] = i[6072];
  assign o[6071] = i[6071];
  assign o[6070] = i[6070];
  assign o[6069] = i[6069];
  assign o[6068] = i[6068];
  assign o[6067] = i[6067];
  assign o[6066] = i[6066];
  assign o[6065] = i[6065];
  assign o[6064] = i[6064];
  assign o[6063] = i[6063];
  assign o[6062] = i[6062];
  assign o[6061] = i[6061];
  assign o[6060] = i[6060];
  assign o[6059] = i[6059];
  assign o[6058] = i[6058];
  assign o[6057] = i[6057];
  assign o[6056] = i[6056];
  assign o[6055] = i[6055];
  assign o[6054] = i[6054];
  assign o[6053] = i[6053];
  assign o[6052] = i[6052];
  assign o[6051] = i[6051];
  assign o[6050] = i[6050];
  assign o[6049] = i[6049];
  assign o[6048] = i[6048];
  assign o[6047] = i[6047];
  assign o[6046] = i[6046];
  assign o[6045] = i[6045];
  assign o[6044] = i[6044];
  assign o[6043] = i[6043];
  assign o[6042] = i[6042];
  assign o[6041] = i[6041];
  assign o[6040] = i[6040];
  assign o[6039] = i[6039];
  assign o[6038] = i[6038];
  assign o[6037] = i[6037];
  assign o[6036] = i[6036];
  assign o[6035] = i[6035];
  assign o[6034] = i[6034];
  assign o[6033] = i[6033];
  assign o[6032] = i[6032];
  assign o[6031] = i[6031];
  assign o[6030] = i[6030];
  assign o[6029] = i[6029];
  assign o[6028] = i[6028];
  assign o[6027] = i[6027];
  assign o[6026] = i[6026];
  assign o[6025] = i[6025];
  assign o[6024] = i[6024];
  assign o[6023] = i[6023];
  assign o[6022] = i[6022];
  assign o[6021] = i[6021];
  assign o[6020] = i[6020];
  assign o[6019] = i[6019];
  assign o[6018] = i[6018];
  assign o[6017] = i[6017];
  assign o[6016] = i[6016];
  assign o[6015] = i[6015];
  assign o[6014] = i[6014];
  assign o[6013] = i[6013];
  assign o[6012] = i[6012];
  assign o[6011] = i[6011];
  assign o[6010] = i[6010];
  assign o[6009] = i[6009];
  assign o[6008] = i[6008];
  assign o[6007] = i[6007];
  assign o[6006] = i[6006];
  assign o[6005] = i[6005];
  assign o[6004] = i[6004];
  assign o[6003] = i[6003];
  assign o[6002] = i[6002];
  assign o[6001] = i[6001];
  assign o[6000] = i[6000];
  assign o[5999] = i[5999];
  assign o[5998] = i[5998];
  assign o[5997] = i[5997];
  assign o[5996] = i[5996];
  assign o[5995] = i[5995];
  assign o[5994] = i[5994];
  assign o[5993] = i[5993];
  assign o[5992] = i[5992];
  assign o[5991] = i[5991];
  assign o[5990] = i[5990];
  assign o[5989] = i[5989];
  assign o[5988] = i[5988];
  assign o[5987] = i[5987];
  assign o[5986] = i[5986];
  assign o[5985] = i[5985];
  assign o[5984] = i[5984];
  assign o[5983] = i[5983];
  assign o[5982] = i[5982];
  assign o[5981] = i[5981];
  assign o[5980] = i[5980];
  assign o[5979] = i[5979];
  assign o[5978] = i[5978];
  assign o[5977] = i[5977];
  assign o[5976] = i[5976];
  assign o[5975] = i[5975];
  assign o[5974] = i[5974];
  assign o[5973] = i[5973];
  assign o[5972] = i[5972];
  assign o[5971] = i[5971];
  assign o[5970] = i[5970];
  assign o[5969] = i[5969];
  assign o[5968] = i[5968];
  assign o[5967] = i[5967];
  assign o[5966] = i[5966];
  assign o[5965] = i[5965];
  assign o[5964] = i[5964];
  assign o[5963] = i[5963];
  assign o[5962] = i[5962];
  assign o[5961] = i[5961];
  assign o[5960] = i[5960];
  assign o[5959] = i[5959];
  assign o[5958] = i[5958];
  assign o[5957] = i[5957];
  assign o[5956] = i[5956];
  assign o[5955] = i[5955];
  assign o[5954] = i[5954];
  assign o[5953] = i[5953];
  assign o[5952] = i[5952];
  assign o[5951] = i[5951];
  assign o[5950] = i[5950];
  assign o[5949] = i[5949];
  assign o[5948] = i[5948];
  assign o[5947] = i[5947];
  assign o[5946] = i[5946];
  assign o[5945] = i[5945];
  assign o[5944] = i[5944];
  assign o[5943] = i[5943];
  assign o[5942] = i[5942];
  assign o[5941] = i[5941];
  assign o[5940] = i[5940];
  assign o[5939] = i[5939];
  assign o[5938] = i[5938];
  assign o[5937] = i[5937];
  assign o[5936] = i[5936];
  assign o[5935] = i[5935];
  assign o[5934] = i[5934];
  assign o[5933] = i[5933];
  assign o[5932] = i[5932];
  assign o[5931] = i[5931];
  assign o[5930] = i[5930];
  assign o[5929] = i[5929];
  assign o[5928] = i[5928];
  assign o[5927] = i[5927];
  assign o[5926] = i[5926];
  assign o[5925] = i[5925];
  assign o[5924] = i[5924];
  assign o[5923] = i[5923];
  assign o[5922] = i[5922];
  assign o[5921] = i[5921];
  assign o[5920] = i[5920];
  assign o[5919] = i[5919];
  assign o[5918] = i[5918];
  assign o[5917] = i[5917];
  assign o[5916] = i[5916];
  assign o[5915] = i[5915];
  assign o[5914] = i[5914];
  assign o[5913] = i[5913];
  assign o[5912] = i[5912];
  assign o[5911] = i[5911];
  assign o[5910] = i[5910];
  assign o[5909] = i[5909];
  assign o[5908] = i[5908];
  assign o[5907] = i[5907];
  assign o[5906] = i[5906];
  assign o[5905] = i[5905];
  assign o[5904] = i[5904];
  assign o[5903] = i[5903];
  assign o[5902] = i[5902];
  assign o[5901] = i[5901];
  assign o[5900] = i[5900];
  assign o[5899] = i[5899];
  assign o[5898] = i[5898];
  assign o[5897] = i[5897];
  assign o[5896] = i[5896];
  assign o[5895] = i[5895];
  assign o[5894] = i[5894];
  assign o[5893] = i[5893];
  assign o[5892] = i[5892];
  assign o[5891] = i[5891];
  assign o[5890] = i[5890];
  assign o[5889] = i[5889];
  assign o[5888] = i[5888];
  assign o[5887] = i[5887];
  assign o[5886] = i[5886];
  assign o[5885] = i[5885];
  assign o[5884] = i[5884];
  assign o[5883] = i[5883];
  assign o[5882] = i[5882];
  assign o[5881] = i[5881];
  assign o[5880] = i[5880];
  assign o[5879] = i[5879];
  assign o[5878] = i[5878];
  assign o[5877] = i[5877];
  assign o[5876] = i[5876];
  assign o[5875] = i[5875];
  assign o[5874] = i[5874];
  assign o[5873] = i[5873];
  assign o[5872] = i[5872];
  assign o[5871] = i[5871];
  assign o[5870] = i[5870];
  assign o[5869] = i[5869];
  assign o[5868] = i[5868];
  assign o[5867] = i[5867];
  assign o[5866] = i[5866];
  assign o[5865] = i[5865];
  assign o[5864] = i[5864];
  assign o[5863] = i[5863];
  assign o[5862] = i[5862];
  assign o[5861] = i[5861];
  assign o[5860] = i[5860];
  assign o[5859] = i[5859];
  assign o[5858] = i[5858];
  assign o[5857] = i[5857];
  assign o[5856] = i[5856];
  assign o[5855] = i[5855];
  assign o[5854] = i[5854];
  assign o[5853] = i[5853];
  assign o[5852] = i[5852];
  assign o[5851] = i[5851];
  assign o[5850] = i[5850];
  assign o[5849] = i[5849];
  assign o[5848] = i[5848];
  assign o[5847] = i[5847];
  assign o[5846] = i[5846];
  assign o[5845] = i[5845];
  assign o[5844] = i[5844];
  assign o[5843] = i[5843];
  assign o[5842] = i[5842];
  assign o[5841] = i[5841];
  assign o[5840] = i[5840];
  assign o[5839] = i[5839];
  assign o[5838] = i[5838];
  assign o[5837] = i[5837];
  assign o[5836] = i[5836];
  assign o[5835] = i[5835];
  assign o[5834] = i[5834];
  assign o[5833] = i[5833];
  assign o[5832] = i[5832];
  assign o[5831] = i[5831];
  assign o[5830] = i[5830];
  assign o[5829] = i[5829];
  assign o[5828] = i[5828];
  assign o[5827] = i[5827];
  assign o[5826] = i[5826];
  assign o[5825] = i[5825];
  assign o[5824] = i[5824];
  assign o[5823] = i[5823];
  assign o[5822] = i[5822];
  assign o[5821] = i[5821];
  assign o[5820] = i[5820];
  assign o[5819] = i[5819];
  assign o[5818] = i[5818];
  assign o[5817] = i[5817];
  assign o[5816] = i[5816];
  assign o[5815] = i[5815];
  assign o[5814] = i[5814];
  assign o[5813] = i[5813];
  assign o[5812] = i[5812];
  assign o[5811] = i[5811];
  assign o[5810] = i[5810];
  assign o[5809] = i[5809];
  assign o[5808] = i[5808];
  assign o[5807] = i[5807];
  assign o[5806] = i[5806];
  assign o[5805] = i[5805];
  assign o[5804] = i[5804];
  assign o[5803] = i[5803];
  assign o[5802] = i[5802];
  assign o[5801] = i[5801];
  assign o[5800] = i[5800];
  assign o[5799] = i[5799];
  assign o[5798] = i[5798];
  assign o[5797] = i[5797];
  assign o[5796] = i[5796];
  assign o[5795] = i[5795];
  assign o[5794] = i[5794];
  assign o[5793] = i[5793];
  assign o[5792] = i[5792];
  assign o[5791] = i[5791];
  assign o[5790] = i[5790];
  assign o[5789] = i[5789];
  assign o[5788] = i[5788];
  assign o[5787] = i[5787];
  assign o[5786] = i[5786];
  assign o[5785] = i[5785];
  assign o[5784] = i[5784];
  assign o[5783] = i[5783];
  assign o[5782] = i[5782];
  assign o[5781] = i[5781];
  assign o[5780] = i[5780];
  assign o[5779] = i[5779];
  assign o[5778] = i[5778];
  assign o[5777] = i[5777];
  assign o[5776] = i[5776];
  assign o[5775] = i[5775];
  assign o[5774] = i[5774];
  assign o[5773] = i[5773];
  assign o[5772] = i[5772];
  assign o[5771] = i[5771];
  assign o[5770] = i[5770];
  assign o[5769] = i[5769];
  assign o[5768] = i[5768];
  assign o[5767] = i[5767];
  assign o[5766] = i[5766];
  assign o[5765] = i[5765];
  assign o[5764] = i[5764];
  assign o[5763] = i[5763];
  assign o[5762] = i[5762];
  assign o[5761] = i[5761];
  assign o[5760] = i[5760];
  assign o[5759] = i[5759];
  assign o[5758] = i[5758];
  assign o[5757] = i[5757];
  assign o[5756] = i[5756];
  assign o[5755] = i[5755];
  assign o[5754] = i[5754];
  assign o[5753] = i[5753];
  assign o[5752] = i[5752];
  assign o[5751] = i[5751];
  assign o[5750] = i[5750];
  assign o[5749] = i[5749];
  assign o[5748] = i[5748];
  assign o[5747] = i[5747];
  assign o[5746] = i[5746];
  assign o[5745] = i[5745];
  assign o[5744] = i[5744];
  assign o[5743] = i[5743];
  assign o[5742] = i[5742];
  assign o[5741] = i[5741];
  assign o[5740] = i[5740];
  assign o[5739] = i[5739];
  assign o[5738] = i[5738];
  assign o[5737] = i[5737];
  assign o[5736] = i[5736];
  assign o[5735] = i[5735];
  assign o[5734] = i[5734];
  assign o[5733] = i[5733];
  assign o[5732] = i[5732];
  assign o[5731] = i[5731];
  assign o[5730] = i[5730];
  assign o[5729] = i[5729];
  assign o[5728] = i[5728];
  assign o[5727] = i[5727];
  assign o[5726] = i[5726];
  assign o[5725] = i[5725];
  assign o[5724] = i[5724];
  assign o[5723] = i[5723];
  assign o[5722] = i[5722];
  assign o[5721] = i[5721];
  assign o[5720] = i[5720];
  assign o[5719] = i[5719];
  assign o[5718] = i[5718];
  assign o[5717] = i[5717];
  assign o[5716] = i[5716];
  assign o[5715] = i[5715];
  assign o[5714] = i[5714];
  assign o[5713] = i[5713];
  assign o[5712] = i[5712];
  assign o[5711] = i[5711];
  assign o[5710] = i[5710];
  assign o[5709] = i[5709];
  assign o[5708] = i[5708];
  assign o[5707] = i[5707];
  assign o[5706] = i[5706];
  assign o[5705] = i[5705];
  assign o[5704] = i[5704];
  assign o[5703] = i[5703];
  assign o[5702] = i[5702];
  assign o[5701] = i[5701];
  assign o[5700] = i[5700];
  assign o[5699] = i[5699];
  assign o[5698] = i[5698];
  assign o[5697] = i[5697];
  assign o[5696] = i[5696];
  assign o[5695] = i[5695];
  assign o[5694] = i[5694];
  assign o[5693] = i[5693];
  assign o[5692] = i[5692];
  assign o[5691] = i[5691];
  assign o[5690] = i[5690];
  assign o[5689] = i[5689];
  assign o[5688] = i[5688];
  assign o[5687] = i[5687];
  assign o[5686] = i[5686];
  assign o[5685] = i[5685];
  assign o[5684] = i[5684];
  assign o[5683] = i[5683];
  assign o[5682] = i[5682];
  assign o[5681] = i[5681];
  assign o[5680] = i[5680];
  assign o[5679] = i[5679];
  assign o[5678] = i[5678];
  assign o[5677] = i[5677];
  assign o[5676] = i[5676];
  assign o[5675] = i[5675];
  assign o[5674] = i[5674];
  assign o[5673] = i[5673];
  assign o[5672] = i[5672];
  assign o[5671] = i[5671];
  assign o[5670] = i[5670];
  assign o[5669] = i[5669];
  assign o[5668] = i[5668];
  assign o[5667] = i[5667];
  assign o[5666] = i[5666];
  assign o[5665] = i[5665];
  assign o[5664] = i[5664];
  assign o[5663] = i[5663];
  assign o[5662] = i[5662];
  assign o[5661] = i[5661];
  assign o[5660] = i[5660];
  assign o[5659] = i[5659];
  assign o[5658] = i[5658];
  assign o[5657] = i[5657];
  assign o[5656] = i[5656];
  assign o[5655] = i[5655];
  assign o[5654] = i[5654];
  assign o[5653] = i[5653];
  assign o[5652] = i[5652];
  assign o[5651] = i[5651];
  assign o[5650] = i[5650];
  assign o[5649] = i[5649];
  assign o[5648] = i[5648];
  assign o[5647] = i[5647];
  assign o[5646] = i[5646];
  assign o[5645] = i[5645];
  assign o[5644] = i[5644];
  assign o[5643] = i[5643];
  assign o[5642] = i[5642];
  assign o[5641] = i[5641];
  assign o[5640] = i[5640];
  assign o[5639] = i[5639];
  assign o[5638] = i[5638];
  assign o[5637] = i[5637];
  assign o[5636] = i[5636];
  assign o[5635] = i[5635];
  assign o[5634] = i[5634];
  assign o[5633] = i[5633];
  assign o[5632] = i[5632];
  assign o[5631] = i[5631];
  assign o[5630] = i[5630];
  assign o[5629] = i[5629];
  assign o[5628] = i[5628];
  assign o[5627] = i[5627];
  assign o[5626] = i[5626];
  assign o[5625] = i[5625];
  assign o[5624] = i[5624];
  assign o[5623] = i[5623];
  assign o[5622] = i[5622];
  assign o[5621] = i[5621];
  assign o[5620] = i[5620];
  assign o[5619] = i[5619];
  assign o[5618] = i[5618];
  assign o[5617] = i[5617];
  assign o[5616] = i[5616];
  assign o[5615] = i[5615];
  assign o[5614] = i[5614];
  assign o[5613] = i[5613];
  assign o[5612] = i[5612];
  assign o[5611] = i[5611];
  assign o[5610] = i[5610];
  assign o[5609] = i[5609];
  assign o[5608] = i[5608];
  assign o[5607] = i[5607];
  assign o[5606] = i[5606];
  assign o[5605] = i[5605];
  assign o[5604] = i[5604];
  assign o[5603] = i[5603];
  assign o[5602] = i[5602];
  assign o[5601] = i[5601];
  assign o[5600] = i[5600];
  assign o[5599] = i[5599];
  assign o[5598] = i[5598];
  assign o[5597] = i[5597];
  assign o[5596] = i[5596];
  assign o[5595] = i[5595];
  assign o[5594] = i[5594];
  assign o[5593] = i[5593];
  assign o[5592] = i[5592];
  assign o[5591] = i[5591];
  assign o[5590] = i[5590];
  assign o[5589] = i[5589];
  assign o[5588] = i[5588];
  assign o[5587] = i[5587];
  assign o[5586] = i[5586];
  assign o[5585] = i[5585];
  assign o[5584] = i[5584];
  assign o[5583] = i[5583];
  assign o[5582] = i[5582];
  assign o[5581] = i[5581];
  assign o[5580] = i[5580];
  assign o[5579] = i[5579];
  assign o[5578] = i[5578];
  assign o[5577] = i[5577];
  assign o[5576] = i[5576];
  assign o[5575] = i[5575];
  assign o[5574] = i[5574];
  assign o[5573] = i[5573];
  assign o[5572] = i[5572];
  assign o[5571] = i[5571];
  assign o[5570] = i[5570];
  assign o[5569] = i[5569];
  assign o[5568] = i[5568];
  assign o[5567] = i[5567];
  assign o[5566] = i[5566];
  assign o[5565] = i[5565];
  assign o[5564] = i[5564];
  assign o[5563] = i[5563];
  assign o[5562] = i[5562];
  assign o[5561] = i[5561];
  assign o[5560] = i[5560];
  assign o[5559] = i[5559];
  assign o[5558] = i[5558];
  assign o[5557] = i[5557];
  assign o[5556] = i[5556];
  assign o[5555] = i[5555];
  assign o[5554] = i[5554];
  assign o[5553] = i[5553];
  assign o[5552] = i[5552];
  assign o[5551] = i[5551];
  assign o[5550] = i[5550];
  assign o[5549] = i[5549];
  assign o[5548] = i[5548];
  assign o[5547] = i[5547];
  assign o[5546] = i[5546];
  assign o[5545] = i[5545];
  assign o[5544] = i[5544];
  assign o[5543] = i[5543];
  assign o[5542] = i[5542];
  assign o[5541] = i[5541];
  assign o[5540] = i[5540];
  assign o[5539] = i[5539];
  assign o[5538] = i[5538];
  assign o[5537] = i[5537];
  assign o[5536] = i[5536];
  assign o[5535] = i[5535];
  assign o[5534] = i[5534];
  assign o[5533] = i[5533];
  assign o[5532] = i[5532];
  assign o[5531] = i[5531];
  assign o[5530] = i[5530];
  assign o[5529] = i[5529];
  assign o[5528] = i[5528];
  assign o[5527] = i[5527];
  assign o[5526] = i[5526];
  assign o[5525] = i[5525];
  assign o[5524] = i[5524];
  assign o[5523] = i[5523];
  assign o[5522] = i[5522];
  assign o[5521] = i[5521];
  assign o[5520] = i[5520];
  assign o[5519] = i[5519];
  assign o[5518] = i[5518];
  assign o[5517] = i[5517];
  assign o[5516] = i[5516];
  assign o[5515] = i[5515];
  assign o[5514] = i[5514];
  assign o[5513] = i[5513];
  assign o[5512] = i[5512];
  assign o[5511] = i[5511];
  assign o[5510] = i[5510];
  assign o[5509] = i[5509];
  assign o[5508] = i[5508];
  assign o[5507] = i[5507];
  assign o[5506] = i[5506];
  assign o[5505] = i[5505];
  assign o[5504] = i[5504];
  assign o[5503] = i[5503];
  assign o[5502] = i[5502];
  assign o[5501] = i[5501];
  assign o[5500] = i[5500];
  assign o[5499] = i[5499];
  assign o[5498] = i[5498];
  assign o[5497] = i[5497];
  assign o[5496] = i[5496];
  assign o[5495] = i[5495];
  assign o[5494] = i[5494];
  assign o[5493] = i[5493];
  assign o[5492] = i[5492];
  assign o[5491] = i[5491];
  assign o[5490] = i[5490];
  assign o[5489] = i[5489];
  assign o[5488] = i[5488];
  assign o[5487] = i[5487];
  assign o[5486] = i[5486];
  assign o[5485] = i[5485];
  assign o[5484] = i[5484];
  assign o[5483] = i[5483];
  assign o[5482] = i[5482];
  assign o[5481] = i[5481];
  assign o[5480] = i[5480];
  assign o[5479] = i[5479];
  assign o[5478] = i[5478];
  assign o[5477] = i[5477];
  assign o[5476] = i[5476];
  assign o[5475] = i[5475];
  assign o[5474] = i[5474];
  assign o[5473] = i[5473];
  assign o[5472] = i[5472];
  assign o[5471] = i[5471];
  assign o[5470] = i[5470];
  assign o[5469] = i[5469];
  assign o[5468] = i[5468];
  assign o[5467] = i[5467];
  assign o[5466] = i[5466];
  assign o[5465] = i[5465];
  assign o[5464] = i[5464];
  assign o[5463] = i[5463];
  assign o[5462] = i[5462];
  assign o[5461] = i[5461];
  assign o[5460] = i[5460];
  assign o[5459] = i[5459];
  assign o[5458] = i[5458];
  assign o[5457] = i[5457];
  assign o[5456] = i[5456];
  assign o[5455] = i[5455];
  assign o[5454] = i[5454];
  assign o[5453] = i[5453];
  assign o[5452] = i[5452];
  assign o[5451] = i[5451];
  assign o[5450] = i[5450];
  assign o[5449] = i[5449];
  assign o[5448] = i[5448];
  assign o[5447] = i[5447];
  assign o[5446] = i[5446];
  assign o[5445] = i[5445];
  assign o[5444] = i[5444];
  assign o[5443] = i[5443];
  assign o[5442] = i[5442];
  assign o[5441] = i[5441];
  assign o[5440] = i[5440];
  assign o[5439] = i[5439];
  assign o[5438] = i[5438];
  assign o[5437] = i[5437];
  assign o[5436] = i[5436];
  assign o[5435] = i[5435];
  assign o[5434] = i[5434];
  assign o[5433] = i[5433];
  assign o[5432] = i[5432];
  assign o[5431] = i[5431];
  assign o[5430] = i[5430];
  assign o[5429] = i[5429];
  assign o[5428] = i[5428];
  assign o[5427] = i[5427];
  assign o[5426] = i[5426];
  assign o[5425] = i[5425];
  assign o[5424] = i[5424];
  assign o[5423] = i[5423];
  assign o[5422] = i[5422];
  assign o[5421] = i[5421];
  assign o[5420] = i[5420];
  assign o[5419] = i[5419];
  assign o[5418] = i[5418];
  assign o[5417] = i[5417];
  assign o[5416] = i[5416];
  assign o[5415] = i[5415];
  assign o[5414] = i[5414];
  assign o[5413] = i[5413];
  assign o[5412] = i[5412];
  assign o[5411] = i[5411];
  assign o[5410] = i[5410];
  assign o[5409] = i[5409];
  assign o[5408] = i[5408];
  assign o[5407] = i[5407];
  assign o[5406] = i[5406];
  assign o[5405] = i[5405];
  assign o[5404] = i[5404];
  assign o[5403] = i[5403];
  assign o[5402] = i[5402];
  assign o[5401] = i[5401];
  assign o[5400] = i[5400];
  assign o[5399] = i[5399];
  assign o[5398] = i[5398];
  assign o[5397] = i[5397];
  assign o[5396] = i[5396];
  assign o[5395] = i[5395];
  assign o[5394] = i[5394];
  assign o[5393] = i[5393];
  assign o[5392] = i[5392];
  assign o[5391] = i[5391];
  assign o[5390] = i[5390];
  assign o[5389] = i[5389];
  assign o[5388] = i[5388];
  assign o[5387] = i[5387];
  assign o[5386] = i[5386];
  assign o[5385] = i[5385];
  assign o[5384] = i[5384];
  assign o[5383] = i[5383];
  assign o[5382] = i[5382];
  assign o[5381] = i[5381];
  assign o[5380] = i[5380];
  assign o[5379] = i[5379];
  assign o[5378] = i[5378];
  assign o[5377] = i[5377];
  assign o[5376] = i[5376];
  assign o[5375] = i[5375];
  assign o[5374] = i[5374];
  assign o[5373] = i[5373];
  assign o[5372] = i[5372];
  assign o[5371] = i[5371];
  assign o[5370] = i[5370];
  assign o[5369] = i[5369];
  assign o[5368] = i[5368];
  assign o[5367] = i[5367];
  assign o[5366] = i[5366];
  assign o[5365] = i[5365];
  assign o[5364] = i[5364];
  assign o[5363] = i[5363];
  assign o[5362] = i[5362];
  assign o[5361] = i[5361];
  assign o[5360] = i[5360];
  assign o[5359] = i[5359];
  assign o[5358] = i[5358];
  assign o[5357] = i[5357];
  assign o[5356] = i[5356];
  assign o[5355] = i[5355];
  assign o[5354] = i[5354];
  assign o[5353] = i[5353];
  assign o[5352] = i[5352];
  assign o[5351] = i[5351];
  assign o[5350] = i[5350];
  assign o[5349] = i[5349];
  assign o[5348] = i[5348];
  assign o[5347] = i[5347];
  assign o[5346] = i[5346];
  assign o[5345] = i[5345];
  assign o[5344] = i[5344];
  assign o[5343] = i[5343];
  assign o[5342] = i[5342];
  assign o[5341] = i[5341];
  assign o[5340] = i[5340];
  assign o[5339] = i[5339];
  assign o[5338] = i[5338];
  assign o[5337] = i[5337];
  assign o[5336] = i[5336];
  assign o[5335] = i[5335];
  assign o[5334] = i[5334];
  assign o[5333] = i[5333];
  assign o[5332] = i[5332];
  assign o[5331] = i[5331];
  assign o[5330] = i[5330];
  assign o[5329] = i[5329];
  assign o[5328] = i[5328];
  assign o[5327] = i[5327];
  assign o[5326] = i[5326];
  assign o[5325] = i[5325];
  assign o[5324] = i[5324];
  assign o[5323] = i[5323];
  assign o[5322] = i[5322];
  assign o[5321] = i[5321];
  assign o[5320] = i[5320];
  assign o[5319] = i[5319];
  assign o[5318] = i[5318];
  assign o[5317] = i[5317];
  assign o[5316] = i[5316];
  assign o[5315] = i[5315];
  assign o[5314] = i[5314];
  assign o[5313] = i[5313];
  assign o[5312] = i[5312];
  assign o[5311] = i[5311];
  assign o[5310] = i[5310];
  assign o[5309] = i[5309];
  assign o[5308] = i[5308];
  assign o[5307] = i[5307];
  assign o[5306] = i[5306];
  assign o[5305] = i[5305];
  assign o[5304] = i[5304];
  assign o[5303] = i[5303];
  assign o[5302] = i[5302];
  assign o[5301] = i[5301];
  assign o[5300] = i[5300];
  assign o[5299] = i[5299];
  assign o[5298] = i[5298];
  assign o[5297] = i[5297];
  assign o[5296] = i[5296];
  assign o[5295] = i[5295];
  assign o[5294] = i[5294];
  assign o[5293] = i[5293];
  assign o[5292] = i[5292];
  assign o[5291] = i[5291];
  assign o[5290] = i[5290];
  assign o[5289] = i[5289];
  assign o[5288] = i[5288];
  assign o[5287] = i[5287];
  assign o[5286] = i[5286];
  assign o[5285] = i[5285];
  assign o[5284] = i[5284];
  assign o[5283] = i[5283];
  assign o[5282] = i[5282];
  assign o[5281] = i[5281];
  assign o[5280] = i[5280];
  assign o[5279] = i[5279];
  assign o[5278] = i[5278];
  assign o[5277] = i[5277];
  assign o[5276] = i[5276];
  assign o[5275] = i[5275];
  assign o[5274] = i[5274];
  assign o[5273] = i[5273];
  assign o[5272] = i[5272];
  assign o[5271] = i[5271];
  assign o[5270] = i[5270];
  assign o[5269] = i[5269];
  assign o[5268] = i[5268];
  assign o[5267] = i[5267];
  assign o[5266] = i[5266];
  assign o[5265] = i[5265];
  assign o[5264] = i[5264];
  assign o[5263] = i[5263];
  assign o[5262] = i[5262];
  assign o[5261] = i[5261];
  assign o[5260] = i[5260];
  assign o[5259] = i[5259];
  assign o[5258] = i[5258];
  assign o[5257] = i[5257];
  assign o[5256] = i[5256];
  assign o[5255] = i[5255];
  assign o[5254] = i[5254];
  assign o[5253] = i[5253];
  assign o[5252] = i[5252];
  assign o[5251] = i[5251];
  assign o[5250] = i[5250];
  assign o[5249] = i[5249];
  assign o[5248] = i[5248];
  assign o[5247] = i[5247];
  assign o[5246] = i[5246];
  assign o[5245] = i[5245];
  assign o[5244] = i[5244];
  assign o[5243] = i[5243];
  assign o[5242] = i[5242];
  assign o[5241] = i[5241];
  assign o[5240] = i[5240];
  assign o[5239] = i[5239];
  assign o[5238] = i[5238];
  assign o[5237] = i[5237];
  assign o[5236] = i[5236];
  assign o[5235] = i[5235];
  assign o[5234] = i[5234];
  assign o[5233] = i[5233];
  assign o[5232] = i[5232];
  assign o[5231] = i[5231];
  assign o[5230] = i[5230];
  assign o[5229] = i[5229];
  assign o[5228] = i[5228];
  assign o[5227] = i[5227];
  assign o[5226] = i[5226];
  assign o[5225] = i[5225];
  assign o[5224] = i[5224];
  assign o[5223] = i[5223];
  assign o[5222] = i[5222];
  assign o[5221] = i[5221];
  assign o[5220] = i[5220];
  assign o[5219] = i[5219];
  assign o[5218] = i[5218];
  assign o[5217] = i[5217];
  assign o[5216] = i[5216];
  assign o[5215] = i[5215];
  assign o[5214] = i[5214];
  assign o[5213] = i[5213];
  assign o[5212] = i[5212];
  assign o[5211] = i[5211];
  assign o[5210] = i[5210];
  assign o[5209] = i[5209];
  assign o[5208] = i[5208];
  assign o[5207] = i[5207];
  assign o[5206] = i[5206];
  assign o[5205] = i[5205];
  assign o[5204] = i[5204];
  assign o[5203] = i[5203];
  assign o[5202] = i[5202];
  assign o[5201] = i[5201];
  assign o[5200] = i[5200];
  assign o[5199] = i[5199];
  assign o[5198] = i[5198];
  assign o[5197] = i[5197];
  assign o[5196] = i[5196];
  assign o[5195] = i[5195];
  assign o[5194] = i[5194];
  assign o[5193] = i[5193];
  assign o[5192] = i[5192];
  assign o[5191] = i[5191];
  assign o[5190] = i[5190];
  assign o[5189] = i[5189];
  assign o[5188] = i[5188];
  assign o[5187] = i[5187];
  assign o[5186] = i[5186];
  assign o[5185] = i[5185];
  assign o[5184] = i[5184];
  assign o[5183] = i[5183];
  assign o[5182] = i[5182];
  assign o[5181] = i[5181];
  assign o[5180] = i[5180];
  assign o[5179] = i[5179];
  assign o[5178] = i[5178];
  assign o[5177] = i[5177];
  assign o[5176] = i[5176];
  assign o[5175] = i[5175];
  assign o[5174] = i[5174];
  assign o[5173] = i[5173];
  assign o[5172] = i[5172];
  assign o[5171] = i[5171];
  assign o[5170] = i[5170];
  assign o[5169] = i[5169];
  assign o[5168] = i[5168];
  assign o[5167] = i[5167];
  assign o[5166] = i[5166];
  assign o[5165] = i[5165];
  assign o[5164] = i[5164];
  assign o[5163] = i[5163];
  assign o[5162] = i[5162];
  assign o[5161] = i[5161];
  assign o[5160] = i[5160];
  assign o[5159] = i[5159];
  assign o[5158] = i[5158];
  assign o[5157] = i[5157];
  assign o[5156] = i[5156];
  assign o[5155] = i[5155];
  assign o[5154] = i[5154];
  assign o[5153] = i[5153];
  assign o[5152] = i[5152];
  assign o[5151] = i[5151];
  assign o[5150] = i[5150];
  assign o[5149] = i[5149];
  assign o[5148] = i[5148];
  assign o[5147] = i[5147];
  assign o[5146] = i[5146];
  assign o[5145] = i[5145];
  assign o[5144] = i[5144];
  assign o[5143] = i[5143];
  assign o[5142] = i[5142];
  assign o[5141] = i[5141];
  assign o[5140] = i[5140];
  assign o[5139] = i[5139];
  assign o[5138] = i[5138];
  assign o[5137] = i[5137];
  assign o[5136] = i[5136];
  assign o[5135] = i[5135];
  assign o[5134] = i[5134];
  assign o[5133] = i[5133];
  assign o[5132] = i[5132];
  assign o[5131] = i[5131];
  assign o[5130] = i[5130];
  assign o[5129] = i[5129];
  assign o[5128] = i[5128];
  assign o[5127] = i[5127];
  assign o[5126] = i[5126];
  assign o[5125] = i[5125];
  assign o[5124] = i[5124];
  assign o[5123] = i[5123];
  assign o[5122] = i[5122];
  assign o[5121] = i[5121];
  assign o[5120] = i[5120];
  assign o[5119] = i[5119];
  assign o[5118] = i[5118];
  assign o[5117] = i[5117];
  assign o[5116] = i[5116];
  assign o[5115] = i[5115];
  assign o[5114] = i[5114];
  assign o[5113] = i[5113];
  assign o[5112] = i[5112];
  assign o[5111] = i[5111];
  assign o[5110] = i[5110];
  assign o[5109] = i[5109];
  assign o[5108] = i[5108];
  assign o[5107] = i[5107];
  assign o[5106] = i[5106];
  assign o[5105] = i[5105];
  assign o[5104] = i[5104];
  assign o[5103] = i[5103];
  assign o[5102] = i[5102];
  assign o[5101] = i[5101];
  assign o[5100] = i[5100];
  assign o[5099] = i[5099];
  assign o[5098] = i[5098];
  assign o[5097] = i[5097];
  assign o[5096] = i[5096];
  assign o[5095] = i[5095];
  assign o[5094] = i[5094];
  assign o[5093] = i[5093];
  assign o[5092] = i[5092];
  assign o[5091] = i[5091];
  assign o[5090] = i[5090];
  assign o[5089] = i[5089];
  assign o[5088] = i[5088];
  assign o[5087] = i[5087];
  assign o[5086] = i[5086];
  assign o[5085] = i[5085];
  assign o[5084] = i[5084];
  assign o[5083] = i[5083];
  assign o[5082] = i[5082];
  assign o[5081] = i[5081];
  assign o[5080] = i[5080];
  assign o[5079] = i[5079];
  assign o[5078] = i[5078];
  assign o[5077] = i[5077];
  assign o[5076] = i[5076];
  assign o[5075] = i[5075];
  assign o[5074] = i[5074];
  assign o[5073] = i[5073];
  assign o[5072] = i[5072];
  assign o[5071] = i[5071];
  assign o[5070] = i[5070];
  assign o[5069] = i[5069];
  assign o[5068] = i[5068];
  assign o[5067] = i[5067];
  assign o[5066] = i[5066];
  assign o[5065] = i[5065];
  assign o[5064] = i[5064];
  assign o[5063] = i[5063];
  assign o[5062] = i[5062];
  assign o[5061] = i[5061];
  assign o[5060] = i[5060];
  assign o[5059] = i[5059];
  assign o[5058] = i[5058];
  assign o[5057] = i[5057];
  assign o[5056] = i[5056];
  assign o[5055] = i[5055];
  assign o[5054] = i[5054];
  assign o[5053] = i[5053];
  assign o[5052] = i[5052];
  assign o[5051] = i[5051];
  assign o[5050] = i[5050];
  assign o[5049] = i[5049];
  assign o[5048] = i[5048];
  assign o[5047] = i[5047];
  assign o[5046] = i[5046];
  assign o[5045] = i[5045];
  assign o[5044] = i[5044];
  assign o[5043] = i[5043];
  assign o[5042] = i[5042];
  assign o[5041] = i[5041];
  assign o[5040] = i[5040];
  assign o[5039] = i[5039];
  assign o[5038] = i[5038];
  assign o[5037] = i[5037];
  assign o[5036] = i[5036];
  assign o[5035] = i[5035];
  assign o[5034] = i[5034];
  assign o[5033] = i[5033];
  assign o[5032] = i[5032];
  assign o[5031] = i[5031];
  assign o[5030] = i[5030];
  assign o[5029] = i[5029];
  assign o[5028] = i[5028];
  assign o[5027] = i[5027];
  assign o[5026] = i[5026];
  assign o[5025] = i[5025];
  assign o[5024] = i[5024];
  assign o[5023] = i[5023];
  assign o[5022] = i[5022];
  assign o[5021] = i[5021];
  assign o[5020] = i[5020];
  assign o[5019] = i[5019];
  assign o[5018] = i[5018];
  assign o[5017] = i[5017];
  assign o[5016] = i[5016];
  assign o[5015] = i[5015];
  assign o[5014] = i[5014];
  assign o[5013] = i[5013];
  assign o[5012] = i[5012];
  assign o[5011] = i[5011];
  assign o[5010] = i[5010];
  assign o[5009] = i[5009];
  assign o[5008] = i[5008];
  assign o[5007] = i[5007];
  assign o[5006] = i[5006];
  assign o[5005] = i[5005];
  assign o[5004] = i[5004];
  assign o[5003] = i[5003];
  assign o[5002] = i[5002];
  assign o[5001] = i[5001];
  assign o[5000] = i[5000];
  assign o[4999] = i[4999];
  assign o[4998] = i[4998];
  assign o[4997] = i[4997];
  assign o[4996] = i[4996];
  assign o[4995] = i[4995];
  assign o[4994] = i[4994];
  assign o[4993] = i[4993];
  assign o[4992] = i[4992];
  assign o[4991] = i[4991];
  assign o[4990] = i[4990];
  assign o[4989] = i[4989];
  assign o[4988] = i[4988];
  assign o[4987] = i[4987];
  assign o[4986] = i[4986];
  assign o[4985] = i[4985];
  assign o[4984] = i[4984];
  assign o[4983] = i[4983];
  assign o[4982] = i[4982];
  assign o[4981] = i[4981];
  assign o[4980] = i[4980];
  assign o[4979] = i[4979];
  assign o[4978] = i[4978];
  assign o[4977] = i[4977];
  assign o[4976] = i[4976];
  assign o[4975] = i[4975];
  assign o[4974] = i[4974];
  assign o[4973] = i[4973];
  assign o[4972] = i[4972];
  assign o[4971] = i[4971];
  assign o[4970] = i[4970];
  assign o[4969] = i[4969];
  assign o[4968] = i[4968];
  assign o[4967] = i[4967];
  assign o[4966] = i[4966];
  assign o[4965] = i[4965];
  assign o[4964] = i[4964];
  assign o[4963] = i[4963];
  assign o[4962] = i[4962];
  assign o[4961] = i[4961];
  assign o[4960] = i[4960];
  assign o[4959] = i[4959];
  assign o[4958] = i[4958];
  assign o[4957] = i[4957];
  assign o[4956] = i[4956];
  assign o[4955] = i[4955];
  assign o[4954] = i[4954];
  assign o[4953] = i[4953];
  assign o[4952] = i[4952];
  assign o[4951] = i[4951];
  assign o[4950] = i[4950];
  assign o[4949] = i[4949];
  assign o[4948] = i[4948];
  assign o[4947] = i[4947];
  assign o[4946] = i[4946];
  assign o[4945] = i[4945];
  assign o[4944] = i[4944];
  assign o[4943] = i[4943];
  assign o[4942] = i[4942];
  assign o[4941] = i[4941];
  assign o[4940] = i[4940];
  assign o[4939] = i[4939];
  assign o[4938] = i[4938];
  assign o[4937] = i[4937];
  assign o[4936] = i[4936];
  assign o[4935] = i[4935];
  assign o[4934] = i[4934];
  assign o[4933] = i[4933];
  assign o[4932] = i[4932];
  assign o[4931] = i[4931];
  assign o[4930] = i[4930];
  assign o[4929] = i[4929];
  assign o[4928] = i[4928];
  assign o[4927] = i[4927];
  assign o[4926] = i[4926];
  assign o[4925] = i[4925];
  assign o[4924] = i[4924];
  assign o[4923] = i[4923];
  assign o[4922] = i[4922];
  assign o[4921] = i[4921];
  assign o[4920] = i[4920];
  assign o[4919] = i[4919];
  assign o[4918] = i[4918];
  assign o[4917] = i[4917];
  assign o[4916] = i[4916];
  assign o[4915] = i[4915];
  assign o[4914] = i[4914];
  assign o[4913] = i[4913];
  assign o[4912] = i[4912];
  assign o[4911] = i[4911];
  assign o[4910] = i[4910];
  assign o[4909] = i[4909];
  assign o[4908] = i[4908];
  assign o[4907] = i[4907];
  assign o[4906] = i[4906];
  assign o[4905] = i[4905];
  assign o[4904] = i[4904];
  assign o[4903] = i[4903];
  assign o[4902] = i[4902];
  assign o[4901] = i[4901];
  assign o[4900] = i[4900];
  assign o[4899] = i[4899];
  assign o[4898] = i[4898];
  assign o[4897] = i[4897];
  assign o[4896] = i[4896];
  assign o[4895] = i[4895];
  assign o[4894] = i[4894];
  assign o[4893] = i[4893];
  assign o[4892] = i[4892];
  assign o[4891] = i[4891];
  assign o[4890] = i[4890];
  assign o[4889] = i[4889];
  assign o[4888] = i[4888];
  assign o[4887] = i[4887];
  assign o[4886] = i[4886];
  assign o[4885] = i[4885];
  assign o[4884] = i[4884];
  assign o[4883] = i[4883];
  assign o[4882] = i[4882];
  assign o[4881] = i[4881];
  assign o[4880] = i[4880];
  assign o[4879] = i[4879];
  assign o[4878] = i[4878];
  assign o[4877] = i[4877];
  assign o[4876] = i[4876];
  assign o[4875] = i[4875];
  assign o[4874] = i[4874];
  assign o[4873] = i[4873];
  assign o[4872] = i[4872];
  assign o[4871] = i[4871];
  assign o[4870] = i[4870];
  assign o[4869] = i[4869];
  assign o[4868] = i[4868];
  assign o[4867] = i[4867];
  assign o[4866] = i[4866];
  assign o[4865] = i[4865];
  assign o[4864] = i[4864];
  assign o[4863] = i[4863];
  assign o[4862] = i[4862];
  assign o[4861] = i[4861];
  assign o[4860] = i[4860];
  assign o[4859] = i[4859];
  assign o[4858] = i[4858];
  assign o[4857] = i[4857];
  assign o[4856] = i[4856];
  assign o[4855] = i[4855];
  assign o[4854] = i[4854];
  assign o[4853] = i[4853];
  assign o[4852] = i[4852];
  assign o[4851] = i[4851];
  assign o[4850] = i[4850];
  assign o[4849] = i[4849];
  assign o[4848] = i[4848];
  assign o[4847] = i[4847];
  assign o[4846] = i[4846];
  assign o[4845] = i[4845];
  assign o[4844] = i[4844];
  assign o[4843] = i[4843];
  assign o[4842] = i[4842];
  assign o[4841] = i[4841];
  assign o[4840] = i[4840];
  assign o[4839] = i[4839];
  assign o[4838] = i[4838];
  assign o[4837] = i[4837];
  assign o[4836] = i[4836];
  assign o[4835] = i[4835];
  assign o[4834] = i[4834];
  assign o[4833] = i[4833];
  assign o[4832] = i[4832];
  assign o[4831] = i[4831];
  assign o[4830] = i[4830];
  assign o[4829] = i[4829];
  assign o[4828] = i[4828];
  assign o[4827] = i[4827];
  assign o[4826] = i[4826];
  assign o[4825] = i[4825];
  assign o[4824] = i[4824];
  assign o[4823] = i[4823];
  assign o[4822] = i[4822];
  assign o[4821] = i[4821];
  assign o[4820] = i[4820];
  assign o[4819] = i[4819];
  assign o[4818] = i[4818];
  assign o[4817] = i[4817];
  assign o[4816] = i[4816];
  assign o[4815] = i[4815];
  assign o[4814] = i[4814];
  assign o[4813] = i[4813];
  assign o[4812] = i[4812];
  assign o[4811] = i[4811];
  assign o[4810] = i[4810];
  assign o[4809] = i[4809];
  assign o[4808] = i[4808];
  assign o[4807] = i[4807];
  assign o[4806] = i[4806];
  assign o[4805] = i[4805];
  assign o[4804] = i[4804];
  assign o[4803] = i[4803];
  assign o[4802] = i[4802];
  assign o[4801] = i[4801];
  assign o[4800] = i[4800];
  assign o[4799] = i[4799];
  assign o[4798] = i[4798];
  assign o[4797] = i[4797];
  assign o[4796] = i[4796];
  assign o[4795] = i[4795];
  assign o[4794] = i[4794];
  assign o[4793] = i[4793];
  assign o[4792] = i[4792];
  assign o[4791] = i[4791];
  assign o[4790] = i[4790];
  assign o[4789] = i[4789];
  assign o[4788] = i[4788];
  assign o[4787] = i[4787];
  assign o[4786] = i[4786];
  assign o[4785] = i[4785];
  assign o[4784] = i[4784];
  assign o[4783] = i[4783];
  assign o[4782] = i[4782];
  assign o[4781] = i[4781];
  assign o[4780] = i[4780];
  assign o[4779] = i[4779];
  assign o[4778] = i[4778];
  assign o[4777] = i[4777];
  assign o[4776] = i[4776];
  assign o[4775] = i[4775];
  assign o[4774] = i[4774];
  assign o[4773] = i[4773];
  assign o[4772] = i[4772];
  assign o[4771] = i[4771];
  assign o[4770] = i[4770];
  assign o[4769] = i[4769];
  assign o[4768] = i[4768];
  assign o[4767] = i[4767];
  assign o[4766] = i[4766];
  assign o[4765] = i[4765];
  assign o[4764] = i[4764];
  assign o[4763] = i[4763];
  assign o[4762] = i[4762];
  assign o[4761] = i[4761];
  assign o[4760] = i[4760];
  assign o[4759] = i[4759];
  assign o[4758] = i[4758];
  assign o[4757] = i[4757];
  assign o[4756] = i[4756];
  assign o[4755] = i[4755];
  assign o[4754] = i[4754];
  assign o[4753] = i[4753];
  assign o[4752] = i[4752];
  assign o[4751] = i[4751];
  assign o[4750] = i[4750];
  assign o[4749] = i[4749];
  assign o[4748] = i[4748];
  assign o[4747] = i[4747];
  assign o[4746] = i[4746];
  assign o[4745] = i[4745];
  assign o[4744] = i[4744];
  assign o[4743] = i[4743];
  assign o[4742] = i[4742];
  assign o[4741] = i[4741];
  assign o[4740] = i[4740];
  assign o[4739] = i[4739];
  assign o[4738] = i[4738];
  assign o[4737] = i[4737];
  assign o[4736] = i[4736];
  assign o[4735] = i[4735];
  assign o[4734] = i[4734];
  assign o[4733] = i[4733];
  assign o[4732] = i[4732];
  assign o[4731] = i[4731];
  assign o[4730] = i[4730];
  assign o[4729] = i[4729];
  assign o[4728] = i[4728];
  assign o[4727] = i[4727];
  assign o[4726] = i[4726];
  assign o[4725] = i[4725];
  assign o[4724] = i[4724];
  assign o[4723] = i[4723];
  assign o[4722] = i[4722];
  assign o[4721] = i[4721];
  assign o[4720] = i[4720];
  assign o[4719] = i[4719];
  assign o[4718] = i[4718];
  assign o[4717] = i[4717];
  assign o[4716] = i[4716];
  assign o[4715] = i[4715];
  assign o[4714] = i[4714];
  assign o[4713] = i[4713];
  assign o[4712] = i[4712];
  assign o[4711] = i[4711];
  assign o[4710] = i[4710];
  assign o[4709] = i[4709];
  assign o[4708] = i[4708];
  assign o[4707] = i[4707];
  assign o[4706] = i[4706];
  assign o[4705] = i[4705];
  assign o[4704] = i[4704];
  assign o[4703] = i[4703];
  assign o[4702] = i[4702];
  assign o[4701] = i[4701];
  assign o[4700] = i[4700];
  assign o[4699] = i[4699];
  assign o[4698] = i[4698];
  assign o[4697] = i[4697];
  assign o[4696] = i[4696];
  assign o[4695] = i[4695];
  assign o[4694] = i[4694];
  assign o[4693] = i[4693];
  assign o[4692] = i[4692];
  assign o[4691] = i[4691];
  assign o[4690] = i[4690];
  assign o[4689] = i[4689];
  assign o[4688] = i[4688];
  assign o[4687] = i[4687];
  assign o[4686] = i[4686];
  assign o[4685] = i[4685];
  assign o[4684] = i[4684];
  assign o[4683] = i[4683];
  assign o[4682] = i[4682];
  assign o[4681] = i[4681];
  assign o[4680] = i[4680];
  assign o[4679] = i[4679];
  assign o[4678] = i[4678];
  assign o[4677] = i[4677];
  assign o[4676] = i[4676];
  assign o[4675] = i[4675];
  assign o[4674] = i[4674];
  assign o[4673] = i[4673];
  assign o[4672] = i[4672];
  assign o[4671] = i[4671];
  assign o[4670] = i[4670];
  assign o[4669] = i[4669];
  assign o[4668] = i[4668];
  assign o[4667] = i[4667];
  assign o[4666] = i[4666];
  assign o[4665] = i[4665];
  assign o[4664] = i[4664];
  assign o[4663] = i[4663];
  assign o[4662] = i[4662];
  assign o[4661] = i[4661];
  assign o[4660] = i[4660];
  assign o[4659] = i[4659];
  assign o[4658] = i[4658];
  assign o[4657] = i[4657];
  assign o[4656] = i[4656];
  assign o[4655] = i[4655];
  assign o[4654] = i[4654];
  assign o[4653] = i[4653];
  assign o[4652] = i[4652];
  assign o[4651] = i[4651];
  assign o[4650] = i[4650];
  assign o[4649] = i[4649];
  assign o[4648] = i[4648];
  assign o[4647] = i[4647];
  assign o[4646] = i[4646];
  assign o[4645] = i[4645];
  assign o[4644] = i[4644];
  assign o[4643] = i[4643];
  assign o[4642] = i[4642];
  assign o[4641] = i[4641];
  assign o[4640] = i[4640];
  assign o[4639] = i[4639];
  assign o[4638] = i[4638];
  assign o[4637] = i[4637];
  assign o[4636] = i[4636];
  assign o[4635] = i[4635];
  assign o[4634] = i[4634];
  assign o[4633] = i[4633];
  assign o[4632] = i[4632];
  assign o[4631] = i[4631];
  assign o[4630] = i[4630];
  assign o[4629] = i[4629];
  assign o[4628] = i[4628];
  assign o[4627] = i[4627];
  assign o[4626] = i[4626];
  assign o[4625] = i[4625];
  assign o[4624] = i[4624];
  assign o[4623] = i[4623];
  assign o[4622] = i[4622];
  assign o[4621] = i[4621];
  assign o[4620] = i[4620];
  assign o[4619] = i[4619];
  assign o[4618] = i[4618];
  assign o[4617] = i[4617];
  assign o[4616] = i[4616];
  assign o[4615] = i[4615];
  assign o[4614] = i[4614];
  assign o[4613] = i[4613];
  assign o[4612] = i[4612];
  assign o[4611] = i[4611];
  assign o[4610] = i[4610];
  assign o[4609] = i[4609];
  assign o[4608] = i[4608];
  assign o[4607] = i[4607];
  assign o[4606] = i[4606];
  assign o[4605] = i[4605];
  assign o[4604] = i[4604];
  assign o[4603] = i[4603];
  assign o[4602] = i[4602];
  assign o[4601] = i[4601];
  assign o[4600] = i[4600];
  assign o[4599] = i[4599];
  assign o[4598] = i[4598];
  assign o[4597] = i[4597];
  assign o[4596] = i[4596];
  assign o[4595] = i[4595];
  assign o[4594] = i[4594];
  assign o[4593] = i[4593];
  assign o[4592] = i[4592];
  assign o[4591] = i[4591];
  assign o[4590] = i[4590];
  assign o[4589] = i[4589];
  assign o[4588] = i[4588];
  assign o[4587] = i[4587];
  assign o[4586] = i[4586];
  assign o[4585] = i[4585];
  assign o[4584] = i[4584];
  assign o[4583] = i[4583];
  assign o[4582] = i[4582];
  assign o[4581] = i[4581];
  assign o[4580] = i[4580];
  assign o[4579] = i[4579];
  assign o[4578] = i[4578];
  assign o[4577] = i[4577];
  assign o[4576] = i[4576];
  assign o[4575] = i[4575];
  assign o[4574] = i[4574];
  assign o[4573] = i[4573];
  assign o[4572] = i[4572];
  assign o[4571] = i[4571];
  assign o[4570] = i[4570];
  assign o[4569] = i[4569];
  assign o[4568] = i[4568];
  assign o[4567] = i[4567];
  assign o[4566] = i[4566];
  assign o[4565] = i[4565];
  assign o[4564] = i[4564];
  assign o[4563] = i[4563];
  assign o[4562] = i[4562];
  assign o[4561] = i[4561];
  assign o[4560] = i[4560];
  assign o[4559] = i[4559];
  assign o[4558] = i[4558];
  assign o[4557] = i[4557];
  assign o[4556] = i[4556];
  assign o[4555] = i[4555];
  assign o[4554] = i[4554];
  assign o[4553] = i[4553];
  assign o[4552] = i[4552];
  assign o[4551] = i[4551];
  assign o[4550] = i[4550];
  assign o[4549] = i[4549];
  assign o[4548] = i[4548];
  assign o[4547] = i[4547];
  assign o[4546] = i[4546];
  assign o[4545] = i[4545];
  assign o[4544] = i[4544];
  assign o[4543] = i[4543];
  assign o[4542] = i[4542];
  assign o[4541] = i[4541];
  assign o[4540] = i[4540];
  assign o[4539] = i[4539];
  assign o[4538] = i[4538];
  assign o[4537] = i[4537];
  assign o[4536] = i[4536];
  assign o[4535] = i[4535];
  assign o[4534] = i[4534];
  assign o[4533] = i[4533];
  assign o[4532] = i[4532];
  assign o[4531] = i[4531];
  assign o[4530] = i[4530];
  assign o[4529] = i[4529];
  assign o[4528] = i[4528];
  assign o[4527] = i[4527];
  assign o[4526] = i[4526];
  assign o[4525] = i[4525];
  assign o[4524] = i[4524];
  assign o[4523] = i[4523];
  assign o[4522] = i[4522];
  assign o[4521] = i[4521];
  assign o[4520] = i[4520];
  assign o[4519] = i[4519];
  assign o[4518] = i[4518];
  assign o[4517] = i[4517];
  assign o[4516] = i[4516];
  assign o[4515] = i[4515];
  assign o[4514] = i[4514];
  assign o[4513] = i[4513];
  assign o[4512] = i[4512];
  assign o[4511] = i[4511];
  assign o[4510] = i[4510];
  assign o[4509] = i[4509];
  assign o[4508] = i[4508];
  assign o[4507] = i[4507];
  assign o[4506] = i[4506];
  assign o[4505] = i[4505];
  assign o[4504] = i[4504];
  assign o[4503] = i[4503];
  assign o[4502] = i[4502];
  assign o[4501] = i[4501];
  assign o[4500] = i[4500];
  assign o[4499] = i[4499];
  assign o[4498] = i[4498];
  assign o[4497] = i[4497];
  assign o[4496] = i[4496];
  assign o[4495] = i[4495];
  assign o[4494] = i[4494];
  assign o[4493] = i[4493];
  assign o[4492] = i[4492];
  assign o[4491] = i[4491];
  assign o[4490] = i[4490];
  assign o[4489] = i[4489];
  assign o[4488] = i[4488];
  assign o[4487] = i[4487];
  assign o[4486] = i[4486];
  assign o[4485] = i[4485];
  assign o[4484] = i[4484];
  assign o[4483] = i[4483];
  assign o[4482] = i[4482];
  assign o[4481] = i[4481];
  assign o[4480] = i[4480];
  assign o[4479] = i[4479];
  assign o[4478] = i[4478];
  assign o[4477] = i[4477];
  assign o[4476] = i[4476];
  assign o[4475] = i[4475];
  assign o[4474] = i[4474];
  assign o[4473] = i[4473];
  assign o[4472] = i[4472];
  assign o[4471] = i[4471];
  assign o[4470] = i[4470];
  assign o[4469] = i[4469];
  assign o[4468] = i[4468];
  assign o[4467] = i[4467];
  assign o[4466] = i[4466];
  assign o[4465] = i[4465];
  assign o[4464] = i[4464];
  assign o[4463] = i[4463];
  assign o[4462] = i[4462];
  assign o[4461] = i[4461];
  assign o[4460] = i[4460];
  assign o[4459] = i[4459];
  assign o[4458] = i[4458];
  assign o[4457] = i[4457];
  assign o[4456] = i[4456];
  assign o[4455] = i[4455];
  assign o[4454] = i[4454];
  assign o[4453] = i[4453];
  assign o[4452] = i[4452];
  assign o[4451] = i[4451];
  assign o[4450] = i[4450];
  assign o[4449] = i[4449];
  assign o[4448] = i[4448];
  assign o[4447] = i[4447];
  assign o[4446] = i[4446];
  assign o[4445] = i[4445];
  assign o[4444] = i[4444];
  assign o[4443] = i[4443];
  assign o[4442] = i[4442];
  assign o[4441] = i[4441];
  assign o[4440] = i[4440];
  assign o[4439] = i[4439];
  assign o[4438] = i[4438];
  assign o[4437] = i[4437];
  assign o[4436] = i[4436];
  assign o[4435] = i[4435];
  assign o[4434] = i[4434];
  assign o[4433] = i[4433];
  assign o[4432] = i[4432];
  assign o[4431] = i[4431];
  assign o[4430] = i[4430];
  assign o[4429] = i[4429];
  assign o[4428] = i[4428];
  assign o[4427] = i[4427];
  assign o[4426] = i[4426];
  assign o[4425] = i[4425];
  assign o[4424] = i[4424];
  assign o[4423] = i[4423];
  assign o[4422] = i[4422];
  assign o[4421] = i[4421];
  assign o[4420] = i[4420];
  assign o[4419] = i[4419];
  assign o[4418] = i[4418];
  assign o[4417] = i[4417];
  assign o[4416] = i[4416];
  assign o[4415] = i[4415];
  assign o[4414] = i[4414];
  assign o[4413] = i[4413];
  assign o[4412] = i[4412];
  assign o[4411] = i[4411];
  assign o[4410] = i[4410];
  assign o[4409] = i[4409];
  assign o[4408] = i[4408];
  assign o[4407] = i[4407];
  assign o[4406] = i[4406];
  assign o[4405] = i[4405];
  assign o[4404] = i[4404];
  assign o[4403] = i[4403];
  assign o[4402] = i[4402];
  assign o[4401] = i[4401];
  assign o[4400] = i[4400];
  assign o[4399] = i[4399];
  assign o[4398] = i[4398];
  assign o[4397] = i[4397];
  assign o[4396] = i[4396];
  assign o[4395] = i[4395];
  assign o[4394] = i[4394];
  assign o[4393] = i[4393];
  assign o[4392] = i[4392];
  assign o[4391] = i[4391];
  assign o[4390] = i[4390];
  assign o[4389] = i[4389];
  assign o[4388] = i[4388];
  assign o[4387] = i[4387];
  assign o[4386] = i[4386];
  assign o[4385] = i[4385];
  assign o[4384] = i[4384];
  assign o[4383] = i[4383];
  assign o[4382] = i[4382];
  assign o[4381] = i[4381];
  assign o[4380] = i[4380];
  assign o[4379] = i[4379];
  assign o[4378] = i[4378];
  assign o[4377] = i[4377];
  assign o[4376] = i[4376];
  assign o[4375] = i[4375];
  assign o[4374] = i[4374];
  assign o[4373] = i[4373];
  assign o[4372] = i[4372];
  assign o[4371] = i[4371];
  assign o[4370] = i[4370];
  assign o[4369] = i[4369];
  assign o[4368] = i[4368];
  assign o[4367] = i[4367];
  assign o[4366] = i[4366];
  assign o[4365] = i[4365];
  assign o[4364] = i[4364];
  assign o[4363] = i[4363];
  assign o[4362] = i[4362];
  assign o[4361] = i[4361];
  assign o[4360] = i[4360];
  assign o[4359] = i[4359];
  assign o[4358] = i[4358];
  assign o[4357] = i[4357];
  assign o[4356] = i[4356];
  assign o[4355] = i[4355];
  assign o[4354] = i[4354];
  assign o[4353] = i[4353];
  assign o[4352] = i[4352];
  assign o[4351] = i[4351];
  assign o[4350] = i[4350];
  assign o[4349] = i[4349];
  assign o[4348] = i[4348];
  assign o[4347] = i[4347];
  assign o[4346] = i[4346];
  assign o[4345] = i[4345];
  assign o[4344] = i[4344];
  assign o[4343] = i[4343];
  assign o[4342] = i[4342];
  assign o[4341] = i[4341];
  assign o[4340] = i[4340];
  assign o[4339] = i[4339];
  assign o[4338] = i[4338];
  assign o[4337] = i[4337];
  assign o[4336] = i[4336];
  assign o[4335] = i[4335];
  assign o[4334] = i[4334];
  assign o[4333] = i[4333];
  assign o[4332] = i[4332];
  assign o[4331] = i[4331];
  assign o[4330] = i[4330];
  assign o[4329] = i[4329];
  assign o[4328] = i[4328];
  assign o[4327] = i[4327];
  assign o[4326] = i[4326];
  assign o[4325] = i[4325];
  assign o[4324] = i[4324];
  assign o[4323] = i[4323];
  assign o[4322] = i[4322];
  assign o[4321] = i[4321];
  assign o[4320] = i[4320];
  assign o[4319] = i[4319];
  assign o[4318] = i[4318];
  assign o[4317] = i[4317];
  assign o[4316] = i[4316];
  assign o[4315] = i[4315];
  assign o[4314] = i[4314];
  assign o[4313] = i[4313];
  assign o[4312] = i[4312];
  assign o[4311] = i[4311];
  assign o[4310] = i[4310];
  assign o[4309] = i[4309];
  assign o[4308] = i[4308];
  assign o[4307] = i[4307];
  assign o[4306] = i[4306];
  assign o[4305] = i[4305];
  assign o[4304] = i[4304];
  assign o[4303] = i[4303];
  assign o[4302] = i[4302];
  assign o[4301] = i[4301];
  assign o[4300] = i[4300];
  assign o[4299] = i[4299];
  assign o[4298] = i[4298];
  assign o[4297] = i[4297];
  assign o[4296] = i[4296];
  assign o[4295] = i[4295];
  assign o[4294] = i[4294];
  assign o[4293] = i[4293];
  assign o[4292] = i[4292];
  assign o[4291] = i[4291];
  assign o[4290] = i[4290];
  assign o[4289] = i[4289];
  assign o[4288] = i[4288];
  assign o[4287] = i[4287];
  assign o[4286] = i[4286];
  assign o[4285] = i[4285];
  assign o[4284] = i[4284];
  assign o[4283] = i[4283];
  assign o[4282] = i[4282];
  assign o[4281] = i[4281];
  assign o[4280] = i[4280];
  assign o[4279] = i[4279];
  assign o[4278] = i[4278];
  assign o[4277] = i[4277];
  assign o[4276] = i[4276];
  assign o[4275] = i[4275];
  assign o[4274] = i[4274];
  assign o[4273] = i[4273];
  assign o[4272] = i[4272];
  assign o[4271] = i[4271];
  assign o[4270] = i[4270];
  assign o[4269] = i[4269];
  assign o[4268] = i[4268];
  assign o[4267] = i[4267];
  assign o[4266] = i[4266];
  assign o[4265] = i[4265];
  assign o[4264] = i[4264];
  assign o[4263] = i[4263];
  assign o[4262] = i[4262];
  assign o[4261] = i[4261];
  assign o[4260] = i[4260];
  assign o[4259] = i[4259];
  assign o[4258] = i[4258];
  assign o[4257] = i[4257];
  assign o[4256] = i[4256];
  assign o[4255] = i[4255];
  assign o[4254] = i[4254];
  assign o[4253] = i[4253];
  assign o[4252] = i[4252];
  assign o[4251] = i[4251];
  assign o[4250] = i[4250];
  assign o[4249] = i[4249];
  assign o[4248] = i[4248];
  assign o[4247] = i[4247];
  assign o[4246] = i[4246];
  assign o[4245] = i[4245];
  assign o[4244] = i[4244];
  assign o[4243] = i[4243];
  assign o[4242] = i[4242];
  assign o[4241] = i[4241];
  assign o[4240] = i[4240];
  assign o[4239] = i[4239];
  assign o[4238] = i[4238];
  assign o[4237] = i[4237];
  assign o[4236] = i[4236];
  assign o[4235] = i[4235];
  assign o[4234] = i[4234];
  assign o[4233] = i[4233];
  assign o[4232] = i[4232];
  assign o[4231] = i[4231];
  assign o[4230] = i[4230];
  assign o[4229] = i[4229];
  assign o[4228] = i[4228];
  assign o[4227] = i[4227];
  assign o[4226] = i[4226];
  assign o[4225] = i[4225];
  assign o[4224] = i[4224];
  assign o[4223] = i[4223];
  assign o[4222] = i[4222];
  assign o[4221] = i[4221];
  assign o[4220] = i[4220];
  assign o[4219] = i[4219];
  assign o[4218] = i[4218];
  assign o[4217] = i[4217];
  assign o[4216] = i[4216];
  assign o[4215] = i[4215];
  assign o[4214] = i[4214];
  assign o[4213] = i[4213];
  assign o[4212] = i[4212];
  assign o[4211] = i[4211];
  assign o[4210] = i[4210];
  assign o[4209] = i[4209];
  assign o[4208] = i[4208];
  assign o[4207] = i[4207];
  assign o[4206] = i[4206];
  assign o[4205] = i[4205];
  assign o[4204] = i[4204];
  assign o[4203] = i[4203];
  assign o[4202] = i[4202];
  assign o[4201] = i[4201];
  assign o[4200] = i[4200];
  assign o[4199] = i[4199];
  assign o[4198] = i[4198];
  assign o[4197] = i[4197];
  assign o[4196] = i[4196];
  assign o[4195] = i[4195];
  assign o[4194] = i[4194];
  assign o[4193] = i[4193];
  assign o[4192] = i[4192];
  assign o[4191] = i[4191];
  assign o[4190] = i[4190];
  assign o[4189] = i[4189];
  assign o[4188] = i[4188];
  assign o[4187] = i[4187];
  assign o[4186] = i[4186];
  assign o[4185] = i[4185];
  assign o[4184] = i[4184];
  assign o[4183] = i[4183];
  assign o[4182] = i[4182];
  assign o[4181] = i[4181];
  assign o[4180] = i[4180];
  assign o[4179] = i[4179];
  assign o[4178] = i[4178];
  assign o[4177] = i[4177];
  assign o[4176] = i[4176];
  assign o[4175] = i[4175];
  assign o[4174] = i[4174];
  assign o[4173] = i[4173];
  assign o[4172] = i[4172];
  assign o[4171] = i[4171];
  assign o[4170] = i[4170];
  assign o[4169] = i[4169];
  assign o[4168] = i[4168];
  assign o[4167] = i[4167];
  assign o[4166] = i[4166];
  assign o[4165] = i[4165];
  assign o[4164] = i[4164];
  assign o[4163] = i[4163];
  assign o[4162] = i[4162];
  assign o[4161] = i[4161];
  assign o[4160] = i[4160];
  assign o[4159] = i[4159];
  assign o[4158] = i[4158];
  assign o[4157] = i[4157];
  assign o[4156] = i[4156];
  assign o[4155] = i[4155];
  assign o[4154] = i[4154];
  assign o[4153] = i[4153];
  assign o[4152] = i[4152];
  assign o[4151] = i[4151];
  assign o[4150] = i[4150];
  assign o[4149] = i[4149];
  assign o[4148] = i[4148];
  assign o[4147] = i[4147];
  assign o[4146] = i[4146];
  assign o[4145] = i[4145];
  assign o[4144] = i[4144];
  assign o[4143] = i[4143];
  assign o[4142] = i[4142];
  assign o[4141] = i[4141];
  assign o[4140] = i[4140];
  assign o[4139] = i[4139];
  assign o[4138] = i[4138];
  assign o[4137] = i[4137];
  assign o[4136] = i[4136];
  assign o[4135] = i[4135];
  assign o[4134] = i[4134];
  assign o[4133] = i[4133];
  assign o[4132] = i[4132];
  assign o[4131] = i[4131];
  assign o[4130] = i[4130];
  assign o[4129] = i[4129];
  assign o[4128] = i[4128];
  assign o[4127] = i[4127];
  assign o[4126] = i[4126];
  assign o[4125] = i[4125];
  assign o[4124] = i[4124];
  assign o[4123] = i[4123];
  assign o[4122] = i[4122];
  assign o[4121] = i[4121];
  assign o[4120] = i[4120];
  assign o[4119] = i[4119];
  assign o[4118] = i[4118];
  assign o[4117] = i[4117];
  assign o[4116] = i[4116];
  assign o[4115] = i[4115];
  assign o[4114] = i[4114];
  assign o[4113] = i[4113];
  assign o[4112] = i[4112];
  assign o[4111] = i[4111];
  assign o[4110] = i[4110];
  assign o[4109] = i[4109];
  assign o[4108] = i[4108];
  assign o[4107] = i[4107];
  assign o[4106] = i[4106];
  assign o[4105] = i[4105];
  assign o[4104] = i[4104];
  assign o[4103] = i[4103];
  assign o[4102] = i[4102];
  assign o[4101] = i[4101];
  assign o[4100] = i[4100];
  assign o[4099] = i[4099];
  assign o[4098] = i[4098];
  assign o[4097] = i[4097];
  assign o[4096] = i[4096];
  assign o[4095] = i[4095];
  assign o[4094] = i[4094];
  assign o[4093] = i[4093];
  assign o[4092] = i[4092];
  assign o[4091] = i[4091];
  assign o[4090] = i[4090];
  assign o[4089] = i[4089];
  assign o[4088] = i[4088];
  assign o[4087] = i[4087];
  assign o[4086] = i[4086];
  assign o[4085] = i[4085];
  assign o[4084] = i[4084];
  assign o[4083] = i[4083];
  assign o[4082] = i[4082];
  assign o[4081] = i[4081];
  assign o[4080] = i[4080];
  assign o[4079] = i[4079];
  assign o[4078] = i[4078];
  assign o[4077] = i[4077];
  assign o[4076] = i[4076];
  assign o[4075] = i[4075];
  assign o[4074] = i[4074];
  assign o[4073] = i[4073];
  assign o[4072] = i[4072];
  assign o[4071] = i[4071];
  assign o[4070] = i[4070];
  assign o[4069] = i[4069];
  assign o[4068] = i[4068];
  assign o[4067] = i[4067];
  assign o[4066] = i[4066];
  assign o[4065] = i[4065];
  assign o[4064] = i[4064];
  assign o[4063] = i[4063];
  assign o[4062] = i[4062];
  assign o[4061] = i[4061];
  assign o[4060] = i[4060];
  assign o[4059] = i[4059];
  assign o[4058] = i[4058];
  assign o[4057] = i[4057];
  assign o[4056] = i[4056];
  assign o[4055] = i[4055];
  assign o[4054] = i[4054];
  assign o[4053] = i[4053];
  assign o[4052] = i[4052];
  assign o[4051] = i[4051];
  assign o[4050] = i[4050];
  assign o[4049] = i[4049];
  assign o[4048] = i[4048];
  assign o[4047] = i[4047];
  assign o[4046] = i[4046];
  assign o[4045] = i[4045];
  assign o[4044] = i[4044];
  assign o[4043] = i[4043];
  assign o[4042] = i[4042];
  assign o[4041] = i[4041];
  assign o[4040] = i[4040];
  assign o[4039] = i[4039];
  assign o[4038] = i[4038];
  assign o[4037] = i[4037];
  assign o[4036] = i[4036];
  assign o[4035] = i[4035];
  assign o[4034] = i[4034];
  assign o[4033] = i[4033];
  assign o[4032] = i[4032];
  assign o[4031] = i[4031];
  assign o[4030] = i[4030];
  assign o[4029] = i[4029];
  assign o[4028] = i[4028];
  assign o[4027] = i[4027];
  assign o[4026] = i[4026];
  assign o[4025] = i[4025];
  assign o[4024] = i[4024];
  assign o[4023] = i[4023];
  assign o[4022] = i[4022];
  assign o[4021] = i[4021];
  assign o[4020] = i[4020];
  assign o[4019] = i[4019];
  assign o[4018] = i[4018];
  assign o[4017] = i[4017];
  assign o[4016] = i[4016];
  assign o[4015] = i[4015];
  assign o[4014] = i[4014];
  assign o[4013] = i[4013];
  assign o[4012] = i[4012];
  assign o[4011] = i[4011];
  assign o[4010] = i[4010];
  assign o[4009] = i[4009];
  assign o[4008] = i[4008];
  assign o[4007] = i[4007];
  assign o[4006] = i[4006];
  assign o[4005] = i[4005];
  assign o[4004] = i[4004];
  assign o[4003] = i[4003];
  assign o[4002] = i[4002];
  assign o[4001] = i[4001];
  assign o[4000] = i[4000];
  assign o[3999] = i[3999];
  assign o[3998] = i[3998];
  assign o[3997] = i[3997];
  assign o[3996] = i[3996];
  assign o[3995] = i[3995];
  assign o[3994] = i[3994];
  assign o[3993] = i[3993];
  assign o[3992] = i[3992];
  assign o[3991] = i[3991];
  assign o[3990] = i[3990];
  assign o[3989] = i[3989];
  assign o[3988] = i[3988];
  assign o[3987] = i[3987];
  assign o[3986] = i[3986];
  assign o[3985] = i[3985];
  assign o[3984] = i[3984];
  assign o[3983] = i[3983];
  assign o[3982] = i[3982];
  assign o[3981] = i[3981];
  assign o[3980] = i[3980];
  assign o[3979] = i[3979];
  assign o[3978] = i[3978];
  assign o[3977] = i[3977];
  assign o[3976] = i[3976];
  assign o[3975] = i[3975];
  assign o[3974] = i[3974];
  assign o[3973] = i[3973];
  assign o[3972] = i[3972];
  assign o[3971] = i[3971];
  assign o[3970] = i[3970];
  assign o[3969] = i[3969];
  assign o[3968] = i[3968];
  assign o[3967] = i[3967];
  assign o[3966] = i[3966];
  assign o[3965] = i[3965];
  assign o[3964] = i[3964];
  assign o[3963] = i[3963];
  assign o[3962] = i[3962];
  assign o[3961] = i[3961];
  assign o[3960] = i[3960];
  assign o[3959] = i[3959];
  assign o[3958] = i[3958];
  assign o[3957] = i[3957];
  assign o[3956] = i[3956];
  assign o[3955] = i[3955];
  assign o[3954] = i[3954];
  assign o[3953] = i[3953];
  assign o[3952] = i[3952];
  assign o[3951] = i[3951];
  assign o[3950] = i[3950];
  assign o[3949] = i[3949];
  assign o[3948] = i[3948];
  assign o[3947] = i[3947];
  assign o[3946] = i[3946];
  assign o[3945] = i[3945];
  assign o[3944] = i[3944];
  assign o[3943] = i[3943];
  assign o[3942] = i[3942];
  assign o[3941] = i[3941];
  assign o[3940] = i[3940];
  assign o[3939] = i[3939];
  assign o[3938] = i[3938];
  assign o[3937] = i[3937];
  assign o[3936] = i[3936];
  assign o[3935] = i[3935];
  assign o[3934] = i[3934];
  assign o[3933] = i[3933];
  assign o[3932] = i[3932];
  assign o[3931] = i[3931];
  assign o[3930] = i[3930];
  assign o[3929] = i[3929];
  assign o[3928] = i[3928];
  assign o[3927] = i[3927];
  assign o[3926] = i[3926];
  assign o[3925] = i[3925];
  assign o[3924] = i[3924];
  assign o[3923] = i[3923];
  assign o[3922] = i[3922];
  assign o[3921] = i[3921];
  assign o[3920] = i[3920];
  assign o[3919] = i[3919];
  assign o[3918] = i[3918];
  assign o[3917] = i[3917];
  assign o[3916] = i[3916];
  assign o[3915] = i[3915];
  assign o[3914] = i[3914];
  assign o[3913] = i[3913];
  assign o[3912] = i[3912];
  assign o[3911] = i[3911];
  assign o[3910] = i[3910];
  assign o[3909] = i[3909];
  assign o[3908] = i[3908];
  assign o[3907] = i[3907];
  assign o[3906] = i[3906];
  assign o[3905] = i[3905];
  assign o[3904] = i[3904];
  assign o[3903] = i[3903];
  assign o[3902] = i[3902];
  assign o[3901] = i[3901];
  assign o[3900] = i[3900];
  assign o[3899] = i[3899];
  assign o[3898] = i[3898];
  assign o[3897] = i[3897];
  assign o[3896] = i[3896];
  assign o[3895] = i[3895];
  assign o[3894] = i[3894];
  assign o[3893] = i[3893];
  assign o[3892] = i[3892];
  assign o[3891] = i[3891];
  assign o[3890] = i[3890];
  assign o[3889] = i[3889];
  assign o[3888] = i[3888];
  assign o[3887] = i[3887];
  assign o[3886] = i[3886];
  assign o[3885] = i[3885];
  assign o[3884] = i[3884];
  assign o[3883] = i[3883];
  assign o[3882] = i[3882];
  assign o[3881] = i[3881];
  assign o[3880] = i[3880];
  assign o[3879] = i[3879];
  assign o[3878] = i[3878];
  assign o[3877] = i[3877];
  assign o[3876] = i[3876];
  assign o[3875] = i[3875];
  assign o[3874] = i[3874];
  assign o[3873] = i[3873];
  assign o[3872] = i[3872];
  assign o[3871] = i[3871];
  assign o[3870] = i[3870];
  assign o[3869] = i[3869];
  assign o[3868] = i[3868];
  assign o[3867] = i[3867];
  assign o[3866] = i[3866];
  assign o[3865] = i[3865];
  assign o[3864] = i[3864];
  assign o[3863] = i[3863];
  assign o[3862] = i[3862];
  assign o[3861] = i[3861];
  assign o[3860] = i[3860];
  assign o[3859] = i[3859];
  assign o[3858] = i[3858];
  assign o[3857] = i[3857];
  assign o[3856] = i[3856];
  assign o[3855] = i[3855];
  assign o[3854] = i[3854];
  assign o[3853] = i[3853];
  assign o[3852] = i[3852];
  assign o[3851] = i[3851];
  assign o[3850] = i[3850];
  assign o[3849] = i[3849];
  assign o[3848] = i[3848];
  assign o[3847] = i[3847];
  assign o[3846] = i[3846];
  assign o[3845] = i[3845];
  assign o[3844] = i[3844];
  assign o[3843] = i[3843];
  assign o[3842] = i[3842];
  assign o[3841] = i[3841];
  assign o[3840] = i[3840];
  assign o[3839] = i[3839];
  assign o[3838] = i[3838];
  assign o[3837] = i[3837];
  assign o[3836] = i[3836];
  assign o[3835] = i[3835];
  assign o[3834] = i[3834];
  assign o[3833] = i[3833];
  assign o[3832] = i[3832];
  assign o[3831] = i[3831];
  assign o[3830] = i[3830];
  assign o[3829] = i[3829];
  assign o[3828] = i[3828];
  assign o[3827] = i[3827];
  assign o[3826] = i[3826];
  assign o[3825] = i[3825];
  assign o[3824] = i[3824];
  assign o[3823] = i[3823];
  assign o[3822] = i[3822];
  assign o[3821] = i[3821];
  assign o[3820] = i[3820];
  assign o[3819] = i[3819];
  assign o[3818] = i[3818];
  assign o[3817] = i[3817];
  assign o[3816] = i[3816];
  assign o[3815] = i[3815];
  assign o[3814] = i[3814];
  assign o[3813] = i[3813];
  assign o[3812] = i[3812];
  assign o[3811] = i[3811];
  assign o[3810] = i[3810];
  assign o[3809] = i[3809];
  assign o[3808] = i[3808];
  assign o[3807] = i[3807];
  assign o[3806] = i[3806];
  assign o[3805] = i[3805];
  assign o[3804] = i[3804];
  assign o[3803] = i[3803];
  assign o[3802] = i[3802];
  assign o[3801] = i[3801];
  assign o[3800] = i[3800];
  assign o[3799] = i[3799];
  assign o[3798] = i[3798];
  assign o[3797] = i[3797];
  assign o[3796] = i[3796];
  assign o[3795] = i[3795];
  assign o[3794] = i[3794];
  assign o[3793] = i[3793];
  assign o[3792] = i[3792];
  assign o[3791] = i[3791];
  assign o[3790] = i[3790];
  assign o[3789] = i[3789];
  assign o[3788] = i[3788];
  assign o[3787] = i[3787];
  assign o[3786] = i[3786];
  assign o[3785] = i[3785];
  assign o[3784] = i[3784];
  assign o[3783] = i[3783];
  assign o[3782] = i[3782];
  assign o[3781] = i[3781];
  assign o[3780] = i[3780];
  assign o[3779] = i[3779];
  assign o[3778] = i[3778];
  assign o[3777] = i[3777];
  assign o[3776] = i[3776];
  assign o[3775] = i[3775];
  assign o[3774] = i[3774];
  assign o[3773] = i[3773];
  assign o[3772] = i[3772];
  assign o[3771] = i[3771];
  assign o[3770] = i[3770];
  assign o[3769] = i[3769];
  assign o[3768] = i[3768];
  assign o[3767] = i[3767];
  assign o[3766] = i[3766];
  assign o[3765] = i[3765];
  assign o[3764] = i[3764];
  assign o[3763] = i[3763];
  assign o[3762] = i[3762];
  assign o[3761] = i[3761];
  assign o[3760] = i[3760];
  assign o[3759] = i[3759];
  assign o[3758] = i[3758];
  assign o[3757] = i[3757];
  assign o[3756] = i[3756];
  assign o[3755] = i[3755];
  assign o[3754] = i[3754];
  assign o[3753] = i[3753];
  assign o[3752] = i[3752];
  assign o[3751] = i[3751];
  assign o[3750] = i[3750];
  assign o[3749] = i[3749];
  assign o[3748] = i[3748];
  assign o[3747] = i[3747];
  assign o[3746] = i[3746];
  assign o[3745] = i[3745];
  assign o[3744] = i[3744];
  assign o[3743] = i[3743];
  assign o[3742] = i[3742];
  assign o[3741] = i[3741];
  assign o[3740] = i[3740];
  assign o[3739] = i[3739];
  assign o[3738] = i[3738];
  assign o[3737] = i[3737];
  assign o[3736] = i[3736];
  assign o[3735] = i[3735];
  assign o[3734] = i[3734];
  assign o[3733] = i[3733];
  assign o[3732] = i[3732];
  assign o[3731] = i[3731];
  assign o[3730] = i[3730];
  assign o[3729] = i[3729];
  assign o[3728] = i[3728];
  assign o[3727] = i[3727];
  assign o[3726] = i[3726];
  assign o[3725] = i[3725];
  assign o[3724] = i[3724];
  assign o[3723] = i[3723];
  assign o[3722] = i[3722];
  assign o[3721] = i[3721];
  assign o[3720] = i[3720];
  assign o[3719] = i[3719];
  assign o[3718] = i[3718];
  assign o[3717] = i[3717];
  assign o[3716] = i[3716];
  assign o[3715] = i[3715];
  assign o[3714] = i[3714];
  assign o[3713] = i[3713];
  assign o[3712] = i[3712];
  assign o[3711] = i[3711];
  assign o[3710] = i[3710];
  assign o[3709] = i[3709];
  assign o[3708] = i[3708];
  assign o[3707] = i[3707];
  assign o[3706] = i[3706];
  assign o[3705] = i[3705];
  assign o[3704] = i[3704];
  assign o[3703] = i[3703];
  assign o[3702] = i[3702];
  assign o[3701] = i[3701];
  assign o[3700] = i[3700];
  assign o[3699] = i[3699];
  assign o[3698] = i[3698];
  assign o[3697] = i[3697];
  assign o[3696] = i[3696];
  assign o[3695] = i[3695];
  assign o[3694] = i[3694];
  assign o[3693] = i[3693];
  assign o[3692] = i[3692];
  assign o[3691] = i[3691];
  assign o[3690] = i[3690];
  assign o[3689] = i[3689];
  assign o[3688] = i[3688];
  assign o[3687] = i[3687];
  assign o[3686] = i[3686];
  assign o[3685] = i[3685];
  assign o[3684] = i[3684];
  assign o[3683] = i[3683];
  assign o[3682] = i[3682];
  assign o[3681] = i[3681];
  assign o[3680] = i[3680];
  assign o[3679] = i[3679];
  assign o[3678] = i[3678];
  assign o[3677] = i[3677];
  assign o[3676] = i[3676];
  assign o[3675] = i[3675];
  assign o[3674] = i[3674];
  assign o[3673] = i[3673];
  assign o[3672] = i[3672];
  assign o[3671] = i[3671];
  assign o[3670] = i[3670];
  assign o[3669] = i[3669];
  assign o[3668] = i[3668];
  assign o[3667] = i[3667];
  assign o[3666] = i[3666];
  assign o[3665] = i[3665];
  assign o[3664] = i[3664];
  assign o[3663] = i[3663];
  assign o[3662] = i[3662];
  assign o[3661] = i[3661];
  assign o[3660] = i[3660];
  assign o[3659] = i[3659];
  assign o[3658] = i[3658];
  assign o[3657] = i[3657];
  assign o[3656] = i[3656];
  assign o[3655] = i[3655];
  assign o[3654] = i[3654];
  assign o[3653] = i[3653];
  assign o[3652] = i[3652];
  assign o[3651] = i[3651];
  assign o[3650] = i[3650];
  assign o[3649] = i[3649];
  assign o[3648] = i[3648];
  assign o[3647] = i[3647];
  assign o[3646] = i[3646];
  assign o[3645] = i[3645];
  assign o[3644] = i[3644];
  assign o[3643] = i[3643];
  assign o[3642] = i[3642];
  assign o[3641] = i[3641];
  assign o[3640] = i[3640];
  assign o[3639] = i[3639];
  assign o[3638] = i[3638];
  assign o[3637] = i[3637];
  assign o[3636] = i[3636];
  assign o[3635] = i[3635];
  assign o[3634] = i[3634];
  assign o[3633] = i[3633];
  assign o[3632] = i[3632];
  assign o[3631] = i[3631];
  assign o[3630] = i[3630];
  assign o[3629] = i[3629];
  assign o[3628] = i[3628];
  assign o[3627] = i[3627];
  assign o[3626] = i[3626];
  assign o[3625] = i[3625];
  assign o[3624] = i[3624];
  assign o[3623] = i[3623];
  assign o[3622] = i[3622];
  assign o[3621] = i[3621];
  assign o[3620] = i[3620];
  assign o[3619] = i[3619];
  assign o[3618] = i[3618];
  assign o[3617] = i[3617];
  assign o[3616] = i[3616];
  assign o[3615] = i[3615];
  assign o[3614] = i[3614];
  assign o[3613] = i[3613];
  assign o[3612] = i[3612];
  assign o[3611] = i[3611];
  assign o[3610] = i[3610];
  assign o[3609] = i[3609];
  assign o[3608] = i[3608];
  assign o[3607] = i[3607];
  assign o[3606] = i[3606];
  assign o[3605] = i[3605];
  assign o[3604] = i[3604];
  assign o[3603] = i[3603];
  assign o[3602] = i[3602];
  assign o[3601] = i[3601];
  assign o[3600] = i[3600];
  assign o[3599] = i[3599];
  assign o[3598] = i[3598];
  assign o[3597] = i[3597];
  assign o[3596] = i[3596];
  assign o[3595] = i[3595];
  assign o[3594] = i[3594];
  assign o[3593] = i[3593];
  assign o[3592] = i[3592];
  assign o[3591] = i[3591];
  assign o[3590] = i[3590];
  assign o[3589] = i[3589];
  assign o[3588] = i[3588];
  assign o[3587] = i[3587];
  assign o[3586] = i[3586];
  assign o[3585] = i[3585];
  assign o[3584] = i[3584];
  assign o[3583] = i[3583];
  assign o[3582] = i[3582];
  assign o[3581] = i[3581];
  assign o[3580] = i[3580];
  assign o[3579] = i[3579];
  assign o[3578] = i[3578];
  assign o[3577] = i[3577];
  assign o[3576] = i[3576];
  assign o[3575] = i[3575];
  assign o[3574] = i[3574];
  assign o[3573] = i[3573];
  assign o[3572] = i[3572];
  assign o[3571] = i[3571];
  assign o[3570] = i[3570];
  assign o[3569] = i[3569];
  assign o[3568] = i[3568];
  assign o[3567] = i[3567];
  assign o[3566] = i[3566];
  assign o[3565] = i[3565];
  assign o[3564] = i[3564];
  assign o[3563] = i[3563];
  assign o[3562] = i[3562];
  assign o[3561] = i[3561];
  assign o[3560] = i[3560];
  assign o[3559] = i[3559];
  assign o[3558] = i[3558];
  assign o[3557] = i[3557];
  assign o[3556] = i[3556];
  assign o[3555] = i[3555];
  assign o[3554] = i[3554];
  assign o[3553] = i[3553];
  assign o[3552] = i[3552];
  assign o[3551] = i[3551];
  assign o[3550] = i[3550];
  assign o[3549] = i[3549];
  assign o[3548] = i[3548];
  assign o[3547] = i[3547];
  assign o[3546] = i[3546];
  assign o[3545] = i[3545];
  assign o[3544] = i[3544];
  assign o[3543] = i[3543];
  assign o[3542] = i[3542];
  assign o[3541] = i[3541];
  assign o[3540] = i[3540];
  assign o[3539] = i[3539];
  assign o[3538] = i[3538];
  assign o[3537] = i[3537];
  assign o[3536] = i[3536];
  assign o[3535] = i[3535];
  assign o[3534] = i[3534];
  assign o[3533] = i[3533];
  assign o[3532] = i[3532];
  assign o[3531] = i[3531];
  assign o[3530] = i[3530];
  assign o[3529] = i[3529];
  assign o[3528] = i[3528];
  assign o[3527] = i[3527];
  assign o[3526] = i[3526];
  assign o[3525] = i[3525];
  assign o[3524] = i[3524];
  assign o[3523] = i[3523];
  assign o[3522] = i[3522];
  assign o[3521] = i[3521];
  assign o[3520] = i[3520];
  assign o[3519] = i[3519];
  assign o[3518] = i[3518];
  assign o[3517] = i[3517];
  assign o[3516] = i[3516];
  assign o[3515] = i[3515];
  assign o[3514] = i[3514];
  assign o[3513] = i[3513];
  assign o[3512] = i[3512];
  assign o[3511] = i[3511];
  assign o[3510] = i[3510];
  assign o[3509] = i[3509];
  assign o[3508] = i[3508];
  assign o[3507] = i[3507];
  assign o[3506] = i[3506];
  assign o[3505] = i[3505];
  assign o[3504] = i[3504];
  assign o[3503] = i[3503];
  assign o[3502] = i[3502];
  assign o[3501] = i[3501];
  assign o[3500] = i[3500];
  assign o[3499] = i[3499];
  assign o[3498] = i[3498];
  assign o[3497] = i[3497];
  assign o[3496] = i[3496];
  assign o[3495] = i[3495];
  assign o[3494] = i[3494];
  assign o[3493] = i[3493];
  assign o[3492] = i[3492];
  assign o[3491] = i[3491];
  assign o[3490] = i[3490];
  assign o[3489] = i[3489];
  assign o[3488] = i[3488];
  assign o[3487] = i[3487];
  assign o[3486] = i[3486];
  assign o[3485] = i[3485];
  assign o[3484] = i[3484];
  assign o[3483] = i[3483];
  assign o[3482] = i[3482];
  assign o[3481] = i[3481];
  assign o[3480] = i[3480];
  assign o[3479] = i[3479];
  assign o[3478] = i[3478];
  assign o[3477] = i[3477];
  assign o[3476] = i[3476];
  assign o[3475] = i[3475];
  assign o[3474] = i[3474];
  assign o[3473] = i[3473];
  assign o[3472] = i[3472];
  assign o[3471] = i[3471];
  assign o[3470] = i[3470];
  assign o[3469] = i[3469];
  assign o[3468] = i[3468];
  assign o[3467] = i[3467];
  assign o[3466] = i[3466];
  assign o[3465] = i[3465];
  assign o[3464] = i[3464];
  assign o[3463] = i[3463];
  assign o[3462] = i[3462];
  assign o[3461] = i[3461];
  assign o[3460] = i[3460];
  assign o[3459] = i[3459];
  assign o[3458] = i[3458];
  assign o[3457] = i[3457];
  assign o[3456] = i[3456];
  assign o[3455] = i[3455];
  assign o[3454] = i[3454];
  assign o[3453] = i[3453];
  assign o[3452] = i[3452];
  assign o[3451] = i[3451];
  assign o[3450] = i[3450];
  assign o[3449] = i[3449];
  assign o[3448] = i[3448];
  assign o[3447] = i[3447];
  assign o[3446] = i[3446];
  assign o[3445] = i[3445];
  assign o[3444] = i[3444];
  assign o[3443] = i[3443];
  assign o[3442] = i[3442];
  assign o[3441] = i[3441];
  assign o[3440] = i[3440];
  assign o[3439] = i[3439];
  assign o[3438] = i[3438];
  assign o[3437] = i[3437];
  assign o[3436] = i[3436];
  assign o[3435] = i[3435];
  assign o[3434] = i[3434];
  assign o[3433] = i[3433];
  assign o[3432] = i[3432];
  assign o[3431] = i[3431];
  assign o[3430] = i[3430];
  assign o[3429] = i[3429];
  assign o[3428] = i[3428];
  assign o[3427] = i[3427];
  assign o[3426] = i[3426];
  assign o[3425] = i[3425];
  assign o[3424] = i[3424];
  assign o[3423] = i[3423];
  assign o[3422] = i[3422];
  assign o[3421] = i[3421];
  assign o[3420] = i[3420];
  assign o[3419] = i[3419];
  assign o[3418] = i[3418];
  assign o[3417] = i[3417];
  assign o[3416] = i[3416];
  assign o[3415] = i[3415];
  assign o[3414] = i[3414];
  assign o[3413] = i[3413];
  assign o[3412] = i[3412];
  assign o[3411] = i[3411];
  assign o[3410] = i[3410];
  assign o[3409] = i[3409];
  assign o[3408] = i[3408];
  assign o[3407] = i[3407];
  assign o[3406] = i[3406];
  assign o[3405] = i[3405];
  assign o[3404] = i[3404];
  assign o[3403] = i[3403];
  assign o[3402] = i[3402];
  assign o[3401] = i[3401];
  assign o[3400] = i[3400];
  assign o[3399] = i[3399];
  assign o[3398] = i[3398];
  assign o[3397] = i[3397];
  assign o[3396] = i[3396];
  assign o[3395] = i[3395];
  assign o[3394] = i[3394];
  assign o[3393] = i[3393];
  assign o[3392] = i[3392];
  assign o[3391] = i[3391];
  assign o[3390] = i[3390];
  assign o[3389] = i[3389];
  assign o[3388] = i[3388];
  assign o[3387] = i[3387];
  assign o[3386] = i[3386];
  assign o[3385] = i[3385];
  assign o[3384] = i[3384];
  assign o[3383] = i[3383];
  assign o[3382] = i[3382];
  assign o[3381] = i[3381];
  assign o[3380] = i[3380];
  assign o[3379] = i[3379];
  assign o[3378] = i[3378];
  assign o[3377] = i[3377];
  assign o[3376] = i[3376];
  assign o[3375] = i[3375];
  assign o[3374] = i[3374];
  assign o[3373] = i[3373];
  assign o[3372] = i[3372];
  assign o[3371] = i[3371];
  assign o[3370] = i[3370];
  assign o[3369] = i[3369];
  assign o[3368] = i[3368];
  assign o[3367] = i[3367];
  assign o[3366] = i[3366];
  assign o[3365] = i[3365];
  assign o[3364] = i[3364];
  assign o[3363] = i[3363];
  assign o[3362] = i[3362];
  assign o[3361] = i[3361];
  assign o[3360] = i[3360];
  assign o[3359] = i[3359];
  assign o[3358] = i[3358];
  assign o[3357] = i[3357];
  assign o[3356] = i[3356];
  assign o[3355] = i[3355];
  assign o[3354] = i[3354];
  assign o[3353] = i[3353];
  assign o[3352] = i[3352];
  assign o[3351] = i[3351];
  assign o[3350] = i[3350];
  assign o[3349] = i[3349];
  assign o[3348] = i[3348];
  assign o[3347] = i[3347];
  assign o[3346] = i[3346];
  assign o[3345] = i[3345];
  assign o[3344] = i[3344];
  assign o[3343] = i[3343];
  assign o[3342] = i[3342];
  assign o[3341] = i[3341];
  assign o[3340] = i[3340];
  assign o[3339] = i[3339];
  assign o[3338] = i[3338];
  assign o[3337] = i[3337];
  assign o[3336] = i[3336];
  assign o[3335] = i[3335];
  assign o[3334] = i[3334];
  assign o[3333] = i[3333];
  assign o[3332] = i[3332];
  assign o[3331] = i[3331];
  assign o[3330] = i[3330];
  assign o[3329] = i[3329];
  assign o[3328] = i[3328];
  assign o[3327] = i[3327];
  assign o[3326] = i[3326];
  assign o[3325] = i[3325];
  assign o[3324] = i[3324];
  assign o[3323] = i[3323];
  assign o[3322] = i[3322];
  assign o[3321] = i[3321];
  assign o[3320] = i[3320];
  assign o[3319] = i[3319];
  assign o[3318] = i[3318];
  assign o[3317] = i[3317];
  assign o[3316] = i[3316];
  assign o[3315] = i[3315];
  assign o[3314] = i[3314];
  assign o[3313] = i[3313];
  assign o[3312] = i[3312];
  assign o[3311] = i[3311];
  assign o[3310] = i[3310];
  assign o[3309] = i[3309];
  assign o[3308] = i[3308];
  assign o[3307] = i[3307];
  assign o[3306] = i[3306];
  assign o[3305] = i[3305];
  assign o[3304] = i[3304];
  assign o[3303] = i[3303];
  assign o[3302] = i[3302];
  assign o[3301] = i[3301];
  assign o[3300] = i[3300];
  assign o[3299] = i[3299];
  assign o[3298] = i[3298];
  assign o[3297] = i[3297];
  assign o[3296] = i[3296];
  assign o[3295] = i[3295];
  assign o[3294] = i[3294];
  assign o[3293] = i[3293];
  assign o[3292] = i[3292];
  assign o[3291] = i[3291];
  assign o[3290] = i[3290];
  assign o[3289] = i[3289];
  assign o[3288] = i[3288];
  assign o[3287] = i[3287];
  assign o[3286] = i[3286];
  assign o[3285] = i[3285];
  assign o[3284] = i[3284];
  assign o[3283] = i[3283];
  assign o[3282] = i[3282];
  assign o[3281] = i[3281];
  assign o[3280] = i[3280];
  assign o[3279] = i[3279];
  assign o[3278] = i[3278];
  assign o[3277] = i[3277];
  assign o[3276] = i[3276];
  assign o[3275] = i[3275];
  assign o[3274] = i[3274];
  assign o[3273] = i[3273];
  assign o[3272] = i[3272];
  assign o[3271] = i[3271];
  assign o[3270] = i[3270];
  assign o[3269] = i[3269];
  assign o[3268] = i[3268];
  assign o[3267] = i[3267];
  assign o[3266] = i[3266];
  assign o[3265] = i[3265];
  assign o[3264] = i[3264];
  assign o[3263] = i[3263];
  assign o[3262] = i[3262];
  assign o[3261] = i[3261];
  assign o[3260] = i[3260];
  assign o[3259] = i[3259];
  assign o[3258] = i[3258];
  assign o[3257] = i[3257];
  assign o[3256] = i[3256];
  assign o[3255] = i[3255];
  assign o[3254] = i[3254];
  assign o[3253] = i[3253];
  assign o[3252] = i[3252];
  assign o[3251] = i[3251];
  assign o[3250] = i[3250];
  assign o[3249] = i[3249];
  assign o[3248] = i[3248];
  assign o[3247] = i[3247];
  assign o[3246] = i[3246];
  assign o[3245] = i[3245];
  assign o[3244] = i[3244];
  assign o[3243] = i[3243];
  assign o[3242] = i[3242];
  assign o[3241] = i[3241];
  assign o[3240] = i[3240];
  assign o[3239] = i[3239];
  assign o[3238] = i[3238];
  assign o[3237] = i[3237];
  assign o[3236] = i[3236];
  assign o[3235] = i[3235];
  assign o[3234] = i[3234];
  assign o[3233] = i[3233];
  assign o[3232] = i[3232];
  assign o[3231] = i[3231];
  assign o[3230] = i[3230];
  assign o[3229] = i[3229];
  assign o[3228] = i[3228];
  assign o[3227] = i[3227];
  assign o[3226] = i[3226];
  assign o[3225] = i[3225];
  assign o[3224] = i[3224];
  assign o[3223] = i[3223];
  assign o[3222] = i[3222];
  assign o[3221] = i[3221];
  assign o[3220] = i[3220];
  assign o[3219] = i[3219];
  assign o[3218] = i[3218];
  assign o[3217] = i[3217];
  assign o[3216] = i[3216];
  assign o[3215] = i[3215];
  assign o[3214] = i[3214];
  assign o[3213] = i[3213];
  assign o[3212] = i[3212];
  assign o[3211] = i[3211];
  assign o[3210] = i[3210];
  assign o[3209] = i[3209];
  assign o[3208] = i[3208];
  assign o[3207] = i[3207];
  assign o[3206] = i[3206];
  assign o[3205] = i[3205];
  assign o[3204] = i[3204];
  assign o[3203] = i[3203];
  assign o[3202] = i[3202];
  assign o[3201] = i[3201];
  assign o[3200] = i[3200];
  assign o[3199] = i[3199];
  assign o[3198] = i[3198];
  assign o[3197] = i[3197];
  assign o[3196] = i[3196];
  assign o[3195] = i[3195];
  assign o[3194] = i[3194];
  assign o[3193] = i[3193];
  assign o[3192] = i[3192];
  assign o[3191] = i[3191];
  assign o[3190] = i[3190];
  assign o[3189] = i[3189];
  assign o[3188] = i[3188];
  assign o[3187] = i[3187];
  assign o[3186] = i[3186];
  assign o[3185] = i[3185];
  assign o[3184] = i[3184];
  assign o[3183] = i[3183];
  assign o[3182] = i[3182];
  assign o[3181] = i[3181];
  assign o[3180] = i[3180];
  assign o[3179] = i[3179];
  assign o[3178] = i[3178];
  assign o[3177] = i[3177];
  assign o[3176] = i[3176];
  assign o[3175] = i[3175];
  assign o[3174] = i[3174];
  assign o[3173] = i[3173];
  assign o[3172] = i[3172];
  assign o[3171] = i[3171];
  assign o[3170] = i[3170];
  assign o[3169] = i[3169];
  assign o[3168] = i[3168];
  assign o[3167] = i[3167];
  assign o[3166] = i[3166];
  assign o[3165] = i[3165];
  assign o[3164] = i[3164];
  assign o[3163] = i[3163];
  assign o[3162] = i[3162];
  assign o[3161] = i[3161];
  assign o[3160] = i[3160];
  assign o[3159] = i[3159];
  assign o[3158] = i[3158];
  assign o[3157] = i[3157];
  assign o[3156] = i[3156];
  assign o[3155] = i[3155];
  assign o[3154] = i[3154];
  assign o[3153] = i[3153];
  assign o[3152] = i[3152];
  assign o[3151] = i[3151];
  assign o[3150] = i[3150];
  assign o[3149] = i[3149];
  assign o[3148] = i[3148];
  assign o[3147] = i[3147];
  assign o[3146] = i[3146];
  assign o[3145] = i[3145];
  assign o[3144] = i[3144];
  assign o[3143] = i[3143];
  assign o[3142] = i[3142];
  assign o[3141] = i[3141];
  assign o[3140] = i[3140];
  assign o[3139] = i[3139];
  assign o[3138] = i[3138];
  assign o[3137] = i[3137];
  assign o[3136] = i[3136];
  assign o[3135] = i[3135];
  assign o[3134] = i[3134];
  assign o[3133] = i[3133];
  assign o[3132] = i[3132];
  assign o[3131] = i[3131];
  assign o[3130] = i[3130];
  assign o[3129] = i[3129];
  assign o[3128] = i[3128];
  assign o[3127] = i[3127];
  assign o[3126] = i[3126];
  assign o[3125] = i[3125];
  assign o[3124] = i[3124];
  assign o[3123] = i[3123];
  assign o[3122] = i[3122];
  assign o[3121] = i[3121];
  assign o[3120] = i[3120];
  assign o[3119] = i[3119];
  assign o[3118] = i[3118];
  assign o[3117] = i[3117];
  assign o[3116] = i[3116];
  assign o[3115] = i[3115];
  assign o[3114] = i[3114];
  assign o[3113] = i[3113];
  assign o[3112] = i[3112];
  assign o[3111] = i[3111];
  assign o[3110] = i[3110];
  assign o[3109] = i[3109];
  assign o[3108] = i[3108];
  assign o[3107] = i[3107];
  assign o[3106] = i[3106];
  assign o[3105] = i[3105];
  assign o[3104] = i[3104];
  assign o[3103] = i[3103];
  assign o[3102] = i[3102];
  assign o[3101] = i[3101];
  assign o[3100] = i[3100];
  assign o[3099] = i[3099];
  assign o[3098] = i[3098];
  assign o[3097] = i[3097];
  assign o[3096] = i[3096];
  assign o[3095] = i[3095];
  assign o[3094] = i[3094];
  assign o[3093] = i[3093];
  assign o[3092] = i[3092];
  assign o[3091] = i[3091];
  assign o[3090] = i[3090];
  assign o[3089] = i[3089];
  assign o[3088] = i[3088];
  assign o[3087] = i[3087];
  assign o[3086] = i[3086];
  assign o[3085] = i[3085];
  assign o[3084] = i[3084];
  assign o[3083] = i[3083];
  assign o[3082] = i[3082];
  assign o[3081] = i[3081];
  assign o[3080] = i[3080];
  assign o[3079] = i[3079];
  assign o[3078] = i[3078];
  assign o[3077] = i[3077];
  assign o[3076] = i[3076];
  assign o[3075] = i[3075];
  assign o[3074] = i[3074];
  assign o[3073] = i[3073];
  assign o[3072] = i[3072];
  assign o[3071] = i[3071];
  assign o[3070] = i[3070];
  assign o[3069] = i[3069];
  assign o[3068] = i[3068];
  assign o[3067] = i[3067];
  assign o[3066] = i[3066];
  assign o[3065] = i[3065];
  assign o[3064] = i[3064];
  assign o[3063] = i[3063];
  assign o[3062] = i[3062];
  assign o[3061] = i[3061];
  assign o[3060] = i[3060];
  assign o[3059] = i[3059];
  assign o[3058] = i[3058];
  assign o[3057] = i[3057];
  assign o[3056] = i[3056];
  assign o[3055] = i[3055];
  assign o[3054] = i[3054];
  assign o[3053] = i[3053];
  assign o[3052] = i[3052];
  assign o[3051] = i[3051];
  assign o[3050] = i[3050];
  assign o[3049] = i[3049];
  assign o[3048] = i[3048];
  assign o[3047] = i[3047];
  assign o[3046] = i[3046];
  assign o[3045] = i[3045];
  assign o[3044] = i[3044];
  assign o[3043] = i[3043];
  assign o[3042] = i[3042];
  assign o[3041] = i[3041];
  assign o[3040] = i[3040];
  assign o[3039] = i[3039];
  assign o[3038] = i[3038];
  assign o[3037] = i[3037];
  assign o[3036] = i[3036];
  assign o[3035] = i[3035];
  assign o[3034] = i[3034];
  assign o[3033] = i[3033];
  assign o[3032] = i[3032];
  assign o[3031] = i[3031];
  assign o[3030] = i[3030];
  assign o[3029] = i[3029];
  assign o[3028] = i[3028];
  assign o[3027] = i[3027];
  assign o[3026] = i[3026];
  assign o[3025] = i[3025];
  assign o[3024] = i[3024];
  assign o[3023] = i[3023];
  assign o[3022] = i[3022];
  assign o[3021] = i[3021];
  assign o[3020] = i[3020];
  assign o[3019] = i[3019];
  assign o[3018] = i[3018];
  assign o[3017] = i[3017];
  assign o[3016] = i[3016];
  assign o[3015] = i[3015];
  assign o[3014] = i[3014];
  assign o[3013] = i[3013];
  assign o[3012] = i[3012];
  assign o[3011] = i[3011];
  assign o[3010] = i[3010];
  assign o[3009] = i[3009];
  assign o[3008] = i[3008];
  assign o[3007] = i[3007];
  assign o[3006] = i[3006];
  assign o[3005] = i[3005];
  assign o[3004] = i[3004];
  assign o[3003] = i[3003];
  assign o[3002] = i[3002];
  assign o[3001] = i[3001];
  assign o[3000] = i[3000];
  assign o[2999] = i[2999];
  assign o[2998] = i[2998];
  assign o[2997] = i[2997];
  assign o[2996] = i[2996];
  assign o[2995] = i[2995];
  assign o[2994] = i[2994];
  assign o[2993] = i[2993];
  assign o[2992] = i[2992];
  assign o[2991] = i[2991];
  assign o[2990] = i[2990];
  assign o[2989] = i[2989];
  assign o[2988] = i[2988];
  assign o[2987] = i[2987];
  assign o[2986] = i[2986];
  assign o[2985] = i[2985];
  assign o[2984] = i[2984];
  assign o[2983] = i[2983];
  assign o[2982] = i[2982];
  assign o[2981] = i[2981];
  assign o[2980] = i[2980];
  assign o[2979] = i[2979];
  assign o[2978] = i[2978];
  assign o[2977] = i[2977];
  assign o[2976] = i[2976];
  assign o[2975] = i[2975];
  assign o[2974] = i[2974];
  assign o[2973] = i[2973];
  assign o[2972] = i[2972];
  assign o[2971] = i[2971];
  assign o[2970] = i[2970];
  assign o[2969] = i[2969];
  assign o[2968] = i[2968];
  assign o[2967] = i[2967];
  assign o[2966] = i[2966];
  assign o[2965] = i[2965];
  assign o[2964] = i[2964];
  assign o[2963] = i[2963];
  assign o[2962] = i[2962];
  assign o[2961] = i[2961];
  assign o[2960] = i[2960];
  assign o[2959] = i[2959];
  assign o[2958] = i[2958];
  assign o[2957] = i[2957];
  assign o[2956] = i[2956];
  assign o[2955] = i[2955];
  assign o[2954] = i[2954];
  assign o[2953] = i[2953];
  assign o[2952] = i[2952];
  assign o[2951] = i[2951];
  assign o[2950] = i[2950];
  assign o[2949] = i[2949];
  assign o[2948] = i[2948];
  assign o[2947] = i[2947];
  assign o[2946] = i[2946];
  assign o[2945] = i[2945];
  assign o[2944] = i[2944];
  assign o[2943] = i[2943];
  assign o[2942] = i[2942];
  assign o[2941] = i[2941];
  assign o[2940] = i[2940];
  assign o[2939] = i[2939];
  assign o[2938] = i[2938];
  assign o[2937] = i[2937];
  assign o[2936] = i[2936];
  assign o[2935] = i[2935];
  assign o[2934] = i[2934];
  assign o[2933] = i[2933];
  assign o[2932] = i[2932];
  assign o[2931] = i[2931];
  assign o[2930] = i[2930];
  assign o[2929] = i[2929];
  assign o[2928] = i[2928];
  assign o[2927] = i[2927];
  assign o[2926] = i[2926];
  assign o[2925] = i[2925];
  assign o[2924] = i[2924];
  assign o[2923] = i[2923];
  assign o[2922] = i[2922];
  assign o[2921] = i[2921];
  assign o[2920] = i[2920];
  assign o[2919] = i[2919];
  assign o[2918] = i[2918];
  assign o[2917] = i[2917];
  assign o[2916] = i[2916];
  assign o[2915] = i[2915];
  assign o[2914] = i[2914];
  assign o[2913] = i[2913];
  assign o[2912] = i[2912];
  assign o[2911] = i[2911];
  assign o[2910] = i[2910];
  assign o[2909] = i[2909];
  assign o[2908] = i[2908];
  assign o[2907] = i[2907];
  assign o[2906] = i[2906];
  assign o[2905] = i[2905];
  assign o[2904] = i[2904];
  assign o[2903] = i[2903];
  assign o[2902] = i[2902];
  assign o[2901] = i[2901];
  assign o[2900] = i[2900];
  assign o[2899] = i[2899];
  assign o[2898] = i[2898];
  assign o[2897] = i[2897];
  assign o[2896] = i[2896];
  assign o[2895] = i[2895];
  assign o[2894] = i[2894];
  assign o[2893] = i[2893];
  assign o[2892] = i[2892];
  assign o[2891] = i[2891];
  assign o[2890] = i[2890];
  assign o[2889] = i[2889];
  assign o[2888] = i[2888];
  assign o[2887] = i[2887];
  assign o[2886] = i[2886];
  assign o[2885] = i[2885];
  assign o[2884] = i[2884];
  assign o[2883] = i[2883];
  assign o[2882] = i[2882];
  assign o[2881] = i[2881];
  assign o[2880] = i[2880];
  assign o[2879] = i[2879];
  assign o[2878] = i[2878];
  assign o[2877] = i[2877];
  assign o[2876] = i[2876];
  assign o[2875] = i[2875];
  assign o[2874] = i[2874];
  assign o[2873] = i[2873];
  assign o[2872] = i[2872];
  assign o[2871] = i[2871];
  assign o[2870] = i[2870];
  assign o[2869] = i[2869];
  assign o[2868] = i[2868];
  assign o[2867] = i[2867];
  assign o[2866] = i[2866];
  assign o[2865] = i[2865];
  assign o[2864] = i[2864];
  assign o[2863] = i[2863];
  assign o[2862] = i[2862];
  assign o[2861] = i[2861];
  assign o[2860] = i[2860];
  assign o[2859] = i[2859];
  assign o[2858] = i[2858];
  assign o[2857] = i[2857];
  assign o[2856] = i[2856];
  assign o[2855] = i[2855];
  assign o[2854] = i[2854];
  assign o[2853] = i[2853];
  assign o[2852] = i[2852];
  assign o[2851] = i[2851];
  assign o[2850] = i[2850];
  assign o[2849] = i[2849];
  assign o[2848] = i[2848];
  assign o[2847] = i[2847];
  assign o[2846] = i[2846];
  assign o[2845] = i[2845];
  assign o[2844] = i[2844];
  assign o[2843] = i[2843];
  assign o[2842] = i[2842];
  assign o[2841] = i[2841];
  assign o[2840] = i[2840];
  assign o[2839] = i[2839];
  assign o[2838] = i[2838];
  assign o[2837] = i[2837];
  assign o[2836] = i[2836];
  assign o[2835] = i[2835];
  assign o[2834] = i[2834];
  assign o[2833] = i[2833];
  assign o[2832] = i[2832];
  assign o[2831] = i[2831];
  assign o[2830] = i[2830];
  assign o[2829] = i[2829];
  assign o[2828] = i[2828];
  assign o[2827] = i[2827];
  assign o[2826] = i[2826];
  assign o[2825] = i[2825];
  assign o[2824] = i[2824];
  assign o[2823] = i[2823];
  assign o[2822] = i[2822];
  assign o[2821] = i[2821];
  assign o[2820] = i[2820];
  assign o[2819] = i[2819];
  assign o[2818] = i[2818];
  assign o[2817] = i[2817];
  assign o[2816] = i[2816];
  assign o[2815] = i[2815];
  assign o[2814] = i[2814];
  assign o[2813] = i[2813];
  assign o[2812] = i[2812];
  assign o[2811] = i[2811];
  assign o[2810] = i[2810];
  assign o[2809] = i[2809];
  assign o[2808] = i[2808];
  assign o[2807] = i[2807];
  assign o[2806] = i[2806];
  assign o[2805] = i[2805];
  assign o[2804] = i[2804];
  assign o[2803] = i[2803];
  assign o[2802] = i[2802];
  assign o[2801] = i[2801];
  assign o[2800] = i[2800];
  assign o[2799] = i[2799];
  assign o[2798] = i[2798];
  assign o[2797] = i[2797];
  assign o[2796] = i[2796];
  assign o[2795] = i[2795];
  assign o[2794] = i[2794];
  assign o[2793] = i[2793];
  assign o[2792] = i[2792];
  assign o[2791] = i[2791];
  assign o[2790] = i[2790];
  assign o[2789] = i[2789];
  assign o[2788] = i[2788];
  assign o[2787] = i[2787];
  assign o[2786] = i[2786];
  assign o[2785] = i[2785];
  assign o[2784] = i[2784];
  assign o[2783] = i[2783];
  assign o[2782] = i[2782];
  assign o[2781] = i[2781];
  assign o[2780] = i[2780];
  assign o[2779] = i[2779];
  assign o[2778] = i[2778];
  assign o[2777] = i[2777];
  assign o[2776] = i[2776];
  assign o[2775] = i[2775];
  assign o[2774] = i[2774];
  assign o[2773] = i[2773];
  assign o[2772] = i[2772];
  assign o[2771] = i[2771];
  assign o[2770] = i[2770];
  assign o[2769] = i[2769];
  assign o[2768] = i[2768];
  assign o[2767] = i[2767];
  assign o[2766] = i[2766];
  assign o[2765] = i[2765];
  assign o[2764] = i[2764];
  assign o[2763] = i[2763];
  assign o[2762] = i[2762];
  assign o[2761] = i[2761];
  assign o[2760] = i[2760];
  assign o[2759] = i[2759];
  assign o[2758] = i[2758];
  assign o[2757] = i[2757];
  assign o[2756] = i[2756];
  assign o[2755] = i[2755];
  assign o[2754] = i[2754];
  assign o[2753] = i[2753];
  assign o[2752] = i[2752];
  assign o[2751] = i[2751];
  assign o[2750] = i[2750];
  assign o[2749] = i[2749];
  assign o[2748] = i[2748];
  assign o[2747] = i[2747];
  assign o[2746] = i[2746];
  assign o[2745] = i[2745];
  assign o[2744] = i[2744];
  assign o[2743] = i[2743];
  assign o[2742] = i[2742];
  assign o[2741] = i[2741];
  assign o[2740] = i[2740];
  assign o[2739] = i[2739];
  assign o[2738] = i[2738];
  assign o[2737] = i[2737];
  assign o[2736] = i[2736];
  assign o[2735] = i[2735];
  assign o[2734] = i[2734];
  assign o[2733] = i[2733];
  assign o[2732] = i[2732];
  assign o[2731] = i[2731];
  assign o[2730] = i[2730];
  assign o[2729] = i[2729];
  assign o[2728] = i[2728];
  assign o[2727] = i[2727];
  assign o[2726] = i[2726];
  assign o[2725] = i[2725];
  assign o[2724] = i[2724];
  assign o[2723] = i[2723];
  assign o[2722] = i[2722];
  assign o[2721] = i[2721];
  assign o[2720] = i[2720];
  assign o[2719] = i[2719];
  assign o[2718] = i[2718];
  assign o[2717] = i[2717];
  assign o[2716] = i[2716];
  assign o[2715] = i[2715];
  assign o[2714] = i[2714];
  assign o[2713] = i[2713];
  assign o[2712] = i[2712];
  assign o[2711] = i[2711];
  assign o[2710] = i[2710];
  assign o[2709] = i[2709];
  assign o[2708] = i[2708];
  assign o[2707] = i[2707];
  assign o[2706] = i[2706];
  assign o[2705] = i[2705];
  assign o[2704] = i[2704];
  assign o[2703] = i[2703];
  assign o[2702] = i[2702];
  assign o[2701] = i[2701];
  assign o[2700] = i[2700];
  assign o[2699] = i[2699];
  assign o[2698] = i[2698];
  assign o[2697] = i[2697];
  assign o[2696] = i[2696];
  assign o[2695] = i[2695];
  assign o[2694] = i[2694];
  assign o[2693] = i[2693];
  assign o[2692] = i[2692];
  assign o[2691] = i[2691];
  assign o[2690] = i[2690];
  assign o[2689] = i[2689];
  assign o[2688] = i[2688];
  assign o[2687] = i[2687];
  assign o[2686] = i[2686];
  assign o[2685] = i[2685];
  assign o[2684] = i[2684];
  assign o[2683] = i[2683];
  assign o[2682] = i[2682];
  assign o[2681] = i[2681];
  assign o[2680] = i[2680];
  assign o[2679] = i[2679];
  assign o[2678] = i[2678];
  assign o[2677] = i[2677];
  assign o[2676] = i[2676];
  assign o[2675] = i[2675];
  assign o[2674] = i[2674];
  assign o[2673] = i[2673];
  assign o[2672] = i[2672];
  assign o[2671] = i[2671];
  assign o[2670] = i[2670];
  assign o[2669] = i[2669];
  assign o[2668] = i[2668];
  assign o[2667] = i[2667];
  assign o[2666] = i[2666];
  assign o[2665] = i[2665];
  assign o[2664] = i[2664];
  assign o[2663] = i[2663];
  assign o[2662] = i[2662];
  assign o[2661] = i[2661];
  assign o[2660] = i[2660];
  assign o[2659] = i[2659];
  assign o[2658] = i[2658];
  assign o[2657] = i[2657];
  assign o[2656] = i[2656];
  assign o[2655] = i[2655];
  assign o[2654] = i[2654];
  assign o[2653] = i[2653];
  assign o[2652] = i[2652];
  assign o[2651] = i[2651];
  assign o[2650] = i[2650];
  assign o[2649] = i[2649];
  assign o[2648] = i[2648];
  assign o[2647] = i[2647];
  assign o[2646] = i[2646];
  assign o[2645] = i[2645];
  assign o[2644] = i[2644];
  assign o[2643] = i[2643];
  assign o[2642] = i[2642];
  assign o[2641] = i[2641];
  assign o[2640] = i[2640];
  assign o[2639] = i[2639];
  assign o[2638] = i[2638];
  assign o[2637] = i[2637];
  assign o[2636] = i[2636];
  assign o[2635] = i[2635];
  assign o[2634] = i[2634];
  assign o[2633] = i[2633];
  assign o[2632] = i[2632];
  assign o[2631] = i[2631];
  assign o[2630] = i[2630];
  assign o[2629] = i[2629];
  assign o[2628] = i[2628];
  assign o[2627] = i[2627];
  assign o[2626] = i[2626];
  assign o[2625] = i[2625];
  assign o[2624] = i[2624];
  assign o[2623] = i[2623];
  assign o[2622] = i[2622];
  assign o[2621] = i[2621];
  assign o[2620] = i[2620];
  assign o[2619] = i[2619];
  assign o[2618] = i[2618];
  assign o[2617] = i[2617];
  assign o[2616] = i[2616];
  assign o[2615] = i[2615];
  assign o[2614] = i[2614];
  assign o[2613] = i[2613];
  assign o[2612] = i[2612];
  assign o[2611] = i[2611];
  assign o[2610] = i[2610];
  assign o[2609] = i[2609];
  assign o[2608] = i[2608];
  assign o[2607] = i[2607];
  assign o[2606] = i[2606];
  assign o[2605] = i[2605];
  assign o[2604] = i[2604];
  assign o[2603] = i[2603];
  assign o[2602] = i[2602];
  assign o[2601] = i[2601];
  assign o[2600] = i[2600];
  assign o[2599] = i[2599];
  assign o[2598] = i[2598];
  assign o[2597] = i[2597];
  assign o[2596] = i[2596];
  assign o[2595] = i[2595];
  assign o[2594] = i[2594];
  assign o[2593] = i[2593];
  assign o[2592] = i[2592];
  assign o[2591] = i[2591];
  assign o[2590] = i[2590];
  assign o[2589] = i[2589];
  assign o[2588] = i[2588];
  assign o[2587] = i[2587];
  assign o[2586] = i[2586];
  assign o[2585] = i[2585];
  assign o[2584] = i[2584];
  assign o[2583] = i[2583];
  assign o[2582] = i[2582];
  assign o[2581] = i[2581];
  assign o[2580] = i[2580];
  assign o[2579] = i[2579];
  assign o[2578] = i[2578];
  assign o[2577] = i[2577];
  assign o[2576] = i[2576];
  assign o[2575] = i[2575];
  assign o[2574] = i[2574];
  assign o[2573] = i[2573];
  assign o[2572] = i[2572];
  assign o[2571] = i[2571];
  assign o[2570] = i[2570];
  assign o[2569] = i[2569];
  assign o[2568] = i[2568];
  assign o[2567] = i[2567];
  assign o[2566] = i[2566];
  assign o[2565] = i[2565];
  assign o[2564] = i[2564];
  assign o[2563] = i[2563];
  assign o[2562] = i[2562];
  assign o[2561] = i[2561];
  assign o[2560] = i[2560];
  assign o[2559] = i[2559];
  assign o[2558] = i[2558];
  assign o[2557] = i[2557];
  assign o[2556] = i[2556];
  assign o[2555] = i[2555];
  assign o[2554] = i[2554];
  assign o[2553] = i[2553];
  assign o[2552] = i[2552];
  assign o[2551] = i[2551];
  assign o[2550] = i[2550];
  assign o[2549] = i[2549];
  assign o[2548] = i[2548];
  assign o[2547] = i[2547];
  assign o[2546] = i[2546];
  assign o[2545] = i[2545];
  assign o[2544] = i[2544];
  assign o[2543] = i[2543];
  assign o[2542] = i[2542];
  assign o[2541] = i[2541];
  assign o[2540] = i[2540];
  assign o[2539] = i[2539];
  assign o[2538] = i[2538];
  assign o[2537] = i[2537];
  assign o[2536] = i[2536];
  assign o[2535] = i[2535];
  assign o[2534] = i[2534];
  assign o[2533] = i[2533];
  assign o[2532] = i[2532];
  assign o[2531] = i[2531];
  assign o[2530] = i[2530];
  assign o[2529] = i[2529];
  assign o[2528] = i[2528];
  assign o[2527] = i[2527];
  assign o[2526] = i[2526];
  assign o[2525] = i[2525];
  assign o[2524] = i[2524];
  assign o[2523] = i[2523];
  assign o[2522] = i[2522];
  assign o[2521] = i[2521];
  assign o[2520] = i[2520];
  assign o[2519] = i[2519];
  assign o[2518] = i[2518];
  assign o[2517] = i[2517];
  assign o[2516] = i[2516];
  assign o[2515] = i[2515];
  assign o[2514] = i[2514];
  assign o[2513] = i[2513];
  assign o[2512] = i[2512];
  assign o[2511] = i[2511];
  assign o[2510] = i[2510];
  assign o[2509] = i[2509];
  assign o[2508] = i[2508];
  assign o[2507] = i[2507];
  assign o[2506] = i[2506];
  assign o[2505] = i[2505];
  assign o[2504] = i[2504];
  assign o[2503] = i[2503];
  assign o[2502] = i[2502];
  assign o[2501] = i[2501];
  assign o[2500] = i[2500];
  assign o[2499] = i[2499];
  assign o[2498] = i[2498];
  assign o[2497] = i[2497];
  assign o[2496] = i[2496];
  assign o[2495] = i[2495];
  assign o[2494] = i[2494];
  assign o[2493] = i[2493];
  assign o[2492] = i[2492];
  assign o[2491] = i[2491];
  assign o[2490] = i[2490];
  assign o[2489] = i[2489];
  assign o[2488] = i[2488];
  assign o[2487] = i[2487];
  assign o[2486] = i[2486];
  assign o[2485] = i[2485];
  assign o[2484] = i[2484];
  assign o[2483] = i[2483];
  assign o[2482] = i[2482];
  assign o[2481] = i[2481];
  assign o[2480] = i[2480];
  assign o[2479] = i[2479];
  assign o[2478] = i[2478];
  assign o[2477] = i[2477];
  assign o[2476] = i[2476];
  assign o[2475] = i[2475];
  assign o[2474] = i[2474];
  assign o[2473] = i[2473];
  assign o[2472] = i[2472];
  assign o[2471] = i[2471];
  assign o[2470] = i[2470];
  assign o[2469] = i[2469];
  assign o[2468] = i[2468];
  assign o[2467] = i[2467];
  assign o[2466] = i[2466];
  assign o[2465] = i[2465];
  assign o[2464] = i[2464];
  assign o[2463] = i[2463];
  assign o[2462] = i[2462];
  assign o[2461] = i[2461];
  assign o[2460] = i[2460];
  assign o[2459] = i[2459];
  assign o[2458] = i[2458];
  assign o[2457] = i[2457];
  assign o[2456] = i[2456];
  assign o[2455] = i[2455];
  assign o[2454] = i[2454];
  assign o[2453] = i[2453];
  assign o[2452] = i[2452];
  assign o[2451] = i[2451];
  assign o[2450] = i[2450];
  assign o[2449] = i[2449];
  assign o[2448] = i[2448];
  assign o[2447] = i[2447];
  assign o[2446] = i[2446];
  assign o[2445] = i[2445];
  assign o[2444] = i[2444];
  assign o[2443] = i[2443];
  assign o[2442] = i[2442];
  assign o[2441] = i[2441];
  assign o[2440] = i[2440];
  assign o[2439] = i[2439];
  assign o[2438] = i[2438];
  assign o[2437] = i[2437];
  assign o[2436] = i[2436];
  assign o[2435] = i[2435];
  assign o[2434] = i[2434];
  assign o[2433] = i[2433];
  assign o[2432] = i[2432];
  assign o[2431] = i[2431];
  assign o[2430] = i[2430];
  assign o[2429] = i[2429];
  assign o[2428] = i[2428];
  assign o[2427] = i[2427];
  assign o[2426] = i[2426];
  assign o[2425] = i[2425];
  assign o[2424] = i[2424];
  assign o[2423] = i[2423];
  assign o[2422] = i[2422];
  assign o[2421] = i[2421];
  assign o[2420] = i[2420];
  assign o[2419] = i[2419];
  assign o[2418] = i[2418];
  assign o[2417] = i[2417];
  assign o[2416] = i[2416];
  assign o[2415] = i[2415];
  assign o[2414] = i[2414];
  assign o[2413] = i[2413];
  assign o[2412] = i[2412];
  assign o[2411] = i[2411];
  assign o[2410] = i[2410];
  assign o[2409] = i[2409];
  assign o[2408] = i[2408];
  assign o[2407] = i[2407];
  assign o[2406] = i[2406];
  assign o[2405] = i[2405];
  assign o[2404] = i[2404];
  assign o[2403] = i[2403];
  assign o[2402] = i[2402];
  assign o[2401] = i[2401];
  assign o[2400] = i[2400];
  assign o[2399] = i[2399];
  assign o[2398] = i[2398];
  assign o[2397] = i[2397];
  assign o[2396] = i[2396];
  assign o[2395] = i[2395];
  assign o[2394] = i[2394];
  assign o[2393] = i[2393];
  assign o[2392] = i[2392];
  assign o[2391] = i[2391];
  assign o[2390] = i[2390];
  assign o[2389] = i[2389];
  assign o[2388] = i[2388];
  assign o[2387] = i[2387];
  assign o[2386] = i[2386];
  assign o[2385] = i[2385];
  assign o[2384] = i[2384];
  assign o[2383] = i[2383];
  assign o[2382] = i[2382];
  assign o[2381] = i[2381];
  assign o[2380] = i[2380];
  assign o[2379] = i[2379];
  assign o[2378] = i[2378];
  assign o[2377] = i[2377];
  assign o[2376] = i[2376];
  assign o[2375] = i[2375];
  assign o[2374] = i[2374];
  assign o[2373] = i[2373];
  assign o[2372] = i[2372];
  assign o[2371] = i[2371];
  assign o[2370] = i[2370];
  assign o[2369] = i[2369];
  assign o[2368] = i[2368];
  assign o[2367] = i[2367];
  assign o[2366] = i[2366];
  assign o[2365] = i[2365];
  assign o[2364] = i[2364];
  assign o[2363] = i[2363];
  assign o[2362] = i[2362];
  assign o[2361] = i[2361];
  assign o[2360] = i[2360];
  assign o[2359] = i[2359];
  assign o[2358] = i[2358];
  assign o[2357] = i[2357];
  assign o[2356] = i[2356];
  assign o[2355] = i[2355];
  assign o[2354] = i[2354];
  assign o[2353] = i[2353];
  assign o[2352] = i[2352];
  assign o[2351] = i[2351];
  assign o[2350] = i[2350];
  assign o[2349] = i[2349];
  assign o[2348] = i[2348];
  assign o[2347] = i[2347];
  assign o[2346] = i[2346];
  assign o[2345] = i[2345];
  assign o[2344] = i[2344];
  assign o[2343] = i[2343];
  assign o[2342] = i[2342];
  assign o[2341] = i[2341];
  assign o[2340] = i[2340];
  assign o[2339] = i[2339];
  assign o[2338] = i[2338];
  assign o[2337] = i[2337];
  assign o[2336] = i[2336];
  assign o[2335] = i[2335];
  assign o[2334] = i[2334];
  assign o[2333] = i[2333];
  assign o[2332] = i[2332];
  assign o[2331] = i[2331];
  assign o[2330] = i[2330];
  assign o[2329] = i[2329];
  assign o[2328] = i[2328];
  assign o[2327] = i[2327];
  assign o[2326] = i[2326];
  assign o[2325] = i[2325];
  assign o[2324] = i[2324];
  assign o[2323] = i[2323];
  assign o[2322] = i[2322];
  assign o[2321] = i[2321];
  assign o[2320] = i[2320];
  assign o[2319] = i[2319];
  assign o[2318] = i[2318];
  assign o[2317] = i[2317];
  assign o[2316] = i[2316];
  assign o[2315] = i[2315];
  assign o[2314] = i[2314];
  assign o[2313] = i[2313];
  assign o[2312] = i[2312];
  assign o[2311] = i[2311];
  assign o[2310] = i[2310];
  assign o[2309] = i[2309];
  assign o[2308] = i[2308];
  assign o[2307] = i[2307];
  assign o[2306] = i[2306];
  assign o[2305] = i[2305];
  assign o[2304] = i[2304];
  assign o[2303] = i[2303];
  assign o[2302] = i[2302];
  assign o[2301] = i[2301];
  assign o[2300] = i[2300];
  assign o[2299] = i[2299];
  assign o[2298] = i[2298];
  assign o[2297] = i[2297];
  assign o[2296] = i[2296];
  assign o[2295] = i[2295];
  assign o[2294] = i[2294];
  assign o[2293] = i[2293];
  assign o[2292] = i[2292];
  assign o[2291] = i[2291];
  assign o[2290] = i[2290];
  assign o[2289] = i[2289];
  assign o[2288] = i[2288];
  assign o[2287] = i[2287];
  assign o[2286] = i[2286];
  assign o[2285] = i[2285];
  assign o[2284] = i[2284];
  assign o[2283] = i[2283];
  assign o[2282] = i[2282];
  assign o[2281] = i[2281];
  assign o[2280] = i[2280];
  assign o[2279] = i[2279];
  assign o[2278] = i[2278];
  assign o[2277] = i[2277];
  assign o[2276] = i[2276];
  assign o[2275] = i[2275];
  assign o[2274] = i[2274];
  assign o[2273] = i[2273];
  assign o[2272] = i[2272];
  assign o[2271] = i[2271];
  assign o[2270] = i[2270];
  assign o[2269] = i[2269];
  assign o[2268] = i[2268];
  assign o[2267] = i[2267];
  assign o[2266] = i[2266];
  assign o[2265] = i[2265];
  assign o[2264] = i[2264];
  assign o[2263] = i[2263];
  assign o[2262] = i[2262];
  assign o[2261] = i[2261];
  assign o[2260] = i[2260];
  assign o[2259] = i[2259];
  assign o[2258] = i[2258];
  assign o[2257] = i[2257];
  assign o[2256] = i[2256];
  assign o[2255] = i[2255];
  assign o[2254] = i[2254];
  assign o[2253] = i[2253];
  assign o[2252] = i[2252];
  assign o[2251] = i[2251];
  assign o[2250] = i[2250];
  assign o[2249] = i[2249];
  assign o[2248] = i[2248];
  assign o[2247] = i[2247];
  assign o[2246] = i[2246];
  assign o[2245] = i[2245];
  assign o[2244] = i[2244];
  assign o[2243] = i[2243];
  assign o[2242] = i[2242];
  assign o[2241] = i[2241];
  assign o[2240] = i[2240];
  assign o[2239] = i[2239];
  assign o[2238] = i[2238];
  assign o[2237] = i[2237];
  assign o[2236] = i[2236];
  assign o[2235] = i[2235];
  assign o[2234] = i[2234];
  assign o[2233] = i[2233];
  assign o[2232] = i[2232];
  assign o[2231] = i[2231];
  assign o[2230] = i[2230];
  assign o[2229] = i[2229];
  assign o[2228] = i[2228];
  assign o[2227] = i[2227];
  assign o[2226] = i[2226];
  assign o[2225] = i[2225];
  assign o[2224] = i[2224];
  assign o[2223] = i[2223];
  assign o[2222] = i[2222];
  assign o[2221] = i[2221];
  assign o[2220] = i[2220];
  assign o[2219] = i[2219];
  assign o[2218] = i[2218];
  assign o[2217] = i[2217];
  assign o[2216] = i[2216];
  assign o[2215] = i[2215];
  assign o[2214] = i[2214];
  assign o[2213] = i[2213];
  assign o[2212] = i[2212];
  assign o[2211] = i[2211];
  assign o[2210] = i[2210];
  assign o[2209] = i[2209];
  assign o[2208] = i[2208];
  assign o[2207] = i[2207];
  assign o[2206] = i[2206];
  assign o[2205] = i[2205];
  assign o[2204] = i[2204];
  assign o[2203] = i[2203];
  assign o[2202] = i[2202];
  assign o[2201] = i[2201];
  assign o[2200] = i[2200];
  assign o[2199] = i[2199];
  assign o[2198] = i[2198];
  assign o[2197] = i[2197];
  assign o[2196] = i[2196];
  assign o[2195] = i[2195];
  assign o[2194] = i[2194];
  assign o[2193] = i[2193];
  assign o[2192] = i[2192];
  assign o[2191] = i[2191];
  assign o[2190] = i[2190];
  assign o[2189] = i[2189];
  assign o[2188] = i[2188];
  assign o[2187] = i[2187];
  assign o[2186] = i[2186];
  assign o[2185] = i[2185];
  assign o[2184] = i[2184];
  assign o[2183] = i[2183];
  assign o[2182] = i[2182];
  assign o[2181] = i[2181];
  assign o[2180] = i[2180];
  assign o[2179] = i[2179];
  assign o[2178] = i[2178];
  assign o[2177] = i[2177];
  assign o[2176] = i[2176];
  assign o[2175] = i[2175];
  assign o[2174] = i[2174];
  assign o[2173] = i[2173];
  assign o[2172] = i[2172];
  assign o[2171] = i[2171];
  assign o[2170] = i[2170];
  assign o[2169] = i[2169];
  assign o[2168] = i[2168];
  assign o[2167] = i[2167];
  assign o[2166] = i[2166];
  assign o[2165] = i[2165];
  assign o[2164] = i[2164];
  assign o[2163] = i[2163];
  assign o[2162] = i[2162];
  assign o[2161] = i[2161];
  assign o[2160] = i[2160];
  assign o[2159] = i[2159];
  assign o[2158] = i[2158];
  assign o[2157] = i[2157];
  assign o[2156] = i[2156];
  assign o[2155] = i[2155];
  assign o[2154] = i[2154];
  assign o[2153] = i[2153];
  assign o[2152] = i[2152];
  assign o[2151] = i[2151];
  assign o[2150] = i[2150];
  assign o[2149] = i[2149];
  assign o[2148] = i[2148];
  assign o[2147] = i[2147];
  assign o[2146] = i[2146];
  assign o[2145] = i[2145];
  assign o[2144] = i[2144];
  assign o[2143] = i[2143];
  assign o[2142] = i[2142];
  assign o[2141] = i[2141];
  assign o[2140] = i[2140];
  assign o[2139] = i[2139];
  assign o[2138] = i[2138];
  assign o[2137] = i[2137];
  assign o[2136] = i[2136];
  assign o[2135] = i[2135];
  assign o[2134] = i[2134];
  assign o[2133] = i[2133];
  assign o[2132] = i[2132];
  assign o[2131] = i[2131];
  assign o[2130] = i[2130];
  assign o[2129] = i[2129];
  assign o[2128] = i[2128];
  assign o[2127] = i[2127];
  assign o[2126] = i[2126];
  assign o[2125] = i[2125];
  assign o[2124] = i[2124];
  assign o[2123] = i[2123];
  assign o[2122] = i[2122];
  assign o[2121] = i[2121];
  assign o[2120] = i[2120];
  assign o[2119] = i[2119];
  assign o[2118] = i[2118];
  assign o[2117] = i[2117];
  assign o[2116] = i[2116];
  assign o[2115] = i[2115];
  assign o[2114] = i[2114];
  assign o[2113] = i[2113];
  assign o[2112] = i[2112];
  assign o[2111] = i[2111];
  assign o[2110] = i[2110];
  assign o[2109] = i[2109];
  assign o[2108] = i[2108];
  assign o[2107] = i[2107];
  assign o[2106] = i[2106];
  assign o[2105] = i[2105];
  assign o[2104] = i[2104];
  assign o[2103] = i[2103];
  assign o[2102] = i[2102];
  assign o[2101] = i[2101];
  assign o[2100] = i[2100];
  assign o[2099] = i[2099];
  assign o[2098] = i[2098];
  assign o[2097] = i[2097];
  assign o[2096] = i[2096];
  assign o[2095] = i[2095];
  assign o[2094] = i[2094];
  assign o[2093] = i[2093];
  assign o[2092] = i[2092];
  assign o[2091] = i[2091];
  assign o[2090] = i[2090];
  assign o[2089] = i[2089];
  assign o[2088] = i[2088];
  assign o[2087] = i[2087];
  assign o[2086] = i[2086];
  assign o[2085] = i[2085];
  assign o[2084] = i[2084];
  assign o[2083] = i[2083];
  assign o[2082] = i[2082];
  assign o[2081] = i[2081];
  assign o[2080] = i[2080];
  assign o[2079] = i[2079];
  assign o[2078] = i[2078];
  assign o[2077] = i[2077];
  assign o[2076] = i[2076];
  assign o[2075] = i[2075];
  assign o[2074] = i[2074];
  assign o[2073] = i[2073];
  assign o[2072] = i[2072];
  assign o[2071] = i[2071];
  assign o[2070] = i[2070];
  assign o[2069] = i[2069];
  assign o[2068] = i[2068];
  assign o[2067] = i[2067];
  assign o[2066] = i[2066];
  assign o[2065] = i[2065];
  assign o[2064] = i[2064];
  assign o[2063] = i[2063];
  assign o[2062] = i[2062];
  assign o[2061] = i[2061];
  assign o[2060] = i[2060];
  assign o[2059] = i[2059];
  assign o[2058] = i[2058];
  assign o[2057] = i[2057];
  assign o[2056] = i[2056];
  assign o[2055] = i[2055];
  assign o[2054] = i[2054];
  assign o[2053] = i[2053];
  assign o[2052] = i[2052];
  assign o[2051] = i[2051];
  assign o[2050] = i[2050];
  assign o[2049] = i[2049];
  assign o[2048] = i[2048];
  assign o[2047] = i[2047];
  assign o[2046] = i[2046];
  assign o[2045] = i[2045];
  assign o[2044] = i[2044];
  assign o[2043] = i[2043];
  assign o[2042] = i[2042];
  assign o[2041] = i[2041];
  assign o[2040] = i[2040];
  assign o[2039] = i[2039];
  assign o[2038] = i[2038];
  assign o[2037] = i[2037];
  assign o[2036] = i[2036];
  assign o[2035] = i[2035];
  assign o[2034] = i[2034];
  assign o[2033] = i[2033];
  assign o[2032] = i[2032];
  assign o[2031] = i[2031];
  assign o[2030] = i[2030];
  assign o[2029] = i[2029];
  assign o[2028] = i[2028];
  assign o[2027] = i[2027];
  assign o[2026] = i[2026];
  assign o[2025] = i[2025];
  assign o[2024] = i[2024];
  assign o[2023] = i[2023];
  assign o[2022] = i[2022];
  assign o[2021] = i[2021];
  assign o[2020] = i[2020];
  assign o[2019] = i[2019];
  assign o[2018] = i[2018];
  assign o[2017] = i[2017];
  assign o[2016] = i[2016];
  assign o[2015] = i[2015];
  assign o[2014] = i[2014];
  assign o[2013] = i[2013];
  assign o[2012] = i[2012];
  assign o[2011] = i[2011];
  assign o[2010] = i[2010];
  assign o[2009] = i[2009];
  assign o[2008] = i[2008];
  assign o[2007] = i[2007];
  assign o[2006] = i[2006];
  assign o[2005] = i[2005];
  assign o[2004] = i[2004];
  assign o[2003] = i[2003];
  assign o[2002] = i[2002];
  assign o[2001] = i[2001];
  assign o[2000] = i[2000];
  assign o[1999] = i[1999];
  assign o[1998] = i[1998];
  assign o[1997] = i[1997];
  assign o[1996] = i[1996];
  assign o[1995] = i[1995];
  assign o[1994] = i[1994];
  assign o[1993] = i[1993];
  assign o[1992] = i[1992];
  assign o[1991] = i[1991];
  assign o[1990] = i[1990];
  assign o[1989] = i[1989];
  assign o[1988] = i[1988];
  assign o[1987] = i[1987];
  assign o[1986] = i[1986];
  assign o[1985] = i[1985];
  assign o[1984] = i[1984];
  assign o[1983] = i[1983];
  assign o[1982] = i[1982];
  assign o[1981] = i[1981];
  assign o[1980] = i[1980];
  assign o[1979] = i[1979];
  assign o[1978] = i[1978];
  assign o[1977] = i[1977];
  assign o[1976] = i[1976];
  assign o[1975] = i[1975];
  assign o[1974] = i[1974];
  assign o[1973] = i[1973];
  assign o[1972] = i[1972];
  assign o[1971] = i[1971];
  assign o[1970] = i[1970];
  assign o[1969] = i[1969];
  assign o[1968] = i[1968];
  assign o[1967] = i[1967];
  assign o[1966] = i[1966];
  assign o[1965] = i[1965];
  assign o[1964] = i[1964];
  assign o[1963] = i[1963];
  assign o[1962] = i[1962];
  assign o[1961] = i[1961];
  assign o[1960] = i[1960];
  assign o[1959] = i[1959];
  assign o[1958] = i[1958];
  assign o[1957] = i[1957];
  assign o[1956] = i[1956];
  assign o[1955] = i[1955];
  assign o[1954] = i[1954];
  assign o[1953] = i[1953];
  assign o[1952] = i[1952];
  assign o[1951] = i[1951];
  assign o[1950] = i[1950];
  assign o[1949] = i[1949];
  assign o[1948] = i[1948];
  assign o[1947] = i[1947];
  assign o[1946] = i[1946];
  assign o[1945] = i[1945];
  assign o[1944] = i[1944];
  assign o[1943] = i[1943];
  assign o[1942] = i[1942];
  assign o[1941] = i[1941];
  assign o[1940] = i[1940];
  assign o[1939] = i[1939];
  assign o[1938] = i[1938];
  assign o[1937] = i[1937];
  assign o[1936] = i[1936];
  assign o[1935] = i[1935];
  assign o[1934] = i[1934];
  assign o[1933] = i[1933];
  assign o[1932] = i[1932];
  assign o[1931] = i[1931];
  assign o[1930] = i[1930];
  assign o[1929] = i[1929];
  assign o[1928] = i[1928];
  assign o[1927] = i[1927];
  assign o[1926] = i[1926];
  assign o[1925] = i[1925];
  assign o[1924] = i[1924];
  assign o[1923] = i[1923];
  assign o[1922] = i[1922];
  assign o[1921] = i[1921];
  assign o[1920] = i[1920];
  assign o[1919] = i[1919];
  assign o[1918] = i[1918];
  assign o[1917] = i[1917];
  assign o[1916] = i[1916];
  assign o[1915] = i[1915];
  assign o[1914] = i[1914];
  assign o[1913] = i[1913];
  assign o[1912] = i[1912];
  assign o[1911] = i[1911];
  assign o[1910] = i[1910];
  assign o[1909] = i[1909];
  assign o[1908] = i[1908];
  assign o[1907] = i[1907];
  assign o[1906] = i[1906];
  assign o[1905] = i[1905];
  assign o[1904] = i[1904];
  assign o[1903] = i[1903];
  assign o[1902] = i[1902];
  assign o[1901] = i[1901];
  assign o[1900] = i[1900];
  assign o[1899] = i[1899];
  assign o[1898] = i[1898];
  assign o[1897] = i[1897];
  assign o[1896] = i[1896];
  assign o[1895] = i[1895];
  assign o[1894] = i[1894];
  assign o[1893] = i[1893];
  assign o[1892] = i[1892];
  assign o[1891] = i[1891];
  assign o[1890] = i[1890];
  assign o[1889] = i[1889];
  assign o[1888] = i[1888];
  assign o[1887] = i[1887];
  assign o[1886] = i[1886];
  assign o[1885] = i[1885];
  assign o[1884] = i[1884];
  assign o[1883] = i[1883];
  assign o[1882] = i[1882];
  assign o[1881] = i[1881];
  assign o[1880] = i[1880];
  assign o[1879] = i[1879];
  assign o[1878] = i[1878];
  assign o[1877] = i[1877];
  assign o[1876] = i[1876];
  assign o[1875] = i[1875];
  assign o[1874] = i[1874];
  assign o[1873] = i[1873];
  assign o[1872] = i[1872];
  assign o[1871] = i[1871];
  assign o[1870] = i[1870];
  assign o[1869] = i[1869];
  assign o[1868] = i[1868];
  assign o[1867] = i[1867];
  assign o[1866] = i[1866];
  assign o[1865] = i[1865];
  assign o[1864] = i[1864];
  assign o[1863] = i[1863];
  assign o[1862] = i[1862];
  assign o[1861] = i[1861];
  assign o[1860] = i[1860];
  assign o[1859] = i[1859];
  assign o[1858] = i[1858];
  assign o[1857] = i[1857];
  assign o[1856] = i[1856];
  assign o[1855] = i[1855];
  assign o[1854] = i[1854];
  assign o[1853] = i[1853];
  assign o[1852] = i[1852];
  assign o[1851] = i[1851];
  assign o[1850] = i[1850];
  assign o[1849] = i[1849];
  assign o[1848] = i[1848];
  assign o[1847] = i[1847];
  assign o[1846] = i[1846];
  assign o[1845] = i[1845];
  assign o[1844] = i[1844];
  assign o[1843] = i[1843];
  assign o[1842] = i[1842];
  assign o[1841] = i[1841];
  assign o[1840] = i[1840];
  assign o[1839] = i[1839];
  assign o[1838] = i[1838];
  assign o[1837] = i[1837];
  assign o[1836] = i[1836];
  assign o[1835] = i[1835];
  assign o[1834] = i[1834];
  assign o[1833] = i[1833];
  assign o[1832] = i[1832];
  assign o[1831] = i[1831];
  assign o[1830] = i[1830];
  assign o[1829] = i[1829];
  assign o[1828] = i[1828];
  assign o[1827] = i[1827];
  assign o[1826] = i[1826];
  assign o[1825] = i[1825];
  assign o[1824] = i[1824];
  assign o[1823] = i[1823];
  assign o[1822] = i[1822];
  assign o[1821] = i[1821];
  assign o[1820] = i[1820];
  assign o[1819] = i[1819];
  assign o[1818] = i[1818];
  assign o[1817] = i[1817];
  assign o[1816] = i[1816];
  assign o[1815] = i[1815];
  assign o[1814] = i[1814];
  assign o[1813] = i[1813];
  assign o[1812] = i[1812];
  assign o[1811] = i[1811];
  assign o[1810] = i[1810];
  assign o[1809] = i[1809];
  assign o[1808] = i[1808];
  assign o[1807] = i[1807];
  assign o[1806] = i[1806];
  assign o[1805] = i[1805];
  assign o[1804] = i[1804];
  assign o[1803] = i[1803];
  assign o[1802] = i[1802];
  assign o[1801] = i[1801];
  assign o[1800] = i[1800];
  assign o[1799] = i[1799];
  assign o[1798] = i[1798];
  assign o[1797] = i[1797];
  assign o[1796] = i[1796];
  assign o[1795] = i[1795];
  assign o[1794] = i[1794];
  assign o[1793] = i[1793];
  assign o[1792] = i[1792];
  assign o[1791] = i[1791];
  assign o[1790] = i[1790];
  assign o[1789] = i[1789];
  assign o[1788] = i[1788];
  assign o[1787] = i[1787];
  assign o[1786] = i[1786];
  assign o[1785] = i[1785];
  assign o[1784] = i[1784];
  assign o[1783] = i[1783];
  assign o[1782] = i[1782];
  assign o[1781] = i[1781];
  assign o[1780] = i[1780];
  assign o[1779] = i[1779];
  assign o[1778] = i[1778];
  assign o[1777] = i[1777];
  assign o[1776] = i[1776];
  assign o[1775] = i[1775];
  assign o[1774] = i[1774];
  assign o[1773] = i[1773];
  assign o[1772] = i[1772];
  assign o[1771] = i[1771];
  assign o[1770] = i[1770];
  assign o[1769] = i[1769];
  assign o[1768] = i[1768];
  assign o[1767] = i[1767];
  assign o[1766] = i[1766];
  assign o[1765] = i[1765];
  assign o[1764] = i[1764];
  assign o[1763] = i[1763];
  assign o[1762] = i[1762];
  assign o[1761] = i[1761];
  assign o[1760] = i[1760];
  assign o[1759] = i[1759];
  assign o[1758] = i[1758];
  assign o[1757] = i[1757];
  assign o[1756] = i[1756];
  assign o[1755] = i[1755];
  assign o[1754] = i[1754];
  assign o[1753] = i[1753];
  assign o[1752] = i[1752];
  assign o[1751] = i[1751];
  assign o[1750] = i[1750];
  assign o[1749] = i[1749];
  assign o[1748] = i[1748];
  assign o[1747] = i[1747];
  assign o[1746] = i[1746];
  assign o[1745] = i[1745];
  assign o[1744] = i[1744];
  assign o[1743] = i[1743];
  assign o[1742] = i[1742];
  assign o[1741] = i[1741];
  assign o[1740] = i[1740];
  assign o[1739] = i[1739];
  assign o[1738] = i[1738];
  assign o[1737] = i[1737];
  assign o[1736] = i[1736];
  assign o[1735] = i[1735];
  assign o[1734] = i[1734];
  assign o[1733] = i[1733];
  assign o[1732] = i[1732];
  assign o[1731] = i[1731];
  assign o[1730] = i[1730];
  assign o[1729] = i[1729];
  assign o[1728] = i[1728];
  assign o[1727] = i[1727];
  assign o[1726] = i[1726];
  assign o[1725] = i[1725];
  assign o[1724] = i[1724];
  assign o[1723] = i[1723];
  assign o[1722] = i[1722];
  assign o[1721] = i[1721];
  assign o[1720] = i[1720];
  assign o[1719] = i[1719];
  assign o[1718] = i[1718];
  assign o[1717] = i[1717];
  assign o[1716] = i[1716];
  assign o[1715] = i[1715];
  assign o[1714] = i[1714];
  assign o[1713] = i[1713];
  assign o[1712] = i[1712];
  assign o[1711] = i[1711];
  assign o[1710] = i[1710];
  assign o[1709] = i[1709];
  assign o[1708] = i[1708];
  assign o[1707] = i[1707];
  assign o[1706] = i[1706];
  assign o[1705] = i[1705];
  assign o[1704] = i[1704];
  assign o[1703] = i[1703];
  assign o[1702] = i[1702];
  assign o[1701] = i[1701];
  assign o[1700] = i[1700];
  assign o[1699] = i[1699];
  assign o[1698] = i[1698];
  assign o[1697] = i[1697];
  assign o[1696] = i[1696];
  assign o[1695] = i[1695];
  assign o[1694] = i[1694];
  assign o[1693] = i[1693];
  assign o[1692] = i[1692];
  assign o[1691] = i[1691];
  assign o[1690] = i[1690];
  assign o[1689] = i[1689];
  assign o[1688] = i[1688];
  assign o[1687] = i[1687];
  assign o[1686] = i[1686];
  assign o[1685] = i[1685];
  assign o[1684] = i[1684];
  assign o[1683] = i[1683];
  assign o[1682] = i[1682];
  assign o[1681] = i[1681];
  assign o[1680] = i[1680];
  assign o[1679] = i[1679];
  assign o[1678] = i[1678];
  assign o[1677] = i[1677];
  assign o[1676] = i[1676];
  assign o[1675] = i[1675];
  assign o[1674] = i[1674];
  assign o[1673] = i[1673];
  assign o[1672] = i[1672];
  assign o[1671] = i[1671];
  assign o[1670] = i[1670];
  assign o[1669] = i[1669];
  assign o[1668] = i[1668];
  assign o[1667] = i[1667];
  assign o[1666] = i[1666];
  assign o[1665] = i[1665];
  assign o[1664] = i[1664];
  assign o[1663] = i[1663];
  assign o[1662] = i[1662];
  assign o[1661] = i[1661];
  assign o[1660] = i[1660];
  assign o[1659] = i[1659];
  assign o[1658] = i[1658];
  assign o[1657] = i[1657];
  assign o[1656] = i[1656];
  assign o[1655] = i[1655];
  assign o[1654] = i[1654];
  assign o[1653] = i[1653];
  assign o[1652] = i[1652];
  assign o[1651] = i[1651];
  assign o[1650] = i[1650];
  assign o[1649] = i[1649];
  assign o[1648] = i[1648];
  assign o[1647] = i[1647];
  assign o[1646] = i[1646];
  assign o[1645] = i[1645];
  assign o[1644] = i[1644];
  assign o[1643] = i[1643];
  assign o[1642] = i[1642];
  assign o[1641] = i[1641];
  assign o[1640] = i[1640];
  assign o[1639] = i[1639];
  assign o[1638] = i[1638];
  assign o[1637] = i[1637];
  assign o[1636] = i[1636];
  assign o[1635] = i[1635];
  assign o[1634] = i[1634];
  assign o[1633] = i[1633];
  assign o[1632] = i[1632];
  assign o[1631] = i[1631];
  assign o[1630] = i[1630];
  assign o[1629] = i[1629];
  assign o[1628] = i[1628];
  assign o[1627] = i[1627];
  assign o[1626] = i[1626];
  assign o[1625] = i[1625];
  assign o[1624] = i[1624];
  assign o[1623] = i[1623];
  assign o[1622] = i[1622];
  assign o[1621] = i[1621];
  assign o[1620] = i[1620];
  assign o[1619] = i[1619];
  assign o[1618] = i[1618];
  assign o[1617] = i[1617];
  assign o[1616] = i[1616];
  assign o[1615] = i[1615];
  assign o[1614] = i[1614];
  assign o[1613] = i[1613];
  assign o[1612] = i[1612];
  assign o[1611] = i[1611];
  assign o[1610] = i[1610];
  assign o[1609] = i[1609];
  assign o[1608] = i[1608];
  assign o[1607] = i[1607];
  assign o[1606] = i[1606];
  assign o[1605] = i[1605];
  assign o[1604] = i[1604];
  assign o[1603] = i[1603];
  assign o[1602] = i[1602];
  assign o[1601] = i[1601];
  assign o[1600] = i[1600];
  assign o[1599] = i[1599];
  assign o[1598] = i[1598];
  assign o[1597] = i[1597];
  assign o[1596] = i[1596];
  assign o[1595] = i[1595];
  assign o[1594] = i[1594];
  assign o[1593] = i[1593];
  assign o[1592] = i[1592];
  assign o[1591] = i[1591];
  assign o[1590] = i[1590];
  assign o[1589] = i[1589];
  assign o[1588] = i[1588];
  assign o[1587] = i[1587];
  assign o[1586] = i[1586];
  assign o[1585] = i[1585];
  assign o[1584] = i[1584];
  assign o[1583] = i[1583];
  assign o[1582] = i[1582];
  assign o[1581] = i[1581];
  assign o[1580] = i[1580];
  assign o[1579] = i[1579];
  assign o[1578] = i[1578];
  assign o[1577] = i[1577];
  assign o[1576] = i[1576];
  assign o[1575] = i[1575];
  assign o[1574] = i[1574];
  assign o[1573] = i[1573];
  assign o[1572] = i[1572];
  assign o[1571] = i[1571];
  assign o[1570] = i[1570];
  assign o[1569] = i[1569];
  assign o[1568] = i[1568];
  assign o[1567] = i[1567];
  assign o[1566] = i[1566];
  assign o[1565] = i[1565];
  assign o[1564] = i[1564];
  assign o[1563] = i[1563];
  assign o[1562] = i[1562];
  assign o[1561] = i[1561];
  assign o[1560] = i[1560];
  assign o[1559] = i[1559];
  assign o[1558] = i[1558];
  assign o[1557] = i[1557];
  assign o[1556] = i[1556];
  assign o[1555] = i[1555];
  assign o[1554] = i[1554];
  assign o[1553] = i[1553];
  assign o[1552] = i[1552];
  assign o[1551] = i[1551];
  assign o[1550] = i[1550];
  assign o[1549] = i[1549];
  assign o[1548] = i[1548];
  assign o[1547] = i[1547];
  assign o[1546] = i[1546];
  assign o[1545] = i[1545];
  assign o[1544] = i[1544];
  assign o[1543] = i[1543];
  assign o[1542] = i[1542];
  assign o[1541] = i[1541];
  assign o[1540] = i[1540];
  assign o[1539] = i[1539];
  assign o[1538] = i[1538];
  assign o[1537] = i[1537];
  assign o[1536] = i[1536];
  assign o[1535] = i[1535];
  assign o[1534] = i[1534];
  assign o[1533] = i[1533];
  assign o[1532] = i[1532];
  assign o[1531] = i[1531];
  assign o[1530] = i[1530];
  assign o[1529] = i[1529];
  assign o[1528] = i[1528];
  assign o[1527] = i[1527];
  assign o[1526] = i[1526];
  assign o[1525] = i[1525];
  assign o[1524] = i[1524];
  assign o[1523] = i[1523];
  assign o[1522] = i[1522];
  assign o[1521] = i[1521];
  assign o[1520] = i[1520];
  assign o[1519] = i[1519];
  assign o[1518] = i[1518];
  assign o[1517] = i[1517];
  assign o[1516] = i[1516];
  assign o[1515] = i[1515];
  assign o[1514] = i[1514];
  assign o[1513] = i[1513];
  assign o[1512] = i[1512];
  assign o[1511] = i[1511];
  assign o[1510] = i[1510];
  assign o[1509] = i[1509];
  assign o[1508] = i[1508];
  assign o[1507] = i[1507];
  assign o[1506] = i[1506];
  assign o[1505] = i[1505];
  assign o[1504] = i[1504];
  assign o[1503] = i[1503];
  assign o[1502] = i[1502];
  assign o[1501] = i[1501];
  assign o[1500] = i[1500];
  assign o[1499] = i[1499];
  assign o[1498] = i[1498];
  assign o[1497] = i[1497];
  assign o[1496] = i[1496];
  assign o[1495] = i[1495];
  assign o[1494] = i[1494];
  assign o[1493] = i[1493];
  assign o[1492] = i[1492];
  assign o[1491] = i[1491];
  assign o[1490] = i[1490];
  assign o[1489] = i[1489];
  assign o[1488] = i[1488];
  assign o[1487] = i[1487];
  assign o[1486] = i[1486];
  assign o[1485] = i[1485];
  assign o[1484] = i[1484];
  assign o[1483] = i[1483];
  assign o[1482] = i[1482];
  assign o[1481] = i[1481];
  assign o[1480] = i[1480];
  assign o[1479] = i[1479];
  assign o[1478] = i[1478];
  assign o[1477] = i[1477];
  assign o[1476] = i[1476];
  assign o[1475] = i[1475];
  assign o[1474] = i[1474];
  assign o[1473] = i[1473];
  assign o[1472] = i[1472];
  assign o[1471] = i[1471];
  assign o[1470] = i[1470];
  assign o[1469] = i[1469];
  assign o[1468] = i[1468];
  assign o[1467] = i[1467];
  assign o[1466] = i[1466];
  assign o[1465] = i[1465];
  assign o[1464] = i[1464];
  assign o[1463] = i[1463];
  assign o[1462] = i[1462];
  assign o[1461] = i[1461];
  assign o[1460] = i[1460];
  assign o[1459] = i[1459];
  assign o[1458] = i[1458];
  assign o[1457] = i[1457];
  assign o[1456] = i[1456];
  assign o[1455] = i[1455];
  assign o[1454] = i[1454];
  assign o[1453] = i[1453];
  assign o[1452] = i[1452];
  assign o[1451] = i[1451];
  assign o[1450] = i[1450];
  assign o[1449] = i[1449];
  assign o[1448] = i[1448];
  assign o[1447] = i[1447];
  assign o[1446] = i[1446];
  assign o[1445] = i[1445];
  assign o[1444] = i[1444];
  assign o[1443] = i[1443];
  assign o[1442] = i[1442];
  assign o[1441] = i[1441];
  assign o[1440] = i[1440];
  assign o[1439] = i[1439];
  assign o[1438] = i[1438];
  assign o[1437] = i[1437];
  assign o[1436] = i[1436];
  assign o[1435] = i[1435];
  assign o[1434] = i[1434];
  assign o[1433] = i[1433];
  assign o[1432] = i[1432];
  assign o[1431] = i[1431];
  assign o[1430] = i[1430];
  assign o[1429] = i[1429];
  assign o[1428] = i[1428];
  assign o[1427] = i[1427];
  assign o[1426] = i[1426];
  assign o[1425] = i[1425];
  assign o[1424] = i[1424];
  assign o[1423] = i[1423];
  assign o[1422] = i[1422];
  assign o[1421] = i[1421];
  assign o[1420] = i[1420];
  assign o[1419] = i[1419];
  assign o[1418] = i[1418];
  assign o[1417] = i[1417];
  assign o[1416] = i[1416];
  assign o[1415] = i[1415];
  assign o[1414] = i[1414];
  assign o[1413] = i[1413];
  assign o[1412] = i[1412];
  assign o[1411] = i[1411];
  assign o[1410] = i[1410];
  assign o[1409] = i[1409];
  assign o[1408] = i[1408];
  assign o[1407] = i[1407];
  assign o[1406] = i[1406];
  assign o[1405] = i[1405];
  assign o[1404] = i[1404];
  assign o[1403] = i[1403];
  assign o[1402] = i[1402];
  assign o[1401] = i[1401];
  assign o[1400] = i[1400];
  assign o[1399] = i[1399];
  assign o[1398] = i[1398];
  assign o[1397] = i[1397];
  assign o[1396] = i[1396];
  assign o[1395] = i[1395];
  assign o[1394] = i[1394];
  assign o[1393] = i[1393];
  assign o[1392] = i[1392];
  assign o[1391] = i[1391];
  assign o[1390] = i[1390];
  assign o[1389] = i[1389];
  assign o[1388] = i[1388];
  assign o[1387] = i[1387];
  assign o[1386] = i[1386];
  assign o[1385] = i[1385];
  assign o[1384] = i[1384];
  assign o[1383] = i[1383];
  assign o[1382] = i[1382];
  assign o[1381] = i[1381];
  assign o[1380] = i[1380];
  assign o[1379] = i[1379];
  assign o[1378] = i[1378];
  assign o[1377] = i[1377];
  assign o[1376] = i[1376];
  assign o[1375] = i[1375];
  assign o[1374] = i[1374];
  assign o[1373] = i[1373];
  assign o[1372] = i[1372];
  assign o[1371] = i[1371];
  assign o[1370] = i[1370];
  assign o[1369] = i[1369];
  assign o[1368] = i[1368];
  assign o[1367] = i[1367];
  assign o[1366] = i[1366];
  assign o[1365] = i[1365];
  assign o[1364] = i[1364];
  assign o[1363] = i[1363];
  assign o[1362] = i[1362];
  assign o[1361] = i[1361];
  assign o[1360] = i[1360];
  assign o[1359] = i[1359];
  assign o[1358] = i[1358];
  assign o[1357] = i[1357];
  assign o[1356] = i[1356];
  assign o[1355] = i[1355];
  assign o[1354] = i[1354];
  assign o[1353] = i[1353];
  assign o[1352] = i[1352];
  assign o[1351] = i[1351];
  assign o[1350] = i[1350];
  assign o[1349] = i[1349];
  assign o[1348] = i[1348];
  assign o[1347] = i[1347];
  assign o[1346] = i[1346];
  assign o[1345] = i[1345];
  assign o[1344] = i[1344];
  assign o[1343] = i[1343];
  assign o[1342] = i[1342];
  assign o[1341] = i[1341];
  assign o[1340] = i[1340];
  assign o[1339] = i[1339];
  assign o[1338] = i[1338];
  assign o[1337] = i[1337];
  assign o[1336] = i[1336];
  assign o[1335] = i[1335];
  assign o[1334] = i[1334];
  assign o[1333] = i[1333];
  assign o[1332] = i[1332];
  assign o[1331] = i[1331];
  assign o[1330] = i[1330];
  assign o[1329] = i[1329];
  assign o[1328] = i[1328];
  assign o[1327] = i[1327];
  assign o[1326] = i[1326];
  assign o[1325] = i[1325];
  assign o[1324] = i[1324];
  assign o[1323] = i[1323];
  assign o[1322] = i[1322];
  assign o[1321] = i[1321];
  assign o[1320] = i[1320];
  assign o[1319] = i[1319];
  assign o[1318] = i[1318];
  assign o[1317] = i[1317];
  assign o[1316] = i[1316];
  assign o[1315] = i[1315];
  assign o[1314] = i[1314];
  assign o[1313] = i[1313];
  assign o[1312] = i[1312];
  assign o[1311] = i[1311];
  assign o[1310] = i[1310];
  assign o[1309] = i[1309];
  assign o[1308] = i[1308];
  assign o[1307] = i[1307];
  assign o[1306] = i[1306];
  assign o[1305] = i[1305];
  assign o[1304] = i[1304];
  assign o[1303] = i[1303];
  assign o[1302] = i[1302];
  assign o[1301] = i[1301];
  assign o[1300] = i[1300];
  assign o[1299] = i[1299];
  assign o[1298] = i[1298];
  assign o[1297] = i[1297];
  assign o[1296] = i[1296];
  assign o[1295] = i[1295];
  assign o[1294] = i[1294];
  assign o[1293] = i[1293];
  assign o[1292] = i[1292];
  assign o[1291] = i[1291];
  assign o[1290] = i[1290];
  assign o[1289] = i[1289];
  assign o[1288] = i[1288];
  assign o[1287] = i[1287];
  assign o[1286] = i[1286];
  assign o[1285] = i[1285];
  assign o[1284] = i[1284];
  assign o[1283] = i[1283];
  assign o[1282] = i[1282];
  assign o[1281] = i[1281];
  assign o[1280] = i[1280];
  assign o[1279] = i[1279];
  assign o[1278] = i[1278];
  assign o[1277] = i[1277];
  assign o[1276] = i[1276];
  assign o[1275] = i[1275];
  assign o[1274] = i[1274];
  assign o[1273] = i[1273];
  assign o[1272] = i[1272];
  assign o[1271] = i[1271];
  assign o[1270] = i[1270];
  assign o[1269] = i[1269];
  assign o[1268] = i[1268];
  assign o[1267] = i[1267];
  assign o[1266] = i[1266];
  assign o[1265] = i[1265];
  assign o[1264] = i[1264];
  assign o[1263] = i[1263];
  assign o[1262] = i[1262];
  assign o[1261] = i[1261];
  assign o[1260] = i[1260];
  assign o[1259] = i[1259];
  assign o[1258] = i[1258];
  assign o[1257] = i[1257];
  assign o[1256] = i[1256];
  assign o[1255] = i[1255];
  assign o[1254] = i[1254];
  assign o[1253] = i[1253];
  assign o[1252] = i[1252];
  assign o[1251] = i[1251];
  assign o[1250] = i[1250];
  assign o[1249] = i[1249];
  assign o[1248] = i[1248];
  assign o[1247] = i[1247];
  assign o[1246] = i[1246];
  assign o[1245] = i[1245];
  assign o[1244] = i[1244];
  assign o[1243] = i[1243];
  assign o[1242] = i[1242];
  assign o[1241] = i[1241];
  assign o[1240] = i[1240];
  assign o[1239] = i[1239];
  assign o[1238] = i[1238];
  assign o[1237] = i[1237];
  assign o[1236] = i[1236];
  assign o[1235] = i[1235];
  assign o[1234] = i[1234];
  assign o[1233] = i[1233];
  assign o[1232] = i[1232];
  assign o[1231] = i[1231];
  assign o[1230] = i[1230];
  assign o[1229] = i[1229];
  assign o[1228] = i[1228];
  assign o[1227] = i[1227];
  assign o[1226] = i[1226];
  assign o[1225] = i[1225];
  assign o[1224] = i[1224];
  assign o[1223] = i[1223];
  assign o[1222] = i[1222];
  assign o[1221] = i[1221];
  assign o[1220] = i[1220];
  assign o[1219] = i[1219];
  assign o[1218] = i[1218];
  assign o[1217] = i[1217];
  assign o[1216] = i[1216];
  assign o[1215] = i[1215];
  assign o[1214] = i[1214];
  assign o[1213] = i[1213];
  assign o[1212] = i[1212];
  assign o[1211] = i[1211];
  assign o[1210] = i[1210];
  assign o[1209] = i[1209];
  assign o[1208] = i[1208];
  assign o[1207] = i[1207];
  assign o[1206] = i[1206];
  assign o[1205] = i[1205];
  assign o[1204] = i[1204];
  assign o[1203] = i[1203];
  assign o[1202] = i[1202];
  assign o[1201] = i[1201];
  assign o[1200] = i[1200];
  assign o[1199] = i[1199];
  assign o[1198] = i[1198];
  assign o[1197] = i[1197];
  assign o[1196] = i[1196];
  assign o[1195] = i[1195];
  assign o[1194] = i[1194];
  assign o[1193] = i[1193];
  assign o[1192] = i[1192];
  assign o[1191] = i[1191];
  assign o[1190] = i[1190];
  assign o[1189] = i[1189];
  assign o[1188] = i[1188];
  assign o[1187] = i[1187];
  assign o[1186] = i[1186];
  assign o[1185] = i[1185];
  assign o[1184] = i[1184];
  assign o[1183] = i[1183];
  assign o[1182] = i[1182];
  assign o[1181] = i[1181];
  assign o[1180] = i[1180];
  assign o[1179] = i[1179];
  assign o[1178] = i[1178];
  assign o[1177] = i[1177];
  assign o[1176] = i[1176];
  assign o[1175] = i[1175];
  assign o[1174] = i[1174];
  assign o[1173] = i[1173];
  assign o[1172] = i[1172];
  assign o[1171] = i[1171];
  assign o[1170] = i[1170];
  assign o[1169] = i[1169];
  assign o[1168] = i[1168];
  assign o[1167] = i[1167];
  assign o[1166] = i[1166];
  assign o[1165] = i[1165];
  assign o[1164] = i[1164];
  assign o[1163] = i[1163];
  assign o[1162] = i[1162];
  assign o[1161] = i[1161];
  assign o[1160] = i[1160];
  assign o[1159] = i[1159];
  assign o[1158] = i[1158];
  assign o[1157] = i[1157];
  assign o[1156] = i[1156];
  assign o[1155] = i[1155];
  assign o[1154] = i[1154];
  assign o[1153] = i[1153];
  assign o[1152] = i[1152];
  assign o[1151] = i[1151];
  assign o[1150] = i[1150];
  assign o[1149] = i[1149];
  assign o[1148] = i[1148];
  assign o[1147] = i[1147];
  assign o[1146] = i[1146];
  assign o[1145] = i[1145];
  assign o[1144] = i[1144];
  assign o[1143] = i[1143];
  assign o[1142] = i[1142];
  assign o[1141] = i[1141];
  assign o[1140] = i[1140];
  assign o[1139] = i[1139];
  assign o[1138] = i[1138];
  assign o[1137] = i[1137];
  assign o[1136] = i[1136];
  assign o[1135] = i[1135];
  assign o[1134] = i[1134];
  assign o[1133] = i[1133];
  assign o[1132] = i[1132];
  assign o[1131] = i[1131];
  assign o[1130] = i[1130];
  assign o[1129] = i[1129];
  assign o[1128] = i[1128];
  assign o[1127] = i[1127];
  assign o[1126] = i[1126];
  assign o[1125] = i[1125];
  assign o[1124] = i[1124];
  assign o[1123] = i[1123];
  assign o[1122] = i[1122];
  assign o[1121] = i[1121];
  assign o[1120] = i[1120];
  assign o[1119] = i[1119];
  assign o[1118] = i[1118];
  assign o[1117] = i[1117];
  assign o[1116] = i[1116];
  assign o[1115] = i[1115];
  assign o[1114] = i[1114];
  assign o[1113] = i[1113];
  assign o[1112] = i[1112];
  assign o[1111] = i[1111];
  assign o[1110] = i[1110];
  assign o[1109] = i[1109];
  assign o[1108] = i[1108];
  assign o[1107] = i[1107];
  assign o[1106] = i[1106];
  assign o[1105] = i[1105];
  assign o[1104] = i[1104];
  assign o[1103] = i[1103];
  assign o[1102] = i[1102];
  assign o[1101] = i[1101];
  assign o[1100] = i[1100];
  assign o[1099] = i[1099];
  assign o[1098] = i[1098];
  assign o[1097] = i[1097];
  assign o[1096] = i[1096];
  assign o[1095] = i[1095];
  assign o[1094] = i[1094];
  assign o[1093] = i[1093];
  assign o[1092] = i[1092];
  assign o[1091] = i[1091];
  assign o[1090] = i[1090];
  assign o[1089] = i[1089];
  assign o[1088] = i[1088];
  assign o[1087] = i[1087];
  assign o[1086] = i[1086];
  assign o[1085] = i[1085];
  assign o[1084] = i[1084];
  assign o[1083] = i[1083];
  assign o[1082] = i[1082];
  assign o[1081] = i[1081];
  assign o[1080] = i[1080];
  assign o[1079] = i[1079];
  assign o[1078] = i[1078];
  assign o[1077] = i[1077];
  assign o[1076] = i[1076];
  assign o[1075] = i[1075];
  assign o[1074] = i[1074];
  assign o[1073] = i[1073];
  assign o[1072] = i[1072];
  assign o[1071] = i[1071];
  assign o[1070] = i[1070];
  assign o[1069] = i[1069];
  assign o[1068] = i[1068];
  assign o[1067] = i[1067];
  assign o[1066] = i[1066];
  assign o[1065] = i[1065];
  assign o[1064] = i[1064];
  assign o[1063] = i[1063];
  assign o[1062] = i[1062];
  assign o[1061] = i[1061];
  assign o[1060] = i[1060];
  assign o[1059] = i[1059];
  assign o[1058] = i[1058];
  assign o[1057] = i[1057];
  assign o[1056] = i[1056];
  assign o[1055] = i[1055];
  assign o[1054] = i[1054];
  assign o[1053] = i[1053];
  assign o[1052] = i[1052];
  assign o[1051] = i[1051];
  assign o[1050] = i[1050];
  assign o[1049] = i[1049];
  assign o[1048] = i[1048];
  assign o[1047] = i[1047];
  assign o[1046] = i[1046];
  assign o[1045] = i[1045];
  assign o[1044] = i[1044];
  assign o[1043] = i[1043];
  assign o[1042] = i[1042];
  assign o[1041] = i[1041];
  assign o[1040] = i[1040];
  assign o[1039] = i[1039];
  assign o[1038] = i[1038];
  assign o[1037] = i[1037];
  assign o[1036] = i[1036];
  assign o[1035] = i[1035];
  assign o[1034] = i[1034];
  assign o[1033] = i[1033];
  assign o[1032] = i[1032];
  assign o[1031] = i[1031];
  assign o[1030] = i[1030];
  assign o[1029] = i[1029];
  assign o[1028] = i[1028];
  assign o[1027] = i[1027];
  assign o[1026] = i[1026];
  assign o[1025] = i[1025];
  assign o[1024] = i[1024];
  assign o[1023] = i[1023];
  assign o[1022] = i[1022];
  assign o[1021] = i[1021];
  assign o[1020] = i[1020];
  assign o[1019] = i[1019];
  assign o[1018] = i[1018];
  assign o[1017] = i[1017];
  assign o[1016] = i[1016];
  assign o[1015] = i[1015];
  assign o[1014] = i[1014];
  assign o[1013] = i[1013];
  assign o[1012] = i[1012];
  assign o[1011] = i[1011];
  assign o[1010] = i[1010];
  assign o[1009] = i[1009];
  assign o[1008] = i[1008];
  assign o[1007] = i[1007];
  assign o[1006] = i[1006];
  assign o[1005] = i[1005];
  assign o[1004] = i[1004];
  assign o[1003] = i[1003];
  assign o[1002] = i[1002];
  assign o[1001] = i[1001];
  assign o[1000] = i[1000];
  assign o[999] = i[999];
  assign o[998] = i[998];
  assign o[997] = i[997];
  assign o[996] = i[996];
  assign o[995] = i[995];
  assign o[994] = i[994];
  assign o[993] = i[993];
  assign o[992] = i[992];
  assign o[991] = i[991];
  assign o[990] = i[990];
  assign o[989] = i[989];
  assign o[988] = i[988];
  assign o[987] = i[987];
  assign o[986] = i[986];
  assign o[985] = i[985];
  assign o[984] = i[984];
  assign o[983] = i[983];
  assign o[982] = i[982];
  assign o[981] = i[981];
  assign o[980] = i[980];
  assign o[979] = i[979];
  assign o[978] = i[978];
  assign o[977] = i[977];
  assign o[976] = i[976];
  assign o[975] = i[975];
  assign o[974] = i[974];
  assign o[973] = i[973];
  assign o[972] = i[972];
  assign o[971] = i[971];
  assign o[970] = i[970];
  assign o[969] = i[969];
  assign o[968] = i[968];
  assign o[967] = i[967];
  assign o[966] = i[966];
  assign o[965] = i[965];
  assign o[964] = i[964];
  assign o[963] = i[963];
  assign o[962] = i[962];
  assign o[961] = i[961];
  assign o[960] = i[960];
  assign o[959] = i[959];
  assign o[958] = i[958];
  assign o[957] = i[957];
  assign o[956] = i[956];
  assign o[955] = i[955];
  assign o[954] = i[954];
  assign o[953] = i[953];
  assign o[952] = i[952];
  assign o[951] = i[951];
  assign o[950] = i[950];
  assign o[949] = i[949];
  assign o[948] = i[948];
  assign o[947] = i[947];
  assign o[946] = i[946];
  assign o[945] = i[945];
  assign o[944] = i[944];
  assign o[943] = i[943];
  assign o[942] = i[942];
  assign o[941] = i[941];
  assign o[940] = i[940];
  assign o[939] = i[939];
  assign o[938] = i[938];
  assign o[937] = i[937];
  assign o[936] = i[936];
  assign o[935] = i[935];
  assign o[934] = i[934];
  assign o[933] = i[933];
  assign o[932] = i[932];
  assign o[931] = i[931];
  assign o[930] = i[930];
  assign o[929] = i[929];
  assign o[928] = i[928];
  assign o[927] = i[927];
  assign o[926] = i[926];
  assign o[925] = i[925];
  assign o[924] = i[924];
  assign o[923] = i[923];
  assign o[922] = i[922];
  assign o[921] = i[921];
  assign o[920] = i[920];
  assign o[919] = i[919];
  assign o[918] = i[918];
  assign o[917] = i[917];
  assign o[916] = i[916];
  assign o[915] = i[915];
  assign o[914] = i[914];
  assign o[913] = i[913];
  assign o[912] = i[912];
  assign o[911] = i[911];
  assign o[910] = i[910];
  assign o[909] = i[909];
  assign o[908] = i[908];
  assign o[907] = i[907];
  assign o[906] = i[906];
  assign o[905] = i[905];
  assign o[904] = i[904];
  assign o[903] = i[903];
  assign o[902] = i[902];
  assign o[901] = i[901];
  assign o[900] = i[900];
  assign o[899] = i[899];
  assign o[898] = i[898];
  assign o[897] = i[897];
  assign o[896] = i[896];
  assign o[895] = i[895];
  assign o[894] = i[894];
  assign o[893] = i[893];
  assign o[892] = i[892];
  assign o[891] = i[891];
  assign o[890] = i[890];
  assign o[889] = i[889];
  assign o[888] = i[888];
  assign o[887] = i[887];
  assign o[886] = i[886];
  assign o[885] = i[885];
  assign o[884] = i[884];
  assign o[883] = i[883];
  assign o[882] = i[882];
  assign o[881] = i[881];
  assign o[880] = i[880];
  assign o[879] = i[879];
  assign o[878] = i[878];
  assign o[877] = i[877];
  assign o[876] = i[876];
  assign o[875] = i[875];
  assign o[874] = i[874];
  assign o[873] = i[873];
  assign o[872] = i[872];
  assign o[871] = i[871];
  assign o[870] = i[870];
  assign o[869] = i[869];
  assign o[868] = i[868];
  assign o[867] = i[867];
  assign o[866] = i[866];
  assign o[865] = i[865];
  assign o[864] = i[864];
  assign o[863] = i[863];
  assign o[862] = i[862];
  assign o[861] = i[861];
  assign o[860] = i[860];
  assign o[859] = i[859];
  assign o[858] = i[858];
  assign o[857] = i[857];
  assign o[856] = i[856];
  assign o[855] = i[855];
  assign o[854] = i[854];
  assign o[853] = i[853];
  assign o[852] = i[852];
  assign o[851] = i[851];
  assign o[850] = i[850];
  assign o[849] = i[849];
  assign o[848] = i[848];
  assign o[847] = i[847];
  assign o[846] = i[846];
  assign o[845] = i[845];
  assign o[844] = i[844];
  assign o[843] = i[843];
  assign o[842] = i[842];
  assign o[841] = i[841];
  assign o[840] = i[840];
  assign o[839] = i[839];
  assign o[838] = i[838];
  assign o[837] = i[837];
  assign o[836] = i[836];
  assign o[835] = i[835];
  assign o[834] = i[834];
  assign o[833] = i[833];
  assign o[832] = i[832];
  assign o[831] = i[831];
  assign o[830] = i[830];
  assign o[829] = i[829];
  assign o[828] = i[828];
  assign o[827] = i[827];
  assign o[826] = i[826];
  assign o[825] = i[825];
  assign o[824] = i[824];
  assign o[823] = i[823];
  assign o[822] = i[822];
  assign o[821] = i[821];
  assign o[820] = i[820];
  assign o[819] = i[819];
  assign o[818] = i[818];
  assign o[817] = i[817];
  assign o[816] = i[816];
  assign o[815] = i[815];
  assign o[814] = i[814];
  assign o[813] = i[813];
  assign o[812] = i[812];
  assign o[811] = i[811];
  assign o[810] = i[810];
  assign o[809] = i[809];
  assign o[808] = i[808];
  assign o[807] = i[807];
  assign o[806] = i[806];
  assign o[805] = i[805];
  assign o[804] = i[804];
  assign o[803] = i[803];
  assign o[802] = i[802];
  assign o[801] = i[801];
  assign o[800] = i[800];
  assign o[799] = i[799];
  assign o[798] = i[798];
  assign o[797] = i[797];
  assign o[796] = i[796];
  assign o[795] = i[795];
  assign o[794] = i[794];
  assign o[793] = i[793];
  assign o[792] = i[792];
  assign o[791] = i[791];
  assign o[790] = i[790];
  assign o[789] = i[789];
  assign o[788] = i[788];
  assign o[787] = i[787];
  assign o[786] = i[786];
  assign o[785] = i[785];
  assign o[784] = i[784];
  assign o[783] = i[783];
  assign o[782] = i[782];
  assign o[781] = i[781];
  assign o[780] = i[780];
  assign o[779] = i[779];
  assign o[778] = i[778];
  assign o[777] = i[777];
  assign o[776] = i[776];
  assign o[775] = i[775];
  assign o[774] = i[774];
  assign o[773] = i[773];
  assign o[772] = i[772];
  assign o[771] = i[771];
  assign o[770] = i[770];
  assign o[769] = i[769];
  assign o[768] = i[768];
  assign o[767] = i[767];
  assign o[766] = i[766];
  assign o[765] = i[765];
  assign o[764] = i[764];
  assign o[763] = i[763];
  assign o[762] = i[762];
  assign o[761] = i[761];
  assign o[760] = i[760];
  assign o[759] = i[759];
  assign o[758] = i[758];
  assign o[757] = i[757];
  assign o[756] = i[756];
  assign o[755] = i[755];
  assign o[754] = i[754];
  assign o[753] = i[753];
  assign o[752] = i[752];
  assign o[751] = i[751];
  assign o[750] = i[750];
  assign o[749] = i[749];
  assign o[748] = i[748];
  assign o[747] = i[747];
  assign o[746] = i[746];
  assign o[745] = i[745];
  assign o[744] = i[744];
  assign o[743] = i[743];
  assign o[742] = i[742];
  assign o[741] = i[741];
  assign o[740] = i[740];
  assign o[739] = i[739];
  assign o[738] = i[738];
  assign o[737] = i[737];
  assign o[736] = i[736];
  assign o[735] = i[735];
  assign o[734] = i[734];
  assign o[733] = i[733];
  assign o[732] = i[732];
  assign o[731] = i[731];
  assign o[730] = i[730];
  assign o[729] = i[729];
  assign o[728] = i[728];
  assign o[727] = i[727];
  assign o[726] = i[726];
  assign o[725] = i[725];
  assign o[724] = i[724];
  assign o[723] = i[723];
  assign o[722] = i[722];
  assign o[721] = i[721];
  assign o[720] = i[720];
  assign o[719] = i[719];
  assign o[718] = i[718];
  assign o[717] = i[717];
  assign o[716] = i[716];
  assign o[715] = i[715];
  assign o[714] = i[714];
  assign o[713] = i[713];
  assign o[712] = i[712];
  assign o[711] = i[711];
  assign o[710] = i[710];
  assign o[709] = i[709];
  assign o[708] = i[708];
  assign o[707] = i[707];
  assign o[706] = i[706];
  assign o[705] = i[705];
  assign o[704] = i[704];
  assign o[703] = i[703];
  assign o[702] = i[702];
  assign o[701] = i[701];
  assign o[700] = i[700];
  assign o[699] = i[699];
  assign o[698] = i[698];
  assign o[697] = i[697];
  assign o[696] = i[696];
  assign o[695] = i[695];
  assign o[694] = i[694];
  assign o[693] = i[693];
  assign o[692] = i[692];
  assign o[691] = i[691];
  assign o[690] = i[690];
  assign o[689] = i[689];
  assign o[688] = i[688];
  assign o[687] = i[687];
  assign o[686] = i[686];
  assign o[685] = i[685];
  assign o[684] = i[684];
  assign o[683] = i[683];
  assign o[682] = i[682];
  assign o[681] = i[681];
  assign o[680] = i[680];
  assign o[679] = i[679];
  assign o[678] = i[678];
  assign o[677] = i[677];
  assign o[676] = i[676];
  assign o[675] = i[675];
  assign o[674] = i[674];
  assign o[673] = i[673];
  assign o[672] = i[672];
  assign o[671] = i[671];
  assign o[670] = i[670];
  assign o[669] = i[669];
  assign o[668] = i[668];
  assign o[667] = i[667];
  assign o[666] = i[666];
  assign o[665] = i[665];
  assign o[664] = i[664];
  assign o[663] = i[663];
  assign o[662] = i[662];
  assign o[661] = i[661];
  assign o[660] = i[660];
  assign o[659] = i[659];
  assign o[658] = i[658];
  assign o[657] = i[657];
  assign o[656] = i[656];
  assign o[655] = i[655];
  assign o[654] = i[654];
  assign o[653] = i[653];
  assign o[652] = i[652];
  assign o[651] = i[651];
  assign o[650] = i[650];
  assign o[649] = i[649];
  assign o[648] = i[648];
  assign o[647] = i[647];
  assign o[646] = i[646];
  assign o[645] = i[645];
  assign o[644] = i[644];
  assign o[643] = i[643];
  assign o[642] = i[642];
  assign o[641] = i[641];
  assign o[640] = i[640];
  assign o[639] = i[639];
  assign o[638] = i[638];
  assign o[637] = i[637];
  assign o[636] = i[636];
  assign o[635] = i[635];
  assign o[634] = i[634];
  assign o[633] = i[633];
  assign o[632] = i[632];
  assign o[631] = i[631];
  assign o[630] = i[630];
  assign o[629] = i[629];
  assign o[628] = i[628];
  assign o[627] = i[627];
  assign o[626] = i[626];
  assign o[625] = i[625];
  assign o[624] = i[624];
  assign o[623] = i[623];
  assign o[622] = i[622];
  assign o[621] = i[621];
  assign o[620] = i[620];
  assign o[619] = i[619];
  assign o[618] = i[618];
  assign o[617] = i[617];
  assign o[616] = i[616];
  assign o[615] = i[615];
  assign o[614] = i[614];
  assign o[613] = i[613];
  assign o[612] = i[612];
  assign o[611] = i[611];
  assign o[610] = i[610];
  assign o[609] = i[609];
  assign o[608] = i[608];
  assign o[607] = i[607];
  assign o[606] = i[606];
  assign o[605] = i[605];
  assign o[604] = i[604];
  assign o[603] = i[603];
  assign o[602] = i[602];
  assign o[601] = i[601];
  assign o[600] = i[600];
  assign o[599] = i[599];
  assign o[598] = i[598];
  assign o[597] = i[597];
  assign o[596] = i[596];
  assign o[595] = i[595];
  assign o[594] = i[594];
  assign o[593] = i[593];
  assign o[592] = i[592];
  assign o[591] = i[591];
  assign o[590] = i[590];
  assign o[589] = i[589];
  assign o[588] = i[588];
  assign o[587] = i[587];
  assign o[586] = i[586];
  assign o[585] = i[585];
  assign o[584] = i[584];
  assign o[583] = i[583];
  assign o[582] = i[582];
  assign o[581] = i[581];
  assign o[580] = i[580];
  assign o[579] = i[579];
  assign o[578] = i[578];
  assign o[577] = i[577];
  assign o[576] = i[576];
  assign o[575] = i[575];
  assign o[574] = i[574];
  assign o[573] = i[573];
  assign o[572] = i[572];
  assign o[571] = i[571];
  assign o[570] = i[570];
  assign o[569] = i[569];
  assign o[568] = i[568];
  assign o[567] = i[567];
  assign o[566] = i[566];
  assign o[565] = i[565];
  assign o[564] = i[564];
  assign o[563] = i[563];
  assign o[562] = i[562];
  assign o[561] = i[561];
  assign o[560] = i[560];
  assign o[559] = i[559];
  assign o[558] = i[558];
  assign o[557] = i[557];
  assign o[556] = i[556];
  assign o[555] = i[555];
  assign o[554] = i[554];
  assign o[553] = i[553];
  assign o[552] = i[552];
  assign o[551] = i[551];
  assign o[550] = i[550];
  assign o[549] = i[549];
  assign o[548] = i[548];
  assign o[547] = i[547];
  assign o[546] = i[546];
  assign o[545] = i[545];
  assign o[544] = i[544];
  assign o[543] = i[543];
  assign o[542] = i[542];
  assign o[541] = i[541];
  assign o[540] = i[540];
  assign o[539] = i[539];
  assign o[538] = i[538];
  assign o[537] = i[537];
  assign o[536] = i[536];
  assign o[535] = i[535];
  assign o[534] = i[534];
  assign o[533] = i[533];
  assign o[532] = i[532];
  assign o[531] = i[531];
  assign o[530] = i[530];
  assign o[529] = i[529];
  assign o[528] = i[528];
  assign o[527] = i[527];
  assign o[526] = i[526];
  assign o[525] = i[525];
  assign o[524] = i[524];
  assign o[523] = i[523];
  assign o[522] = i[522];
  assign o[521] = i[521];
  assign o[520] = i[520];
  assign o[519] = i[519];
  assign o[518] = i[518];
  assign o[517] = i[517];
  assign o[516] = i[516];
  assign o[515] = i[515];
  assign o[514] = i[514];
  assign o[513] = i[513];
  assign o[512] = i[512];
  assign o[511] = i[511];
  assign o[510] = i[510];
  assign o[509] = i[509];
  assign o[508] = i[508];
  assign o[507] = i[507];
  assign o[506] = i[506];
  assign o[505] = i[505];
  assign o[504] = i[504];
  assign o[503] = i[503];
  assign o[502] = i[502];
  assign o[501] = i[501];
  assign o[500] = i[500];
  assign o[499] = i[499];
  assign o[498] = i[498];
  assign o[497] = i[497];
  assign o[496] = i[496];
  assign o[495] = i[495];
  assign o[494] = i[494];
  assign o[493] = i[493];
  assign o[492] = i[492];
  assign o[491] = i[491];
  assign o[490] = i[490];
  assign o[489] = i[489];
  assign o[488] = i[488];
  assign o[487] = i[487];
  assign o[486] = i[486];
  assign o[485] = i[485];
  assign o[484] = i[484];
  assign o[483] = i[483];
  assign o[482] = i[482];
  assign o[481] = i[481];
  assign o[480] = i[480];
  assign o[479] = i[479];
  assign o[478] = i[478];
  assign o[477] = i[477];
  assign o[476] = i[476];
  assign o[475] = i[475];
  assign o[474] = i[474];
  assign o[473] = i[473];
  assign o[472] = i[472];
  assign o[471] = i[471];
  assign o[470] = i[470];
  assign o[469] = i[469];
  assign o[468] = i[468];
  assign o[467] = i[467];
  assign o[466] = i[466];
  assign o[465] = i[465];
  assign o[464] = i[464];
  assign o[463] = i[463];
  assign o[462] = i[462];
  assign o[461] = i[461];
  assign o[460] = i[460];
  assign o[459] = i[459];
  assign o[458] = i[458];
  assign o[457] = i[457];
  assign o[456] = i[456];
  assign o[455] = i[455];
  assign o[454] = i[454];
  assign o[453] = i[453];
  assign o[452] = i[452];
  assign o[451] = i[451];
  assign o[450] = i[450];
  assign o[449] = i[449];
  assign o[448] = i[448];
  assign o[447] = i[447];
  assign o[446] = i[446];
  assign o[445] = i[445];
  assign o[444] = i[444];
  assign o[443] = i[443];
  assign o[442] = i[442];
  assign o[441] = i[441];
  assign o[440] = i[440];
  assign o[439] = i[439];
  assign o[438] = i[438];
  assign o[437] = i[437];
  assign o[436] = i[436];
  assign o[435] = i[435];
  assign o[434] = i[434];
  assign o[433] = i[433];
  assign o[432] = i[432];
  assign o[431] = i[431];
  assign o[430] = i[430];
  assign o[429] = i[429];
  assign o[428] = i[428];
  assign o[427] = i[427];
  assign o[426] = i[426];
  assign o[425] = i[425];
  assign o[424] = i[424];
  assign o[423] = i[423];
  assign o[422] = i[422];
  assign o[421] = i[421];
  assign o[420] = i[420];
  assign o[419] = i[419];
  assign o[418] = i[418];
  assign o[417] = i[417];
  assign o[416] = i[416];
  assign o[415] = i[415];
  assign o[414] = i[414];
  assign o[413] = i[413];
  assign o[412] = i[412];
  assign o[411] = i[411];
  assign o[410] = i[410];
  assign o[409] = i[409];
  assign o[408] = i[408];
  assign o[407] = i[407];
  assign o[406] = i[406];
  assign o[405] = i[405];
  assign o[404] = i[404];
  assign o[403] = i[403];
  assign o[402] = i[402];
  assign o[401] = i[401];
  assign o[400] = i[400];
  assign o[399] = i[399];
  assign o[398] = i[398];
  assign o[397] = i[397];
  assign o[396] = i[396];
  assign o[395] = i[395];
  assign o[394] = i[394];
  assign o[393] = i[393];
  assign o[392] = i[392];
  assign o[391] = i[391];
  assign o[390] = i[390];
  assign o[389] = i[389];
  assign o[388] = i[388];
  assign o[387] = i[387];
  assign o[386] = i[386];
  assign o[385] = i[385];
  assign o[384] = i[384];
  assign o[383] = i[383];
  assign o[382] = i[382];
  assign o[381] = i[381];
  assign o[380] = i[380];
  assign o[379] = i[379];
  assign o[378] = i[378];
  assign o[377] = i[377];
  assign o[376] = i[376];
  assign o[375] = i[375];
  assign o[374] = i[374];
  assign o[373] = i[373];
  assign o[372] = i[372];
  assign o[371] = i[371];
  assign o[370] = i[370];
  assign o[369] = i[369];
  assign o[368] = i[368];
  assign o[367] = i[367];
  assign o[366] = i[366];
  assign o[365] = i[365];
  assign o[364] = i[364];
  assign o[363] = i[363];
  assign o[362] = i[362];
  assign o[361] = i[361];
  assign o[360] = i[360];
  assign o[359] = i[359];
  assign o[358] = i[358];
  assign o[357] = i[357];
  assign o[356] = i[356];
  assign o[355] = i[355];
  assign o[354] = i[354];
  assign o[353] = i[353];
  assign o[352] = i[352];
  assign o[351] = i[351];
  assign o[350] = i[350];
  assign o[349] = i[349];
  assign o[348] = i[348];
  assign o[347] = i[347];
  assign o[346] = i[346];
  assign o[345] = i[345];
  assign o[344] = i[344];
  assign o[343] = i[343];
  assign o[342] = i[342];
  assign o[341] = i[341];
  assign o[340] = i[340];
  assign o[339] = i[339];
  assign o[338] = i[338];
  assign o[337] = i[337];
  assign o[336] = i[336];
  assign o[335] = i[335];
  assign o[334] = i[334];
  assign o[333] = i[333];
  assign o[332] = i[332];
  assign o[331] = i[331];
  assign o[330] = i[330];
  assign o[329] = i[329];
  assign o[328] = i[328];
  assign o[327] = i[327];
  assign o[326] = i[326];
  assign o[325] = i[325];
  assign o[324] = i[324];
  assign o[323] = i[323];
  assign o[322] = i[322];
  assign o[321] = i[321];
  assign o[320] = i[320];
  assign o[319] = i[319];
  assign o[318] = i[318];
  assign o[317] = i[317];
  assign o[316] = i[316];
  assign o[315] = i[315];
  assign o[314] = i[314];
  assign o[313] = i[313];
  assign o[312] = i[312];
  assign o[311] = i[311];
  assign o[310] = i[310];
  assign o[309] = i[309];
  assign o[308] = i[308];
  assign o[307] = i[307];
  assign o[306] = i[306];
  assign o[305] = i[305];
  assign o[304] = i[304];
  assign o[303] = i[303];
  assign o[302] = i[302];
  assign o[301] = i[301];
  assign o[300] = i[300];
  assign o[299] = i[299];
  assign o[298] = i[298];
  assign o[297] = i[297];
  assign o[296] = i[296];
  assign o[295] = i[295];
  assign o[294] = i[294];
  assign o[293] = i[293];
  assign o[292] = i[292];
  assign o[291] = i[291];
  assign o[290] = i[290];
  assign o[289] = i[289];
  assign o[288] = i[288];
  assign o[287] = i[287];
  assign o[286] = i[286];
  assign o[285] = i[285];
  assign o[284] = i[284];
  assign o[283] = i[283];
  assign o[282] = i[282];
  assign o[281] = i[281];
  assign o[280] = i[280];
  assign o[279] = i[279];
  assign o[278] = i[278];
  assign o[277] = i[277];
  assign o[276] = i[276];
  assign o[275] = i[275];
  assign o[274] = i[274];
  assign o[273] = i[273];
  assign o[272] = i[272];
  assign o[271] = i[271];
  assign o[270] = i[270];
  assign o[269] = i[269];
  assign o[268] = i[268];
  assign o[267] = i[267];
  assign o[266] = i[266];
  assign o[265] = i[265];
  assign o[264] = i[264];
  assign o[263] = i[263];
  assign o[262] = i[262];
  assign o[261] = i[261];
  assign o[260] = i[260];
  assign o[259] = i[259];
  assign o[258] = i[258];
  assign o[257] = i[257];
  assign o[256] = i[256];
  assign o[255] = i[255];
  assign o[254] = i[254];
  assign o[253] = i[253];
  assign o[252] = i[252];
  assign o[251] = i[251];
  assign o[250] = i[250];
  assign o[249] = i[249];
  assign o[248] = i[248];
  assign o[247] = i[247];
  assign o[246] = i[246];
  assign o[245] = i[245];
  assign o[244] = i[244];
  assign o[243] = i[243];
  assign o[242] = i[242];
  assign o[241] = i[241];
  assign o[240] = i[240];
  assign o[239] = i[239];
  assign o[238] = i[238];
  assign o[237] = i[237];
  assign o[236] = i[236];
  assign o[235] = i[235];
  assign o[234] = i[234];
  assign o[233] = i[233];
  assign o[232] = i[232];
  assign o[231] = i[231];
  assign o[230] = i[230];
  assign o[229] = i[229];
  assign o[228] = i[228];
  assign o[227] = i[227];
  assign o[226] = i[226];
  assign o[225] = i[225];
  assign o[224] = i[224];
  assign o[223] = i[223];
  assign o[222] = i[222];
  assign o[221] = i[221];
  assign o[220] = i[220];
  assign o[219] = i[219];
  assign o[218] = i[218];
  assign o[217] = i[217];
  assign o[216] = i[216];
  assign o[215] = i[215];
  assign o[214] = i[214];
  assign o[213] = i[213];
  assign o[212] = i[212];
  assign o[211] = i[211];
  assign o[210] = i[210];
  assign o[209] = i[209];
  assign o[208] = i[208];
  assign o[207] = i[207];
  assign o[206] = i[206];
  assign o[205] = i[205];
  assign o[204] = i[204];
  assign o[203] = i[203];
  assign o[202] = i[202];
  assign o[201] = i[201];
  assign o[200] = i[200];
  assign o[199] = i[199];
  assign o[198] = i[198];
  assign o[197] = i[197];
  assign o[196] = i[196];
  assign o[195] = i[195];
  assign o[194] = i[194];
  assign o[193] = i[193];
  assign o[192] = i[192];
  assign o[191] = i[191];
  assign o[190] = i[190];
  assign o[189] = i[189];
  assign o[188] = i[188];
  assign o[187] = i[187];
  assign o[186] = i[186];
  assign o[185] = i[185];
  assign o[184] = i[184];
  assign o[183] = i[183];
  assign o[182] = i[182];
  assign o[181] = i[181];
  assign o[180] = i[180];
  assign o[179] = i[179];
  assign o[178] = i[178];
  assign o[177] = i[177];
  assign o[176] = i[176];
  assign o[175] = i[175];
  assign o[174] = i[174];
  assign o[173] = i[173];
  assign o[172] = i[172];
  assign o[171] = i[171];
  assign o[170] = i[170];
  assign o[169] = i[169];
  assign o[168] = i[168];
  assign o[167] = i[167];
  assign o[166] = i[166];
  assign o[165] = i[165];
  assign o[164] = i[164];
  assign o[163] = i[163];
  assign o[162] = i[162];
  assign o[161] = i[161];
  assign o[160] = i[160];
  assign o[159] = i[159];
  assign o[158] = i[158];
  assign o[157] = i[157];
  assign o[156] = i[156];
  assign o[155] = i[155];
  assign o[154] = i[154];
  assign o[153] = i[153];
  assign o[152] = i[152];
  assign o[151] = i[151];
  assign o[150] = i[150];
  assign o[149] = i[149];
  assign o[148] = i[148];
  assign o[147] = i[147];
  assign o[146] = i[146];
  assign o[145] = i[145];
  assign o[144] = i[144];
  assign o[143] = i[143];
  assign o[142] = i[142];
  assign o[141] = i[141];
  assign o[140] = i[140];
  assign o[139] = i[139];
  assign o[138] = i[138];
  assign o[137] = i[137];
  assign o[136] = i[136];
  assign o[135] = i[135];
  assign o[134] = i[134];
  assign o[133] = i[133];
  assign o[132] = i[132];
  assign o[131] = i[131];
  assign o[130] = i[130];
  assign o[129] = i[129];
  assign o[128] = i[128];
  assign o[127] = i[127];
  assign o[126] = i[126];
  assign o[125] = i[125];
  assign o[124] = i[124];
  assign o[123] = i[123];
  assign o[122] = i[122];
  assign o[121] = i[121];
  assign o[120] = i[120];
  assign o[119] = i[119];
  assign o[118] = i[118];
  assign o[117] = i[117];
  assign o[116] = i[116];
  assign o[115] = i[115];
  assign o[114] = i[114];
  assign o[113] = i[113];
  assign o[112] = i[112];
  assign o[111] = i[111];
  assign o[110] = i[110];
  assign o[109] = i[109];
  assign o[108] = i[108];
  assign o[107] = i[107];
  assign o[106] = i[106];
  assign o[105] = i[105];
  assign o[104] = i[104];
  assign o[103] = i[103];
  assign o[102] = i[102];
  assign o[101] = i[101];
  assign o[100] = i[100];
  assign o[99] = i[99];
  assign o[98] = i[98];
  assign o[97] = i[97];
  assign o[96] = i[96];
  assign o[95] = i[95];
  assign o[94] = i[94];
  assign o[93] = i[93];
  assign o[92] = i[92];
  assign o[91] = i[91];
  assign o[90] = i[90];
  assign o[89] = i[89];
  assign o[88] = i[88];
  assign o[87] = i[87];
  assign o[86] = i[86];
  assign o[85] = i[85];
  assign o[84] = i[84];
  assign o[83] = i[83];
  assign o[82] = i[82];
  assign o[81] = i[81];
  assign o[80] = i[80];
  assign o[79] = i[79];
  assign o[78] = i[78];
  assign o[77] = i[77];
  assign o[76] = i[76];
  assign o[75] = i[75];
  assign o[74] = i[74];
  assign o[73] = i[73];
  assign o[72] = i[72];
  assign o[71] = i[71];
  assign o[70] = i[70];
  assign o[69] = i[69];
  assign o[68] = i[68];
  assign o[67] = i[67];
  assign o[66] = i[66];
  assign o[65] = i[65];
  assign o[64] = i[64];
  assign o[63] = i[63];
  assign o[62] = i[62];
  assign o[61] = i[61];
  assign o[60] = i[60];
  assign o[59] = i[59];
  assign o[58] = i[58];
  assign o[57] = i[57];
  assign o[56] = i[56];
  assign o[55] = i[55];
  assign o[54] = i[54];
  assign o[53] = i[53];
  assign o[52] = i[52];
  assign o[51] = i[51];
  assign o[50] = i[50];
  assign o[49] = i[49];
  assign o[48] = i[48];
  assign o[47] = i[47];
  assign o[46] = i[46];
  assign o[45] = i[45];
  assign o[44] = i[44];
  assign o[43] = i[43];
  assign o[42] = i[42];
  assign o[41] = i[41];
  assign o[40] = i[40];
  assign o[39] = i[39];
  assign o[38] = i[38];
  assign o[37] = i[37];
  assign o[36] = i[36];
  assign o[35] = i[35];
  assign o[34] = i[34];
  assign o[33] = i[33];
  assign o[32] = i[32];
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule

