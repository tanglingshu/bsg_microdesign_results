

module top
(
  i,
  sel_oi_one_hot_i,
  o
);

  input [16383:0] i;
  input [16383:0] sel_oi_one_hot_i;
  output [16383:0] o;

  bsg_crossbar_o_by_i
  wrapper
  (
    .i(i),
    .sel_oi_one_hot_i(sel_oi_one_hot_i),
    .o(o)
  );


endmodule



module bsg_mux_one_hot_width_p128_els_p128
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [16383:0] data_i;
  input [127:0] sel_one_hot_i;
  output [127:0] data_o;
  wire [127:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
  N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,
  N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,
  N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,
  N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,
  N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,
  N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,
  N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,
  N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,
  N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,
  N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,
  N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,
  N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,
  N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,
  N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,
  N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,
  N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,
  N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
  N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,
  N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,
  N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,
  N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,
  N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,
  N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,
  N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,
  N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,
  N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,
  N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,
  N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,
  N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,
  N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,
  N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,
  N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,
  N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,
  N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,
  N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,
  N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,
  N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,
  N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,
  N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,
  N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,
  N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,
  N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,
  N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,
  N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,
  N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,
  N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,
  N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,
  N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,
  N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,
  N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,
  N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,
  N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,
  N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,
  N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,
  N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,
  N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,
  N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,
  N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,
  N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,
  N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,
  N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,
  N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,
  N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,
  N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,
  N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,
  N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,
  N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,
  N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,
  N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,
  N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,
  N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,
  N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,
  N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,
  N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,
  N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,
  N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,
  N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,
  N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,
  N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,
  N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,
  N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,
  N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,
  N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144,
  N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,
  N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,N2170,
  N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,N2184,
  N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197,
  N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,N2210,
  N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,N2224,
  N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,
  N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,
  N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,N2264,
  N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,
  N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290,
  N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302,N2303,N2304,
  N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,
  N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,
  N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,
  N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,
  N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2369,N2370,
  N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382,N2383,N2384,
  N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,N2394,N2395,N2396,N2397,
  N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407,N2408,N2409,N2410,
  N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422,N2423,N2424,
  N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,
  N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447,N2448,N2449,N2450,
  N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,N2460,N2461,N2462,N2463,N2464,
  N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,N2474,N2475,N2476,N2477,
  N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,N2488,N2489,N2490,
  N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,N2500,N2501,N2502,N2503,N2504,
  N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,N2514,N2515,N2516,N2517,
  N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528,N2529,N2530,
  N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539,N2540,N2541,N2542,N2543,N2544,
  N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2554,N2555,N2556,N2557,
  N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,N2567,N2568,N2569,N2570,
  N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579,N2580,N2581,N2582,N2583,N2584,
  N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,N2594,N2595,N2596,N2597,
  N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,N2609,N2610,
  N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,N2620,N2621,N2622,N2623,N2624,
  N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2637,
  N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,N2649,N2650,
  N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662,N2663,N2664,
  N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,
  N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,N2687,N2688,N2689,N2690,
  N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2704,
  N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,N2714,N2715,N2716,N2717,
  N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,N2727,N2728,N2729,N2730,
  N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,
  N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,N2754,N2755,N2756,N2757,
  N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,N2767,N2768,N2769,N2770,
  N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2779,N2780,N2781,N2782,N2783,N2784,
  N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793,N2794,N2795,N2796,N2797,
  N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,N2807,N2808,N2809,N2810,
  N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,N2819,N2820,N2821,N2822,N2823,N2824,
  N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,N2834,N2835,N2836,N2837,
  N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,N2847,N2848,N2849,N2850,
  N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,N2859,N2860,N2861,N2862,N2863,N2864,
  N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877,
  N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,N2887,N2888,N2889,N2890,
  N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,N2899,N2900,N2901,N2902,N2903,N2904,
  N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,N2917,
  N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,N2930,
  N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,N2939,N2940,N2941,N2942,N2943,N2944,
  N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952,N2953,N2954,N2955,N2956,N2957,
  N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2965,N2966,N2967,N2968,N2969,N2970,
  N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980,N2981,N2982,N2983,N2984,
  N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,
  N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,N3010,
  N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022,N3023,N3024,
  N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3036,N3037,
  N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,N3050,
  N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3062,N3063,N3064,
  N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,N3076,N3077,
  N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,N3090,
  N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,N3101,N3102,N3103,N3104,
  N3105,N3106,N3107,N3108,N3109,N3110,N3111,N3112,N3113,N3114,N3115,N3116,N3117,
  N3118,N3119,N3120,N3121,N3122,N3123,N3124,N3125,N3126,N3127,N3128,N3129,N3130,
  N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,N3139,N3140,N3141,N3142,N3143,N3144,
  N3145,N3146,N3147,N3148,N3149,N3150,N3151,N3152,N3153,N3154,N3155,N3156,N3157,
  N3158,N3159,N3160,N3161,N3162,N3163,N3164,N3165,N3166,N3167,N3168,N3169,N3170,
  N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,N3179,N3180,N3181,N3182,N3183,N3184,
  N3185,N3186,N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194,N3195,N3196,N3197,
  N3198,N3199,N3200,N3201,N3202,N3203,N3204,N3205,N3206,N3207,N3208,N3209,N3210,
  N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,N3220,N3221,N3222,N3223,N3224,
  N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,
  N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,N3249,N3250,
  N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,N3260,N3261,N3262,N3263,N3264,
  N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,
  N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,N3290,
  N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,N3300,N3301,N3302,N3303,N3304,
  N3305,N3306,N3307,N3308,N3309,N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,
  N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,N3330,
  N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,N3339,N3340,N3341,N3342,N3343,N3344,
  N3345,N3346,N3347,N3348,N3349,N3350,N3351,N3352,N3353,N3354,N3355,N3356,N3357,
  N3358,N3359,N3360,N3361,N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,N3370,
  N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,N3379,N3380,N3381,N3382,N3383,N3384,
  N3385,N3386,N3387,N3388,N3389,N3390,N3391,N3392,N3393,N3394,N3395,N3396,N3397,
  N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3408,N3409,N3410,
  N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,N3419,N3420,N3421,N3422,N3423,N3424,
  N3425,N3426,N3427,N3428,N3429,N3430,N3431,N3432,N3433,N3434,N3435,N3436,N3437,
  N3438,N3439,N3440,N3441,N3442,N3443,N3444,N3445,N3446,N3447,N3448,N3449,N3450,
  N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,N3459,N3460,N3461,N3462,N3463,N3464,
  N3465,N3466,N3467,N3468,N3469,N3470,N3471,N3472,N3473,N3474,N3475,N3476,N3477,
  N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,N3487,N3488,N3489,N3490,
  N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,N3499,N3500,N3501,N3502,N3503,N3504,
  N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,N3513,N3514,N3515,N3516,N3517,
  N3518,N3519,N3520,N3521,N3522,N3523,N3524,N3525,N3526,N3527,N3528,N3529,N3530,
  N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,N3539,N3540,N3541,N3542,N3543,N3544,
  N3545,N3546,N3547,N3548,N3549,N3550,N3551,N3552,N3553,N3554,N3555,N3556,N3557,
  N3558,N3559,N3560,N3561,N3562,N3563,N3564,N3565,N3566,N3567,N3568,N3569,N3570,
  N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,N3579,N3580,N3581,N3582,N3583,N3584,
  N3585,N3586,N3587,N3588,N3589,N3590,N3591,N3592,N3593,N3594,N3595,N3596,N3597,
  N3598,N3599,N3600,N3601,N3602,N3603,N3604,N3605,N3606,N3607,N3608,N3609,N3610,
  N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,N3619,N3620,N3621,N3622,N3623,N3624,
  N3625,N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3636,N3637,
  N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3646,N3647,N3648,N3649,N3650,
  N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,N3659,N3660,N3661,N3662,N3663,N3664,
  N3665,N3666,N3667,N3668,N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3676,N3677,
  N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685,N3686,N3687,N3688,N3689,N3690,
  N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,N3699,N3700,N3701,N3702,N3703,N3704,
  N3705,N3706,N3707,N3708,N3709,N3710,N3711,N3712,N3713,N3714,N3715,N3716,N3717,
  N3718,N3719,N3720,N3721,N3722,N3723,N3724,N3725,N3726,N3727,N3728,N3729,N3730,
  N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,N3739,N3740,N3741,N3742,N3743,N3744,
  N3745,N3746,N3747,N3748,N3749,N3750,N3751,N3752,N3753,N3754,N3755,N3756,N3757,
  N3758,N3759,N3760,N3761,N3762,N3763,N3764,N3765,N3766,N3767,N3768,N3769,N3770,
  N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,N3779,N3780,N3781,N3782,N3783,N3784,
  N3785,N3786,N3787,N3788,N3789,N3790,N3791,N3792,N3793,N3794,N3795,N3796,N3797,
  N3798,N3799,N3800,N3801,N3802,N3803,N3804,N3805,N3806,N3807,N3808,N3809,N3810,
  N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,N3819,N3820,N3821,N3822,N3823,N3824,
  N3825,N3826,N3827,N3828,N3829,N3830,N3831,N3832,N3833,N3834,N3835,N3836,N3837,
  N3838,N3839,N3840,N3841,N3842,N3843,N3844,N3845,N3846,N3847,N3848,N3849,N3850,
  N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,N3859,N3860,N3861,N3862,N3863,N3864,
  N3865,N3866,N3867,N3868,N3869,N3870,N3871,N3872,N3873,N3874,N3875,N3876,N3877,
  N3878,N3879,N3880,N3881,N3882,N3883,N3884,N3885,N3886,N3887,N3888,N3889,N3890,
  N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,N3899,N3900,N3901,N3902,N3903,N3904,
  N3905,N3906,N3907,N3908,N3909,N3910,N3911,N3912,N3913,N3914,N3915,N3916,N3917,
  N3918,N3919,N3920,N3921,N3922,N3923,N3924,N3925,N3926,N3927,N3928,N3929,N3930,
  N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,N3939,N3940,N3941,N3942,N3943,N3944,
  N3945,N3946,N3947,N3948,N3949,N3950,N3951,N3952,N3953,N3954,N3955,N3956,N3957,
  N3958,N3959,N3960,N3961,N3962,N3963,N3964,N3965,N3966,N3967,N3968,N3969,N3970,
  N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978,N3979,N3980,N3981,N3982,N3983,N3984,
  N3985,N3986,N3987,N3988,N3989,N3990,N3991,N3992,N3993,N3994,N3995,N3996,N3997,
  N3998,N3999,N4000,N4001,N4002,N4003,N4004,N4005,N4006,N4007,N4008,N4009,N4010,
  N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,N4019,N4020,N4021,N4022,N4023,N4024,
  N4025,N4026,N4027,N4028,N4029,N4030,N4031,N4032,N4033,N4034,N4035,N4036,N4037,
  N4038,N4039,N4040,N4041,N4042,N4043,N4044,N4045,N4046,N4047,N4048,N4049,N4050,
  N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,N4059,N4060,N4061,N4062,N4063,N4064,
  N4065,N4066,N4067,N4068,N4069,N4070,N4071,N4072,N4073,N4074,N4075,N4076,N4077,
  N4078,N4079,N4080,N4081,N4082,N4083,N4084,N4085,N4086,N4087,N4088,N4089,N4090,
  N4091,N4092,N4093,N4094,N4095,N4096,N4097,N4098,N4099,N4100,N4101,N4102,N4103,N4104,
  N4105,N4106,N4107,N4108,N4109,N4110,N4111,N4112,N4113,N4114,N4115,N4116,N4117,
  N4118,N4119,N4120,N4121,N4122,N4123,N4124,N4125,N4126,N4127,N4128,N4129,N4130,
  N4131,N4132,N4133,N4134,N4135,N4136,N4137,N4138,N4139,N4140,N4141,N4142,N4143,N4144,
  N4145,N4146,N4147,N4148,N4149,N4150,N4151,N4152,N4153,N4154,N4155,N4156,N4157,
  N4158,N4159,N4160,N4161,N4162,N4163,N4164,N4165,N4166,N4167,N4168,N4169,N4170,
  N4171,N4172,N4173,N4174,N4175,N4176,N4177,N4178,N4179,N4180,N4181,N4182,N4183,N4184,
  N4185,N4186,N4187,N4188,N4189,N4190,N4191,N4192,N4193,N4194,N4195,N4196,N4197,
  N4198,N4199,N4200,N4201,N4202,N4203,N4204,N4205,N4206,N4207,N4208,N4209,N4210,
  N4211,N4212,N4213,N4214,N4215,N4216,N4217,N4218,N4219,N4220,N4221,N4222,N4223,N4224,
  N4225,N4226,N4227,N4228,N4229,N4230,N4231,N4232,N4233,N4234,N4235,N4236,N4237,
  N4238,N4239,N4240,N4241,N4242,N4243,N4244,N4245,N4246,N4247,N4248,N4249,N4250,
  N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,N4259,N4260,N4261,N4262,N4263,N4264,
  N4265,N4266,N4267,N4268,N4269,N4270,N4271,N4272,N4273,N4274,N4275,N4276,N4277,
  N4278,N4279,N4280,N4281,N4282,N4283,N4284,N4285,N4286,N4287,N4288,N4289,N4290,
  N4291,N4292,N4293,N4294,N4295,N4296,N4297,N4298,N4299,N4300,N4301,N4302,N4303,N4304,
  N4305,N4306,N4307,N4308,N4309,N4310,N4311,N4312,N4313,N4314,N4315,N4316,N4317,
  N4318,N4319,N4320,N4321,N4322,N4323,N4324,N4325,N4326,N4327,N4328,N4329,N4330,
  N4331,N4332,N4333,N4334,N4335,N4336,N4337,N4338,N4339,N4340,N4341,N4342,N4343,N4344,
  N4345,N4346,N4347,N4348,N4349,N4350,N4351,N4352,N4353,N4354,N4355,N4356,N4357,
  N4358,N4359,N4360,N4361,N4362,N4363,N4364,N4365,N4366,N4367,N4368,N4369,N4370,
  N4371,N4372,N4373,N4374,N4375,N4376,N4377,N4378,N4379,N4380,N4381,N4382,N4383,N4384,
  N4385,N4386,N4387,N4388,N4389,N4390,N4391,N4392,N4393,N4394,N4395,N4396,N4397,
  N4398,N4399,N4400,N4401,N4402,N4403,N4404,N4405,N4406,N4407,N4408,N4409,N4410,
  N4411,N4412,N4413,N4414,N4415,N4416,N4417,N4418,N4419,N4420,N4421,N4422,N4423,N4424,
  N4425,N4426,N4427,N4428,N4429,N4430,N4431,N4432,N4433,N4434,N4435,N4436,N4437,
  N4438,N4439,N4440,N4441,N4442,N4443,N4444,N4445,N4446,N4447,N4448,N4449,N4450,
  N4451,N4452,N4453,N4454,N4455,N4456,N4457,N4458,N4459,N4460,N4461,N4462,N4463,N4464,
  N4465,N4466,N4467,N4468,N4469,N4470,N4471,N4472,N4473,N4474,N4475,N4476,N4477,
  N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,N4487,N4488,N4489,N4490,
  N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,N4499,N4500,N4501,N4502,N4503,N4504,
  N4505,N4506,N4507,N4508,N4509,N4510,N4511,N4512,N4513,N4514,N4515,N4516,N4517,
  N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,N4527,N4528,N4529,N4530,
  N4531,N4532,N4533,N4534,N4535,N4536,N4537,N4538,N4539,N4540,N4541,N4542,N4543,N4544,
  N4545,N4546,N4547,N4548,N4549,N4550,N4551,N4552,N4553,N4554,N4555,N4556,N4557,
  N4558,N4559,N4560,N4561,N4562,N4563,N4564,N4565,N4566,N4567,N4568,N4569,N4570,
  N4571,N4572,N4573,N4574,N4575,N4576,N4577,N4578,N4579,N4580,N4581,N4582,N4583,N4584,
  N4585,N4586,N4587,N4588,N4589,N4590,N4591,N4592,N4593,N4594,N4595,N4596,N4597,
  N4598,N4599,N4600,N4601,N4602,N4603,N4604,N4605,N4606,N4607,N4608,N4609,N4610,
  N4611,N4612,N4613,N4614,N4615,N4616,N4617,N4618,N4619,N4620,N4621,N4622,N4623,N4624,
  N4625,N4626,N4627,N4628,N4629,N4630,N4631,N4632,N4633,N4634,N4635,N4636,N4637,
  N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,N4647,N4648,N4649,N4650,
  N4651,N4652,N4653,N4654,N4655,N4656,N4657,N4658,N4659,N4660,N4661,N4662,N4663,N4664,
  N4665,N4666,N4667,N4668,N4669,N4670,N4671,N4672,N4673,N4674,N4675,N4676,N4677,
  N4678,N4679,N4680,N4681,N4682,N4683,N4684,N4685,N4686,N4687,N4688,N4689,N4690,
  N4691,N4692,N4693,N4694,N4695,N4696,N4697,N4698,N4699,N4700,N4701,N4702,N4703,N4704,
  N4705,N4706,N4707,N4708,N4709,N4710,N4711,N4712,N4713,N4714,N4715,N4716,N4717,
  N4718,N4719,N4720,N4721,N4722,N4723,N4724,N4725,N4726,N4727,N4728,N4729,N4730,
  N4731,N4732,N4733,N4734,N4735,N4736,N4737,N4738,N4739,N4740,N4741,N4742,N4743,N4744,
  N4745,N4746,N4747,N4748,N4749,N4750,N4751,N4752,N4753,N4754,N4755,N4756,N4757,
  N4758,N4759,N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,N4768,N4769,N4770,
  N4771,N4772,N4773,N4774,N4775,N4776,N4777,N4778,N4779,N4780,N4781,N4782,N4783,N4784,
  N4785,N4786,N4787,N4788,N4789,N4790,N4791,N4792,N4793,N4794,N4795,N4796,N4797,
  N4798,N4799,N4800,N4801,N4802,N4803,N4804,N4805,N4806,N4807,N4808,N4809,N4810,
  N4811,N4812,N4813,N4814,N4815,N4816,N4817,N4818,N4819,N4820,N4821,N4822,N4823,N4824,
  N4825,N4826,N4827,N4828,N4829,N4830,N4831,N4832,N4833,N4834,N4835,N4836,N4837,
  N4838,N4839,N4840,N4841,N4842,N4843,N4844,N4845,N4846,N4847,N4848,N4849,N4850,
  N4851,N4852,N4853,N4854,N4855,N4856,N4857,N4858,N4859,N4860,N4861,N4862,N4863,N4864,
  N4865,N4866,N4867,N4868,N4869,N4870,N4871,N4872,N4873,N4874,N4875,N4876,N4877,
  N4878,N4879,N4880,N4881,N4882,N4883,N4884,N4885,N4886,N4887,N4888,N4889,N4890,
  N4891,N4892,N4893,N4894,N4895,N4896,N4897,N4898,N4899,N4900,N4901,N4902,N4903,N4904,
  N4905,N4906,N4907,N4908,N4909,N4910,N4911,N4912,N4913,N4914,N4915,N4916,N4917,
  N4918,N4919,N4920,N4921,N4922,N4923,N4924,N4925,N4926,N4927,N4928,N4929,N4930,
  N4931,N4932,N4933,N4934,N4935,N4936,N4937,N4938,N4939,N4940,N4941,N4942,N4943,N4944,
  N4945,N4946,N4947,N4948,N4949,N4950,N4951,N4952,N4953,N4954,N4955,N4956,N4957,
  N4958,N4959,N4960,N4961,N4962,N4963,N4964,N4965,N4966,N4967,N4968,N4969,N4970,
  N4971,N4972,N4973,N4974,N4975,N4976,N4977,N4978,N4979,N4980,N4981,N4982,N4983,N4984,
  N4985,N4986,N4987,N4988,N4989,N4990,N4991,N4992,N4993,N4994,N4995,N4996,N4997,
  N4998,N4999,N5000,N5001,N5002,N5003,N5004,N5005,N5006,N5007,N5008,N5009,N5010,
  N5011,N5012,N5013,N5014,N5015,N5016,N5017,N5018,N5019,N5020,N5021,N5022,N5023,N5024,
  N5025,N5026,N5027,N5028,N5029,N5030,N5031,N5032,N5033,N5034,N5035,N5036,N5037,
  N5038,N5039,N5040,N5041,N5042,N5043,N5044,N5045,N5046,N5047,N5048,N5049,N5050,
  N5051,N5052,N5053,N5054,N5055,N5056,N5057,N5058,N5059,N5060,N5061,N5062,N5063,N5064,
  N5065,N5066,N5067,N5068,N5069,N5070,N5071,N5072,N5073,N5074,N5075,N5076,N5077,
  N5078,N5079,N5080,N5081,N5082,N5083,N5084,N5085,N5086,N5087,N5088,N5089,N5090,
  N5091,N5092,N5093,N5094,N5095,N5096,N5097,N5098,N5099,N5100,N5101,N5102,N5103,N5104,
  N5105,N5106,N5107,N5108,N5109,N5110,N5111,N5112,N5113,N5114,N5115,N5116,N5117,
  N5118,N5119,N5120,N5121,N5122,N5123,N5124,N5125,N5126,N5127,N5128,N5129,N5130,
  N5131,N5132,N5133,N5134,N5135,N5136,N5137,N5138,N5139,N5140,N5141,N5142,N5143,N5144,
  N5145,N5146,N5147,N5148,N5149,N5150,N5151,N5152,N5153,N5154,N5155,N5156,N5157,
  N5158,N5159,N5160,N5161,N5162,N5163,N5164,N5165,N5166,N5167,N5168,N5169,N5170,
  N5171,N5172,N5173,N5174,N5175,N5176,N5177,N5178,N5179,N5180,N5181,N5182,N5183,N5184,
  N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,N5193,N5194,N5195,N5196,N5197,
  N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,N5207,N5208,N5209,N5210,
  N5211,N5212,N5213,N5214,N5215,N5216,N5217,N5218,N5219,N5220,N5221,N5222,N5223,N5224,
  N5225,N5226,N5227,N5228,N5229,N5230,N5231,N5232,N5233,N5234,N5235,N5236,N5237,
  N5238,N5239,N5240,N5241,N5242,N5243,N5244,N5245,N5246,N5247,N5248,N5249,N5250,
  N5251,N5252,N5253,N5254,N5255,N5256,N5257,N5258,N5259,N5260,N5261,N5262,N5263,N5264,
  N5265,N5266,N5267,N5268,N5269,N5270,N5271,N5272,N5273,N5274,N5275,N5276,N5277,
  N5278,N5279,N5280,N5281,N5282,N5283,N5284,N5285,N5286,N5287,N5288,N5289,N5290,
  N5291,N5292,N5293,N5294,N5295,N5296,N5297,N5298,N5299,N5300,N5301,N5302,N5303,N5304,
  N5305,N5306,N5307,N5308,N5309,N5310,N5311,N5312,N5313,N5314,N5315,N5316,N5317,
  N5318,N5319,N5320,N5321,N5322,N5323,N5324,N5325,N5326,N5327,N5328,N5329,N5330,
  N5331,N5332,N5333,N5334,N5335,N5336,N5337,N5338,N5339,N5340,N5341,N5342,N5343,N5344,
  N5345,N5346,N5347,N5348,N5349,N5350,N5351,N5352,N5353,N5354,N5355,N5356,N5357,
  N5358,N5359,N5360,N5361,N5362,N5363,N5364,N5365,N5366,N5367,N5368,N5369,N5370,
  N5371,N5372,N5373,N5374,N5375,N5376,N5377,N5378,N5379,N5380,N5381,N5382,N5383,N5384,
  N5385,N5386,N5387,N5388,N5389,N5390,N5391,N5392,N5393,N5394,N5395,N5396,N5397,
  N5398,N5399,N5400,N5401,N5402,N5403,N5404,N5405,N5406,N5407,N5408,N5409,N5410,
  N5411,N5412,N5413,N5414,N5415,N5416,N5417,N5418,N5419,N5420,N5421,N5422,N5423,N5424,
  N5425,N5426,N5427,N5428,N5429,N5430,N5431,N5432,N5433,N5434,N5435,N5436,N5437,
  N5438,N5439,N5440,N5441,N5442,N5443,N5444,N5445,N5446,N5447,N5448,N5449,N5450,
  N5451,N5452,N5453,N5454,N5455,N5456,N5457,N5458,N5459,N5460,N5461,N5462,N5463,N5464,
  N5465,N5466,N5467,N5468,N5469,N5470,N5471,N5472,N5473,N5474,N5475,N5476,N5477,
  N5478,N5479,N5480,N5481,N5482,N5483,N5484,N5485,N5486,N5487,N5488,N5489,N5490,
  N5491,N5492,N5493,N5494,N5495,N5496,N5497,N5498,N5499,N5500,N5501,N5502,N5503,N5504,
  N5505,N5506,N5507,N5508,N5509,N5510,N5511,N5512,N5513,N5514,N5515,N5516,N5517,
  N5518,N5519,N5520,N5521,N5522,N5523,N5524,N5525,N5526,N5527,N5528,N5529,N5530,
  N5531,N5532,N5533,N5534,N5535,N5536,N5537,N5538,N5539,N5540,N5541,N5542,N5543,N5544,
  N5545,N5546,N5547,N5548,N5549,N5550,N5551,N5552,N5553,N5554,N5555,N5556,N5557,
  N5558,N5559,N5560,N5561,N5562,N5563,N5564,N5565,N5566,N5567,N5568,N5569,N5570,
  N5571,N5572,N5573,N5574,N5575,N5576,N5577,N5578,N5579,N5580,N5581,N5582,N5583,N5584,
  N5585,N5586,N5587,N5588,N5589,N5590,N5591,N5592,N5593,N5594,N5595,N5596,N5597,
  N5598,N5599,N5600,N5601,N5602,N5603,N5604,N5605,N5606,N5607,N5608,N5609,N5610,
  N5611,N5612,N5613,N5614,N5615,N5616,N5617,N5618,N5619,N5620,N5621,N5622,N5623,N5624,
  N5625,N5626,N5627,N5628,N5629,N5630,N5631,N5632,N5633,N5634,N5635,N5636,N5637,
  N5638,N5639,N5640,N5641,N5642,N5643,N5644,N5645,N5646,N5647,N5648,N5649,N5650,
  N5651,N5652,N5653,N5654,N5655,N5656,N5657,N5658,N5659,N5660,N5661,N5662,N5663,N5664,
  N5665,N5666,N5667,N5668,N5669,N5670,N5671,N5672,N5673,N5674,N5675,N5676,N5677,
  N5678,N5679,N5680,N5681,N5682,N5683,N5684,N5685,N5686,N5687,N5688,N5689,N5690,
  N5691,N5692,N5693,N5694,N5695,N5696,N5697,N5698,N5699,N5700,N5701,N5702,N5703,N5704,
  N5705,N5706,N5707,N5708,N5709,N5710,N5711,N5712,N5713,N5714,N5715,N5716,N5717,
  N5718,N5719,N5720,N5721,N5722,N5723,N5724,N5725,N5726,N5727,N5728,N5729,N5730,
  N5731,N5732,N5733,N5734,N5735,N5736,N5737,N5738,N5739,N5740,N5741,N5742,N5743,N5744,
  N5745,N5746,N5747,N5748,N5749,N5750,N5751,N5752,N5753,N5754,N5755,N5756,N5757,
  N5758,N5759,N5760,N5761,N5762,N5763,N5764,N5765,N5766,N5767,N5768,N5769,N5770,
  N5771,N5772,N5773,N5774,N5775,N5776,N5777,N5778,N5779,N5780,N5781,N5782,N5783,N5784,
  N5785,N5786,N5787,N5788,N5789,N5790,N5791,N5792,N5793,N5794,N5795,N5796,N5797,
  N5798,N5799,N5800,N5801,N5802,N5803,N5804,N5805,N5806,N5807,N5808,N5809,N5810,
  N5811,N5812,N5813,N5814,N5815,N5816,N5817,N5818,N5819,N5820,N5821,N5822,N5823,N5824,
  N5825,N5826,N5827,N5828,N5829,N5830,N5831,N5832,N5833,N5834,N5835,N5836,N5837,
  N5838,N5839,N5840,N5841,N5842,N5843,N5844,N5845,N5846,N5847,N5848,N5849,N5850,
  N5851,N5852,N5853,N5854,N5855,N5856,N5857,N5858,N5859,N5860,N5861,N5862,N5863,N5864,
  N5865,N5866,N5867,N5868,N5869,N5870,N5871,N5872,N5873,N5874,N5875,N5876,N5877,
  N5878,N5879,N5880,N5881,N5882,N5883,N5884,N5885,N5886,N5887,N5888,N5889,N5890,
  N5891,N5892,N5893,N5894,N5895,N5896,N5897,N5898,N5899,N5900,N5901,N5902,N5903,N5904,
  N5905,N5906,N5907,N5908,N5909,N5910,N5911,N5912,N5913,N5914,N5915,N5916,N5917,
  N5918,N5919,N5920,N5921,N5922,N5923,N5924,N5925,N5926,N5927,N5928,N5929,N5930,
  N5931,N5932,N5933,N5934,N5935,N5936,N5937,N5938,N5939,N5940,N5941,N5942,N5943,N5944,
  N5945,N5946,N5947,N5948,N5949,N5950,N5951,N5952,N5953,N5954,N5955,N5956,N5957,
  N5958,N5959,N5960,N5961,N5962,N5963,N5964,N5965,N5966,N5967,N5968,N5969,N5970,
  N5971,N5972,N5973,N5974,N5975,N5976,N5977,N5978,N5979,N5980,N5981,N5982,N5983,N5984,
  N5985,N5986,N5987,N5988,N5989,N5990,N5991,N5992,N5993,N5994,N5995,N5996,N5997,
  N5998,N5999,N6000,N6001,N6002,N6003,N6004,N6005,N6006,N6007,N6008,N6009,N6010,
  N6011,N6012,N6013,N6014,N6015,N6016,N6017,N6018,N6019,N6020,N6021,N6022,N6023,N6024,
  N6025,N6026,N6027,N6028,N6029,N6030,N6031,N6032,N6033,N6034,N6035,N6036,N6037,
  N6038,N6039,N6040,N6041,N6042,N6043,N6044,N6045,N6046,N6047,N6048,N6049,N6050,
  N6051,N6052,N6053,N6054,N6055,N6056,N6057,N6058,N6059,N6060,N6061,N6062,N6063,N6064,
  N6065,N6066,N6067,N6068,N6069,N6070,N6071,N6072,N6073,N6074,N6075,N6076,N6077,
  N6078,N6079,N6080,N6081,N6082,N6083,N6084,N6085,N6086,N6087,N6088,N6089,N6090,
  N6091,N6092,N6093,N6094,N6095,N6096,N6097,N6098,N6099,N6100,N6101,N6102,N6103,N6104,
  N6105,N6106,N6107,N6108,N6109,N6110,N6111,N6112,N6113,N6114,N6115,N6116,N6117,
  N6118,N6119,N6120,N6121,N6122,N6123,N6124,N6125,N6126,N6127,N6128,N6129,N6130,
  N6131,N6132,N6133,N6134,N6135,N6136,N6137,N6138,N6139,N6140,N6141,N6142,N6143,N6144,
  N6145,N6146,N6147,N6148,N6149,N6150,N6151,N6152,N6153,N6154,N6155,N6156,N6157,
  N6158,N6159,N6160,N6161,N6162,N6163,N6164,N6165,N6166,N6167,N6168,N6169,N6170,
  N6171,N6172,N6173,N6174,N6175,N6176,N6177,N6178,N6179,N6180,N6181,N6182,N6183,N6184,
  N6185,N6186,N6187,N6188,N6189,N6190,N6191,N6192,N6193,N6194,N6195,N6196,N6197,
  N6198,N6199,N6200,N6201,N6202,N6203,N6204,N6205,N6206,N6207,N6208,N6209,N6210,
  N6211,N6212,N6213,N6214,N6215,N6216,N6217,N6218,N6219,N6220,N6221,N6222,N6223,N6224,
  N6225,N6226,N6227,N6228,N6229,N6230,N6231,N6232,N6233,N6234,N6235,N6236,N6237,
  N6238,N6239,N6240,N6241,N6242,N6243,N6244,N6245,N6246,N6247,N6248,N6249,N6250,
  N6251,N6252,N6253,N6254,N6255,N6256,N6257,N6258,N6259,N6260,N6261,N6262,N6263,N6264,
  N6265,N6266,N6267,N6268,N6269,N6270,N6271,N6272,N6273,N6274,N6275,N6276,N6277,
  N6278,N6279,N6280,N6281,N6282,N6283,N6284,N6285,N6286,N6287,N6288,N6289,N6290,
  N6291,N6292,N6293,N6294,N6295,N6296,N6297,N6298,N6299,N6300,N6301,N6302,N6303,N6304,
  N6305,N6306,N6307,N6308,N6309,N6310,N6311,N6312,N6313,N6314,N6315,N6316,N6317,
  N6318,N6319,N6320,N6321,N6322,N6323,N6324,N6325,N6326,N6327,N6328,N6329,N6330,
  N6331,N6332,N6333,N6334,N6335,N6336,N6337,N6338,N6339,N6340,N6341,N6342,N6343,N6344,
  N6345,N6346,N6347,N6348,N6349,N6350,N6351,N6352,N6353,N6354,N6355,N6356,N6357,
  N6358,N6359,N6360,N6361,N6362,N6363,N6364,N6365,N6366,N6367,N6368,N6369,N6370,
  N6371,N6372,N6373,N6374,N6375,N6376,N6377,N6378,N6379,N6380,N6381,N6382,N6383,N6384,
  N6385,N6386,N6387,N6388,N6389,N6390,N6391,N6392,N6393,N6394,N6395,N6396,N6397,
  N6398,N6399,N6400,N6401,N6402,N6403,N6404,N6405,N6406,N6407,N6408,N6409,N6410,
  N6411,N6412,N6413,N6414,N6415,N6416,N6417,N6418,N6419,N6420,N6421,N6422,N6423,N6424,
  N6425,N6426,N6427,N6428,N6429,N6430,N6431,N6432,N6433,N6434,N6435,N6436,N6437,
  N6438,N6439,N6440,N6441,N6442,N6443,N6444,N6445,N6446,N6447,N6448,N6449,N6450,
  N6451,N6452,N6453,N6454,N6455,N6456,N6457,N6458,N6459,N6460,N6461,N6462,N6463,N6464,
  N6465,N6466,N6467,N6468,N6469,N6470,N6471,N6472,N6473,N6474,N6475,N6476,N6477,
  N6478,N6479,N6480,N6481,N6482,N6483,N6484,N6485,N6486,N6487,N6488,N6489,N6490,
  N6491,N6492,N6493,N6494,N6495,N6496,N6497,N6498,N6499,N6500,N6501,N6502,N6503,N6504,
  N6505,N6506,N6507,N6508,N6509,N6510,N6511,N6512,N6513,N6514,N6515,N6516,N6517,
  N6518,N6519,N6520,N6521,N6522,N6523,N6524,N6525,N6526,N6527,N6528,N6529,N6530,
  N6531,N6532,N6533,N6534,N6535,N6536,N6537,N6538,N6539,N6540,N6541,N6542,N6543,N6544,
  N6545,N6546,N6547,N6548,N6549,N6550,N6551,N6552,N6553,N6554,N6555,N6556,N6557,
  N6558,N6559,N6560,N6561,N6562,N6563,N6564,N6565,N6566,N6567,N6568,N6569,N6570,
  N6571,N6572,N6573,N6574,N6575,N6576,N6577,N6578,N6579,N6580,N6581,N6582,N6583,N6584,
  N6585,N6586,N6587,N6588,N6589,N6590,N6591,N6592,N6593,N6594,N6595,N6596,N6597,
  N6598,N6599,N6600,N6601,N6602,N6603,N6604,N6605,N6606,N6607,N6608,N6609,N6610,
  N6611,N6612,N6613,N6614,N6615,N6616,N6617,N6618,N6619,N6620,N6621,N6622,N6623,N6624,
  N6625,N6626,N6627,N6628,N6629,N6630,N6631,N6632,N6633,N6634,N6635,N6636,N6637,
  N6638,N6639,N6640,N6641,N6642,N6643,N6644,N6645,N6646,N6647,N6648,N6649,N6650,
  N6651,N6652,N6653,N6654,N6655,N6656,N6657,N6658,N6659,N6660,N6661,N6662,N6663,N6664,
  N6665,N6666,N6667,N6668,N6669,N6670,N6671,N6672,N6673,N6674,N6675,N6676,N6677,
  N6678,N6679,N6680,N6681,N6682,N6683,N6684,N6685,N6686,N6687,N6688,N6689,N6690,
  N6691,N6692,N6693,N6694,N6695,N6696,N6697,N6698,N6699,N6700,N6701,N6702,N6703,N6704,
  N6705,N6706,N6707,N6708,N6709,N6710,N6711,N6712,N6713,N6714,N6715,N6716,N6717,
  N6718,N6719,N6720,N6721,N6722,N6723,N6724,N6725,N6726,N6727,N6728,N6729,N6730,
  N6731,N6732,N6733,N6734,N6735,N6736,N6737,N6738,N6739,N6740,N6741,N6742,N6743,N6744,
  N6745,N6746,N6747,N6748,N6749,N6750,N6751,N6752,N6753,N6754,N6755,N6756,N6757,
  N6758,N6759,N6760,N6761,N6762,N6763,N6764,N6765,N6766,N6767,N6768,N6769,N6770,
  N6771,N6772,N6773,N6774,N6775,N6776,N6777,N6778,N6779,N6780,N6781,N6782,N6783,N6784,
  N6785,N6786,N6787,N6788,N6789,N6790,N6791,N6792,N6793,N6794,N6795,N6796,N6797,
  N6798,N6799,N6800,N6801,N6802,N6803,N6804,N6805,N6806,N6807,N6808,N6809,N6810,
  N6811,N6812,N6813,N6814,N6815,N6816,N6817,N6818,N6819,N6820,N6821,N6822,N6823,N6824,
  N6825,N6826,N6827,N6828,N6829,N6830,N6831,N6832,N6833,N6834,N6835,N6836,N6837,
  N6838,N6839,N6840,N6841,N6842,N6843,N6844,N6845,N6846,N6847,N6848,N6849,N6850,
  N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6858,N6859,N6860,N6861,N6862,N6863,N6864,
  N6865,N6866,N6867,N6868,N6869,N6870,N6871,N6872,N6873,N6874,N6875,N6876,N6877,
  N6878,N6879,N6880,N6881,N6882,N6883,N6884,N6885,N6886,N6887,N6888,N6889,N6890,
  N6891,N6892,N6893,N6894,N6895,N6896,N6897,N6898,N6899,N6900,N6901,N6902,N6903,N6904,
  N6905,N6906,N6907,N6908,N6909,N6910,N6911,N6912,N6913,N6914,N6915,N6916,N6917,
  N6918,N6919,N6920,N6921,N6922,N6923,N6924,N6925,N6926,N6927,N6928,N6929,N6930,
  N6931,N6932,N6933,N6934,N6935,N6936,N6937,N6938,N6939,N6940,N6941,N6942,N6943,N6944,
  N6945,N6946,N6947,N6948,N6949,N6950,N6951,N6952,N6953,N6954,N6955,N6956,N6957,
  N6958,N6959,N6960,N6961,N6962,N6963,N6964,N6965,N6966,N6967,N6968,N6969,N6970,
  N6971,N6972,N6973,N6974,N6975,N6976,N6977,N6978,N6979,N6980,N6981,N6982,N6983,N6984,
  N6985,N6986,N6987,N6988,N6989,N6990,N6991,N6992,N6993,N6994,N6995,N6996,N6997,
  N6998,N6999,N7000,N7001,N7002,N7003,N7004,N7005,N7006,N7007,N7008,N7009,N7010,
  N7011,N7012,N7013,N7014,N7015,N7016,N7017,N7018,N7019,N7020,N7021,N7022,N7023,N7024,
  N7025,N7026,N7027,N7028,N7029,N7030,N7031,N7032,N7033,N7034,N7035,N7036,N7037,
  N7038,N7039,N7040,N7041,N7042,N7043,N7044,N7045,N7046,N7047,N7048,N7049,N7050,
  N7051,N7052,N7053,N7054,N7055,N7056,N7057,N7058,N7059,N7060,N7061,N7062,N7063,N7064,
  N7065,N7066,N7067,N7068,N7069,N7070,N7071,N7072,N7073,N7074,N7075,N7076,N7077,
  N7078,N7079,N7080,N7081,N7082,N7083,N7084,N7085,N7086,N7087,N7088,N7089,N7090,
  N7091,N7092,N7093,N7094,N7095,N7096,N7097,N7098,N7099,N7100,N7101,N7102,N7103,N7104,
  N7105,N7106,N7107,N7108,N7109,N7110,N7111,N7112,N7113,N7114,N7115,N7116,N7117,
  N7118,N7119,N7120,N7121,N7122,N7123,N7124,N7125,N7126,N7127,N7128,N7129,N7130,
  N7131,N7132,N7133,N7134,N7135,N7136,N7137,N7138,N7139,N7140,N7141,N7142,N7143,N7144,
  N7145,N7146,N7147,N7148,N7149,N7150,N7151,N7152,N7153,N7154,N7155,N7156,N7157,
  N7158,N7159,N7160,N7161,N7162,N7163,N7164,N7165,N7166,N7167,N7168,N7169,N7170,
  N7171,N7172,N7173,N7174,N7175,N7176,N7177,N7178,N7179,N7180,N7181,N7182,N7183,N7184,
  N7185,N7186,N7187,N7188,N7189,N7190,N7191,N7192,N7193,N7194,N7195,N7196,N7197,
  N7198,N7199,N7200,N7201,N7202,N7203,N7204,N7205,N7206,N7207,N7208,N7209,N7210,
  N7211,N7212,N7213,N7214,N7215,N7216,N7217,N7218,N7219,N7220,N7221,N7222,N7223,N7224,
  N7225,N7226,N7227,N7228,N7229,N7230,N7231,N7232,N7233,N7234,N7235,N7236,N7237,
  N7238,N7239,N7240,N7241,N7242,N7243,N7244,N7245,N7246,N7247,N7248,N7249,N7250,
  N7251,N7252,N7253,N7254,N7255,N7256,N7257,N7258,N7259,N7260,N7261,N7262,N7263,N7264,
  N7265,N7266,N7267,N7268,N7269,N7270,N7271,N7272,N7273,N7274,N7275,N7276,N7277,
  N7278,N7279,N7280,N7281,N7282,N7283,N7284,N7285,N7286,N7287,N7288,N7289,N7290,
  N7291,N7292,N7293,N7294,N7295,N7296,N7297,N7298,N7299,N7300,N7301,N7302,N7303,N7304,
  N7305,N7306,N7307,N7308,N7309,N7310,N7311,N7312,N7313,N7314,N7315,N7316,N7317,
  N7318,N7319,N7320,N7321,N7322,N7323,N7324,N7325,N7326,N7327,N7328,N7329,N7330,
  N7331,N7332,N7333,N7334,N7335,N7336,N7337,N7338,N7339,N7340,N7341,N7342,N7343,N7344,
  N7345,N7346,N7347,N7348,N7349,N7350,N7351,N7352,N7353,N7354,N7355,N7356,N7357,
  N7358,N7359,N7360,N7361,N7362,N7363,N7364,N7365,N7366,N7367,N7368,N7369,N7370,
  N7371,N7372,N7373,N7374,N7375,N7376,N7377,N7378,N7379,N7380,N7381,N7382,N7383,N7384,
  N7385,N7386,N7387,N7388,N7389,N7390,N7391,N7392,N7393,N7394,N7395,N7396,N7397,
  N7398,N7399,N7400,N7401,N7402,N7403,N7404,N7405,N7406,N7407,N7408,N7409,N7410,
  N7411,N7412,N7413,N7414,N7415,N7416,N7417,N7418,N7419,N7420,N7421,N7422,N7423,N7424,
  N7425,N7426,N7427,N7428,N7429,N7430,N7431,N7432,N7433,N7434,N7435,N7436,N7437,
  N7438,N7439,N7440,N7441,N7442,N7443,N7444,N7445,N7446,N7447,N7448,N7449,N7450,
  N7451,N7452,N7453,N7454,N7455,N7456,N7457,N7458,N7459,N7460,N7461,N7462,N7463,N7464,
  N7465,N7466,N7467,N7468,N7469,N7470,N7471,N7472,N7473,N7474,N7475,N7476,N7477,
  N7478,N7479,N7480,N7481,N7482,N7483,N7484,N7485,N7486,N7487,N7488,N7489,N7490,
  N7491,N7492,N7493,N7494,N7495,N7496,N7497,N7498,N7499,N7500,N7501,N7502,N7503,N7504,
  N7505,N7506,N7507,N7508,N7509,N7510,N7511,N7512,N7513,N7514,N7515,N7516,N7517,
  N7518,N7519,N7520,N7521,N7522,N7523,N7524,N7525,N7526,N7527,N7528,N7529,N7530,
  N7531,N7532,N7533,N7534,N7535,N7536,N7537,N7538,N7539,N7540,N7541,N7542,N7543,N7544,
  N7545,N7546,N7547,N7548,N7549,N7550,N7551,N7552,N7553,N7554,N7555,N7556,N7557,
  N7558,N7559,N7560,N7561,N7562,N7563,N7564,N7565,N7566,N7567,N7568,N7569,N7570,
  N7571,N7572,N7573,N7574,N7575,N7576,N7577,N7578,N7579,N7580,N7581,N7582,N7583,N7584,
  N7585,N7586,N7587,N7588,N7589,N7590,N7591,N7592,N7593,N7594,N7595,N7596,N7597,
  N7598,N7599,N7600,N7601,N7602,N7603,N7604,N7605,N7606,N7607,N7608,N7609,N7610,
  N7611,N7612,N7613,N7614,N7615,N7616,N7617,N7618,N7619,N7620,N7621,N7622,N7623,N7624,
  N7625,N7626,N7627,N7628,N7629,N7630,N7631,N7632,N7633,N7634,N7635,N7636,N7637,
  N7638,N7639,N7640,N7641,N7642,N7643,N7644,N7645,N7646,N7647,N7648,N7649,N7650,
  N7651,N7652,N7653,N7654,N7655,N7656,N7657,N7658,N7659,N7660,N7661,N7662,N7663,N7664,
  N7665,N7666,N7667,N7668,N7669,N7670,N7671,N7672,N7673,N7674,N7675,N7676,N7677,
  N7678,N7679,N7680,N7681,N7682,N7683,N7684,N7685,N7686,N7687,N7688,N7689,N7690,
  N7691,N7692,N7693,N7694,N7695,N7696,N7697,N7698,N7699,N7700,N7701,N7702,N7703,N7704,
  N7705,N7706,N7707,N7708,N7709,N7710,N7711,N7712,N7713,N7714,N7715,N7716,N7717,
  N7718,N7719,N7720,N7721,N7722,N7723,N7724,N7725,N7726,N7727,N7728,N7729,N7730,
  N7731,N7732,N7733,N7734,N7735,N7736,N7737,N7738,N7739,N7740,N7741,N7742,N7743,N7744,
  N7745,N7746,N7747,N7748,N7749,N7750,N7751,N7752,N7753,N7754,N7755,N7756,N7757,
  N7758,N7759,N7760,N7761,N7762,N7763,N7764,N7765,N7766,N7767,N7768,N7769,N7770,
  N7771,N7772,N7773,N7774,N7775,N7776,N7777,N7778,N7779,N7780,N7781,N7782,N7783,N7784,
  N7785,N7786,N7787,N7788,N7789,N7790,N7791,N7792,N7793,N7794,N7795,N7796,N7797,
  N7798,N7799,N7800,N7801,N7802,N7803,N7804,N7805,N7806,N7807,N7808,N7809,N7810,
  N7811,N7812,N7813,N7814,N7815,N7816,N7817,N7818,N7819,N7820,N7821,N7822,N7823,N7824,
  N7825,N7826,N7827,N7828,N7829,N7830,N7831,N7832,N7833,N7834,N7835,N7836,N7837,
  N7838,N7839,N7840,N7841,N7842,N7843,N7844,N7845,N7846,N7847,N7848,N7849,N7850,
  N7851,N7852,N7853,N7854,N7855,N7856,N7857,N7858,N7859,N7860,N7861,N7862,N7863,N7864,
  N7865,N7866,N7867,N7868,N7869,N7870,N7871,N7872,N7873,N7874,N7875,N7876,N7877,
  N7878,N7879,N7880,N7881,N7882,N7883,N7884,N7885,N7886,N7887,N7888,N7889,N7890,
  N7891,N7892,N7893,N7894,N7895,N7896,N7897,N7898,N7899,N7900,N7901,N7902,N7903,N7904,
  N7905,N7906,N7907,N7908,N7909,N7910,N7911,N7912,N7913,N7914,N7915,N7916,N7917,
  N7918,N7919,N7920,N7921,N7922,N7923,N7924,N7925,N7926,N7927,N7928,N7929,N7930,
  N7931,N7932,N7933,N7934,N7935,N7936,N7937,N7938,N7939,N7940,N7941,N7942,N7943,N7944,
  N7945,N7946,N7947,N7948,N7949,N7950,N7951,N7952,N7953,N7954,N7955,N7956,N7957,
  N7958,N7959,N7960,N7961,N7962,N7963,N7964,N7965,N7966,N7967,N7968,N7969,N7970,
  N7971,N7972,N7973,N7974,N7975,N7976,N7977,N7978,N7979,N7980,N7981,N7982,N7983,N7984,
  N7985,N7986,N7987,N7988,N7989,N7990,N7991,N7992,N7993,N7994,N7995,N7996,N7997,
  N7998,N7999,N8000,N8001,N8002,N8003,N8004,N8005,N8006,N8007,N8008,N8009,N8010,
  N8011,N8012,N8013,N8014,N8015,N8016,N8017,N8018,N8019,N8020,N8021,N8022,N8023,N8024,
  N8025,N8026,N8027,N8028,N8029,N8030,N8031,N8032,N8033,N8034,N8035,N8036,N8037,
  N8038,N8039,N8040,N8041,N8042,N8043,N8044,N8045,N8046,N8047,N8048,N8049,N8050,
  N8051,N8052,N8053,N8054,N8055,N8056,N8057,N8058,N8059,N8060,N8061,N8062,N8063,N8064,
  N8065,N8066,N8067,N8068,N8069,N8070,N8071,N8072,N8073,N8074,N8075,N8076,N8077,
  N8078,N8079,N8080,N8081,N8082,N8083,N8084,N8085,N8086,N8087,N8088,N8089,N8090,
  N8091,N8092,N8093,N8094,N8095,N8096,N8097,N8098,N8099,N8100,N8101,N8102,N8103,N8104,
  N8105,N8106,N8107,N8108,N8109,N8110,N8111,N8112,N8113,N8114,N8115,N8116,N8117,
  N8118,N8119,N8120,N8121,N8122,N8123,N8124,N8125,N8126,N8127,N8128,N8129,N8130,
  N8131,N8132,N8133,N8134,N8135,N8136,N8137,N8138,N8139,N8140,N8141,N8142,N8143,N8144,
  N8145,N8146,N8147,N8148,N8149,N8150,N8151,N8152,N8153,N8154,N8155,N8156,N8157,
  N8158,N8159,N8160,N8161,N8162,N8163,N8164,N8165,N8166,N8167,N8168,N8169,N8170,
  N8171,N8172,N8173,N8174,N8175,N8176,N8177,N8178,N8179,N8180,N8181,N8182,N8183,N8184,
  N8185,N8186,N8187,N8188,N8189,N8190,N8191,N8192,N8193,N8194,N8195,N8196,N8197,
  N8198,N8199,N8200,N8201,N8202,N8203,N8204,N8205,N8206,N8207,N8208,N8209,N8210,
  N8211,N8212,N8213,N8214,N8215,N8216,N8217,N8218,N8219,N8220,N8221,N8222,N8223,N8224,
  N8225,N8226,N8227,N8228,N8229,N8230,N8231,N8232,N8233,N8234,N8235,N8236,N8237,
  N8238,N8239,N8240,N8241,N8242,N8243,N8244,N8245,N8246,N8247,N8248,N8249,N8250,
  N8251,N8252,N8253,N8254,N8255,N8256,N8257,N8258,N8259,N8260,N8261,N8262,N8263,N8264,
  N8265,N8266,N8267,N8268,N8269,N8270,N8271,N8272,N8273,N8274,N8275,N8276,N8277,
  N8278,N8279,N8280,N8281,N8282,N8283,N8284,N8285,N8286,N8287,N8288,N8289,N8290,
  N8291,N8292,N8293,N8294,N8295,N8296,N8297,N8298,N8299,N8300,N8301,N8302,N8303,N8304,
  N8305,N8306,N8307,N8308,N8309,N8310,N8311,N8312,N8313,N8314,N8315,N8316,N8317,
  N8318,N8319,N8320,N8321,N8322,N8323,N8324,N8325,N8326,N8327,N8328,N8329,N8330,
  N8331,N8332,N8333,N8334,N8335,N8336,N8337,N8338,N8339,N8340,N8341,N8342,N8343,N8344,
  N8345,N8346,N8347,N8348,N8349,N8350,N8351,N8352,N8353,N8354,N8355,N8356,N8357,
  N8358,N8359,N8360,N8361,N8362,N8363,N8364,N8365,N8366,N8367,N8368,N8369,N8370,
  N8371,N8372,N8373,N8374,N8375,N8376,N8377,N8378,N8379,N8380,N8381,N8382,N8383,N8384,
  N8385,N8386,N8387,N8388,N8389,N8390,N8391,N8392,N8393,N8394,N8395,N8396,N8397,
  N8398,N8399,N8400,N8401,N8402,N8403,N8404,N8405,N8406,N8407,N8408,N8409,N8410,
  N8411,N8412,N8413,N8414,N8415,N8416,N8417,N8418,N8419,N8420,N8421,N8422,N8423,N8424,
  N8425,N8426,N8427,N8428,N8429,N8430,N8431,N8432,N8433,N8434,N8435,N8436,N8437,
  N8438,N8439,N8440,N8441,N8442,N8443,N8444,N8445,N8446,N8447,N8448,N8449,N8450,
  N8451,N8452,N8453,N8454,N8455,N8456,N8457,N8458,N8459,N8460,N8461,N8462,N8463,N8464,
  N8465,N8466,N8467,N8468,N8469,N8470,N8471,N8472,N8473,N8474,N8475,N8476,N8477,
  N8478,N8479,N8480,N8481,N8482,N8483,N8484,N8485,N8486,N8487,N8488,N8489,N8490,
  N8491,N8492,N8493,N8494,N8495,N8496,N8497,N8498,N8499,N8500,N8501,N8502,N8503,N8504,
  N8505,N8506,N8507,N8508,N8509,N8510,N8511,N8512,N8513,N8514,N8515,N8516,N8517,
  N8518,N8519,N8520,N8521,N8522,N8523,N8524,N8525,N8526,N8527,N8528,N8529,N8530,
  N8531,N8532,N8533,N8534,N8535,N8536,N8537,N8538,N8539,N8540,N8541,N8542,N8543,N8544,
  N8545,N8546,N8547,N8548,N8549,N8550,N8551,N8552,N8553,N8554,N8555,N8556,N8557,
  N8558,N8559,N8560,N8561,N8562,N8563,N8564,N8565,N8566,N8567,N8568,N8569,N8570,
  N8571,N8572,N8573,N8574,N8575,N8576,N8577,N8578,N8579,N8580,N8581,N8582,N8583,N8584,
  N8585,N8586,N8587,N8588,N8589,N8590,N8591,N8592,N8593,N8594,N8595,N8596,N8597,
  N8598,N8599,N8600,N8601,N8602,N8603,N8604,N8605,N8606,N8607,N8608,N8609,N8610,
  N8611,N8612,N8613,N8614,N8615,N8616,N8617,N8618,N8619,N8620,N8621,N8622,N8623,N8624,
  N8625,N8626,N8627,N8628,N8629,N8630,N8631,N8632,N8633,N8634,N8635,N8636,N8637,
  N8638,N8639,N8640,N8641,N8642,N8643,N8644,N8645,N8646,N8647,N8648,N8649,N8650,
  N8651,N8652,N8653,N8654,N8655,N8656,N8657,N8658,N8659,N8660,N8661,N8662,N8663,N8664,
  N8665,N8666,N8667,N8668,N8669,N8670,N8671,N8672,N8673,N8674,N8675,N8676,N8677,
  N8678,N8679,N8680,N8681,N8682,N8683,N8684,N8685,N8686,N8687,N8688,N8689,N8690,
  N8691,N8692,N8693,N8694,N8695,N8696,N8697,N8698,N8699,N8700,N8701,N8702,N8703,N8704,
  N8705,N8706,N8707,N8708,N8709,N8710,N8711,N8712,N8713,N8714,N8715,N8716,N8717,
  N8718,N8719,N8720,N8721,N8722,N8723,N8724,N8725,N8726,N8727,N8728,N8729,N8730,
  N8731,N8732,N8733,N8734,N8735,N8736,N8737,N8738,N8739,N8740,N8741,N8742,N8743,N8744,
  N8745,N8746,N8747,N8748,N8749,N8750,N8751,N8752,N8753,N8754,N8755,N8756,N8757,
  N8758,N8759,N8760,N8761,N8762,N8763,N8764,N8765,N8766,N8767,N8768,N8769,N8770,
  N8771,N8772,N8773,N8774,N8775,N8776,N8777,N8778,N8779,N8780,N8781,N8782,N8783,N8784,
  N8785,N8786,N8787,N8788,N8789,N8790,N8791,N8792,N8793,N8794,N8795,N8796,N8797,
  N8798,N8799,N8800,N8801,N8802,N8803,N8804,N8805,N8806,N8807,N8808,N8809,N8810,
  N8811,N8812,N8813,N8814,N8815,N8816,N8817,N8818,N8819,N8820,N8821,N8822,N8823,N8824,
  N8825,N8826,N8827,N8828,N8829,N8830,N8831,N8832,N8833,N8834,N8835,N8836,N8837,
  N8838,N8839,N8840,N8841,N8842,N8843,N8844,N8845,N8846,N8847,N8848,N8849,N8850,
  N8851,N8852,N8853,N8854,N8855,N8856,N8857,N8858,N8859,N8860,N8861,N8862,N8863,N8864,
  N8865,N8866,N8867,N8868,N8869,N8870,N8871,N8872,N8873,N8874,N8875,N8876,N8877,
  N8878,N8879,N8880,N8881,N8882,N8883,N8884,N8885,N8886,N8887,N8888,N8889,N8890,
  N8891,N8892,N8893,N8894,N8895,N8896,N8897,N8898,N8899,N8900,N8901,N8902,N8903,N8904,
  N8905,N8906,N8907,N8908,N8909,N8910,N8911,N8912,N8913,N8914,N8915,N8916,N8917,
  N8918,N8919,N8920,N8921,N8922,N8923,N8924,N8925,N8926,N8927,N8928,N8929,N8930,
  N8931,N8932,N8933,N8934,N8935,N8936,N8937,N8938,N8939,N8940,N8941,N8942,N8943,N8944,
  N8945,N8946,N8947,N8948,N8949,N8950,N8951,N8952,N8953,N8954,N8955,N8956,N8957,
  N8958,N8959,N8960,N8961,N8962,N8963,N8964,N8965,N8966,N8967,N8968,N8969,N8970,
  N8971,N8972,N8973,N8974,N8975,N8976,N8977,N8978,N8979,N8980,N8981,N8982,N8983,N8984,
  N8985,N8986,N8987,N8988,N8989,N8990,N8991,N8992,N8993,N8994,N8995,N8996,N8997,
  N8998,N8999,N9000,N9001,N9002,N9003,N9004,N9005,N9006,N9007,N9008,N9009,N9010,
  N9011,N9012,N9013,N9014,N9015,N9016,N9017,N9018,N9019,N9020,N9021,N9022,N9023,N9024,
  N9025,N9026,N9027,N9028,N9029,N9030,N9031,N9032,N9033,N9034,N9035,N9036,N9037,
  N9038,N9039,N9040,N9041,N9042,N9043,N9044,N9045,N9046,N9047,N9048,N9049,N9050,
  N9051,N9052,N9053,N9054,N9055,N9056,N9057,N9058,N9059,N9060,N9061,N9062,N9063,N9064,
  N9065,N9066,N9067,N9068,N9069,N9070,N9071,N9072,N9073,N9074,N9075,N9076,N9077,
  N9078,N9079,N9080,N9081,N9082,N9083,N9084,N9085,N9086,N9087,N9088,N9089,N9090,
  N9091,N9092,N9093,N9094,N9095,N9096,N9097,N9098,N9099,N9100,N9101,N9102,N9103,N9104,
  N9105,N9106,N9107,N9108,N9109,N9110,N9111,N9112,N9113,N9114,N9115,N9116,N9117,
  N9118,N9119,N9120,N9121,N9122,N9123,N9124,N9125,N9126,N9127,N9128,N9129,N9130,
  N9131,N9132,N9133,N9134,N9135,N9136,N9137,N9138,N9139,N9140,N9141,N9142,N9143,N9144,
  N9145,N9146,N9147,N9148,N9149,N9150,N9151,N9152,N9153,N9154,N9155,N9156,N9157,
  N9158,N9159,N9160,N9161,N9162,N9163,N9164,N9165,N9166,N9167,N9168,N9169,N9170,
  N9171,N9172,N9173,N9174,N9175,N9176,N9177,N9178,N9179,N9180,N9181,N9182,N9183,N9184,
  N9185,N9186,N9187,N9188,N9189,N9190,N9191,N9192,N9193,N9194,N9195,N9196,N9197,
  N9198,N9199,N9200,N9201,N9202,N9203,N9204,N9205,N9206,N9207,N9208,N9209,N9210,
  N9211,N9212,N9213,N9214,N9215,N9216,N9217,N9218,N9219,N9220,N9221,N9222,N9223,N9224,
  N9225,N9226,N9227,N9228,N9229,N9230,N9231,N9232,N9233,N9234,N9235,N9236,N9237,
  N9238,N9239,N9240,N9241,N9242,N9243,N9244,N9245,N9246,N9247,N9248,N9249,N9250,
  N9251,N9252,N9253,N9254,N9255,N9256,N9257,N9258,N9259,N9260,N9261,N9262,N9263,N9264,
  N9265,N9266,N9267,N9268,N9269,N9270,N9271,N9272,N9273,N9274,N9275,N9276,N9277,
  N9278,N9279,N9280,N9281,N9282,N9283,N9284,N9285,N9286,N9287,N9288,N9289,N9290,
  N9291,N9292,N9293,N9294,N9295,N9296,N9297,N9298,N9299,N9300,N9301,N9302,N9303,N9304,
  N9305,N9306,N9307,N9308,N9309,N9310,N9311,N9312,N9313,N9314,N9315,N9316,N9317,
  N9318,N9319,N9320,N9321,N9322,N9323,N9324,N9325,N9326,N9327,N9328,N9329,N9330,
  N9331,N9332,N9333,N9334,N9335,N9336,N9337,N9338,N9339,N9340,N9341,N9342,N9343,N9344,
  N9345,N9346,N9347,N9348,N9349,N9350,N9351,N9352,N9353,N9354,N9355,N9356,N9357,
  N9358,N9359,N9360,N9361,N9362,N9363,N9364,N9365,N9366,N9367,N9368,N9369,N9370,
  N9371,N9372,N9373,N9374,N9375,N9376,N9377,N9378,N9379,N9380,N9381,N9382,N9383,N9384,
  N9385,N9386,N9387,N9388,N9389,N9390,N9391,N9392,N9393,N9394,N9395,N9396,N9397,
  N9398,N9399,N9400,N9401,N9402,N9403,N9404,N9405,N9406,N9407,N9408,N9409,N9410,
  N9411,N9412,N9413,N9414,N9415,N9416,N9417,N9418,N9419,N9420,N9421,N9422,N9423,N9424,
  N9425,N9426,N9427,N9428,N9429,N9430,N9431,N9432,N9433,N9434,N9435,N9436,N9437,
  N9438,N9439,N9440,N9441,N9442,N9443,N9444,N9445,N9446,N9447,N9448,N9449,N9450,
  N9451,N9452,N9453,N9454,N9455,N9456,N9457,N9458,N9459,N9460,N9461,N9462,N9463,N9464,
  N9465,N9466,N9467,N9468,N9469,N9470,N9471,N9472,N9473,N9474,N9475,N9476,N9477,
  N9478,N9479,N9480,N9481,N9482,N9483,N9484,N9485,N9486,N9487,N9488,N9489,N9490,
  N9491,N9492,N9493,N9494,N9495,N9496,N9497,N9498,N9499,N9500,N9501,N9502,N9503,N9504,
  N9505,N9506,N9507,N9508,N9509,N9510,N9511,N9512,N9513,N9514,N9515,N9516,N9517,
  N9518,N9519,N9520,N9521,N9522,N9523,N9524,N9525,N9526,N9527,N9528,N9529,N9530,
  N9531,N9532,N9533,N9534,N9535,N9536,N9537,N9538,N9539,N9540,N9541,N9542,N9543,N9544,
  N9545,N9546,N9547,N9548,N9549,N9550,N9551,N9552,N9553,N9554,N9555,N9556,N9557,
  N9558,N9559,N9560,N9561,N9562,N9563,N9564,N9565,N9566,N9567,N9568,N9569,N9570,
  N9571,N9572,N9573,N9574,N9575,N9576,N9577,N9578,N9579,N9580,N9581,N9582,N9583,N9584,
  N9585,N9586,N9587,N9588,N9589,N9590,N9591,N9592,N9593,N9594,N9595,N9596,N9597,
  N9598,N9599,N9600,N9601,N9602,N9603,N9604,N9605,N9606,N9607,N9608,N9609,N9610,
  N9611,N9612,N9613,N9614,N9615,N9616,N9617,N9618,N9619,N9620,N9621,N9622,N9623,N9624,
  N9625,N9626,N9627,N9628,N9629,N9630,N9631,N9632,N9633,N9634,N9635,N9636,N9637,
  N9638,N9639,N9640,N9641,N9642,N9643,N9644,N9645,N9646,N9647,N9648,N9649,N9650,
  N9651,N9652,N9653,N9654,N9655,N9656,N9657,N9658,N9659,N9660,N9661,N9662,N9663,N9664,
  N9665,N9666,N9667,N9668,N9669,N9670,N9671,N9672,N9673,N9674,N9675,N9676,N9677,
  N9678,N9679,N9680,N9681,N9682,N9683,N9684,N9685,N9686,N9687,N9688,N9689,N9690,
  N9691,N9692,N9693,N9694,N9695,N9696,N9697,N9698,N9699,N9700,N9701,N9702,N9703,N9704,
  N9705,N9706,N9707,N9708,N9709,N9710,N9711,N9712,N9713,N9714,N9715,N9716,N9717,
  N9718,N9719,N9720,N9721,N9722,N9723,N9724,N9725,N9726,N9727,N9728,N9729,N9730,
  N9731,N9732,N9733,N9734,N9735,N9736,N9737,N9738,N9739,N9740,N9741,N9742,N9743,N9744,
  N9745,N9746,N9747,N9748,N9749,N9750,N9751,N9752,N9753,N9754,N9755,N9756,N9757,
  N9758,N9759,N9760,N9761,N9762,N9763,N9764,N9765,N9766,N9767,N9768,N9769,N9770,
  N9771,N9772,N9773,N9774,N9775,N9776,N9777,N9778,N9779,N9780,N9781,N9782,N9783,N9784,
  N9785,N9786,N9787,N9788,N9789,N9790,N9791,N9792,N9793,N9794,N9795,N9796,N9797,
  N9798,N9799,N9800,N9801,N9802,N9803,N9804,N9805,N9806,N9807,N9808,N9809,N9810,
  N9811,N9812,N9813,N9814,N9815,N9816,N9817,N9818,N9819,N9820,N9821,N9822,N9823,N9824,
  N9825,N9826,N9827,N9828,N9829,N9830,N9831,N9832,N9833,N9834,N9835,N9836,N9837,
  N9838,N9839,N9840,N9841,N9842,N9843,N9844,N9845,N9846,N9847,N9848,N9849,N9850,
  N9851,N9852,N9853,N9854,N9855,N9856,N9857,N9858,N9859,N9860,N9861,N9862,N9863,N9864,
  N9865,N9866,N9867,N9868,N9869,N9870,N9871,N9872,N9873,N9874,N9875,N9876,N9877,
  N9878,N9879,N9880,N9881,N9882,N9883,N9884,N9885,N9886,N9887,N9888,N9889,N9890,
  N9891,N9892,N9893,N9894,N9895,N9896,N9897,N9898,N9899,N9900,N9901,N9902,N9903,N9904,
  N9905,N9906,N9907,N9908,N9909,N9910,N9911,N9912,N9913,N9914,N9915,N9916,N9917,
  N9918,N9919,N9920,N9921,N9922,N9923,N9924,N9925,N9926,N9927,N9928,N9929,N9930,
  N9931,N9932,N9933,N9934,N9935,N9936,N9937,N9938,N9939,N9940,N9941,N9942,N9943,N9944,
  N9945,N9946,N9947,N9948,N9949,N9950,N9951,N9952,N9953,N9954,N9955,N9956,N9957,
  N9958,N9959,N9960,N9961,N9962,N9963,N9964,N9965,N9966,N9967,N9968,N9969,N9970,
  N9971,N9972,N9973,N9974,N9975,N9976,N9977,N9978,N9979,N9980,N9981,N9982,N9983,N9984,
  N9985,N9986,N9987,N9988,N9989,N9990,N9991,N9992,N9993,N9994,N9995,N9996,N9997,
  N9998,N9999,N10000,N10001,N10002,N10003,N10004,N10005,N10006,N10007,N10008,N10009,
  N10010,N10011,N10012,N10013,N10014,N10015,N10016,N10017,N10018,N10019,N10020,
  N10021,N10022,N10023,N10024,N10025,N10026,N10027,N10028,N10029,N10030,N10031,
  N10032,N10033,N10034,N10035,N10036,N10037,N10038,N10039,N10040,N10041,N10042,N10043,
  N10044,N10045,N10046,N10047,N10048,N10049,N10050,N10051,N10052,N10053,N10054,
  N10055,N10056,N10057,N10058,N10059,N10060,N10061,N10062,N10063,N10064,N10065,N10066,
  N10067,N10068,N10069,N10070,N10071,N10072,N10073,N10074,N10075,N10076,N10077,
  N10078,N10079,N10080,N10081,N10082,N10083,N10084,N10085,N10086,N10087,N10088,N10089,
  N10090,N10091,N10092,N10093,N10094,N10095,N10096,N10097,N10098,N10099,N10100,
  N10101,N10102,N10103,N10104,N10105,N10106,N10107,N10108,N10109,N10110,N10111,
  N10112,N10113,N10114,N10115,N10116,N10117,N10118,N10119,N10120,N10121,N10122,N10123,
  N10124,N10125,N10126,N10127,N10128,N10129,N10130,N10131,N10132,N10133,N10134,
  N10135,N10136,N10137,N10138,N10139,N10140,N10141,N10142,N10143,N10144,N10145,N10146,
  N10147,N10148,N10149,N10150,N10151,N10152,N10153,N10154,N10155,N10156,N10157,
  N10158,N10159,N10160,N10161,N10162,N10163,N10164,N10165,N10166,N10167,N10168,N10169,
  N10170,N10171,N10172,N10173,N10174,N10175,N10176,N10177,N10178,N10179,N10180,
  N10181,N10182,N10183,N10184,N10185,N10186,N10187,N10188,N10189,N10190,N10191,
  N10192,N10193,N10194,N10195,N10196,N10197,N10198,N10199,N10200,N10201,N10202,N10203,
  N10204,N10205,N10206,N10207,N10208,N10209,N10210,N10211,N10212,N10213,N10214,
  N10215,N10216,N10217,N10218,N10219,N10220,N10221,N10222,N10223,N10224,N10225,N10226,
  N10227,N10228,N10229,N10230,N10231,N10232,N10233,N10234,N10235,N10236,N10237,
  N10238,N10239,N10240,N10241,N10242,N10243,N10244,N10245,N10246,N10247,N10248,N10249,
  N10250,N10251,N10252,N10253,N10254,N10255,N10256,N10257,N10258,N10259,N10260,
  N10261,N10262,N10263,N10264,N10265,N10266,N10267,N10268,N10269,N10270,N10271,
  N10272,N10273,N10274,N10275,N10276,N10277,N10278,N10279,N10280,N10281,N10282,N10283,
  N10284,N10285,N10286,N10287,N10288,N10289,N10290,N10291,N10292,N10293,N10294,
  N10295,N10296,N10297,N10298,N10299,N10300,N10301,N10302,N10303,N10304,N10305,N10306,
  N10307,N10308,N10309,N10310,N10311,N10312,N10313,N10314,N10315,N10316,N10317,
  N10318,N10319,N10320,N10321,N10322,N10323,N10324,N10325,N10326,N10327,N10328,N10329,
  N10330,N10331,N10332,N10333,N10334,N10335,N10336,N10337,N10338,N10339,N10340,
  N10341,N10342,N10343,N10344,N10345,N10346,N10347,N10348,N10349,N10350,N10351,
  N10352,N10353,N10354,N10355,N10356,N10357,N10358,N10359,N10360,N10361,N10362,N10363,
  N10364,N10365,N10366,N10367,N10368,N10369,N10370,N10371,N10372,N10373,N10374,
  N10375,N10376,N10377,N10378,N10379,N10380,N10381,N10382,N10383,N10384,N10385,N10386,
  N10387,N10388,N10389,N10390,N10391,N10392,N10393,N10394,N10395,N10396,N10397,
  N10398,N10399,N10400,N10401,N10402,N10403,N10404,N10405,N10406,N10407,N10408,N10409,
  N10410,N10411,N10412,N10413,N10414,N10415,N10416,N10417,N10418,N10419,N10420,
  N10421,N10422,N10423,N10424,N10425,N10426,N10427,N10428,N10429,N10430,N10431,
  N10432,N10433,N10434,N10435,N10436,N10437,N10438,N10439,N10440,N10441,N10442,N10443,
  N10444,N10445,N10446,N10447,N10448,N10449,N10450,N10451,N10452,N10453,N10454,
  N10455,N10456,N10457,N10458,N10459,N10460,N10461,N10462,N10463,N10464,N10465,N10466,
  N10467,N10468,N10469,N10470,N10471,N10472,N10473,N10474,N10475,N10476,N10477,
  N10478,N10479,N10480,N10481,N10482,N10483,N10484,N10485,N10486,N10487,N10488,N10489,
  N10490,N10491,N10492,N10493,N10494,N10495,N10496,N10497,N10498,N10499,N10500,
  N10501,N10502,N10503,N10504,N10505,N10506,N10507,N10508,N10509,N10510,N10511,
  N10512,N10513,N10514,N10515,N10516,N10517,N10518,N10519,N10520,N10521,N10522,N10523,
  N10524,N10525,N10526,N10527,N10528,N10529,N10530,N10531,N10532,N10533,N10534,
  N10535,N10536,N10537,N10538,N10539,N10540,N10541,N10542,N10543,N10544,N10545,N10546,
  N10547,N10548,N10549,N10550,N10551,N10552,N10553,N10554,N10555,N10556,N10557,
  N10558,N10559,N10560,N10561,N10562,N10563,N10564,N10565,N10566,N10567,N10568,N10569,
  N10570,N10571,N10572,N10573,N10574,N10575,N10576,N10577,N10578,N10579,N10580,
  N10581,N10582,N10583,N10584,N10585,N10586,N10587,N10588,N10589,N10590,N10591,
  N10592,N10593,N10594,N10595,N10596,N10597,N10598,N10599,N10600,N10601,N10602,N10603,
  N10604,N10605,N10606,N10607,N10608,N10609,N10610,N10611,N10612,N10613,N10614,
  N10615,N10616,N10617,N10618,N10619,N10620,N10621,N10622,N10623,N10624,N10625,N10626,
  N10627,N10628,N10629,N10630,N10631,N10632,N10633,N10634,N10635,N10636,N10637,
  N10638,N10639,N10640,N10641,N10642,N10643,N10644,N10645,N10646,N10647,N10648,N10649,
  N10650,N10651,N10652,N10653,N10654,N10655,N10656,N10657,N10658,N10659,N10660,
  N10661,N10662,N10663,N10664,N10665,N10666,N10667,N10668,N10669,N10670,N10671,
  N10672,N10673,N10674,N10675,N10676,N10677,N10678,N10679,N10680,N10681,N10682,N10683,
  N10684,N10685,N10686,N10687,N10688,N10689,N10690,N10691,N10692,N10693,N10694,
  N10695,N10696,N10697,N10698,N10699,N10700,N10701,N10702,N10703,N10704,N10705,N10706,
  N10707,N10708,N10709,N10710,N10711,N10712,N10713,N10714,N10715,N10716,N10717,
  N10718,N10719,N10720,N10721,N10722,N10723,N10724,N10725,N10726,N10727,N10728,N10729,
  N10730,N10731,N10732,N10733,N10734,N10735,N10736,N10737,N10738,N10739,N10740,
  N10741,N10742,N10743,N10744,N10745,N10746,N10747,N10748,N10749,N10750,N10751,
  N10752,N10753,N10754,N10755,N10756,N10757,N10758,N10759,N10760,N10761,N10762,N10763,
  N10764,N10765,N10766,N10767,N10768,N10769,N10770,N10771,N10772,N10773,N10774,
  N10775,N10776,N10777,N10778,N10779,N10780,N10781,N10782,N10783,N10784,N10785,N10786,
  N10787,N10788,N10789,N10790,N10791,N10792,N10793,N10794,N10795,N10796,N10797,
  N10798,N10799,N10800,N10801,N10802,N10803,N10804,N10805,N10806,N10807,N10808,N10809,
  N10810,N10811,N10812,N10813,N10814,N10815,N10816,N10817,N10818,N10819,N10820,
  N10821,N10822,N10823,N10824,N10825,N10826,N10827,N10828,N10829,N10830,N10831,
  N10832,N10833,N10834,N10835,N10836,N10837,N10838,N10839,N10840,N10841,N10842,N10843,
  N10844,N10845,N10846,N10847,N10848,N10849,N10850,N10851,N10852,N10853,N10854,
  N10855,N10856,N10857,N10858,N10859,N10860,N10861,N10862,N10863,N10864,N10865,N10866,
  N10867,N10868,N10869,N10870,N10871,N10872,N10873,N10874,N10875,N10876,N10877,
  N10878,N10879,N10880,N10881,N10882,N10883,N10884,N10885,N10886,N10887,N10888,N10889,
  N10890,N10891,N10892,N10893,N10894,N10895,N10896,N10897,N10898,N10899,N10900,
  N10901,N10902,N10903,N10904,N10905,N10906,N10907,N10908,N10909,N10910,N10911,
  N10912,N10913,N10914,N10915,N10916,N10917,N10918,N10919,N10920,N10921,N10922,N10923,
  N10924,N10925,N10926,N10927,N10928,N10929,N10930,N10931,N10932,N10933,N10934,
  N10935,N10936,N10937,N10938,N10939,N10940,N10941,N10942,N10943,N10944,N10945,N10946,
  N10947,N10948,N10949,N10950,N10951,N10952,N10953,N10954,N10955,N10956,N10957,
  N10958,N10959,N10960,N10961,N10962,N10963,N10964,N10965,N10966,N10967,N10968,N10969,
  N10970,N10971,N10972,N10973,N10974,N10975,N10976,N10977,N10978,N10979,N10980,
  N10981,N10982,N10983,N10984,N10985,N10986,N10987,N10988,N10989,N10990,N10991,
  N10992,N10993,N10994,N10995,N10996,N10997,N10998,N10999,N11000,N11001,N11002,N11003,
  N11004,N11005,N11006,N11007,N11008,N11009,N11010,N11011,N11012,N11013,N11014,
  N11015,N11016,N11017,N11018,N11019,N11020,N11021,N11022,N11023,N11024,N11025,N11026,
  N11027,N11028,N11029,N11030,N11031,N11032,N11033,N11034,N11035,N11036,N11037,
  N11038,N11039,N11040,N11041,N11042,N11043,N11044,N11045,N11046,N11047,N11048,N11049,
  N11050,N11051,N11052,N11053,N11054,N11055,N11056,N11057,N11058,N11059,N11060,
  N11061,N11062,N11063,N11064,N11065,N11066,N11067,N11068,N11069,N11070,N11071,
  N11072,N11073,N11074,N11075,N11076,N11077,N11078,N11079,N11080,N11081,N11082,N11083,
  N11084,N11085,N11086,N11087,N11088,N11089,N11090,N11091,N11092,N11093,N11094,
  N11095,N11096,N11097,N11098,N11099,N11100,N11101,N11102,N11103,N11104,N11105,N11106,
  N11107,N11108,N11109,N11110,N11111,N11112,N11113,N11114,N11115,N11116,N11117,
  N11118,N11119,N11120,N11121,N11122,N11123,N11124,N11125,N11126,N11127,N11128,N11129,
  N11130,N11131,N11132,N11133,N11134,N11135,N11136,N11137,N11138,N11139,N11140,
  N11141,N11142,N11143,N11144,N11145,N11146,N11147,N11148,N11149,N11150,N11151,
  N11152,N11153,N11154,N11155,N11156,N11157,N11158,N11159,N11160,N11161,N11162,N11163,
  N11164,N11165,N11166,N11167,N11168,N11169,N11170,N11171,N11172,N11173,N11174,
  N11175,N11176,N11177,N11178,N11179,N11180,N11181,N11182,N11183,N11184,N11185,N11186,
  N11187,N11188,N11189,N11190,N11191,N11192,N11193,N11194,N11195,N11196,N11197,
  N11198,N11199,N11200,N11201,N11202,N11203,N11204,N11205,N11206,N11207,N11208,N11209,
  N11210,N11211,N11212,N11213,N11214,N11215,N11216,N11217,N11218,N11219,N11220,
  N11221,N11222,N11223,N11224,N11225,N11226,N11227,N11228,N11229,N11230,N11231,
  N11232,N11233,N11234,N11235,N11236,N11237,N11238,N11239,N11240,N11241,N11242,N11243,
  N11244,N11245,N11246,N11247,N11248,N11249,N11250,N11251,N11252,N11253,N11254,
  N11255,N11256,N11257,N11258,N11259,N11260,N11261,N11262,N11263,N11264,N11265,N11266,
  N11267,N11268,N11269,N11270,N11271,N11272,N11273,N11274,N11275,N11276,N11277,
  N11278,N11279,N11280,N11281,N11282,N11283,N11284,N11285,N11286,N11287,N11288,N11289,
  N11290,N11291,N11292,N11293,N11294,N11295,N11296,N11297,N11298,N11299,N11300,
  N11301,N11302,N11303,N11304,N11305,N11306,N11307,N11308,N11309,N11310,N11311,
  N11312,N11313,N11314,N11315,N11316,N11317,N11318,N11319,N11320,N11321,N11322,N11323,
  N11324,N11325,N11326,N11327,N11328,N11329,N11330,N11331,N11332,N11333,N11334,
  N11335,N11336,N11337,N11338,N11339,N11340,N11341,N11342,N11343,N11344,N11345,N11346,
  N11347,N11348,N11349,N11350,N11351,N11352,N11353,N11354,N11355,N11356,N11357,
  N11358,N11359,N11360,N11361,N11362,N11363,N11364,N11365,N11366,N11367,N11368,N11369,
  N11370,N11371,N11372,N11373,N11374,N11375,N11376,N11377,N11378,N11379,N11380,
  N11381,N11382,N11383,N11384,N11385,N11386,N11387,N11388,N11389,N11390,N11391,
  N11392,N11393,N11394,N11395,N11396,N11397,N11398,N11399,N11400,N11401,N11402,N11403,
  N11404,N11405,N11406,N11407,N11408,N11409,N11410,N11411,N11412,N11413,N11414,
  N11415,N11416,N11417,N11418,N11419,N11420,N11421,N11422,N11423,N11424,N11425,N11426,
  N11427,N11428,N11429,N11430,N11431,N11432,N11433,N11434,N11435,N11436,N11437,
  N11438,N11439,N11440,N11441,N11442,N11443,N11444,N11445,N11446,N11447,N11448,N11449,
  N11450,N11451,N11452,N11453,N11454,N11455,N11456,N11457,N11458,N11459,N11460,
  N11461,N11462,N11463,N11464,N11465,N11466,N11467,N11468,N11469,N11470,N11471,
  N11472,N11473,N11474,N11475,N11476,N11477,N11478,N11479,N11480,N11481,N11482,N11483,
  N11484,N11485,N11486,N11487,N11488,N11489,N11490,N11491,N11492,N11493,N11494,
  N11495,N11496,N11497,N11498,N11499,N11500,N11501,N11502,N11503,N11504,N11505,N11506,
  N11507,N11508,N11509,N11510,N11511,N11512,N11513,N11514,N11515,N11516,N11517,
  N11518,N11519,N11520,N11521,N11522,N11523,N11524,N11525,N11526,N11527,N11528,N11529,
  N11530,N11531,N11532,N11533,N11534,N11535,N11536,N11537,N11538,N11539,N11540,
  N11541,N11542,N11543,N11544,N11545,N11546,N11547,N11548,N11549,N11550,N11551,
  N11552,N11553,N11554,N11555,N11556,N11557,N11558,N11559,N11560,N11561,N11562,N11563,
  N11564,N11565,N11566,N11567,N11568,N11569,N11570,N11571,N11572,N11573,N11574,
  N11575,N11576,N11577,N11578,N11579,N11580,N11581,N11582,N11583,N11584,N11585,N11586,
  N11587,N11588,N11589,N11590,N11591,N11592,N11593,N11594,N11595,N11596,N11597,
  N11598,N11599,N11600,N11601,N11602,N11603,N11604,N11605,N11606,N11607,N11608,N11609,
  N11610,N11611,N11612,N11613,N11614,N11615,N11616,N11617,N11618,N11619,N11620,
  N11621,N11622,N11623,N11624,N11625,N11626,N11627,N11628,N11629,N11630,N11631,
  N11632,N11633,N11634,N11635,N11636,N11637,N11638,N11639,N11640,N11641,N11642,N11643,
  N11644,N11645,N11646,N11647,N11648,N11649,N11650,N11651,N11652,N11653,N11654,
  N11655,N11656,N11657,N11658,N11659,N11660,N11661,N11662,N11663,N11664,N11665,N11666,
  N11667,N11668,N11669,N11670,N11671,N11672,N11673,N11674,N11675,N11676,N11677,
  N11678,N11679,N11680,N11681,N11682,N11683,N11684,N11685,N11686,N11687,N11688,N11689,
  N11690,N11691,N11692,N11693,N11694,N11695,N11696,N11697,N11698,N11699,N11700,
  N11701,N11702,N11703,N11704,N11705,N11706,N11707,N11708,N11709,N11710,N11711,
  N11712,N11713,N11714,N11715,N11716,N11717,N11718,N11719,N11720,N11721,N11722,N11723,
  N11724,N11725,N11726,N11727,N11728,N11729,N11730,N11731,N11732,N11733,N11734,
  N11735,N11736,N11737,N11738,N11739,N11740,N11741,N11742,N11743,N11744,N11745,N11746,
  N11747,N11748,N11749,N11750,N11751,N11752,N11753,N11754,N11755,N11756,N11757,
  N11758,N11759,N11760,N11761,N11762,N11763,N11764,N11765,N11766,N11767,N11768,N11769,
  N11770,N11771,N11772,N11773,N11774,N11775,N11776,N11777,N11778,N11779,N11780,
  N11781,N11782,N11783,N11784,N11785,N11786,N11787,N11788,N11789,N11790,N11791,
  N11792,N11793,N11794,N11795,N11796,N11797,N11798,N11799,N11800,N11801,N11802,N11803,
  N11804,N11805,N11806,N11807,N11808,N11809,N11810,N11811,N11812,N11813,N11814,
  N11815,N11816,N11817,N11818,N11819,N11820,N11821,N11822,N11823,N11824,N11825,N11826,
  N11827,N11828,N11829,N11830,N11831,N11832,N11833,N11834,N11835,N11836,N11837,
  N11838,N11839,N11840,N11841,N11842,N11843,N11844,N11845,N11846,N11847,N11848,N11849,
  N11850,N11851,N11852,N11853,N11854,N11855,N11856,N11857,N11858,N11859,N11860,
  N11861,N11862,N11863,N11864,N11865,N11866,N11867,N11868,N11869,N11870,N11871,
  N11872,N11873,N11874,N11875,N11876,N11877,N11878,N11879,N11880,N11881,N11882,N11883,
  N11884,N11885,N11886,N11887,N11888,N11889,N11890,N11891,N11892,N11893,N11894,
  N11895,N11896,N11897,N11898,N11899,N11900,N11901,N11902,N11903,N11904,N11905,N11906,
  N11907,N11908,N11909,N11910,N11911,N11912,N11913,N11914,N11915,N11916,N11917,
  N11918,N11919,N11920,N11921,N11922,N11923,N11924,N11925,N11926,N11927,N11928,N11929,
  N11930,N11931,N11932,N11933,N11934,N11935,N11936,N11937,N11938,N11939,N11940,
  N11941,N11942,N11943,N11944,N11945,N11946,N11947,N11948,N11949,N11950,N11951,
  N11952,N11953,N11954,N11955,N11956,N11957,N11958,N11959,N11960,N11961,N11962,N11963,
  N11964,N11965,N11966,N11967,N11968,N11969,N11970,N11971,N11972,N11973,N11974,
  N11975,N11976,N11977,N11978,N11979,N11980,N11981,N11982,N11983,N11984,N11985,N11986,
  N11987,N11988,N11989,N11990,N11991,N11992,N11993,N11994,N11995,N11996,N11997,
  N11998,N11999,N12000,N12001,N12002,N12003,N12004,N12005,N12006,N12007,N12008,N12009,
  N12010,N12011,N12012,N12013,N12014,N12015,N12016,N12017,N12018,N12019,N12020,
  N12021,N12022,N12023,N12024,N12025,N12026,N12027,N12028,N12029,N12030,N12031,
  N12032,N12033,N12034,N12035,N12036,N12037,N12038,N12039,N12040,N12041,N12042,N12043,
  N12044,N12045,N12046,N12047,N12048,N12049,N12050,N12051,N12052,N12053,N12054,
  N12055,N12056,N12057,N12058,N12059,N12060,N12061,N12062,N12063,N12064,N12065,N12066,
  N12067,N12068,N12069,N12070,N12071,N12072,N12073,N12074,N12075,N12076,N12077,
  N12078,N12079,N12080,N12081,N12082,N12083,N12084,N12085,N12086,N12087,N12088,N12089,
  N12090,N12091,N12092,N12093,N12094,N12095,N12096,N12097,N12098,N12099,N12100,
  N12101,N12102,N12103,N12104,N12105,N12106,N12107,N12108,N12109,N12110,N12111,
  N12112,N12113,N12114,N12115,N12116,N12117,N12118,N12119,N12120,N12121,N12122,N12123,
  N12124,N12125,N12126,N12127,N12128,N12129,N12130,N12131,N12132,N12133,N12134,
  N12135,N12136,N12137,N12138,N12139,N12140,N12141,N12142,N12143,N12144,N12145,N12146,
  N12147,N12148,N12149,N12150,N12151,N12152,N12153,N12154,N12155,N12156,N12157,
  N12158,N12159,N12160,N12161,N12162,N12163,N12164,N12165,N12166,N12167,N12168,N12169,
  N12170,N12171,N12172,N12173,N12174,N12175,N12176,N12177,N12178,N12179,N12180,
  N12181,N12182,N12183,N12184,N12185,N12186,N12187,N12188,N12189,N12190,N12191,
  N12192,N12193,N12194,N12195,N12196,N12197,N12198,N12199,N12200,N12201,N12202,N12203,
  N12204,N12205,N12206,N12207,N12208,N12209,N12210,N12211,N12212,N12213,N12214,
  N12215,N12216,N12217,N12218,N12219,N12220,N12221,N12222,N12223,N12224,N12225,N12226,
  N12227,N12228,N12229,N12230,N12231,N12232,N12233,N12234,N12235,N12236,N12237,
  N12238,N12239,N12240,N12241,N12242,N12243,N12244,N12245,N12246,N12247,N12248,N12249,
  N12250,N12251,N12252,N12253,N12254,N12255,N12256,N12257,N12258,N12259,N12260,
  N12261,N12262,N12263,N12264,N12265,N12266,N12267,N12268,N12269,N12270,N12271,
  N12272,N12273,N12274,N12275,N12276,N12277,N12278,N12279,N12280,N12281,N12282,N12283,
  N12284,N12285,N12286,N12287,N12288,N12289,N12290,N12291,N12292,N12293,N12294,
  N12295,N12296,N12297,N12298,N12299,N12300,N12301,N12302,N12303,N12304,N12305,N12306,
  N12307,N12308,N12309,N12310,N12311,N12312,N12313,N12314,N12315,N12316,N12317,
  N12318,N12319,N12320,N12321,N12322,N12323,N12324,N12325,N12326,N12327,N12328,N12329,
  N12330,N12331,N12332,N12333,N12334,N12335,N12336,N12337,N12338,N12339,N12340,
  N12341,N12342,N12343,N12344,N12345,N12346,N12347,N12348,N12349,N12350,N12351,
  N12352,N12353,N12354,N12355,N12356,N12357,N12358,N12359,N12360,N12361,N12362,N12363,
  N12364,N12365,N12366,N12367,N12368,N12369,N12370,N12371,N12372,N12373,N12374,
  N12375,N12376,N12377,N12378,N12379,N12380,N12381,N12382,N12383,N12384,N12385,N12386,
  N12387,N12388,N12389,N12390,N12391,N12392,N12393,N12394,N12395,N12396,N12397,
  N12398,N12399,N12400,N12401,N12402,N12403,N12404,N12405,N12406,N12407,N12408,N12409,
  N12410,N12411,N12412,N12413,N12414,N12415,N12416,N12417,N12418,N12419,N12420,
  N12421,N12422,N12423,N12424,N12425,N12426,N12427,N12428,N12429,N12430,N12431,
  N12432,N12433,N12434,N12435,N12436,N12437,N12438,N12439,N12440,N12441,N12442,N12443,
  N12444,N12445,N12446,N12447,N12448,N12449,N12450,N12451,N12452,N12453,N12454,
  N12455,N12456,N12457,N12458,N12459,N12460,N12461,N12462,N12463,N12464,N12465,N12466,
  N12467,N12468,N12469,N12470,N12471,N12472,N12473,N12474,N12475,N12476,N12477,
  N12478,N12479,N12480,N12481,N12482,N12483,N12484,N12485,N12486,N12487,N12488,N12489,
  N12490,N12491,N12492,N12493,N12494,N12495,N12496,N12497,N12498,N12499,N12500,
  N12501,N12502,N12503,N12504,N12505,N12506,N12507,N12508,N12509,N12510,N12511,
  N12512,N12513,N12514,N12515,N12516,N12517,N12518,N12519,N12520,N12521,N12522,N12523,
  N12524,N12525,N12526,N12527,N12528,N12529,N12530,N12531,N12532,N12533,N12534,
  N12535,N12536,N12537,N12538,N12539,N12540,N12541,N12542,N12543,N12544,N12545,N12546,
  N12547,N12548,N12549,N12550,N12551,N12552,N12553,N12554,N12555,N12556,N12557,
  N12558,N12559,N12560,N12561,N12562,N12563,N12564,N12565,N12566,N12567,N12568,N12569,
  N12570,N12571,N12572,N12573,N12574,N12575,N12576,N12577,N12578,N12579,N12580,
  N12581,N12582,N12583,N12584,N12585,N12586,N12587,N12588,N12589,N12590,N12591,
  N12592,N12593,N12594,N12595,N12596,N12597,N12598,N12599,N12600,N12601,N12602,N12603,
  N12604,N12605,N12606,N12607,N12608,N12609,N12610,N12611,N12612,N12613,N12614,
  N12615,N12616,N12617,N12618,N12619,N12620,N12621,N12622,N12623,N12624,N12625,N12626,
  N12627,N12628,N12629,N12630,N12631,N12632,N12633,N12634,N12635,N12636,N12637,
  N12638,N12639,N12640,N12641,N12642,N12643,N12644,N12645,N12646,N12647,N12648,N12649,
  N12650,N12651,N12652,N12653,N12654,N12655,N12656,N12657,N12658,N12659,N12660,
  N12661,N12662,N12663,N12664,N12665,N12666,N12667,N12668,N12669,N12670,N12671,
  N12672,N12673,N12674,N12675,N12676,N12677,N12678,N12679,N12680,N12681,N12682,N12683,
  N12684,N12685,N12686,N12687,N12688,N12689,N12690,N12691,N12692,N12693,N12694,
  N12695,N12696,N12697,N12698,N12699,N12700,N12701,N12702,N12703,N12704,N12705,N12706,
  N12707,N12708,N12709,N12710,N12711,N12712,N12713,N12714,N12715,N12716,N12717,
  N12718,N12719,N12720,N12721,N12722,N12723,N12724,N12725,N12726,N12727,N12728,N12729,
  N12730,N12731,N12732,N12733,N12734,N12735,N12736,N12737,N12738,N12739,N12740,
  N12741,N12742,N12743,N12744,N12745,N12746,N12747,N12748,N12749,N12750,N12751,
  N12752,N12753,N12754,N12755,N12756,N12757,N12758,N12759,N12760,N12761,N12762,N12763,
  N12764,N12765,N12766,N12767,N12768,N12769,N12770,N12771,N12772,N12773,N12774,
  N12775,N12776,N12777,N12778,N12779,N12780,N12781,N12782,N12783,N12784,N12785,N12786,
  N12787,N12788,N12789,N12790,N12791,N12792,N12793,N12794,N12795,N12796,N12797,
  N12798,N12799,N12800,N12801,N12802,N12803,N12804,N12805,N12806,N12807,N12808,N12809,
  N12810,N12811,N12812,N12813,N12814,N12815,N12816,N12817,N12818,N12819,N12820,
  N12821,N12822,N12823,N12824,N12825,N12826,N12827,N12828,N12829,N12830,N12831,
  N12832,N12833,N12834,N12835,N12836,N12837,N12838,N12839,N12840,N12841,N12842,N12843,
  N12844,N12845,N12846,N12847,N12848,N12849,N12850,N12851,N12852,N12853,N12854,
  N12855,N12856,N12857,N12858,N12859,N12860,N12861,N12862,N12863,N12864,N12865,N12866,
  N12867,N12868,N12869,N12870,N12871,N12872,N12873,N12874,N12875,N12876,N12877,
  N12878,N12879,N12880,N12881,N12882,N12883,N12884,N12885,N12886,N12887,N12888,N12889,
  N12890,N12891,N12892,N12893,N12894,N12895,N12896,N12897,N12898,N12899,N12900,
  N12901,N12902,N12903,N12904,N12905,N12906,N12907,N12908,N12909,N12910,N12911,
  N12912,N12913,N12914,N12915,N12916,N12917,N12918,N12919,N12920,N12921,N12922,N12923,
  N12924,N12925,N12926,N12927,N12928,N12929,N12930,N12931,N12932,N12933,N12934,
  N12935,N12936,N12937,N12938,N12939,N12940,N12941,N12942,N12943,N12944,N12945,N12946,
  N12947,N12948,N12949,N12950,N12951,N12952,N12953,N12954,N12955,N12956,N12957,
  N12958,N12959,N12960,N12961,N12962,N12963,N12964,N12965,N12966,N12967,N12968,N12969,
  N12970,N12971,N12972,N12973,N12974,N12975,N12976,N12977,N12978,N12979,N12980,
  N12981,N12982,N12983,N12984,N12985,N12986,N12987,N12988,N12989,N12990,N12991,
  N12992,N12993,N12994,N12995,N12996,N12997,N12998,N12999,N13000,N13001,N13002,N13003,
  N13004,N13005,N13006,N13007,N13008,N13009,N13010,N13011,N13012,N13013,N13014,
  N13015,N13016,N13017,N13018,N13019,N13020,N13021,N13022,N13023,N13024,N13025,N13026,
  N13027,N13028,N13029,N13030,N13031,N13032,N13033,N13034,N13035,N13036,N13037,
  N13038,N13039,N13040,N13041,N13042,N13043,N13044,N13045,N13046,N13047,N13048,N13049,
  N13050,N13051,N13052,N13053,N13054,N13055,N13056,N13057,N13058,N13059,N13060,
  N13061,N13062,N13063,N13064,N13065,N13066,N13067,N13068,N13069,N13070,N13071,
  N13072,N13073,N13074,N13075,N13076,N13077,N13078,N13079,N13080,N13081,N13082,N13083,
  N13084,N13085,N13086,N13087,N13088,N13089,N13090,N13091,N13092,N13093,N13094,
  N13095,N13096,N13097,N13098,N13099,N13100,N13101,N13102,N13103,N13104,N13105,N13106,
  N13107,N13108,N13109,N13110,N13111,N13112,N13113,N13114,N13115,N13116,N13117,
  N13118,N13119,N13120,N13121,N13122,N13123,N13124,N13125,N13126,N13127,N13128,N13129,
  N13130,N13131,N13132,N13133,N13134,N13135,N13136,N13137,N13138,N13139,N13140,
  N13141,N13142,N13143,N13144,N13145,N13146,N13147,N13148,N13149,N13150,N13151,
  N13152,N13153,N13154,N13155,N13156,N13157,N13158,N13159,N13160,N13161,N13162,N13163,
  N13164,N13165,N13166,N13167,N13168,N13169,N13170,N13171,N13172,N13173,N13174,
  N13175,N13176,N13177,N13178,N13179,N13180,N13181,N13182,N13183,N13184,N13185,N13186,
  N13187,N13188,N13189,N13190,N13191,N13192,N13193,N13194,N13195,N13196,N13197,
  N13198,N13199,N13200,N13201,N13202,N13203,N13204,N13205,N13206,N13207,N13208,N13209,
  N13210,N13211,N13212,N13213,N13214,N13215,N13216,N13217,N13218,N13219,N13220,
  N13221,N13222,N13223,N13224,N13225,N13226,N13227,N13228,N13229,N13230,N13231,
  N13232,N13233,N13234,N13235,N13236,N13237,N13238,N13239,N13240,N13241,N13242,N13243,
  N13244,N13245,N13246,N13247,N13248,N13249,N13250,N13251,N13252,N13253,N13254,
  N13255,N13256,N13257,N13258,N13259,N13260,N13261,N13262,N13263,N13264,N13265,N13266,
  N13267,N13268,N13269,N13270,N13271,N13272,N13273,N13274,N13275,N13276,N13277,
  N13278,N13279,N13280,N13281,N13282,N13283,N13284,N13285,N13286,N13287,N13288,N13289,
  N13290,N13291,N13292,N13293,N13294,N13295,N13296,N13297,N13298,N13299,N13300,
  N13301,N13302,N13303,N13304,N13305,N13306,N13307,N13308,N13309,N13310,N13311,
  N13312,N13313,N13314,N13315,N13316,N13317,N13318,N13319,N13320,N13321,N13322,N13323,
  N13324,N13325,N13326,N13327,N13328,N13329,N13330,N13331,N13332,N13333,N13334,
  N13335,N13336,N13337,N13338,N13339,N13340,N13341,N13342,N13343,N13344,N13345,N13346,
  N13347,N13348,N13349,N13350,N13351,N13352,N13353,N13354,N13355,N13356,N13357,
  N13358,N13359,N13360,N13361,N13362,N13363,N13364,N13365,N13366,N13367,N13368,N13369,
  N13370,N13371,N13372,N13373,N13374,N13375,N13376,N13377,N13378,N13379,N13380,
  N13381,N13382,N13383,N13384,N13385,N13386,N13387,N13388,N13389,N13390,N13391,
  N13392,N13393,N13394,N13395,N13396,N13397,N13398,N13399,N13400,N13401,N13402,N13403,
  N13404,N13405,N13406,N13407,N13408,N13409,N13410,N13411,N13412,N13413,N13414,
  N13415,N13416,N13417,N13418,N13419,N13420,N13421,N13422,N13423,N13424,N13425,N13426,
  N13427,N13428,N13429,N13430,N13431,N13432,N13433,N13434,N13435,N13436,N13437,
  N13438,N13439,N13440,N13441,N13442,N13443,N13444,N13445,N13446,N13447,N13448,N13449,
  N13450,N13451,N13452,N13453,N13454,N13455,N13456,N13457,N13458,N13459,N13460,
  N13461,N13462,N13463,N13464,N13465,N13466,N13467,N13468,N13469,N13470,N13471,
  N13472,N13473,N13474,N13475,N13476,N13477,N13478,N13479,N13480,N13481,N13482,N13483,
  N13484,N13485,N13486,N13487,N13488,N13489,N13490,N13491,N13492,N13493,N13494,
  N13495,N13496,N13497,N13498,N13499,N13500,N13501,N13502,N13503,N13504,N13505,N13506,
  N13507,N13508,N13509,N13510,N13511,N13512,N13513,N13514,N13515,N13516,N13517,
  N13518,N13519,N13520,N13521,N13522,N13523,N13524,N13525,N13526,N13527,N13528,N13529,
  N13530,N13531,N13532,N13533,N13534,N13535,N13536,N13537,N13538,N13539,N13540,
  N13541,N13542,N13543,N13544,N13545,N13546,N13547,N13548,N13549,N13550,N13551,
  N13552,N13553,N13554,N13555,N13556,N13557,N13558,N13559,N13560,N13561,N13562,N13563,
  N13564,N13565,N13566,N13567,N13568,N13569,N13570,N13571,N13572,N13573,N13574,
  N13575,N13576,N13577,N13578,N13579,N13580,N13581,N13582,N13583,N13584,N13585,N13586,
  N13587,N13588,N13589,N13590,N13591,N13592,N13593,N13594,N13595,N13596,N13597,
  N13598,N13599,N13600,N13601,N13602,N13603,N13604,N13605,N13606,N13607,N13608,N13609,
  N13610,N13611,N13612,N13613,N13614,N13615,N13616,N13617,N13618,N13619,N13620,
  N13621,N13622,N13623,N13624,N13625,N13626,N13627,N13628,N13629,N13630,N13631,
  N13632,N13633,N13634,N13635,N13636,N13637,N13638,N13639,N13640,N13641,N13642,N13643,
  N13644,N13645,N13646,N13647,N13648,N13649,N13650,N13651,N13652,N13653,N13654,
  N13655,N13656,N13657,N13658,N13659,N13660,N13661,N13662,N13663,N13664,N13665,N13666,
  N13667,N13668,N13669,N13670,N13671,N13672,N13673,N13674,N13675,N13676,N13677,
  N13678,N13679,N13680,N13681,N13682,N13683,N13684,N13685,N13686,N13687,N13688,N13689,
  N13690,N13691,N13692,N13693,N13694,N13695,N13696,N13697,N13698,N13699,N13700,
  N13701,N13702,N13703,N13704,N13705,N13706,N13707,N13708,N13709,N13710,N13711,
  N13712,N13713,N13714,N13715,N13716,N13717,N13718,N13719,N13720,N13721,N13722,N13723,
  N13724,N13725,N13726,N13727,N13728,N13729,N13730,N13731,N13732,N13733,N13734,
  N13735,N13736,N13737,N13738,N13739,N13740,N13741,N13742,N13743,N13744,N13745,N13746,
  N13747,N13748,N13749,N13750,N13751,N13752,N13753,N13754,N13755,N13756,N13757,
  N13758,N13759,N13760,N13761,N13762,N13763,N13764,N13765,N13766,N13767,N13768,N13769,
  N13770,N13771,N13772,N13773,N13774,N13775,N13776,N13777,N13778,N13779,N13780,
  N13781,N13782,N13783,N13784,N13785,N13786,N13787,N13788,N13789,N13790,N13791,
  N13792,N13793,N13794,N13795,N13796,N13797,N13798,N13799,N13800,N13801,N13802,N13803,
  N13804,N13805,N13806,N13807,N13808,N13809,N13810,N13811,N13812,N13813,N13814,
  N13815,N13816,N13817,N13818,N13819,N13820,N13821,N13822,N13823,N13824,N13825,N13826,
  N13827,N13828,N13829,N13830,N13831,N13832,N13833,N13834,N13835,N13836,N13837,
  N13838,N13839,N13840,N13841,N13842,N13843,N13844,N13845,N13846,N13847,N13848,N13849,
  N13850,N13851,N13852,N13853,N13854,N13855,N13856,N13857,N13858,N13859,N13860,
  N13861,N13862,N13863,N13864,N13865,N13866,N13867,N13868,N13869,N13870,N13871,
  N13872,N13873,N13874,N13875,N13876,N13877,N13878,N13879,N13880,N13881,N13882,N13883,
  N13884,N13885,N13886,N13887,N13888,N13889,N13890,N13891,N13892,N13893,N13894,
  N13895,N13896,N13897,N13898,N13899,N13900,N13901,N13902,N13903,N13904,N13905,N13906,
  N13907,N13908,N13909,N13910,N13911,N13912,N13913,N13914,N13915,N13916,N13917,
  N13918,N13919,N13920,N13921,N13922,N13923,N13924,N13925,N13926,N13927,N13928,N13929,
  N13930,N13931,N13932,N13933,N13934,N13935,N13936,N13937,N13938,N13939,N13940,
  N13941,N13942,N13943,N13944,N13945,N13946,N13947,N13948,N13949,N13950,N13951,
  N13952,N13953,N13954,N13955,N13956,N13957,N13958,N13959,N13960,N13961,N13962,N13963,
  N13964,N13965,N13966,N13967,N13968,N13969,N13970,N13971,N13972,N13973,N13974,
  N13975,N13976,N13977,N13978,N13979,N13980,N13981,N13982,N13983,N13984,N13985,N13986,
  N13987,N13988,N13989,N13990,N13991,N13992,N13993,N13994,N13995,N13996,N13997,
  N13998,N13999,N14000,N14001,N14002,N14003,N14004,N14005,N14006,N14007,N14008,N14009,
  N14010,N14011,N14012,N14013,N14014,N14015,N14016,N14017,N14018,N14019,N14020,
  N14021,N14022,N14023,N14024,N14025,N14026,N14027,N14028,N14029,N14030,N14031,
  N14032,N14033,N14034,N14035,N14036,N14037,N14038,N14039,N14040,N14041,N14042,N14043,
  N14044,N14045,N14046,N14047,N14048,N14049,N14050,N14051,N14052,N14053,N14054,
  N14055,N14056,N14057,N14058,N14059,N14060,N14061,N14062,N14063,N14064,N14065,N14066,
  N14067,N14068,N14069,N14070,N14071,N14072,N14073,N14074,N14075,N14076,N14077,
  N14078,N14079,N14080,N14081,N14082,N14083,N14084,N14085,N14086,N14087,N14088,N14089,
  N14090,N14091,N14092,N14093,N14094,N14095,N14096,N14097,N14098,N14099,N14100,
  N14101,N14102,N14103,N14104,N14105,N14106,N14107,N14108,N14109,N14110,N14111,
  N14112,N14113,N14114,N14115,N14116,N14117,N14118,N14119,N14120,N14121,N14122,N14123,
  N14124,N14125,N14126,N14127,N14128,N14129,N14130,N14131,N14132,N14133,N14134,
  N14135,N14136,N14137,N14138,N14139,N14140,N14141,N14142,N14143,N14144,N14145,N14146,
  N14147,N14148,N14149,N14150,N14151,N14152,N14153,N14154,N14155,N14156,N14157,
  N14158,N14159,N14160,N14161,N14162,N14163,N14164,N14165,N14166,N14167,N14168,N14169,
  N14170,N14171,N14172,N14173,N14174,N14175,N14176,N14177,N14178,N14179,N14180,
  N14181,N14182,N14183,N14184,N14185,N14186,N14187,N14188,N14189,N14190,N14191,
  N14192,N14193,N14194,N14195,N14196,N14197,N14198,N14199,N14200,N14201,N14202,N14203,
  N14204,N14205,N14206,N14207,N14208,N14209,N14210,N14211,N14212,N14213,N14214,
  N14215,N14216,N14217,N14218,N14219,N14220,N14221,N14222,N14223,N14224,N14225,N14226,
  N14227,N14228,N14229,N14230,N14231,N14232,N14233,N14234,N14235,N14236,N14237,
  N14238,N14239,N14240,N14241,N14242,N14243,N14244,N14245,N14246,N14247,N14248,N14249,
  N14250,N14251,N14252,N14253,N14254,N14255,N14256,N14257,N14258,N14259,N14260,
  N14261,N14262,N14263,N14264,N14265,N14266,N14267,N14268,N14269,N14270,N14271,
  N14272,N14273,N14274,N14275,N14276,N14277,N14278,N14279,N14280,N14281,N14282,N14283,
  N14284,N14285,N14286,N14287,N14288,N14289,N14290,N14291,N14292,N14293,N14294,
  N14295,N14296,N14297,N14298,N14299,N14300,N14301,N14302,N14303,N14304,N14305,N14306,
  N14307,N14308,N14309,N14310,N14311,N14312,N14313,N14314,N14315,N14316,N14317,
  N14318,N14319,N14320,N14321,N14322,N14323,N14324,N14325,N14326,N14327,N14328,N14329,
  N14330,N14331,N14332,N14333,N14334,N14335,N14336,N14337,N14338,N14339,N14340,
  N14341,N14342,N14343,N14344,N14345,N14346,N14347,N14348,N14349,N14350,N14351,
  N14352,N14353,N14354,N14355,N14356,N14357,N14358,N14359,N14360,N14361,N14362,N14363,
  N14364,N14365,N14366,N14367,N14368,N14369,N14370,N14371,N14372,N14373,N14374,
  N14375,N14376,N14377,N14378,N14379,N14380,N14381,N14382,N14383,N14384,N14385,N14386,
  N14387,N14388,N14389,N14390,N14391,N14392,N14393,N14394,N14395,N14396,N14397,
  N14398,N14399,N14400,N14401,N14402,N14403,N14404,N14405,N14406,N14407,N14408,N14409,
  N14410,N14411,N14412,N14413,N14414,N14415,N14416,N14417,N14418,N14419,N14420,
  N14421,N14422,N14423,N14424,N14425,N14426,N14427,N14428,N14429,N14430,N14431,
  N14432,N14433,N14434,N14435,N14436,N14437,N14438,N14439,N14440,N14441,N14442,N14443,
  N14444,N14445,N14446,N14447,N14448,N14449,N14450,N14451,N14452,N14453,N14454,
  N14455,N14456,N14457,N14458,N14459,N14460,N14461,N14462,N14463,N14464,N14465,N14466,
  N14467,N14468,N14469,N14470,N14471,N14472,N14473,N14474,N14475,N14476,N14477,
  N14478,N14479,N14480,N14481,N14482,N14483,N14484,N14485,N14486,N14487,N14488,N14489,
  N14490,N14491,N14492,N14493,N14494,N14495,N14496,N14497,N14498,N14499,N14500,
  N14501,N14502,N14503,N14504,N14505,N14506,N14507,N14508,N14509,N14510,N14511,
  N14512,N14513,N14514,N14515,N14516,N14517,N14518,N14519,N14520,N14521,N14522,N14523,
  N14524,N14525,N14526,N14527,N14528,N14529,N14530,N14531,N14532,N14533,N14534,
  N14535,N14536,N14537,N14538,N14539,N14540,N14541,N14542,N14543,N14544,N14545,N14546,
  N14547,N14548,N14549,N14550,N14551,N14552,N14553,N14554,N14555,N14556,N14557,
  N14558,N14559,N14560,N14561,N14562,N14563,N14564,N14565,N14566,N14567,N14568,N14569,
  N14570,N14571,N14572,N14573,N14574,N14575,N14576,N14577,N14578,N14579,N14580,
  N14581,N14582,N14583,N14584,N14585,N14586,N14587,N14588,N14589,N14590,N14591,
  N14592,N14593,N14594,N14595,N14596,N14597,N14598,N14599,N14600,N14601,N14602,N14603,
  N14604,N14605,N14606,N14607,N14608,N14609,N14610,N14611,N14612,N14613,N14614,
  N14615,N14616,N14617,N14618,N14619,N14620,N14621,N14622,N14623,N14624,N14625,N14626,
  N14627,N14628,N14629,N14630,N14631,N14632,N14633,N14634,N14635,N14636,N14637,
  N14638,N14639,N14640,N14641,N14642,N14643,N14644,N14645,N14646,N14647,N14648,N14649,
  N14650,N14651,N14652,N14653,N14654,N14655,N14656,N14657,N14658,N14659,N14660,
  N14661,N14662,N14663,N14664,N14665,N14666,N14667,N14668,N14669,N14670,N14671,
  N14672,N14673,N14674,N14675,N14676,N14677,N14678,N14679,N14680,N14681,N14682,N14683,
  N14684,N14685,N14686,N14687,N14688,N14689,N14690,N14691,N14692,N14693,N14694,
  N14695,N14696,N14697,N14698,N14699,N14700,N14701,N14702,N14703,N14704,N14705,N14706,
  N14707,N14708,N14709,N14710,N14711,N14712,N14713,N14714,N14715,N14716,N14717,
  N14718,N14719,N14720,N14721,N14722,N14723,N14724,N14725,N14726,N14727,N14728,N14729,
  N14730,N14731,N14732,N14733,N14734,N14735,N14736,N14737,N14738,N14739,N14740,
  N14741,N14742,N14743,N14744,N14745,N14746,N14747,N14748,N14749,N14750,N14751,
  N14752,N14753,N14754,N14755,N14756,N14757,N14758,N14759,N14760,N14761,N14762,N14763,
  N14764,N14765,N14766,N14767,N14768,N14769,N14770,N14771,N14772,N14773,N14774,
  N14775,N14776,N14777,N14778,N14779,N14780,N14781,N14782,N14783,N14784,N14785,N14786,
  N14787,N14788,N14789,N14790,N14791,N14792,N14793,N14794,N14795,N14796,N14797,
  N14798,N14799,N14800,N14801,N14802,N14803,N14804,N14805,N14806,N14807,N14808,N14809,
  N14810,N14811,N14812,N14813,N14814,N14815,N14816,N14817,N14818,N14819,N14820,
  N14821,N14822,N14823,N14824,N14825,N14826,N14827,N14828,N14829,N14830,N14831,
  N14832,N14833,N14834,N14835,N14836,N14837,N14838,N14839,N14840,N14841,N14842,N14843,
  N14844,N14845,N14846,N14847,N14848,N14849,N14850,N14851,N14852,N14853,N14854,
  N14855,N14856,N14857,N14858,N14859,N14860,N14861,N14862,N14863,N14864,N14865,N14866,
  N14867,N14868,N14869,N14870,N14871,N14872,N14873,N14874,N14875,N14876,N14877,
  N14878,N14879,N14880,N14881,N14882,N14883,N14884,N14885,N14886,N14887,N14888,N14889,
  N14890,N14891,N14892,N14893,N14894,N14895,N14896,N14897,N14898,N14899,N14900,
  N14901,N14902,N14903,N14904,N14905,N14906,N14907,N14908,N14909,N14910,N14911,
  N14912,N14913,N14914,N14915,N14916,N14917,N14918,N14919,N14920,N14921,N14922,N14923,
  N14924,N14925,N14926,N14927,N14928,N14929,N14930,N14931,N14932,N14933,N14934,
  N14935,N14936,N14937,N14938,N14939,N14940,N14941,N14942,N14943,N14944,N14945,N14946,
  N14947,N14948,N14949,N14950,N14951,N14952,N14953,N14954,N14955,N14956,N14957,
  N14958,N14959,N14960,N14961,N14962,N14963,N14964,N14965,N14966,N14967,N14968,N14969,
  N14970,N14971,N14972,N14973,N14974,N14975,N14976,N14977,N14978,N14979,N14980,
  N14981,N14982,N14983,N14984,N14985,N14986,N14987,N14988,N14989,N14990,N14991,
  N14992,N14993,N14994,N14995,N14996,N14997,N14998,N14999,N15000,N15001,N15002,N15003,
  N15004,N15005,N15006,N15007,N15008,N15009,N15010,N15011,N15012,N15013,N15014,
  N15015,N15016,N15017,N15018,N15019,N15020,N15021,N15022,N15023,N15024,N15025,N15026,
  N15027,N15028,N15029,N15030,N15031,N15032,N15033,N15034,N15035,N15036,N15037,
  N15038,N15039,N15040,N15041,N15042,N15043,N15044,N15045,N15046,N15047,N15048,N15049,
  N15050,N15051,N15052,N15053,N15054,N15055,N15056,N15057,N15058,N15059,N15060,
  N15061,N15062,N15063,N15064,N15065,N15066,N15067,N15068,N15069,N15070,N15071,
  N15072,N15073,N15074,N15075,N15076,N15077,N15078,N15079,N15080,N15081,N15082,N15083,
  N15084,N15085,N15086,N15087,N15088,N15089,N15090,N15091,N15092,N15093,N15094,
  N15095,N15096,N15097,N15098,N15099,N15100,N15101,N15102,N15103,N15104,N15105,N15106,
  N15107,N15108,N15109,N15110,N15111,N15112,N15113,N15114,N15115,N15116,N15117,
  N15118,N15119,N15120,N15121,N15122,N15123,N15124,N15125,N15126,N15127,N15128,N15129,
  N15130,N15131,N15132,N15133,N15134,N15135,N15136,N15137,N15138,N15139,N15140,
  N15141,N15142,N15143,N15144,N15145,N15146,N15147,N15148,N15149,N15150,N15151,
  N15152,N15153,N15154,N15155,N15156,N15157,N15158,N15159,N15160,N15161,N15162,N15163,
  N15164,N15165,N15166,N15167,N15168,N15169,N15170,N15171,N15172,N15173,N15174,
  N15175,N15176,N15177,N15178,N15179,N15180,N15181,N15182,N15183,N15184,N15185,N15186,
  N15187,N15188,N15189,N15190,N15191,N15192,N15193,N15194,N15195,N15196,N15197,
  N15198,N15199,N15200,N15201,N15202,N15203,N15204,N15205,N15206,N15207,N15208,N15209,
  N15210,N15211,N15212,N15213,N15214,N15215,N15216,N15217,N15218,N15219,N15220,
  N15221,N15222,N15223,N15224,N15225,N15226,N15227,N15228,N15229,N15230,N15231,
  N15232,N15233,N15234,N15235,N15236,N15237,N15238,N15239,N15240,N15241,N15242,N15243,
  N15244,N15245,N15246,N15247,N15248,N15249,N15250,N15251,N15252,N15253,N15254,
  N15255,N15256,N15257,N15258,N15259,N15260,N15261,N15262,N15263,N15264,N15265,N15266,
  N15267,N15268,N15269,N15270,N15271,N15272,N15273,N15274,N15275,N15276,N15277,
  N15278,N15279,N15280,N15281,N15282,N15283,N15284,N15285,N15286,N15287,N15288,N15289,
  N15290,N15291,N15292,N15293,N15294,N15295,N15296,N15297,N15298,N15299,N15300,
  N15301,N15302,N15303,N15304,N15305,N15306,N15307,N15308,N15309,N15310,N15311,
  N15312,N15313,N15314,N15315,N15316,N15317,N15318,N15319,N15320,N15321,N15322,N15323,
  N15324,N15325,N15326,N15327,N15328,N15329,N15330,N15331,N15332,N15333,N15334,
  N15335,N15336,N15337,N15338,N15339,N15340,N15341,N15342,N15343,N15344,N15345,N15346,
  N15347,N15348,N15349,N15350,N15351,N15352,N15353,N15354,N15355,N15356,N15357,
  N15358,N15359,N15360,N15361,N15362,N15363,N15364,N15365,N15366,N15367,N15368,N15369,
  N15370,N15371,N15372,N15373,N15374,N15375,N15376,N15377,N15378,N15379,N15380,
  N15381,N15382,N15383,N15384,N15385,N15386,N15387,N15388,N15389,N15390,N15391,
  N15392,N15393,N15394,N15395,N15396,N15397,N15398,N15399,N15400,N15401,N15402,N15403,
  N15404,N15405,N15406,N15407,N15408,N15409,N15410,N15411,N15412,N15413,N15414,
  N15415,N15416,N15417,N15418,N15419,N15420,N15421,N15422,N15423,N15424,N15425,N15426,
  N15427,N15428,N15429,N15430,N15431,N15432,N15433,N15434,N15435,N15436,N15437,
  N15438,N15439,N15440,N15441,N15442,N15443,N15444,N15445,N15446,N15447,N15448,N15449,
  N15450,N15451,N15452,N15453,N15454,N15455,N15456,N15457,N15458,N15459,N15460,
  N15461,N15462,N15463,N15464,N15465,N15466,N15467,N15468,N15469,N15470,N15471,
  N15472,N15473,N15474,N15475,N15476,N15477,N15478,N15479,N15480,N15481,N15482,N15483,
  N15484,N15485,N15486,N15487,N15488,N15489,N15490,N15491,N15492,N15493,N15494,
  N15495,N15496,N15497,N15498,N15499,N15500,N15501,N15502,N15503,N15504,N15505,N15506,
  N15507,N15508,N15509,N15510,N15511,N15512,N15513,N15514,N15515,N15516,N15517,
  N15518,N15519,N15520,N15521,N15522,N15523,N15524,N15525,N15526,N15527,N15528,N15529,
  N15530,N15531,N15532,N15533,N15534,N15535,N15536,N15537,N15538,N15539,N15540,
  N15541,N15542,N15543,N15544,N15545,N15546,N15547,N15548,N15549,N15550,N15551,
  N15552,N15553,N15554,N15555,N15556,N15557,N15558,N15559,N15560,N15561,N15562,N15563,
  N15564,N15565,N15566,N15567,N15568,N15569,N15570,N15571,N15572,N15573,N15574,
  N15575,N15576,N15577,N15578,N15579,N15580,N15581,N15582,N15583,N15584,N15585,N15586,
  N15587,N15588,N15589,N15590,N15591,N15592,N15593,N15594,N15595,N15596,N15597,
  N15598,N15599,N15600,N15601,N15602,N15603,N15604,N15605,N15606,N15607,N15608,N15609,
  N15610,N15611,N15612,N15613,N15614,N15615,N15616,N15617,N15618,N15619,N15620,
  N15621,N15622,N15623,N15624,N15625,N15626,N15627,N15628,N15629,N15630,N15631,
  N15632,N15633,N15634,N15635,N15636,N15637,N15638,N15639,N15640,N15641,N15642,N15643,
  N15644,N15645,N15646,N15647,N15648,N15649,N15650,N15651,N15652,N15653,N15654,
  N15655,N15656,N15657,N15658,N15659,N15660,N15661,N15662,N15663,N15664,N15665,N15666,
  N15667,N15668,N15669,N15670,N15671,N15672,N15673,N15674,N15675,N15676,N15677,
  N15678,N15679,N15680,N15681,N15682,N15683,N15684,N15685,N15686,N15687,N15688,N15689,
  N15690,N15691,N15692,N15693,N15694,N15695,N15696,N15697,N15698,N15699,N15700,
  N15701,N15702,N15703,N15704,N15705,N15706,N15707,N15708,N15709,N15710,N15711,
  N15712,N15713,N15714,N15715,N15716,N15717,N15718,N15719,N15720,N15721,N15722,N15723,
  N15724,N15725,N15726,N15727,N15728,N15729,N15730,N15731,N15732,N15733,N15734,
  N15735,N15736,N15737,N15738,N15739,N15740,N15741,N15742,N15743,N15744,N15745,N15746,
  N15747,N15748,N15749,N15750,N15751,N15752,N15753,N15754,N15755,N15756,N15757,
  N15758,N15759,N15760,N15761,N15762,N15763,N15764,N15765,N15766,N15767,N15768,N15769,
  N15770,N15771,N15772,N15773,N15774,N15775,N15776,N15777,N15778,N15779,N15780,
  N15781,N15782,N15783,N15784,N15785,N15786,N15787,N15788,N15789,N15790,N15791,
  N15792,N15793,N15794,N15795,N15796,N15797,N15798,N15799,N15800,N15801,N15802,N15803,
  N15804,N15805,N15806,N15807,N15808,N15809,N15810,N15811,N15812,N15813,N15814,
  N15815,N15816,N15817,N15818,N15819,N15820,N15821,N15822,N15823,N15824,N15825,N15826,
  N15827,N15828,N15829,N15830,N15831,N15832,N15833,N15834,N15835,N15836,N15837,
  N15838,N15839,N15840,N15841,N15842,N15843,N15844,N15845,N15846,N15847,N15848,N15849,
  N15850,N15851,N15852,N15853,N15854,N15855,N15856,N15857,N15858,N15859,N15860,
  N15861,N15862,N15863,N15864,N15865,N15866,N15867,N15868,N15869,N15870,N15871,
  N15872,N15873,N15874,N15875,N15876,N15877,N15878,N15879,N15880,N15881,N15882,N15883,
  N15884,N15885,N15886,N15887,N15888,N15889,N15890,N15891,N15892,N15893,N15894,
  N15895,N15896,N15897,N15898,N15899,N15900,N15901,N15902,N15903,N15904,N15905,N15906,
  N15907,N15908,N15909,N15910,N15911,N15912,N15913,N15914,N15915,N15916,N15917,
  N15918,N15919,N15920,N15921,N15922,N15923,N15924,N15925,N15926,N15927,N15928,N15929,
  N15930,N15931,N15932,N15933,N15934,N15935,N15936,N15937,N15938,N15939,N15940,
  N15941,N15942,N15943,N15944,N15945,N15946,N15947,N15948,N15949,N15950,N15951,
  N15952,N15953,N15954,N15955,N15956,N15957,N15958,N15959,N15960,N15961,N15962,N15963,
  N15964,N15965,N15966,N15967,N15968,N15969,N15970,N15971,N15972,N15973,N15974,
  N15975,N15976,N15977,N15978,N15979,N15980,N15981,N15982,N15983,N15984,N15985,N15986,
  N15987,N15988,N15989,N15990,N15991,N15992,N15993,N15994,N15995,N15996,N15997,
  N15998,N15999,N16000,N16001,N16002,N16003,N16004,N16005,N16006,N16007,N16008,N16009,
  N16010,N16011,N16012,N16013,N16014,N16015,N16016,N16017,N16018,N16019,N16020,
  N16021,N16022,N16023,N16024,N16025,N16026,N16027,N16028,N16029,N16030,N16031,
  N16032,N16033,N16034,N16035,N16036,N16037,N16038,N16039,N16040,N16041,N16042,N16043,
  N16044,N16045,N16046,N16047,N16048,N16049,N16050,N16051,N16052,N16053,N16054,
  N16055,N16056,N16057,N16058,N16059,N16060,N16061,N16062,N16063,N16064,N16065,N16066,
  N16067,N16068,N16069,N16070,N16071,N16072,N16073,N16074,N16075,N16076,N16077,
  N16078,N16079,N16080,N16081,N16082,N16083,N16084,N16085,N16086,N16087,N16088,N16089,
  N16090,N16091,N16092,N16093,N16094,N16095,N16096,N16097,N16098,N16099,N16100,
  N16101,N16102,N16103,N16104,N16105,N16106,N16107,N16108,N16109,N16110,N16111,
  N16112,N16113,N16114,N16115,N16116,N16117,N16118,N16119,N16120,N16121,N16122,N16123,
  N16124,N16125,N16126,N16127;
  wire [16383:0] data_masked;
  assign data_masked[127] = data_i[127] & sel_one_hot_i[0];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[0];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[0];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[0];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[0];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[0];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[0];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[0];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[0];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[0];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[0];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[0];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[0];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[0];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[0];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[0];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[0];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[0];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[0];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[0];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[0];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[0];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[0];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[0];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[0];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[0];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[0];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[0];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[0];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[0];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[0];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[0];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[0];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[0];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[0];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[0];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[0];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[0];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[0];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[0];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[0];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[0];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[0];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[0];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[0];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[0];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[0];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[0];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[0];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[0];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[0];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[0];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[0];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[0];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[0];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[0];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[0];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[0];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[0];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[0];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[0];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[0];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[1];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[1];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[1];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[1];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[1];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[1];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[1];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[1];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[1];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[1];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[1];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[1];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[1];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[1];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[1];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[1];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[1];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[1];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[1];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[1];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[1];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[1];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[1];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[1];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[1];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[1];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[1];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[1];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[1];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[1];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[1];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[1];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[1];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[1];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[1];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[1];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[1];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[1];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[1];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[1];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[1];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[1];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[1];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[1];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[1];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[1];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[1];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[1];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[1];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[1];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[1];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[1];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[1];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[1];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[1];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[1];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[1];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[1];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[1];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[1];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[1];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[1];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[1];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[1];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[1];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[1];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[1];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[1];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[1];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[1];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[1];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[1];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[1];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[1];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[1];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[1];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[1];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[1];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[1];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[1];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[1];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[1];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[1];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[1];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[1];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[1];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[1];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[1];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[1];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[1];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[1];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[1];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[1];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[1];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[1];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[1];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[1];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[1];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[1];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[1];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[1];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[1];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[1];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[1];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[1];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[1];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[1];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[1];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[1];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[1];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[1];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[1];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[1];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[1];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[1];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[1];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[1];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[1];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[1];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[1];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[1];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[1];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[1];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[1];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[1];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[1];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[1];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[2];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[2];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[2];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[2];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[2];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[2];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[2];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[2];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[2];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[2];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[2];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[2];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[2];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[2];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[2];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[2];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[2];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[2];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[2];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[2];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[2];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[2];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[2];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[2];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[2];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[2];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[2];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[2];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[2];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[2];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[2];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[2];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[2];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[2];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[2];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[2];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[2];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[2];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[2];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[2];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[2];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[2];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[2];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[2];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[2];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[2];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[2];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[2];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[2];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[2];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[2];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[2];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[2];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[2];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[2];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[2];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[2];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[2];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[2];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[2];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[2];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[2];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[2];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[2];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[2];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[2];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[2];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[2];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[2];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[2];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[2];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[2];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[2];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[2];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[2];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[2];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[2];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[2];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[2];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[2];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[2];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[2];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[2];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[2];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[2];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[2];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[2];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[2];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[2];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[2];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[2];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[2];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[2];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[2];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[2];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[2];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[2];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[2];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[2];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[2];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[2];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[2];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[2];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[2];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[2];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[2];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[2];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[2];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[2];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[2];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[2];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[2];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[2];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[2];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[2];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[2];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[2];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[2];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[2];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[2];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[2];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[2];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[2];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[2];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[2];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[2];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[2];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[2];
  assign data_masked[511] = data_i[511] & sel_one_hot_i[3];
  assign data_masked[510] = data_i[510] & sel_one_hot_i[3];
  assign data_masked[509] = data_i[509] & sel_one_hot_i[3];
  assign data_masked[508] = data_i[508] & sel_one_hot_i[3];
  assign data_masked[507] = data_i[507] & sel_one_hot_i[3];
  assign data_masked[506] = data_i[506] & sel_one_hot_i[3];
  assign data_masked[505] = data_i[505] & sel_one_hot_i[3];
  assign data_masked[504] = data_i[504] & sel_one_hot_i[3];
  assign data_masked[503] = data_i[503] & sel_one_hot_i[3];
  assign data_masked[502] = data_i[502] & sel_one_hot_i[3];
  assign data_masked[501] = data_i[501] & sel_one_hot_i[3];
  assign data_masked[500] = data_i[500] & sel_one_hot_i[3];
  assign data_masked[499] = data_i[499] & sel_one_hot_i[3];
  assign data_masked[498] = data_i[498] & sel_one_hot_i[3];
  assign data_masked[497] = data_i[497] & sel_one_hot_i[3];
  assign data_masked[496] = data_i[496] & sel_one_hot_i[3];
  assign data_masked[495] = data_i[495] & sel_one_hot_i[3];
  assign data_masked[494] = data_i[494] & sel_one_hot_i[3];
  assign data_masked[493] = data_i[493] & sel_one_hot_i[3];
  assign data_masked[492] = data_i[492] & sel_one_hot_i[3];
  assign data_masked[491] = data_i[491] & sel_one_hot_i[3];
  assign data_masked[490] = data_i[490] & sel_one_hot_i[3];
  assign data_masked[489] = data_i[489] & sel_one_hot_i[3];
  assign data_masked[488] = data_i[488] & sel_one_hot_i[3];
  assign data_masked[487] = data_i[487] & sel_one_hot_i[3];
  assign data_masked[486] = data_i[486] & sel_one_hot_i[3];
  assign data_masked[485] = data_i[485] & sel_one_hot_i[3];
  assign data_masked[484] = data_i[484] & sel_one_hot_i[3];
  assign data_masked[483] = data_i[483] & sel_one_hot_i[3];
  assign data_masked[482] = data_i[482] & sel_one_hot_i[3];
  assign data_masked[481] = data_i[481] & sel_one_hot_i[3];
  assign data_masked[480] = data_i[480] & sel_one_hot_i[3];
  assign data_masked[479] = data_i[479] & sel_one_hot_i[3];
  assign data_masked[478] = data_i[478] & sel_one_hot_i[3];
  assign data_masked[477] = data_i[477] & sel_one_hot_i[3];
  assign data_masked[476] = data_i[476] & sel_one_hot_i[3];
  assign data_masked[475] = data_i[475] & sel_one_hot_i[3];
  assign data_masked[474] = data_i[474] & sel_one_hot_i[3];
  assign data_masked[473] = data_i[473] & sel_one_hot_i[3];
  assign data_masked[472] = data_i[472] & sel_one_hot_i[3];
  assign data_masked[471] = data_i[471] & sel_one_hot_i[3];
  assign data_masked[470] = data_i[470] & sel_one_hot_i[3];
  assign data_masked[469] = data_i[469] & sel_one_hot_i[3];
  assign data_masked[468] = data_i[468] & sel_one_hot_i[3];
  assign data_masked[467] = data_i[467] & sel_one_hot_i[3];
  assign data_masked[466] = data_i[466] & sel_one_hot_i[3];
  assign data_masked[465] = data_i[465] & sel_one_hot_i[3];
  assign data_masked[464] = data_i[464] & sel_one_hot_i[3];
  assign data_masked[463] = data_i[463] & sel_one_hot_i[3];
  assign data_masked[462] = data_i[462] & sel_one_hot_i[3];
  assign data_masked[461] = data_i[461] & sel_one_hot_i[3];
  assign data_masked[460] = data_i[460] & sel_one_hot_i[3];
  assign data_masked[459] = data_i[459] & sel_one_hot_i[3];
  assign data_masked[458] = data_i[458] & sel_one_hot_i[3];
  assign data_masked[457] = data_i[457] & sel_one_hot_i[3];
  assign data_masked[456] = data_i[456] & sel_one_hot_i[3];
  assign data_masked[455] = data_i[455] & sel_one_hot_i[3];
  assign data_masked[454] = data_i[454] & sel_one_hot_i[3];
  assign data_masked[453] = data_i[453] & sel_one_hot_i[3];
  assign data_masked[452] = data_i[452] & sel_one_hot_i[3];
  assign data_masked[451] = data_i[451] & sel_one_hot_i[3];
  assign data_masked[450] = data_i[450] & sel_one_hot_i[3];
  assign data_masked[449] = data_i[449] & sel_one_hot_i[3];
  assign data_masked[448] = data_i[448] & sel_one_hot_i[3];
  assign data_masked[447] = data_i[447] & sel_one_hot_i[3];
  assign data_masked[446] = data_i[446] & sel_one_hot_i[3];
  assign data_masked[445] = data_i[445] & sel_one_hot_i[3];
  assign data_masked[444] = data_i[444] & sel_one_hot_i[3];
  assign data_masked[443] = data_i[443] & sel_one_hot_i[3];
  assign data_masked[442] = data_i[442] & sel_one_hot_i[3];
  assign data_masked[441] = data_i[441] & sel_one_hot_i[3];
  assign data_masked[440] = data_i[440] & sel_one_hot_i[3];
  assign data_masked[439] = data_i[439] & sel_one_hot_i[3];
  assign data_masked[438] = data_i[438] & sel_one_hot_i[3];
  assign data_masked[437] = data_i[437] & sel_one_hot_i[3];
  assign data_masked[436] = data_i[436] & sel_one_hot_i[3];
  assign data_masked[435] = data_i[435] & sel_one_hot_i[3];
  assign data_masked[434] = data_i[434] & sel_one_hot_i[3];
  assign data_masked[433] = data_i[433] & sel_one_hot_i[3];
  assign data_masked[432] = data_i[432] & sel_one_hot_i[3];
  assign data_masked[431] = data_i[431] & sel_one_hot_i[3];
  assign data_masked[430] = data_i[430] & sel_one_hot_i[3];
  assign data_masked[429] = data_i[429] & sel_one_hot_i[3];
  assign data_masked[428] = data_i[428] & sel_one_hot_i[3];
  assign data_masked[427] = data_i[427] & sel_one_hot_i[3];
  assign data_masked[426] = data_i[426] & sel_one_hot_i[3];
  assign data_masked[425] = data_i[425] & sel_one_hot_i[3];
  assign data_masked[424] = data_i[424] & sel_one_hot_i[3];
  assign data_masked[423] = data_i[423] & sel_one_hot_i[3];
  assign data_masked[422] = data_i[422] & sel_one_hot_i[3];
  assign data_masked[421] = data_i[421] & sel_one_hot_i[3];
  assign data_masked[420] = data_i[420] & sel_one_hot_i[3];
  assign data_masked[419] = data_i[419] & sel_one_hot_i[3];
  assign data_masked[418] = data_i[418] & sel_one_hot_i[3];
  assign data_masked[417] = data_i[417] & sel_one_hot_i[3];
  assign data_masked[416] = data_i[416] & sel_one_hot_i[3];
  assign data_masked[415] = data_i[415] & sel_one_hot_i[3];
  assign data_masked[414] = data_i[414] & sel_one_hot_i[3];
  assign data_masked[413] = data_i[413] & sel_one_hot_i[3];
  assign data_masked[412] = data_i[412] & sel_one_hot_i[3];
  assign data_masked[411] = data_i[411] & sel_one_hot_i[3];
  assign data_masked[410] = data_i[410] & sel_one_hot_i[3];
  assign data_masked[409] = data_i[409] & sel_one_hot_i[3];
  assign data_masked[408] = data_i[408] & sel_one_hot_i[3];
  assign data_masked[407] = data_i[407] & sel_one_hot_i[3];
  assign data_masked[406] = data_i[406] & sel_one_hot_i[3];
  assign data_masked[405] = data_i[405] & sel_one_hot_i[3];
  assign data_masked[404] = data_i[404] & sel_one_hot_i[3];
  assign data_masked[403] = data_i[403] & sel_one_hot_i[3];
  assign data_masked[402] = data_i[402] & sel_one_hot_i[3];
  assign data_masked[401] = data_i[401] & sel_one_hot_i[3];
  assign data_masked[400] = data_i[400] & sel_one_hot_i[3];
  assign data_masked[399] = data_i[399] & sel_one_hot_i[3];
  assign data_masked[398] = data_i[398] & sel_one_hot_i[3];
  assign data_masked[397] = data_i[397] & sel_one_hot_i[3];
  assign data_masked[396] = data_i[396] & sel_one_hot_i[3];
  assign data_masked[395] = data_i[395] & sel_one_hot_i[3];
  assign data_masked[394] = data_i[394] & sel_one_hot_i[3];
  assign data_masked[393] = data_i[393] & sel_one_hot_i[3];
  assign data_masked[392] = data_i[392] & sel_one_hot_i[3];
  assign data_masked[391] = data_i[391] & sel_one_hot_i[3];
  assign data_masked[390] = data_i[390] & sel_one_hot_i[3];
  assign data_masked[389] = data_i[389] & sel_one_hot_i[3];
  assign data_masked[388] = data_i[388] & sel_one_hot_i[3];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[3];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[3];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[3];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[3];
  assign data_masked[639] = data_i[639] & sel_one_hot_i[4];
  assign data_masked[638] = data_i[638] & sel_one_hot_i[4];
  assign data_masked[637] = data_i[637] & sel_one_hot_i[4];
  assign data_masked[636] = data_i[636] & sel_one_hot_i[4];
  assign data_masked[635] = data_i[635] & sel_one_hot_i[4];
  assign data_masked[634] = data_i[634] & sel_one_hot_i[4];
  assign data_masked[633] = data_i[633] & sel_one_hot_i[4];
  assign data_masked[632] = data_i[632] & sel_one_hot_i[4];
  assign data_masked[631] = data_i[631] & sel_one_hot_i[4];
  assign data_masked[630] = data_i[630] & sel_one_hot_i[4];
  assign data_masked[629] = data_i[629] & sel_one_hot_i[4];
  assign data_masked[628] = data_i[628] & sel_one_hot_i[4];
  assign data_masked[627] = data_i[627] & sel_one_hot_i[4];
  assign data_masked[626] = data_i[626] & sel_one_hot_i[4];
  assign data_masked[625] = data_i[625] & sel_one_hot_i[4];
  assign data_masked[624] = data_i[624] & sel_one_hot_i[4];
  assign data_masked[623] = data_i[623] & sel_one_hot_i[4];
  assign data_masked[622] = data_i[622] & sel_one_hot_i[4];
  assign data_masked[621] = data_i[621] & sel_one_hot_i[4];
  assign data_masked[620] = data_i[620] & sel_one_hot_i[4];
  assign data_masked[619] = data_i[619] & sel_one_hot_i[4];
  assign data_masked[618] = data_i[618] & sel_one_hot_i[4];
  assign data_masked[617] = data_i[617] & sel_one_hot_i[4];
  assign data_masked[616] = data_i[616] & sel_one_hot_i[4];
  assign data_masked[615] = data_i[615] & sel_one_hot_i[4];
  assign data_masked[614] = data_i[614] & sel_one_hot_i[4];
  assign data_masked[613] = data_i[613] & sel_one_hot_i[4];
  assign data_masked[612] = data_i[612] & sel_one_hot_i[4];
  assign data_masked[611] = data_i[611] & sel_one_hot_i[4];
  assign data_masked[610] = data_i[610] & sel_one_hot_i[4];
  assign data_masked[609] = data_i[609] & sel_one_hot_i[4];
  assign data_masked[608] = data_i[608] & sel_one_hot_i[4];
  assign data_masked[607] = data_i[607] & sel_one_hot_i[4];
  assign data_masked[606] = data_i[606] & sel_one_hot_i[4];
  assign data_masked[605] = data_i[605] & sel_one_hot_i[4];
  assign data_masked[604] = data_i[604] & sel_one_hot_i[4];
  assign data_masked[603] = data_i[603] & sel_one_hot_i[4];
  assign data_masked[602] = data_i[602] & sel_one_hot_i[4];
  assign data_masked[601] = data_i[601] & sel_one_hot_i[4];
  assign data_masked[600] = data_i[600] & sel_one_hot_i[4];
  assign data_masked[599] = data_i[599] & sel_one_hot_i[4];
  assign data_masked[598] = data_i[598] & sel_one_hot_i[4];
  assign data_masked[597] = data_i[597] & sel_one_hot_i[4];
  assign data_masked[596] = data_i[596] & sel_one_hot_i[4];
  assign data_masked[595] = data_i[595] & sel_one_hot_i[4];
  assign data_masked[594] = data_i[594] & sel_one_hot_i[4];
  assign data_masked[593] = data_i[593] & sel_one_hot_i[4];
  assign data_masked[592] = data_i[592] & sel_one_hot_i[4];
  assign data_masked[591] = data_i[591] & sel_one_hot_i[4];
  assign data_masked[590] = data_i[590] & sel_one_hot_i[4];
  assign data_masked[589] = data_i[589] & sel_one_hot_i[4];
  assign data_masked[588] = data_i[588] & sel_one_hot_i[4];
  assign data_masked[587] = data_i[587] & sel_one_hot_i[4];
  assign data_masked[586] = data_i[586] & sel_one_hot_i[4];
  assign data_masked[585] = data_i[585] & sel_one_hot_i[4];
  assign data_masked[584] = data_i[584] & sel_one_hot_i[4];
  assign data_masked[583] = data_i[583] & sel_one_hot_i[4];
  assign data_masked[582] = data_i[582] & sel_one_hot_i[4];
  assign data_masked[581] = data_i[581] & sel_one_hot_i[4];
  assign data_masked[580] = data_i[580] & sel_one_hot_i[4];
  assign data_masked[579] = data_i[579] & sel_one_hot_i[4];
  assign data_masked[578] = data_i[578] & sel_one_hot_i[4];
  assign data_masked[577] = data_i[577] & sel_one_hot_i[4];
  assign data_masked[576] = data_i[576] & sel_one_hot_i[4];
  assign data_masked[575] = data_i[575] & sel_one_hot_i[4];
  assign data_masked[574] = data_i[574] & sel_one_hot_i[4];
  assign data_masked[573] = data_i[573] & sel_one_hot_i[4];
  assign data_masked[572] = data_i[572] & sel_one_hot_i[4];
  assign data_masked[571] = data_i[571] & sel_one_hot_i[4];
  assign data_masked[570] = data_i[570] & sel_one_hot_i[4];
  assign data_masked[569] = data_i[569] & sel_one_hot_i[4];
  assign data_masked[568] = data_i[568] & sel_one_hot_i[4];
  assign data_masked[567] = data_i[567] & sel_one_hot_i[4];
  assign data_masked[566] = data_i[566] & sel_one_hot_i[4];
  assign data_masked[565] = data_i[565] & sel_one_hot_i[4];
  assign data_masked[564] = data_i[564] & sel_one_hot_i[4];
  assign data_masked[563] = data_i[563] & sel_one_hot_i[4];
  assign data_masked[562] = data_i[562] & sel_one_hot_i[4];
  assign data_masked[561] = data_i[561] & sel_one_hot_i[4];
  assign data_masked[560] = data_i[560] & sel_one_hot_i[4];
  assign data_masked[559] = data_i[559] & sel_one_hot_i[4];
  assign data_masked[558] = data_i[558] & sel_one_hot_i[4];
  assign data_masked[557] = data_i[557] & sel_one_hot_i[4];
  assign data_masked[556] = data_i[556] & sel_one_hot_i[4];
  assign data_masked[555] = data_i[555] & sel_one_hot_i[4];
  assign data_masked[554] = data_i[554] & sel_one_hot_i[4];
  assign data_masked[553] = data_i[553] & sel_one_hot_i[4];
  assign data_masked[552] = data_i[552] & sel_one_hot_i[4];
  assign data_masked[551] = data_i[551] & sel_one_hot_i[4];
  assign data_masked[550] = data_i[550] & sel_one_hot_i[4];
  assign data_masked[549] = data_i[549] & sel_one_hot_i[4];
  assign data_masked[548] = data_i[548] & sel_one_hot_i[4];
  assign data_masked[547] = data_i[547] & sel_one_hot_i[4];
  assign data_masked[546] = data_i[546] & sel_one_hot_i[4];
  assign data_masked[545] = data_i[545] & sel_one_hot_i[4];
  assign data_masked[544] = data_i[544] & sel_one_hot_i[4];
  assign data_masked[543] = data_i[543] & sel_one_hot_i[4];
  assign data_masked[542] = data_i[542] & sel_one_hot_i[4];
  assign data_masked[541] = data_i[541] & sel_one_hot_i[4];
  assign data_masked[540] = data_i[540] & sel_one_hot_i[4];
  assign data_masked[539] = data_i[539] & sel_one_hot_i[4];
  assign data_masked[538] = data_i[538] & sel_one_hot_i[4];
  assign data_masked[537] = data_i[537] & sel_one_hot_i[4];
  assign data_masked[536] = data_i[536] & sel_one_hot_i[4];
  assign data_masked[535] = data_i[535] & sel_one_hot_i[4];
  assign data_masked[534] = data_i[534] & sel_one_hot_i[4];
  assign data_masked[533] = data_i[533] & sel_one_hot_i[4];
  assign data_masked[532] = data_i[532] & sel_one_hot_i[4];
  assign data_masked[531] = data_i[531] & sel_one_hot_i[4];
  assign data_masked[530] = data_i[530] & sel_one_hot_i[4];
  assign data_masked[529] = data_i[529] & sel_one_hot_i[4];
  assign data_masked[528] = data_i[528] & sel_one_hot_i[4];
  assign data_masked[527] = data_i[527] & sel_one_hot_i[4];
  assign data_masked[526] = data_i[526] & sel_one_hot_i[4];
  assign data_masked[525] = data_i[525] & sel_one_hot_i[4];
  assign data_masked[524] = data_i[524] & sel_one_hot_i[4];
  assign data_masked[523] = data_i[523] & sel_one_hot_i[4];
  assign data_masked[522] = data_i[522] & sel_one_hot_i[4];
  assign data_masked[521] = data_i[521] & sel_one_hot_i[4];
  assign data_masked[520] = data_i[520] & sel_one_hot_i[4];
  assign data_masked[519] = data_i[519] & sel_one_hot_i[4];
  assign data_masked[518] = data_i[518] & sel_one_hot_i[4];
  assign data_masked[517] = data_i[517] & sel_one_hot_i[4];
  assign data_masked[516] = data_i[516] & sel_one_hot_i[4];
  assign data_masked[515] = data_i[515] & sel_one_hot_i[4];
  assign data_masked[514] = data_i[514] & sel_one_hot_i[4];
  assign data_masked[513] = data_i[513] & sel_one_hot_i[4];
  assign data_masked[512] = data_i[512] & sel_one_hot_i[4];
  assign data_masked[767] = data_i[767] & sel_one_hot_i[5];
  assign data_masked[766] = data_i[766] & sel_one_hot_i[5];
  assign data_masked[765] = data_i[765] & sel_one_hot_i[5];
  assign data_masked[764] = data_i[764] & sel_one_hot_i[5];
  assign data_masked[763] = data_i[763] & sel_one_hot_i[5];
  assign data_masked[762] = data_i[762] & sel_one_hot_i[5];
  assign data_masked[761] = data_i[761] & sel_one_hot_i[5];
  assign data_masked[760] = data_i[760] & sel_one_hot_i[5];
  assign data_masked[759] = data_i[759] & sel_one_hot_i[5];
  assign data_masked[758] = data_i[758] & sel_one_hot_i[5];
  assign data_masked[757] = data_i[757] & sel_one_hot_i[5];
  assign data_masked[756] = data_i[756] & sel_one_hot_i[5];
  assign data_masked[755] = data_i[755] & sel_one_hot_i[5];
  assign data_masked[754] = data_i[754] & sel_one_hot_i[5];
  assign data_masked[753] = data_i[753] & sel_one_hot_i[5];
  assign data_masked[752] = data_i[752] & sel_one_hot_i[5];
  assign data_masked[751] = data_i[751] & sel_one_hot_i[5];
  assign data_masked[750] = data_i[750] & sel_one_hot_i[5];
  assign data_masked[749] = data_i[749] & sel_one_hot_i[5];
  assign data_masked[748] = data_i[748] & sel_one_hot_i[5];
  assign data_masked[747] = data_i[747] & sel_one_hot_i[5];
  assign data_masked[746] = data_i[746] & sel_one_hot_i[5];
  assign data_masked[745] = data_i[745] & sel_one_hot_i[5];
  assign data_masked[744] = data_i[744] & sel_one_hot_i[5];
  assign data_masked[743] = data_i[743] & sel_one_hot_i[5];
  assign data_masked[742] = data_i[742] & sel_one_hot_i[5];
  assign data_masked[741] = data_i[741] & sel_one_hot_i[5];
  assign data_masked[740] = data_i[740] & sel_one_hot_i[5];
  assign data_masked[739] = data_i[739] & sel_one_hot_i[5];
  assign data_masked[738] = data_i[738] & sel_one_hot_i[5];
  assign data_masked[737] = data_i[737] & sel_one_hot_i[5];
  assign data_masked[736] = data_i[736] & sel_one_hot_i[5];
  assign data_masked[735] = data_i[735] & sel_one_hot_i[5];
  assign data_masked[734] = data_i[734] & sel_one_hot_i[5];
  assign data_masked[733] = data_i[733] & sel_one_hot_i[5];
  assign data_masked[732] = data_i[732] & sel_one_hot_i[5];
  assign data_masked[731] = data_i[731] & sel_one_hot_i[5];
  assign data_masked[730] = data_i[730] & sel_one_hot_i[5];
  assign data_masked[729] = data_i[729] & sel_one_hot_i[5];
  assign data_masked[728] = data_i[728] & sel_one_hot_i[5];
  assign data_masked[727] = data_i[727] & sel_one_hot_i[5];
  assign data_masked[726] = data_i[726] & sel_one_hot_i[5];
  assign data_masked[725] = data_i[725] & sel_one_hot_i[5];
  assign data_masked[724] = data_i[724] & sel_one_hot_i[5];
  assign data_masked[723] = data_i[723] & sel_one_hot_i[5];
  assign data_masked[722] = data_i[722] & sel_one_hot_i[5];
  assign data_masked[721] = data_i[721] & sel_one_hot_i[5];
  assign data_masked[720] = data_i[720] & sel_one_hot_i[5];
  assign data_masked[719] = data_i[719] & sel_one_hot_i[5];
  assign data_masked[718] = data_i[718] & sel_one_hot_i[5];
  assign data_masked[717] = data_i[717] & sel_one_hot_i[5];
  assign data_masked[716] = data_i[716] & sel_one_hot_i[5];
  assign data_masked[715] = data_i[715] & sel_one_hot_i[5];
  assign data_masked[714] = data_i[714] & sel_one_hot_i[5];
  assign data_masked[713] = data_i[713] & sel_one_hot_i[5];
  assign data_masked[712] = data_i[712] & sel_one_hot_i[5];
  assign data_masked[711] = data_i[711] & sel_one_hot_i[5];
  assign data_masked[710] = data_i[710] & sel_one_hot_i[5];
  assign data_masked[709] = data_i[709] & sel_one_hot_i[5];
  assign data_masked[708] = data_i[708] & sel_one_hot_i[5];
  assign data_masked[707] = data_i[707] & sel_one_hot_i[5];
  assign data_masked[706] = data_i[706] & sel_one_hot_i[5];
  assign data_masked[705] = data_i[705] & sel_one_hot_i[5];
  assign data_masked[704] = data_i[704] & sel_one_hot_i[5];
  assign data_masked[703] = data_i[703] & sel_one_hot_i[5];
  assign data_masked[702] = data_i[702] & sel_one_hot_i[5];
  assign data_masked[701] = data_i[701] & sel_one_hot_i[5];
  assign data_masked[700] = data_i[700] & sel_one_hot_i[5];
  assign data_masked[699] = data_i[699] & sel_one_hot_i[5];
  assign data_masked[698] = data_i[698] & sel_one_hot_i[5];
  assign data_masked[697] = data_i[697] & sel_one_hot_i[5];
  assign data_masked[696] = data_i[696] & sel_one_hot_i[5];
  assign data_masked[695] = data_i[695] & sel_one_hot_i[5];
  assign data_masked[694] = data_i[694] & sel_one_hot_i[5];
  assign data_masked[693] = data_i[693] & sel_one_hot_i[5];
  assign data_masked[692] = data_i[692] & sel_one_hot_i[5];
  assign data_masked[691] = data_i[691] & sel_one_hot_i[5];
  assign data_masked[690] = data_i[690] & sel_one_hot_i[5];
  assign data_masked[689] = data_i[689] & sel_one_hot_i[5];
  assign data_masked[688] = data_i[688] & sel_one_hot_i[5];
  assign data_masked[687] = data_i[687] & sel_one_hot_i[5];
  assign data_masked[686] = data_i[686] & sel_one_hot_i[5];
  assign data_masked[685] = data_i[685] & sel_one_hot_i[5];
  assign data_masked[684] = data_i[684] & sel_one_hot_i[5];
  assign data_masked[683] = data_i[683] & sel_one_hot_i[5];
  assign data_masked[682] = data_i[682] & sel_one_hot_i[5];
  assign data_masked[681] = data_i[681] & sel_one_hot_i[5];
  assign data_masked[680] = data_i[680] & sel_one_hot_i[5];
  assign data_masked[679] = data_i[679] & sel_one_hot_i[5];
  assign data_masked[678] = data_i[678] & sel_one_hot_i[5];
  assign data_masked[677] = data_i[677] & sel_one_hot_i[5];
  assign data_masked[676] = data_i[676] & sel_one_hot_i[5];
  assign data_masked[675] = data_i[675] & sel_one_hot_i[5];
  assign data_masked[674] = data_i[674] & sel_one_hot_i[5];
  assign data_masked[673] = data_i[673] & sel_one_hot_i[5];
  assign data_masked[672] = data_i[672] & sel_one_hot_i[5];
  assign data_masked[671] = data_i[671] & sel_one_hot_i[5];
  assign data_masked[670] = data_i[670] & sel_one_hot_i[5];
  assign data_masked[669] = data_i[669] & sel_one_hot_i[5];
  assign data_masked[668] = data_i[668] & sel_one_hot_i[5];
  assign data_masked[667] = data_i[667] & sel_one_hot_i[5];
  assign data_masked[666] = data_i[666] & sel_one_hot_i[5];
  assign data_masked[665] = data_i[665] & sel_one_hot_i[5];
  assign data_masked[664] = data_i[664] & sel_one_hot_i[5];
  assign data_masked[663] = data_i[663] & sel_one_hot_i[5];
  assign data_masked[662] = data_i[662] & sel_one_hot_i[5];
  assign data_masked[661] = data_i[661] & sel_one_hot_i[5];
  assign data_masked[660] = data_i[660] & sel_one_hot_i[5];
  assign data_masked[659] = data_i[659] & sel_one_hot_i[5];
  assign data_masked[658] = data_i[658] & sel_one_hot_i[5];
  assign data_masked[657] = data_i[657] & sel_one_hot_i[5];
  assign data_masked[656] = data_i[656] & sel_one_hot_i[5];
  assign data_masked[655] = data_i[655] & sel_one_hot_i[5];
  assign data_masked[654] = data_i[654] & sel_one_hot_i[5];
  assign data_masked[653] = data_i[653] & sel_one_hot_i[5];
  assign data_masked[652] = data_i[652] & sel_one_hot_i[5];
  assign data_masked[651] = data_i[651] & sel_one_hot_i[5];
  assign data_masked[650] = data_i[650] & sel_one_hot_i[5];
  assign data_masked[649] = data_i[649] & sel_one_hot_i[5];
  assign data_masked[648] = data_i[648] & sel_one_hot_i[5];
  assign data_masked[647] = data_i[647] & sel_one_hot_i[5];
  assign data_masked[646] = data_i[646] & sel_one_hot_i[5];
  assign data_masked[645] = data_i[645] & sel_one_hot_i[5];
  assign data_masked[644] = data_i[644] & sel_one_hot_i[5];
  assign data_masked[643] = data_i[643] & sel_one_hot_i[5];
  assign data_masked[642] = data_i[642] & sel_one_hot_i[5];
  assign data_masked[641] = data_i[641] & sel_one_hot_i[5];
  assign data_masked[640] = data_i[640] & sel_one_hot_i[5];
  assign data_masked[895] = data_i[895] & sel_one_hot_i[6];
  assign data_masked[894] = data_i[894] & sel_one_hot_i[6];
  assign data_masked[893] = data_i[893] & sel_one_hot_i[6];
  assign data_masked[892] = data_i[892] & sel_one_hot_i[6];
  assign data_masked[891] = data_i[891] & sel_one_hot_i[6];
  assign data_masked[890] = data_i[890] & sel_one_hot_i[6];
  assign data_masked[889] = data_i[889] & sel_one_hot_i[6];
  assign data_masked[888] = data_i[888] & sel_one_hot_i[6];
  assign data_masked[887] = data_i[887] & sel_one_hot_i[6];
  assign data_masked[886] = data_i[886] & sel_one_hot_i[6];
  assign data_masked[885] = data_i[885] & sel_one_hot_i[6];
  assign data_masked[884] = data_i[884] & sel_one_hot_i[6];
  assign data_masked[883] = data_i[883] & sel_one_hot_i[6];
  assign data_masked[882] = data_i[882] & sel_one_hot_i[6];
  assign data_masked[881] = data_i[881] & sel_one_hot_i[6];
  assign data_masked[880] = data_i[880] & sel_one_hot_i[6];
  assign data_masked[879] = data_i[879] & sel_one_hot_i[6];
  assign data_masked[878] = data_i[878] & sel_one_hot_i[6];
  assign data_masked[877] = data_i[877] & sel_one_hot_i[6];
  assign data_masked[876] = data_i[876] & sel_one_hot_i[6];
  assign data_masked[875] = data_i[875] & sel_one_hot_i[6];
  assign data_masked[874] = data_i[874] & sel_one_hot_i[6];
  assign data_masked[873] = data_i[873] & sel_one_hot_i[6];
  assign data_masked[872] = data_i[872] & sel_one_hot_i[6];
  assign data_masked[871] = data_i[871] & sel_one_hot_i[6];
  assign data_masked[870] = data_i[870] & sel_one_hot_i[6];
  assign data_masked[869] = data_i[869] & sel_one_hot_i[6];
  assign data_masked[868] = data_i[868] & sel_one_hot_i[6];
  assign data_masked[867] = data_i[867] & sel_one_hot_i[6];
  assign data_masked[866] = data_i[866] & sel_one_hot_i[6];
  assign data_masked[865] = data_i[865] & sel_one_hot_i[6];
  assign data_masked[864] = data_i[864] & sel_one_hot_i[6];
  assign data_masked[863] = data_i[863] & sel_one_hot_i[6];
  assign data_masked[862] = data_i[862] & sel_one_hot_i[6];
  assign data_masked[861] = data_i[861] & sel_one_hot_i[6];
  assign data_masked[860] = data_i[860] & sel_one_hot_i[6];
  assign data_masked[859] = data_i[859] & sel_one_hot_i[6];
  assign data_masked[858] = data_i[858] & sel_one_hot_i[6];
  assign data_masked[857] = data_i[857] & sel_one_hot_i[6];
  assign data_masked[856] = data_i[856] & sel_one_hot_i[6];
  assign data_masked[855] = data_i[855] & sel_one_hot_i[6];
  assign data_masked[854] = data_i[854] & sel_one_hot_i[6];
  assign data_masked[853] = data_i[853] & sel_one_hot_i[6];
  assign data_masked[852] = data_i[852] & sel_one_hot_i[6];
  assign data_masked[851] = data_i[851] & sel_one_hot_i[6];
  assign data_masked[850] = data_i[850] & sel_one_hot_i[6];
  assign data_masked[849] = data_i[849] & sel_one_hot_i[6];
  assign data_masked[848] = data_i[848] & sel_one_hot_i[6];
  assign data_masked[847] = data_i[847] & sel_one_hot_i[6];
  assign data_masked[846] = data_i[846] & sel_one_hot_i[6];
  assign data_masked[845] = data_i[845] & sel_one_hot_i[6];
  assign data_masked[844] = data_i[844] & sel_one_hot_i[6];
  assign data_masked[843] = data_i[843] & sel_one_hot_i[6];
  assign data_masked[842] = data_i[842] & sel_one_hot_i[6];
  assign data_masked[841] = data_i[841] & sel_one_hot_i[6];
  assign data_masked[840] = data_i[840] & sel_one_hot_i[6];
  assign data_masked[839] = data_i[839] & sel_one_hot_i[6];
  assign data_masked[838] = data_i[838] & sel_one_hot_i[6];
  assign data_masked[837] = data_i[837] & sel_one_hot_i[6];
  assign data_masked[836] = data_i[836] & sel_one_hot_i[6];
  assign data_masked[835] = data_i[835] & sel_one_hot_i[6];
  assign data_masked[834] = data_i[834] & sel_one_hot_i[6];
  assign data_masked[833] = data_i[833] & sel_one_hot_i[6];
  assign data_masked[832] = data_i[832] & sel_one_hot_i[6];
  assign data_masked[831] = data_i[831] & sel_one_hot_i[6];
  assign data_masked[830] = data_i[830] & sel_one_hot_i[6];
  assign data_masked[829] = data_i[829] & sel_one_hot_i[6];
  assign data_masked[828] = data_i[828] & sel_one_hot_i[6];
  assign data_masked[827] = data_i[827] & sel_one_hot_i[6];
  assign data_masked[826] = data_i[826] & sel_one_hot_i[6];
  assign data_masked[825] = data_i[825] & sel_one_hot_i[6];
  assign data_masked[824] = data_i[824] & sel_one_hot_i[6];
  assign data_masked[823] = data_i[823] & sel_one_hot_i[6];
  assign data_masked[822] = data_i[822] & sel_one_hot_i[6];
  assign data_masked[821] = data_i[821] & sel_one_hot_i[6];
  assign data_masked[820] = data_i[820] & sel_one_hot_i[6];
  assign data_masked[819] = data_i[819] & sel_one_hot_i[6];
  assign data_masked[818] = data_i[818] & sel_one_hot_i[6];
  assign data_masked[817] = data_i[817] & sel_one_hot_i[6];
  assign data_masked[816] = data_i[816] & sel_one_hot_i[6];
  assign data_masked[815] = data_i[815] & sel_one_hot_i[6];
  assign data_masked[814] = data_i[814] & sel_one_hot_i[6];
  assign data_masked[813] = data_i[813] & sel_one_hot_i[6];
  assign data_masked[812] = data_i[812] & sel_one_hot_i[6];
  assign data_masked[811] = data_i[811] & sel_one_hot_i[6];
  assign data_masked[810] = data_i[810] & sel_one_hot_i[6];
  assign data_masked[809] = data_i[809] & sel_one_hot_i[6];
  assign data_masked[808] = data_i[808] & sel_one_hot_i[6];
  assign data_masked[807] = data_i[807] & sel_one_hot_i[6];
  assign data_masked[806] = data_i[806] & sel_one_hot_i[6];
  assign data_masked[805] = data_i[805] & sel_one_hot_i[6];
  assign data_masked[804] = data_i[804] & sel_one_hot_i[6];
  assign data_masked[803] = data_i[803] & sel_one_hot_i[6];
  assign data_masked[802] = data_i[802] & sel_one_hot_i[6];
  assign data_masked[801] = data_i[801] & sel_one_hot_i[6];
  assign data_masked[800] = data_i[800] & sel_one_hot_i[6];
  assign data_masked[799] = data_i[799] & sel_one_hot_i[6];
  assign data_masked[798] = data_i[798] & sel_one_hot_i[6];
  assign data_masked[797] = data_i[797] & sel_one_hot_i[6];
  assign data_masked[796] = data_i[796] & sel_one_hot_i[6];
  assign data_masked[795] = data_i[795] & sel_one_hot_i[6];
  assign data_masked[794] = data_i[794] & sel_one_hot_i[6];
  assign data_masked[793] = data_i[793] & sel_one_hot_i[6];
  assign data_masked[792] = data_i[792] & sel_one_hot_i[6];
  assign data_masked[791] = data_i[791] & sel_one_hot_i[6];
  assign data_masked[790] = data_i[790] & sel_one_hot_i[6];
  assign data_masked[789] = data_i[789] & sel_one_hot_i[6];
  assign data_masked[788] = data_i[788] & sel_one_hot_i[6];
  assign data_masked[787] = data_i[787] & sel_one_hot_i[6];
  assign data_masked[786] = data_i[786] & sel_one_hot_i[6];
  assign data_masked[785] = data_i[785] & sel_one_hot_i[6];
  assign data_masked[784] = data_i[784] & sel_one_hot_i[6];
  assign data_masked[783] = data_i[783] & sel_one_hot_i[6];
  assign data_masked[782] = data_i[782] & sel_one_hot_i[6];
  assign data_masked[781] = data_i[781] & sel_one_hot_i[6];
  assign data_masked[780] = data_i[780] & sel_one_hot_i[6];
  assign data_masked[779] = data_i[779] & sel_one_hot_i[6];
  assign data_masked[778] = data_i[778] & sel_one_hot_i[6];
  assign data_masked[777] = data_i[777] & sel_one_hot_i[6];
  assign data_masked[776] = data_i[776] & sel_one_hot_i[6];
  assign data_masked[775] = data_i[775] & sel_one_hot_i[6];
  assign data_masked[774] = data_i[774] & sel_one_hot_i[6];
  assign data_masked[773] = data_i[773] & sel_one_hot_i[6];
  assign data_masked[772] = data_i[772] & sel_one_hot_i[6];
  assign data_masked[771] = data_i[771] & sel_one_hot_i[6];
  assign data_masked[770] = data_i[770] & sel_one_hot_i[6];
  assign data_masked[769] = data_i[769] & sel_one_hot_i[6];
  assign data_masked[768] = data_i[768] & sel_one_hot_i[6];
  assign data_masked[1023] = data_i[1023] & sel_one_hot_i[7];
  assign data_masked[1022] = data_i[1022] & sel_one_hot_i[7];
  assign data_masked[1021] = data_i[1021] & sel_one_hot_i[7];
  assign data_masked[1020] = data_i[1020] & sel_one_hot_i[7];
  assign data_masked[1019] = data_i[1019] & sel_one_hot_i[7];
  assign data_masked[1018] = data_i[1018] & sel_one_hot_i[7];
  assign data_masked[1017] = data_i[1017] & sel_one_hot_i[7];
  assign data_masked[1016] = data_i[1016] & sel_one_hot_i[7];
  assign data_masked[1015] = data_i[1015] & sel_one_hot_i[7];
  assign data_masked[1014] = data_i[1014] & sel_one_hot_i[7];
  assign data_masked[1013] = data_i[1013] & sel_one_hot_i[7];
  assign data_masked[1012] = data_i[1012] & sel_one_hot_i[7];
  assign data_masked[1011] = data_i[1011] & sel_one_hot_i[7];
  assign data_masked[1010] = data_i[1010] & sel_one_hot_i[7];
  assign data_masked[1009] = data_i[1009] & sel_one_hot_i[7];
  assign data_masked[1008] = data_i[1008] & sel_one_hot_i[7];
  assign data_masked[1007] = data_i[1007] & sel_one_hot_i[7];
  assign data_masked[1006] = data_i[1006] & sel_one_hot_i[7];
  assign data_masked[1005] = data_i[1005] & sel_one_hot_i[7];
  assign data_masked[1004] = data_i[1004] & sel_one_hot_i[7];
  assign data_masked[1003] = data_i[1003] & sel_one_hot_i[7];
  assign data_masked[1002] = data_i[1002] & sel_one_hot_i[7];
  assign data_masked[1001] = data_i[1001] & sel_one_hot_i[7];
  assign data_masked[1000] = data_i[1000] & sel_one_hot_i[7];
  assign data_masked[999] = data_i[999] & sel_one_hot_i[7];
  assign data_masked[998] = data_i[998] & sel_one_hot_i[7];
  assign data_masked[997] = data_i[997] & sel_one_hot_i[7];
  assign data_masked[996] = data_i[996] & sel_one_hot_i[7];
  assign data_masked[995] = data_i[995] & sel_one_hot_i[7];
  assign data_masked[994] = data_i[994] & sel_one_hot_i[7];
  assign data_masked[993] = data_i[993] & sel_one_hot_i[7];
  assign data_masked[992] = data_i[992] & sel_one_hot_i[7];
  assign data_masked[991] = data_i[991] & sel_one_hot_i[7];
  assign data_masked[990] = data_i[990] & sel_one_hot_i[7];
  assign data_masked[989] = data_i[989] & sel_one_hot_i[7];
  assign data_masked[988] = data_i[988] & sel_one_hot_i[7];
  assign data_masked[987] = data_i[987] & sel_one_hot_i[7];
  assign data_masked[986] = data_i[986] & sel_one_hot_i[7];
  assign data_masked[985] = data_i[985] & sel_one_hot_i[7];
  assign data_masked[984] = data_i[984] & sel_one_hot_i[7];
  assign data_masked[983] = data_i[983] & sel_one_hot_i[7];
  assign data_masked[982] = data_i[982] & sel_one_hot_i[7];
  assign data_masked[981] = data_i[981] & sel_one_hot_i[7];
  assign data_masked[980] = data_i[980] & sel_one_hot_i[7];
  assign data_masked[979] = data_i[979] & sel_one_hot_i[7];
  assign data_masked[978] = data_i[978] & sel_one_hot_i[7];
  assign data_masked[977] = data_i[977] & sel_one_hot_i[7];
  assign data_masked[976] = data_i[976] & sel_one_hot_i[7];
  assign data_masked[975] = data_i[975] & sel_one_hot_i[7];
  assign data_masked[974] = data_i[974] & sel_one_hot_i[7];
  assign data_masked[973] = data_i[973] & sel_one_hot_i[7];
  assign data_masked[972] = data_i[972] & sel_one_hot_i[7];
  assign data_masked[971] = data_i[971] & sel_one_hot_i[7];
  assign data_masked[970] = data_i[970] & sel_one_hot_i[7];
  assign data_masked[969] = data_i[969] & sel_one_hot_i[7];
  assign data_masked[968] = data_i[968] & sel_one_hot_i[7];
  assign data_masked[967] = data_i[967] & sel_one_hot_i[7];
  assign data_masked[966] = data_i[966] & sel_one_hot_i[7];
  assign data_masked[965] = data_i[965] & sel_one_hot_i[7];
  assign data_masked[964] = data_i[964] & sel_one_hot_i[7];
  assign data_masked[963] = data_i[963] & sel_one_hot_i[7];
  assign data_masked[962] = data_i[962] & sel_one_hot_i[7];
  assign data_masked[961] = data_i[961] & sel_one_hot_i[7];
  assign data_masked[960] = data_i[960] & sel_one_hot_i[7];
  assign data_masked[959] = data_i[959] & sel_one_hot_i[7];
  assign data_masked[958] = data_i[958] & sel_one_hot_i[7];
  assign data_masked[957] = data_i[957] & sel_one_hot_i[7];
  assign data_masked[956] = data_i[956] & sel_one_hot_i[7];
  assign data_masked[955] = data_i[955] & sel_one_hot_i[7];
  assign data_masked[954] = data_i[954] & sel_one_hot_i[7];
  assign data_masked[953] = data_i[953] & sel_one_hot_i[7];
  assign data_masked[952] = data_i[952] & sel_one_hot_i[7];
  assign data_masked[951] = data_i[951] & sel_one_hot_i[7];
  assign data_masked[950] = data_i[950] & sel_one_hot_i[7];
  assign data_masked[949] = data_i[949] & sel_one_hot_i[7];
  assign data_masked[948] = data_i[948] & sel_one_hot_i[7];
  assign data_masked[947] = data_i[947] & sel_one_hot_i[7];
  assign data_masked[946] = data_i[946] & sel_one_hot_i[7];
  assign data_masked[945] = data_i[945] & sel_one_hot_i[7];
  assign data_masked[944] = data_i[944] & sel_one_hot_i[7];
  assign data_masked[943] = data_i[943] & sel_one_hot_i[7];
  assign data_masked[942] = data_i[942] & sel_one_hot_i[7];
  assign data_masked[941] = data_i[941] & sel_one_hot_i[7];
  assign data_masked[940] = data_i[940] & sel_one_hot_i[7];
  assign data_masked[939] = data_i[939] & sel_one_hot_i[7];
  assign data_masked[938] = data_i[938] & sel_one_hot_i[7];
  assign data_masked[937] = data_i[937] & sel_one_hot_i[7];
  assign data_masked[936] = data_i[936] & sel_one_hot_i[7];
  assign data_masked[935] = data_i[935] & sel_one_hot_i[7];
  assign data_masked[934] = data_i[934] & sel_one_hot_i[7];
  assign data_masked[933] = data_i[933] & sel_one_hot_i[7];
  assign data_masked[932] = data_i[932] & sel_one_hot_i[7];
  assign data_masked[931] = data_i[931] & sel_one_hot_i[7];
  assign data_masked[930] = data_i[930] & sel_one_hot_i[7];
  assign data_masked[929] = data_i[929] & sel_one_hot_i[7];
  assign data_masked[928] = data_i[928] & sel_one_hot_i[7];
  assign data_masked[927] = data_i[927] & sel_one_hot_i[7];
  assign data_masked[926] = data_i[926] & sel_one_hot_i[7];
  assign data_masked[925] = data_i[925] & sel_one_hot_i[7];
  assign data_masked[924] = data_i[924] & sel_one_hot_i[7];
  assign data_masked[923] = data_i[923] & sel_one_hot_i[7];
  assign data_masked[922] = data_i[922] & sel_one_hot_i[7];
  assign data_masked[921] = data_i[921] & sel_one_hot_i[7];
  assign data_masked[920] = data_i[920] & sel_one_hot_i[7];
  assign data_masked[919] = data_i[919] & sel_one_hot_i[7];
  assign data_masked[918] = data_i[918] & sel_one_hot_i[7];
  assign data_masked[917] = data_i[917] & sel_one_hot_i[7];
  assign data_masked[916] = data_i[916] & sel_one_hot_i[7];
  assign data_masked[915] = data_i[915] & sel_one_hot_i[7];
  assign data_masked[914] = data_i[914] & sel_one_hot_i[7];
  assign data_masked[913] = data_i[913] & sel_one_hot_i[7];
  assign data_masked[912] = data_i[912] & sel_one_hot_i[7];
  assign data_masked[911] = data_i[911] & sel_one_hot_i[7];
  assign data_masked[910] = data_i[910] & sel_one_hot_i[7];
  assign data_masked[909] = data_i[909] & sel_one_hot_i[7];
  assign data_masked[908] = data_i[908] & sel_one_hot_i[7];
  assign data_masked[907] = data_i[907] & sel_one_hot_i[7];
  assign data_masked[906] = data_i[906] & sel_one_hot_i[7];
  assign data_masked[905] = data_i[905] & sel_one_hot_i[7];
  assign data_masked[904] = data_i[904] & sel_one_hot_i[7];
  assign data_masked[903] = data_i[903] & sel_one_hot_i[7];
  assign data_masked[902] = data_i[902] & sel_one_hot_i[7];
  assign data_masked[901] = data_i[901] & sel_one_hot_i[7];
  assign data_masked[900] = data_i[900] & sel_one_hot_i[7];
  assign data_masked[899] = data_i[899] & sel_one_hot_i[7];
  assign data_masked[898] = data_i[898] & sel_one_hot_i[7];
  assign data_masked[897] = data_i[897] & sel_one_hot_i[7];
  assign data_masked[896] = data_i[896] & sel_one_hot_i[7];
  assign data_masked[1151] = data_i[1151] & sel_one_hot_i[8];
  assign data_masked[1150] = data_i[1150] & sel_one_hot_i[8];
  assign data_masked[1149] = data_i[1149] & sel_one_hot_i[8];
  assign data_masked[1148] = data_i[1148] & sel_one_hot_i[8];
  assign data_masked[1147] = data_i[1147] & sel_one_hot_i[8];
  assign data_masked[1146] = data_i[1146] & sel_one_hot_i[8];
  assign data_masked[1145] = data_i[1145] & sel_one_hot_i[8];
  assign data_masked[1144] = data_i[1144] & sel_one_hot_i[8];
  assign data_masked[1143] = data_i[1143] & sel_one_hot_i[8];
  assign data_masked[1142] = data_i[1142] & sel_one_hot_i[8];
  assign data_masked[1141] = data_i[1141] & sel_one_hot_i[8];
  assign data_masked[1140] = data_i[1140] & sel_one_hot_i[8];
  assign data_masked[1139] = data_i[1139] & sel_one_hot_i[8];
  assign data_masked[1138] = data_i[1138] & sel_one_hot_i[8];
  assign data_masked[1137] = data_i[1137] & sel_one_hot_i[8];
  assign data_masked[1136] = data_i[1136] & sel_one_hot_i[8];
  assign data_masked[1135] = data_i[1135] & sel_one_hot_i[8];
  assign data_masked[1134] = data_i[1134] & sel_one_hot_i[8];
  assign data_masked[1133] = data_i[1133] & sel_one_hot_i[8];
  assign data_masked[1132] = data_i[1132] & sel_one_hot_i[8];
  assign data_masked[1131] = data_i[1131] & sel_one_hot_i[8];
  assign data_masked[1130] = data_i[1130] & sel_one_hot_i[8];
  assign data_masked[1129] = data_i[1129] & sel_one_hot_i[8];
  assign data_masked[1128] = data_i[1128] & sel_one_hot_i[8];
  assign data_masked[1127] = data_i[1127] & sel_one_hot_i[8];
  assign data_masked[1126] = data_i[1126] & sel_one_hot_i[8];
  assign data_masked[1125] = data_i[1125] & sel_one_hot_i[8];
  assign data_masked[1124] = data_i[1124] & sel_one_hot_i[8];
  assign data_masked[1123] = data_i[1123] & sel_one_hot_i[8];
  assign data_masked[1122] = data_i[1122] & sel_one_hot_i[8];
  assign data_masked[1121] = data_i[1121] & sel_one_hot_i[8];
  assign data_masked[1120] = data_i[1120] & sel_one_hot_i[8];
  assign data_masked[1119] = data_i[1119] & sel_one_hot_i[8];
  assign data_masked[1118] = data_i[1118] & sel_one_hot_i[8];
  assign data_masked[1117] = data_i[1117] & sel_one_hot_i[8];
  assign data_masked[1116] = data_i[1116] & sel_one_hot_i[8];
  assign data_masked[1115] = data_i[1115] & sel_one_hot_i[8];
  assign data_masked[1114] = data_i[1114] & sel_one_hot_i[8];
  assign data_masked[1113] = data_i[1113] & sel_one_hot_i[8];
  assign data_masked[1112] = data_i[1112] & sel_one_hot_i[8];
  assign data_masked[1111] = data_i[1111] & sel_one_hot_i[8];
  assign data_masked[1110] = data_i[1110] & sel_one_hot_i[8];
  assign data_masked[1109] = data_i[1109] & sel_one_hot_i[8];
  assign data_masked[1108] = data_i[1108] & sel_one_hot_i[8];
  assign data_masked[1107] = data_i[1107] & sel_one_hot_i[8];
  assign data_masked[1106] = data_i[1106] & sel_one_hot_i[8];
  assign data_masked[1105] = data_i[1105] & sel_one_hot_i[8];
  assign data_masked[1104] = data_i[1104] & sel_one_hot_i[8];
  assign data_masked[1103] = data_i[1103] & sel_one_hot_i[8];
  assign data_masked[1102] = data_i[1102] & sel_one_hot_i[8];
  assign data_masked[1101] = data_i[1101] & sel_one_hot_i[8];
  assign data_masked[1100] = data_i[1100] & sel_one_hot_i[8];
  assign data_masked[1099] = data_i[1099] & sel_one_hot_i[8];
  assign data_masked[1098] = data_i[1098] & sel_one_hot_i[8];
  assign data_masked[1097] = data_i[1097] & sel_one_hot_i[8];
  assign data_masked[1096] = data_i[1096] & sel_one_hot_i[8];
  assign data_masked[1095] = data_i[1095] & sel_one_hot_i[8];
  assign data_masked[1094] = data_i[1094] & sel_one_hot_i[8];
  assign data_masked[1093] = data_i[1093] & sel_one_hot_i[8];
  assign data_masked[1092] = data_i[1092] & sel_one_hot_i[8];
  assign data_masked[1091] = data_i[1091] & sel_one_hot_i[8];
  assign data_masked[1090] = data_i[1090] & sel_one_hot_i[8];
  assign data_masked[1089] = data_i[1089] & sel_one_hot_i[8];
  assign data_masked[1088] = data_i[1088] & sel_one_hot_i[8];
  assign data_masked[1087] = data_i[1087] & sel_one_hot_i[8];
  assign data_masked[1086] = data_i[1086] & sel_one_hot_i[8];
  assign data_masked[1085] = data_i[1085] & sel_one_hot_i[8];
  assign data_masked[1084] = data_i[1084] & sel_one_hot_i[8];
  assign data_masked[1083] = data_i[1083] & sel_one_hot_i[8];
  assign data_masked[1082] = data_i[1082] & sel_one_hot_i[8];
  assign data_masked[1081] = data_i[1081] & sel_one_hot_i[8];
  assign data_masked[1080] = data_i[1080] & sel_one_hot_i[8];
  assign data_masked[1079] = data_i[1079] & sel_one_hot_i[8];
  assign data_masked[1078] = data_i[1078] & sel_one_hot_i[8];
  assign data_masked[1077] = data_i[1077] & sel_one_hot_i[8];
  assign data_masked[1076] = data_i[1076] & sel_one_hot_i[8];
  assign data_masked[1075] = data_i[1075] & sel_one_hot_i[8];
  assign data_masked[1074] = data_i[1074] & sel_one_hot_i[8];
  assign data_masked[1073] = data_i[1073] & sel_one_hot_i[8];
  assign data_masked[1072] = data_i[1072] & sel_one_hot_i[8];
  assign data_masked[1071] = data_i[1071] & sel_one_hot_i[8];
  assign data_masked[1070] = data_i[1070] & sel_one_hot_i[8];
  assign data_masked[1069] = data_i[1069] & sel_one_hot_i[8];
  assign data_masked[1068] = data_i[1068] & sel_one_hot_i[8];
  assign data_masked[1067] = data_i[1067] & sel_one_hot_i[8];
  assign data_masked[1066] = data_i[1066] & sel_one_hot_i[8];
  assign data_masked[1065] = data_i[1065] & sel_one_hot_i[8];
  assign data_masked[1064] = data_i[1064] & sel_one_hot_i[8];
  assign data_masked[1063] = data_i[1063] & sel_one_hot_i[8];
  assign data_masked[1062] = data_i[1062] & sel_one_hot_i[8];
  assign data_masked[1061] = data_i[1061] & sel_one_hot_i[8];
  assign data_masked[1060] = data_i[1060] & sel_one_hot_i[8];
  assign data_masked[1059] = data_i[1059] & sel_one_hot_i[8];
  assign data_masked[1058] = data_i[1058] & sel_one_hot_i[8];
  assign data_masked[1057] = data_i[1057] & sel_one_hot_i[8];
  assign data_masked[1056] = data_i[1056] & sel_one_hot_i[8];
  assign data_masked[1055] = data_i[1055] & sel_one_hot_i[8];
  assign data_masked[1054] = data_i[1054] & sel_one_hot_i[8];
  assign data_masked[1053] = data_i[1053] & sel_one_hot_i[8];
  assign data_masked[1052] = data_i[1052] & sel_one_hot_i[8];
  assign data_masked[1051] = data_i[1051] & sel_one_hot_i[8];
  assign data_masked[1050] = data_i[1050] & sel_one_hot_i[8];
  assign data_masked[1049] = data_i[1049] & sel_one_hot_i[8];
  assign data_masked[1048] = data_i[1048] & sel_one_hot_i[8];
  assign data_masked[1047] = data_i[1047] & sel_one_hot_i[8];
  assign data_masked[1046] = data_i[1046] & sel_one_hot_i[8];
  assign data_masked[1045] = data_i[1045] & sel_one_hot_i[8];
  assign data_masked[1044] = data_i[1044] & sel_one_hot_i[8];
  assign data_masked[1043] = data_i[1043] & sel_one_hot_i[8];
  assign data_masked[1042] = data_i[1042] & sel_one_hot_i[8];
  assign data_masked[1041] = data_i[1041] & sel_one_hot_i[8];
  assign data_masked[1040] = data_i[1040] & sel_one_hot_i[8];
  assign data_masked[1039] = data_i[1039] & sel_one_hot_i[8];
  assign data_masked[1038] = data_i[1038] & sel_one_hot_i[8];
  assign data_masked[1037] = data_i[1037] & sel_one_hot_i[8];
  assign data_masked[1036] = data_i[1036] & sel_one_hot_i[8];
  assign data_masked[1035] = data_i[1035] & sel_one_hot_i[8];
  assign data_masked[1034] = data_i[1034] & sel_one_hot_i[8];
  assign data_masked[1033] = data_i[1033] & sel_one_hot_i[8];
  assign data_masked[1032] = data_i[1032] & sel_one_hot_i[8];
  assign data_masked[1031] = data_i[1031] & sel_one_hot_i[8];
  assign data_masked[1030] = data_i[1030] & sel_one_hot_i[8];
  assign data_masked[1029] = data_i[1029] & sel_one_hot_i[8];
  assign data_masked[1028] = data_i[1028] & sel_one_hot_i[8];
  assign data_masked[1027] = data_i[1027] & sel_one_hot_i[8];
  assign data_masked[1026] = data_i[1026] & sel_one_hot_i[8];
  assign data_masked[1025] = data_i[1025] & sel_one_hot_i[8];
  assign data_masked[1024] = data_i[1024] & sel_one_hot_i[8];
  assign data_masked[1279] = data_i[1279] & sel_one_hot_i[9];
  assign data_masked[1278] = data_i[1278] & sel_one_hot_i[9];
  assign data_masked[1277] = data_i[1277] & sel_one_hot_i[9];
  assign data_masked[1276] = data_i[1276] & sel_one_hot_i[9];
  assign data_masked[1275] = data_i[1275] & sel_one_hot_i[9];
  assign data_masked[1274] = data_i[1274] & sel_one_hot_i[9];
  assign data_masked[1273] = data_i[1273] & sel_one_hot_i[9];
  assign data_masked[1272] = data_i[1272] & sel_one_hot_i[9];
  assign data_masked[1271] = data_i[1271] & sel_one_hot_i[9];
  assign data_masked[1270] = data_i[1270] & sel_one_hot_i[9];
  assign data_masked[1269] = data_i[1269] & sel_one_hot_i[9];
  assign data_masked[1268] = data_i[1268] & sel_one_hot_i[9];
  assign data_masked[1267] = data_i[1267] & sel_one_hot_i[9];
  assign data_masked[1266] = data_i[1266] & sel_one_hot_i[9];
  assign data_masked[1265] = data_i[1265] & sel_one_hot_i[9];
  assign data_masked[1264] = data_i[1264] & sel_one_hot_i[9];
  assign data_masked[1263] = data_i[1263] & sel_one_hot_i[9];
  assign data_masked[1262] = data_i[1262] & sel_one_hot_i[9];
  assign data_masked[1261] = data_i[1261] & sel_one_hot_i[9];
  assign data_masked[1260] = data_i[1260] & sel_one_hot_i[9];
  assign data_masked[1259] = data_i[1259] & sel_one_hot_i[9];
  assign data_masked[1258] = data_i[1258] & sel_one_hot_i[9];
  assign data_masked[1257] = data_i[1257] & sel_one_hot_i[9];
  assign data_masked[1256] = data_i[1256] & sel_one_hot_i[9];
  assign data_masked[1255] = data_i[1255] & sel_one_hot_i[9];
  assign data_masked[1254] = data_i[1254] & sel_one_hot_i[9];
  assign data_masked[1253] = data_i[1253] & sel_one_hot_i[9];
  assign data_masked[1252] = data_i[1252] & sel_one_hot_i[9];
  assign data_masked[1251] = data_i[1251] & sel_one_hot_i[9];
  assign data_masked[1250] = data_i[1250] & sel_one_hot_i[9];
  assign data_masked[1249] = data_i[1249] & sel_one_hot_i[9];
  assign data_masked[1248] = data_i[1248] & sel_one_hot_i[9];
  assign data_masked[1247] = data_i[1247] & sel_one_hot_i[9];
  assign data_masked[1246] = data_i[1246] & sel_one_hot_i[9];
  assign data_masked[1245] = data_i[1245] & sel_one_hot_i[9];
  assign data_masked[1244] = data_i[1244] & sel_one_hot_i[9];
  assign data_masked[1243] = data_i[1243] & sel_one_hot_i[9];
  assign data_masked[1242] = data_i[1242] & sel_one_hot_i[9];
  assign data_masked[1241] = data_i[1241] & sel_one_hot_i[9];
  assign data_masked[1240] = data_i[1240] & sel_one_hot_i[9];
  assign data_masked[1239] = data_i[1239] & sel_one_hot_i[9];
  assign data_masked[1238] = data_i[1238] & sel_one_hot_i[9];
  assign data_masked[1237] = data_i[1237] & sel_one_hot_i[9];
  assign data_masked[1236] = data_i[1236] & sel_one_hot_i[9];
  assign data_masked[1235] = data_i[1235] & sel_one_hot_i[9];
  assign data_masked[1234] = data_i[1234] & sel_one_hot_i[9];
  assign data_masked[1233] = data_i[1233] & sel_one_hot_i[9];
  assign data_masked[1232] = data_i[1232] & sel_one_hot_i[9];
  assign data_masked[1231] = data_i[1231] & sel_one_hot_i[9];
  assign data_masked[1230] = data_i[1230] & sel_one_hot_i[9];
  assign data_masked[1229] = data_i[1229] & sel_one_hot_i[9];
  assign data_masked[1228] = data_i[1228] & sel_one_hot_i[9];
  assign data_masked[1227] = data_i[1227] & sel_one_hot_i[9];
  assign data_masked[1226] = data_i[1226] & sel_one_hot_i[9];
  assign data_masked[1225] = data_i[1225] & sel_one_hot_i[9];
  assign data_masked[1224] = data_i[1224] & sel_one_hot_i[9];
  assign data_masked[1223] = data_i[1223] & sel_one_hot_i[9];
  assign data_masked[1222] = data_i[1222] & sel_one_hot_i[9];
  assign data_masked[1221] = data_i[1221] & sel_one_hot_i[9];
  assign data_masked[1220] = data_i[1220] & sel_one_hot_i[9];
  assign data_masked[1219] = data_i[1219] & sel_one_hot_i[9];
  assign data_masked[1218] = data_i[1218] & sel_one_hot_i[9];
  assign data_masked[1217] = data_i[1217] & sel_one_hot_i[9];
  assign data_masked[1216] = data_i[1216] & sel_one_hot_i[9];
  assign data_masked[1215] = data_i[1215] & sel_one_hot_i[9];
  assign data_masked[1214] = data_i[1214] & sel_one_hot_i[9];
  assign data_masked[1213] = data_i[1213] & sel_one_hot_i[9];
  assign data_masked[1212] = data_i[1212] & sel_one_hot_i[9];
  assign data_masked[1211] = data_i[1211] & sel_one_hot_i[9];
  assign data_masked[1210] = data_i[1210] & sel_one_hot_i[9];
  assign data_masked[1209] = data_i[1209] & sel_one_hot_i[9];
  assign data_masked[1208] = data_i[1208] & sel_one_hot_i[9];
  assign data_masked[1207] = data_i[1207] & sel_one_hot_i[9];
  assign data_masked[1206] = data_i[1206] & sel_one_hot_i[9];
  assign data_masked[1205] = data_i[1205] & sel_one_hot_i[9];
  assign data_masked[1204] = data_i[1204] & sel_one_hot_i[9];
  assign data_masked[1203] = data_i[1203] & sel_one_hot_i[9];
  assign data_masked[1202] = data_i[1202] & sel_one_hot_i[9];
  assign data_masked[1201] = data_i[1201] & sel_one_hot_i[9];
  assign data_masked[1200] = data_i[1200] & sel_one_hot_i[9];
  assign data_masked[1199] = data_i[1199] & sel_one_hot_i[9];
  assign data_masked[1198] = data_i[1198] & sel_one_hot_i[9];
  assign data_masked[1197] = data_i[1197] & sel_one_hot_i[9];
  assign data_masked[1196] = data_i[1196] & sel_one_hot_i[9];
  assign data_masked[1195] = data_i[1195] & sel_one_hot_i[9];
  assign data_masked[1194] = data_i[1194] & sel_one_hot_i[9];
  assign data_masked[1193] = data_i[1193] & sel_one_hot_i[9];
  assign data_masked[1192] = data_i[1192] & sel_one_hot_i[9];
  assign data_masked[1191] = data_i[1191] & sel_one_hot_i[9];
  assign data_masked[1190] = data_i[1190] & sel_one_hot_i[9];
  assign data_masked[1189] = data_i[1189] & sel_one_hot_i[9];
  assign data_masked[1188] = data_i[1188] & sel_one_hot_i[9];
  assign data_masked[1187] = data_i[1187] & sel_one_hot_i[9];
  assign data_masked[1186] = data_i[1186] & sel_one_hot_i[9];
  assign data_masked[1185] = data_i[1185] & sel_one_hot_i[9];
  assign data_masked[1184] = data_i[1184] & sel_one_hot_i[9];
  assign data_masked[1183] = data_i[1183] & sel_one_hot_i[9];
  assign data_masked[1182] = data_i[1182] & sel_one_hot_i[9];
  assign data_masked[1181] = data_i[1181] & sel_one_hot_i[9];
  assign data_masked[1180] = data_i[1180] & sel_one_hot_i[9];
  assign data_masked[1179] = data_i[1179] & sel_one_hot_i[9];
  assign data_masked[1178] = data_i[1178] & sel_one_hot_i[9];
  assign data_masked[1177] = data_i[1177] & sel_one_hot_i[9];
  assign data_masked[1176] = data_i[1176] & sel_one_hot_i[9];
  assign data_masked[1175] = data_i[1175] & sel_one_hot_i[9];
  assign data_masked[1174] = data_i[1174] & sel_one_hot_i[9];
  assign data_masked[1173] = data_i[1173] & sel_one_hot_i[9];
  assign data_masked[1172] = data_i[1172] & sel_one_hot_i[9];
  assign data_masked[1171] = data_i[1171] & sel_one_hot_i[9];
  assign data_masked[1170] = data_i[1170] & sel_one_hot_i[9];
  assign data_masked[1169] = data_i[1169] & sel_one_hot_i[9];
  assign data_masked[1168] = data_i[1168] & sel_one_hot_i[9];
  assign data_masked[1167] = data_i[1167] & sel_one_hot_i[9];
  assign data_masked[1166] = data_i[1166] & sel_one_hot_i[9];
  assign data_masked[1165] = data_i[1165] & sel_one_hot_i[9];
  assign data_masked[1164] = data_i[1164] & sel_one_hot_i[9];
  assign data_masked[1163] = data_i[1163] & sel_one_hot_i[9];
  assign data_masked[1162] = data_i[1162] & sel_one_hot_i[9];
  assign data_masked[1161] = data_i[1161] & sel_one_hot_i[9];
  assign data_masked[1160] = data_i[1160] & sel_one_hot_i[9];
  assign data_masked[1159] = data_i[1159] & sel_one_hot_i[9];
  assign data_masked[1158] = data_i[1158] & sel_one_hot_i[9];
  assign data_masked[1157] = data_i[1157] & sel_one_hot_i[9];
  assign data_masked[1156] = data_i[1156] & sel_one_hot_i[9];
  assign data_masked[1155] = data_i[1155] & sel_one_hot_i[9];
  assign data_masked[1154] = data_i[1154] & sel_one_hot_i[9];
  assign data_masked[1153] = data_i[1153] & sel_one_hot_i[9];
  assign data_masked[1152] = data_i[1152] & sel_one_hot_i[9];
  assign data_masked[1407] = data_i[1407] & sel_one_hot_i[10];
  assign data_masked[1406] = data_i[1406] & sel_one_hot_i[10];
  assign data_masked[1405] = data_i[1405] & sel_one_hot_i[10];
  assign data_masked[1404] = data_i[1404] & sel_one_hot_i[10];
  assign data_masked[1403] = data_i[1403] & sel_one_hot_i[10];
  assign data_masked[1402] = data_i[1402] & sel_one_hot_i[10];
  assign data_masked[1401] = data_i[1401] & sel_one_hot_i[10];
  assign data_masked[1400] = data_i[1400] & sel_one_hot_i[10];
  assign data_masked[1399] = data_i[1399] & sel_one_hot_i[10];
  assign data_masked[1398] = data_i[1398] & sel_one_hot_i[10];
  assign data_masked[1397] = data_i[1397] & sel_one_hot_i[10];
  assign data_masked[1396] = data_i[1396] & sel_one_hot_i[10];
  assign data_masked[1395] = data_i[1395] & sel_one_hot_i[10];
  assign data_masked[1394] = data_i[1394] & sel_one_hot_i[10];
  assign data_masked[1393] = data_i[1393] & sel_one_hot_i[10];
  assign data_masked[1392] = data_i[1392] & sel_one_hot_i[10];
  assign data_masked[1391] = data_i[1391] & sel_one_hot_i[10];
  assign data_masked[1390] = data_i[1390] & sel_one_hot_i[10];
  assign data_masked[1389] = data_i[1389] & sel_one_hot_i[10];
  assign data_masked[1388] = data_i[1388] & sel_one_hot_i[10];
  assign data_masked[1387] = data_i[1387] & sel_one_hot_i[10];
  assign data_masked[1386] = data_i[1386] & sel_one_hot_i[10];
  assign data_masked[1385] = data_i[1385] & sel_one_hot_i[10];
  assign data_masked[1384] = data_i[1384] & sel_one_hot_i[10];
  assign data_masked[1383] = data_i[1383] & sel_one_hot_i[10];
  assign data_masked[1382] = data_i[1382] & sel_one_hot_i[10];
  assign data_masked[1381] = data_i[1381] & sel_one_hot_i[10];
  assign data_masked[1380] = data_i[1380] & sel_one_hot_i[10];
  assign data_masked[1379] = data_i[1379] & sel_one_hot_i[10];
  assign data_masked[1378] = data_i[1378] & sel_one_hot_i[10];
  assign data_masked[1377] = data_i[1377] & sel_one_hot_i[10];
  assign data_masked[1376] = data_i[1376] & sel_one_hot_i[10];
  assign data_masked[1375] = data_i[1375] & sel_one_hot_i[10];
  assign data_masked[1374] = data_i[1374] & sel_one_hot_i[10];
  assign data_masked[1373] = data_i[1373] & sel_one_hot_i[10];
  assign data_masked[1372] = data_i[1372] & sel_one_hot_i[10];
  assign data_masked[1371] = data_i[1371] & sel_one_hot_i[10];
  assign data_masked[1370] = data_i[1370] & sel_one_hot_i[10];
  assign data_masked[1369] = data_i[1369] & sel_one_hot_i[10];
  assign data_masked[1368] = data_i[1368] & sel_one_hot_i[10];
  assign data_masked[1367] = data_i[1367] & sel_one_hot_i[10];
  assign data_masked[1366] = data_i[1366] & sel_one_hot_i[10];
  assign data_masked[1365] = data_i[1365] & sel_one_hot_i[10];
  assign data_masked[1364] = data_i[1364] & sel_one_hot_i[10];
  assign data_masked[1363] = data_i[1363] & sel_one_hot_i[10];
  assign data_masked[1362] = data_i[1362] & sel_one_hot_i[10];
  assign data_masked[1361] = data_i[1361] & sel_one_hot_i[10];
  assign data_masked[1360] = data_i[1360] & sel_one_hot_i[10];
  assign data_masked[1359] = data_i[1359] & sel_one_hot_i[10];
  assign data_masked[1358] = data_i[1358] & sel_one_hot_i[10];
  assign data_masked[1357] = data_i[1357] & sel_one_hot_i[10];
  assign data_masked[1356] = data_i[1356] & sel_one_hot_i[10];
  assign data_masked[1355] = data_i[1355] & sel_one_hot_i[10];
  assign data_masked[1354] = data_i[1354] & sel_one_hot_i[10];
  assign data_masked[1353] = data_i[1353] & sel_one_hot_i[10];
  assign data_masked[1352] = data_i[1352] & sel_one_hot_i[10];
  assign data_masked[1351] = data_i[1351] & sel_one_hot_i[10];
  assign data_masked[1350] = data_i[1350] & sel_one_hot_i[10];
  assign data_masked[1349] = data_i[1349] & sel_one_hot_i[10];
  assign data_masked[1348] = data_i[1348] & sel_one_hot_i[10];
  assign data_masked[1347] = data_i[1347] & sel_one_hot_i[10];
  assign data_masked[1346] = data_i[1346] & sel_one_hot_i[10];
  assign data_masked[1345] = data_i[1345] & sel_one_hot_i[10];
  assign data_masked[1344] = data_i[1344] & sel_one_hot_i[10];
  assign data_masked[1343] = data_i[1343] & sel_one_hot_i[10];
  assign data_masked[1342] = data_i[1342] & sel_one_hot_i[10];
  assign data_masked[1341] = data_i[1341] & sel_one_hot_i[10];
  assign data_masked[1340] = data_i[1340] & sel_one_hot_i[10];
  assign data_masked[1339] = data_i[1339] & sel_one_hot_i[10];
  assign data_masked[1338] = data_i[1338] & sel_one_hot_i[10];
  assign data_masked[1337] = data_i[1337] & sel_one_hot_i[10];
  assign data_masked[1336] = data_i[1336] & sel_one_hot_i[10];
  assign data_masked[1335] = data_i[1335] & sel_one_hot_i[10];
  assign data_masked[1334] = data_i[1334] & sel_one_hot_i[10];
  assign data_masked[1333] = data_i[1333] & sel_one_hot_i[10];
  assign data_masked[1332] = data_i[1332] & sel_one_hot_i[10];
  assign data_masked[1331] = data_i[1331] & sel_one_hot_i[10];
  assign data_masked[1330] = data_i[1330] & sel_one_hot_i[10];
  assign data_masked[1329] = data_i[1329] & sel_one_hot_i[10];
  assign data_masked[1328] = data_i[1328] & sel_one_hot_i[10];
  assign data_masked[1327] = data_i[1327] & sel_one_hot_i[10];
  assign data_masked[1326] = data_i[1326] & sel_one_hot_i[10];
  assign data_masked[1325] = data_i[1325] & sel_one_hot_i[10];
  assign data_masked[1324] = data_i[1324] & sel_one_hot_i[10];
  assign data_masked[1323] = data_i[1323] & sel_one_hot_i[10];
  assign data_masked[1322] = data_i[1322] & sel_one_hot_i[10];
  assign data_masked[1321] = data_i[1321] & sel_one_hot_i[10];
  assign data_masked[1320] = data_i[1320] & sel_one_hot_i[10];
  assign data_masked[1319] = data_i[1319] & sel_one_hot_i[10];
  assign data_masked[1318] = data_i[1318] & sel_one_hot_i[10];
  assign data_masked[1317] = data_i[1317] & sel_one_hot_i[10];
  assign data_masked[1316] = data_i[1316] & sel_one_hot_i[10];
  assign data_masked[1315] = data_i[1315] & sel_one_hot_i[10];
  assign data_masked[1314] = data_i[1314] & sel_one_hot_i[10];
  assign data_masked[1313] = data_i[1313] & sel_one_hot_i[10];
  assign data_masked[1312] = data_i[1312] & sel_one_hot_i[10];
  assign data_masked[1311] = data_i[1311] & sel_one_hot_i[10];
  assign data_masked[1310] = data_i[1310] & sel_one_hot_i[10];
  assign data_masked[1309] = data_i[1309] & sel_one_hot_i[10];
  assign data_masked[1308] = data_i[1308] & sel_one_hot_i[10];
  assign data_masked[1307] = data_i[1307] & sel_one_hot_i[10];
  assign data_masked[1306] = data_i[1306] & sel_one_hot_i[10];
  assign data_masked[1305] = data_i[1305] & sel_one_hot_i[10];
  assign data_masked[1304] = data_i[1304] & sel_one_hot_i[10];
  assign data_masked[1303] = data_i[1303] & sel_one_hot_i[10];
  assign data_masked[1302] = data_i[1302] & sel_one_hot_i[10];
  assign data_masked[1301] = data_i[1301] & sel_one_hot_i[10];
  assign data_masked[1300] = data_i[1300] & sel_one_hot_i[10];
  assign data_masked[1299] = data_i[1299] & sel_one_hot_i[10];
  assign data_masked[1298] = data_i[1298] & sel_one_hot_i[10];
  assign data_masked[1297] = data_i[1297] & sel_one_hot_i[10];
  assign data_masked[1296] = data_i[1296] & sel_one_hot_i[10];
  assign data_masked[1295] = data_i[1295] & sel_one_hot_i[10];
  assign data_masked[1294] = data_i[1294] & sel_one_hot_i[10];
  assign data_masked[1293] = data_i[1293] & sel_one_hot_i[10];
  assign data_masked[1292] = data_i[1292] & sel_one_hot_i[10];
  assign data_masked[1291] = data_i[1291] & sel_one_hot_i[10];
  assign data_masked[1290] = data_i[1290] & sel_one_hot_i[10];
  assign data_masked[1289] = data_i[1289] & sel_one_hot_i[10];
  assign data_masked[1288] = data_i[1288] & sel_one_hot_i[10];
  assign data_masked[1287] = data_i[1287] & sel_one_hot_i[10];
  assign data_masked[1286] = data_i[1286] & sel_one_hot_i[10];
  assign data_masked[1285] = data_i[1285] & sel_one_hot_i[10];
  assign data_masked[1284] = data_i[1284] & sel_one_hot_i[10];
  assign data_masked[1283] = data_i[1283] & sel_one_hot_i[10];
  assign data_masked[1282] = data_i[1282] & sel_one_hot_i[10];
  assign data_masked[1281] = data_i[1281] & sel_one_hot_i[10];
  assign data_masked[1280] = data_i[1280] & sel_one_hot_i[10];
  assign data_masked[1535] = data_i[1535] & sel_one_hot_i[11];
  assign data_masked[1534] = data_i[1534] & sel_one_hot_i[11];
  assign data_masked[1533] = data_i[1533] & sel_one_hot_i[11];
  assign data_masked[1532] = data_i[1532] & sel_one_hot_i[11];
  assign data_masked[1531] = data_i[1531] & sel_one_hot_i[11];
  assign data_masked[1530] = data_i[1530] & sel_one_hot_i[11];
  assign data_masked[1529] = data_i[1529] & sel_one_hot_i[11];
  assign data_masked[1528] = data_i[1528] & sel_one_hot_i[11];
  assign data_masked[1527] = data_i[1527] & sel_one_hot_i[11];
  assign data_masked[1526] = data_i[1526] & sel_one_hot_i[11];
  assign data_masked[1525] = data_i[1525] & sel_one_hot_i[11];
  assign data_masked[1524] = data_i[1524] & sel_one_hot_i[11];
  assign data_masked[1523] = data_i[1523] & sel_one_hot_i[11];
  assign data_masked[1522] = data_i[1522] & sel_one_hot_i[11];
  assign data_masked[1521] = data_i[1521] & sel_one_hot_i[11];
  assign data_masked[1520] = data_i[1520] & sel_one_hot_i[11];
  assign data_masked[1519] = data_i[1519] & sel_one_hot_i[11];
  assign data_masked[1518] = data_i[1518] & sel_one_hot_i[11];
  assign data_masked[1517] = data_i[1517] & sel_one_hot_i[11];
  assign data_masked[1516] = data_i[1516] & sel_one_hot_i[11];
  assign data_masked[1515] = data_i[1515] & sel_one_hot_i[11];
  assign data_masked[1514] = data_i[1514] & sel_one_hot_i[11];
  assign data_masked[1513] = data_i[1513] & sel_one_hot_i[11];
  assign data_masked[1512] = data_i[1512] & sel_one_hot_i[11];
  assign data_masked[1511] = data_i[1511] & sel_one_hot_i[11];
  assign data_masked[1510] = data_i[1510] & sel_one_hot_i[11];
  assign data_masked[1509] = data_i[1509] & sel_one_hot_i[11];
  assign data_masked[1508] = data_i[1508] & sel_one_hot_i[11];
  assign data_masked[1507] = data_i[1507] & sel_one_hot_i[11];
  assign data_masked[1506] = data_i[1506] & sel_one_hot_i[11];
  assign data_masked[1505] = data_i[1505] & sel_one_hot_i[11];
  assign data_masked[1504] = data_i[1504] & sel_one_hot_i[11];
  assign data_masked[1503] = data_i[1503] & sel_one_hot_i[11];
  assign data_masked[1502] = data_i[1502] & sel_one_hot_i[11];
  assign data_masked[1501] = data_i[1501] & sel_one_hot_i[11];
  assign data_masked[1500] = data_i[1500] & sel_one_hot_i[11];
  assign data_masked[1499] = data_i[1499] & sel_one_hot_i[11];
  assign data_masked[1498] = data_i[1498] & sel_one_hot_i[11];
  assign data_masked[1497] = data_i[1497] & sel_one_hot_i[11];
  assign data_masked[1496] = data_i[1496] & sel_one_hot_i[11];
  assign data_masked[1495] = data_i[1495] & sel_one_hot_i[11];
  assign data_masked[1494] = data_i[1494] & sel_one_hot_i[11];
  assign data_masked[1493] = data_i[1493] & sel_one_hot_i[11];
  assign data_masked[1492] = data_i[1492] & sel_one_hot_i[11];
  assign data_masked[1491] = data_i[1491] & sel_one_hot_i[11];
  assign data_masked[1490] = data_i[1490] & sel_one_hot_i[11];
  assign data_masked[1489] = data_i[1489] & sel_one_hot_i[11];
  assign data_masked[1488] = data_i[1488] & sel_one_hot_i[11];
  assign data_masked[1487] = data_i[1487] & sel_one_hot_i[11];
  assign data_masked[1486] = data_i[1486] & sel_one_hot_i[11];
  assign data_masked[1485] = data_i[1485] & sel_one_hot_i[11];
  assign data_masked[1484] = data_i[1484] & sel_one_hot_i[11];
  assign data_masked[1483] = data_i[1483] & sel_one_hot_i[11];
  assign data_masked[1482] = data_i[1482] & sel_one_hot_i[11];
  assign data_masked[1481] = data_i[1481] & sel_one_hot_i[11];
  assign data_masked[1480] = data_i[1480] & sel_one_hot_i[11];
  assign data_masked[1479] = data_i[1479] & sel_one_hot_i[11];
  assign data_masked[1478] = data_i[1478] & sel_one_hot_i[11];
  assign data_masked[1477] = data_i[1477] & sel_one_hot_i[11];
  assign data_masked[1476] = data_i[1476] & sel_one_hot_i[11];
  assign data_masked[1475] = data_i[1475] & sel_one_hot_i[11];
  assign data_masked[1474] = data_i[1474] & sel_one_hot_i[11];
  assign data_masked[1473] = data_i[1473] & sel_one_hot_i[11];
  assign data_masked[1472] = data_i[1472] & sel_one_hot_i[11];
  assign data_masked[1471] = data_i[1471] & sel_one_hot_i[11];
  assign data_masked[1470] = data_i[1470] & sel_one_hot_i[11];
  assign data_masked[1469] = data_i[1469] & sel_one_hot_i[11];
  assign data_masked[1468] = data_i[1468] & sel_one_hot_i[11];
  assign data_masked[1467] = data_i[1467] & sel_one_hot_i[11];
  assign data_masked[1466] = data_i[1466] & sel_one_hot_i[11];
  assign data_masked[1465] = data_i[1465] & sel_one_hot_i[11];
  assign data_masked[1464] = data_i[1464] & sel_one_hot_i[11];
  assign data_masked[1463] = data_i[1463] & sel_one_hot_i[11];
  assign data_masked[1462] = data_i[1462] & sel_one_hot_i[11];
  assign data_masked[1461] = data_i[1461] & sel_one_hot_i[11];
  assign data_masked[1460] = data_i[1460] & sel_one_hot_i[11];
  assign data_masked[1459] = data_i[1459] & sel_one_hot_i[11];
  assign data_masked[1458] = data_i[1458] & sel_one_hot_i[11];
  assign data_masked[1457] = data_i[1457] & sel_one_hot_i[11];
  assign data_masked[1456] = data_i[1456] & sel_one_hot_i[11];
  assign data_masked[1455] = data_i[1455] & sel_one_hot_i[11];
  assign data_masked[1454] = data_i[1454] & sel_one_hot_i[11];
  assign data_masked[1453] = data_i[1453] & sel_one_hot_i[11];
  assign data_masked[1452] = data_i[1452] & sel_one_hot_i[11];
  assign data_masked[1451] = data_i[1451] & sel_one_hot_i[11];
  assign data_masked[1450] = data_i[1450] & sel_one_hot_i[11];
  assign data_masked[1449] = data_i[1449] & sel_one_hot_i[11];
  assign data_masked[1448] = data_i[1448] & sel_one_hot_i[11];
  assign data_masked[1447] = data_i[1447] & sel_one_hot_i[11];
  assign data_masked[1446] = data_i[1446] & sel_one_hot_i[11];
  assign data_masked[1445] = data_i[1445] & sel_one_hot_i[11];
  assign data_masked[1444] = data_i[1444] & sel_one_hot_i[11];
  assign data_masked[1443] = data_i[1443] & sel_one_hot_i[11];
  assign data_masked[1442] = data_i[1442] & sel_one_hot_i[11];
  assign data_masked[1441] = data_i[1441] & sel_one_hot_i[11];
  assign data_masked[1440] = data_i[1440] & sel_one_hot_i[11];
  assign data_masked[1439] = data_i[1439] & sel_one_hot_i[11];
  assign data_masked[1438] = data_i[1438] & sel_one_hot_i[11];
  assign data_masked[1437] = data_i[1437] & sel_one_hot_i[11];
  assign data_masked[1436] = data_i[1436] & sel_one_hot_i[11];
  assign data_masked[1435] = data_i[1435] & sel_one_hot_i[11];
  assign data_masked[1434] = data_i[1434] & sel_one_hot_i[11];
  assign data_masked[1433] = data_i[1433] & sel_one_hot_i[11];
  assign data_masked[1432] = data_i[1432] & sel_one_hot_i[11];
  assign data_masked[1431] = data_i[1431] & sel_one_hot_i[11];
  assign data_masked[1430] = data_i[1430] & sel_one_hot_i[11];
  assign data_masked[1429] = data_i[1429] & sel_one_hot_i[11];
  assign data_masked[1428] = data_i[1428] & sel_one_hot_i[11];
  assign data_masked[1427] = data_i[1427] & sel_one_hot_i[11];
  assign data_masked[1426] = data_i[1426] & sel_one_hot_i[11];
  assign data_masked[1425] = data_i[1425] & sel_one_hot_i[11];
  assign data_masked[1424] = data_i[1424] & sel_one_hot_i[11];
  assign data_masked[1423] = data_i[1423] & sel_one_hot_i[11];
  assign data_masked[1422] = data_i[1422] & sel_one_hot_i[11];
  assign data_masked[1421] = data_i[1421] & sel_one_hot_i[11];
  assign data_masked[1420] = data_i[1420] & sel_one_hot_i[11];
  assign data_masked[1419] = data_i[1419] & sel_one_hot_i[11];
  assign data_masked[1418] = data_i[1418] & sel_one_hot_i[11];
  assign data_masked[1417] = data_i[1417] & sel_one_hot_i[11];
  assign data_masked[1416] = data_i[1416] & sel_one_hot_i[11];
  assign data_masked[1415] = data_i[1415] & sel_one_hot_i[11];
  assign data_masked[1414] = data_i[1414] & sel_one_hot_i[11];
  assign data_masked[1413] = data_i[1413] & sel_one_hot_i[11];
  assign data_masked[1412] = data_i[1412] & sel_one_hot_i[11];
  assign data_masked[1411] = data_i[1411] & sel_one_hot_i[11];
  assign data_masked[1410] = data_i[1410] & sel_one_hot_i[11];
  assign data_masked[1409] = data_i[1409] & sel_one_hot_i[11];
  assign data_masked[1408] = data_i[1408] & sel_one_hot_i[11];
  assign data_masked[1663] = data_i[1663] & sel_one_hot_i[12];
  assign data_masked[1662] = data_i[1662] & sel_one_hot_i[12];
  assign data_masked[1661] = data_i[1661] & sel_one_hot_i[12];
  assign data_masked[1660] = data_i[1660] & sel_one_hot_i[12];
  assign data_masked[1659] = data_i[1659] & sel_one_hot_i[12];
  assign data_masked[1658] = data_i[1658] & sel_one_hot_i[12];
  assign data_masked[1657] = data_i[1657] & sel_one_hot_i[12];
  assign data_masked[1656] = data_i[1656] & sel_one_hot_i[12];
  assign data_masked[1655] = data_i[1655] & sel_one_hot_i[12];
  assign data_masked[1654] = data_i[1654] & sel_one_hot_i[12];
  assign data_masked[1653] = data_i[1653] & sel_one_hot_i[12];
  assign data_masked[1652] = data_i[1652] & sel_one_hot_i[12];
  assign data_masked[1651] = data_i[1651] & sel_one_hot_i[12];
  assign data_masked[1650] = data_i[1650] & sel_one_hot_i[12];
  assign data_masked[1649] = data_i[1649] & sel_one_hot_i[12];
  assign data_masked[1648] = data_i[1648] & sel_one_hot_i[12];
  assign data_masked[1647] = data_i[1647] & sel_one_hot_i[12];
  assign data_masked[1646] = data_i[1646] & sel_one_hot_i[12];
  assign data_masked[1645] = data_i[1645] & sel_one_hot_i[12];
  assign data_masked[1644] = data_i[1644] & sel_one_hot_i[12];
  assign data_masked[1643] = data_i[1643] & sel_one_hot_i[12];
  assign data_masked[1642] = data_i[1642] & sel_one_hot_i[12];
  assign data_masked[1641] = data_i[1641] & sel_one_hot_i[12];
  assign data_masked[1640] = data_i[1640] & sel_one_hot_i[12];
  assign data_masked[1639] = data_i[1639] & sel_one_hot_i[12];
  assign data_masked[1638] = data_i[1638] & sel_one_hot_i[12];
  assign data_masked[1637] = data_i[1637] & sel_one_hot_i[12];
  assign data_masked[1636] = data_i[1636] & sel_one_hot_i[12];
  assign data_masked[1635] = data_i[1635] & sel_one_hot_i[12];
  assign data_masked[1634] = data_i[1634] & sel_one_hot_i[12];
  assign data_masked[1633] = data_i[1633] & sel_one_hot_i[12];
  assign data_masked[1632] = data_i[1632] & sel_one_hot_i[12];
  assign data_masked[1631] = data_i[1631] & sel_one_hot_i[12];
  assign data_masked[1630] = data_i[1630] & sel_one_hot_i[12];
  assign data_masked[1629] = data_i[1629] & sel_one_hot_i[12];
  assign data_masked[1628] = data_i[1628] & sel_one_hot_i[12];
  assign data_masked[1627] = data_i[1627] & sel_one_hot_i[12];
  assign data_masked[1626] = data_i[1626] & sel_one_hot_i[12];
  assign data_masked[1625] = data_i[1625] & sel_one_hot_i[12];
  assign data_masked[1624] = data_i[1624] & sel_one_hot_i[12];
  assign data_masked[1623] = data_i[1623] & sel_one_hot_i[12];
  assign data_masked[1622] = data_i[1622] & sel_one_hot_i[12];
  assign data_masked[1621] = data_i[1621] & sel_one_hot_i[12];
  assign data_masked[1620] = data_i[1620] & sel_one_hot_i[12];
  assign data_masked[1619] = data_i[1619] & sel_one_hot_i[12];
  assign data_masked[1618] = data_i[1618] & sel_one_hot_i[12];
  assign data_masked[1617] = data_i[1617] & sel_one_hot_i[12];
  assign data_masked[1616] = data_i[1616] & sel_one_hot_i[12];
  assign data_masked[1615] = data_i[1615] & sel_one_hot_i[12];
  assign data_masked[1614] = data_i[1614] & sel_one_hot_i[12];
  assign data_masked[1613] = data_i[1613] & sel_one_hot_i[12];
  assign data_masked[1612] = data_i[1612] & sel_one_hot_i[12];
  assign data_masked[1611] = data_i[1611] & sel_one_hot_i[12];
  assign data_masked[1610] = data_i[1610] & sel_one_hot_i[12];
  assign data_masked[1609] = data_i[1609] & sel_one_hot_i[12];
  assign data_masked[1608] = data_i[1608] & sel_one_hot_i[12];
  assign data_masked[1607] = data_i[1607] & sel_one_hot_i[12];
  assign data_masked[1606] = data_i[1606] & sel_one_hot_i[12];
  assign data_masked[1605] = data_i[1605] & sel_one_hot_i[12];
  assign data_masked[1604] = data_i[1604] & sel_one_hot_i[12];
  assign data_masked[1603] = data_i[1603] & sel_one_hot_i[12];
  assign data_masked[1602] = data_i[1602] & sel_one_hot_i[12];
  assign data_masked[1601] = data_i[1601] & sel_one_hot_i[12];
  assign data_masked[1600] = data_i[1600] & sel_one_hot_i[12];
  assign data_masked[1599] = data_i[1599] & sel_one_hot_i[12];
  assign data_masked[1598] = data_i[1598] & sel_one_hot_i[12];
  assign data_masked[1597] = data_i[1597] & sel_one_hot_i[12];
  assign data_masked[1596] = data_i[1596] & sel_one_hot_i[12];
  assign data_masked[1595] = data_i[1595] & sel_one_hot_i[12];
  assign data_masked[1594] = data_i[1594] & sel_one_hot_i[12];
  assign data_masked[1593] = data_i[1593] & sel_one_hot_i[12];
  assign data_masked[1592] = data_i[1592] & sel_one_hot_i[12];
  assign data_masked[1591] = data_i[1591] & sel_one_hot_i[12];
  assign data_masked[1590] = data_i[1590] & sel_one_hot_i[12];
  assign data_masked[1589] = data_i[1589] & sel_one_hot_i[12];
  assign data_masked[1588] = data_i[1588] & sel_one_hot_i[12];
  assign data_masked[1587] = data_i[1587] & sel_one_hot_i[12];
  assign data_masked[1586] = data_i[1586] & sel_one_hot_i[12];
  assign data_masked[1585] = data_i[1585] & sel_one_hot_i[12];
  assign data_masked[1584] = data_i[1584] & sel_one_hot_i[12];
  assign data_masked[1583] = data_i[1583] & sel_one_hot_i[12];
  assign data_masked[1582] = data_i[1582] & sel_one_hot_i[12];
  assign data_masked[1581] = data_i[1581] & sel_one_hot_i[12];
  assign data_masked[1580] = data_i[1580] & sel_one_hot_i[12];
  assign data_masked[1579] = data_i[1579] & sel_one_hot_i[12];
  assign data_masked[1578] = data_i[1578] & sel_one_hot_i[12];
  assign data_masked[1577] = data_i[1577] & sel_one_hot_i[12];
  assign data_masked[1576] = data_i[1576] & sel_one_hot_i[12];
  assign data_masked[1575] = data_i[1575] & sel_one_hot_i[12];
  assign data_masked[1574] = data_i[1574] & sel_one_hot_i[12];
  assign data_masked[1573] = data_i[1573] & sel_one_hot_i[12];
  assign data_masked[1572] = data_i[1572] & sel_one_hot_i[12];
  assign data_masked[1571] = data_i[1571] & sel_one_hot_i[12];
  assign data_masked[1570] = data_i[1570] & sel_one_hot_i[12];
  assign data_masked[1569] = data_i[1569] & sel_one_hot_i[12];
  assign data_masked[1568] = data_i[1568] & sel_one_hot_i[12];
  assign data_masked[1567] = data_i[1567] & sel_one_hot_i[12];
  assign data_masked[1566] = data_i[1566] & sel_one_hot_i[12];
  assign data_masked[1565] = data_i[1565] & sel_one_hot_i[12];
  assign data_masked[1564] = data_i[1564] & sel_one_hot_i[12];
  assign data_masked[1563] = data_i[1563] & sel_one_hot_i[12];
  assign data_masked[1562] = data_i[1562] & sel_one_hot_i[12];
  assign data_masked[1561] = data_i[1561] & sel_one_hot_i[12];
  assign data_masked[1560] = data_i[1560] & sel_one_hot_i[12];
  assign data_masked[1559] = data_i[1559] & sel_one_hot_i[12];
  assign data_masked[1558] = data_i[1558] & sel_one_hot_i[12];
  assign data_masked[1557] = data_i[1557] & sel_one_hot_i[12];
  assign data_masked[1556] = data_i[1556] & sel_one_hot_i[12];
  assign data_masked[1555] = data_i[1555] & sel_one_hot_i[12];
  assign data_masked[1554] = data_i[1554] & sel_one_hot_i[12];
  assign data_masked[1553] = data_i[1553] & sel_one_hot_i[12];
  assign data_masked[1552] = data_i[1552] & sel_one_hot_i[12];
  assign data_masked[1551] = data_i[1551] & sel_one_hot_i[12];
  assign data_masked[1550] = data_i[1550] & sel_one_hot_i[12];
  assign data_masked[1549] = data_i[1549] & sel_one_hot_i[12];
  assign data_masked[1548] = data_i[1548] & sel_one_hot_i[12];
  assign data_masked[1547] = data_i[1547] & sel_one_hot_i[12];
  assign data_masked[1546] = data_i[1546] & sel_one_hot_i[12];
  assign data_masked[1545] = data_i[1545] & sel_one_hot_i[12];
  assign data_masked[1544] = data_i[1544] & sel_one_hot_i[12];
  assign data_masked[1543] = data_i[1543] & sel_one_hot_i[12];
  assign data_masked[1542] = data_i[1542] & sel_one_hot_i[12];
  assign data_masked[1541] = data_i[1541] & sel_one_hot_i[12];
  assign data_masked[1540] = data_i[1540] & sel_one_hot_i[12];
  assign data_masked[1539] = data_i[1539] & sel_one_hot_i[12];
  assign data_masked[1538] = data_i[1538] & sel_one_hot_i[12];
  assign data_masked[1537] = data_i[1537] & sel_one_hot_i[12];
  assign data_masked[1536] = data_i[1536] & sel_one_hot_i[12];
  assign data_masked[1791] = data_i[1791] & sel_one_hot_i[13];
  assign data_masked[1790] = data_i[1790] & sel_one_hot_i[13];
  assign data_masked[1789] = data_i[1789] & sel_one_hot_i[13];
  assign data_masked[1788] = data_i[1788] & sel_one_hot_i[13];
  assign data_masked[1787] = data_i[1787] & sel_one_hot_i[13];
  assign data_masked[1786] = data_i[1786] & sel_one_hot_i[13];
  assign data_masked[1785] = data_i[1785] & sel_one_hot_i[13];
  assign data_masked[1784] = data_i[1784] & sel_one_hot_i[13];
  assign data_masked[1783] = data_i[1783] & sel_one_hot_i[13];
  assign data_masked[1782] = data_i[1782] & sel_one_hot_i[13];
  assign data_masked[1781] = data_i[1781] & sel_one_hot_i[13];
  assign data_masked[1780] = data_i[1780] & sel_one_hot_i[13];
  assign data_masked[1779] = data_i[1779] & sel_one_hot_i[13];
  assign data_masked[1778] = data_i[1778] & sel_one_hot_i[13];
  assign data_masked[1777] = data_i[1777] & sel_one_hot_i[13];
  assign data_masked[1776] = data_i[1776] & sel_one_hot_i[13];
  assign data_masked[1775] = data_i[1775] & sel_one_hot_i[13];
  assign data_masked[1774] = data_i[1774] & sel_one_hot_i[13];
  assign data_masked[1773] = data_i[1773] & sel_one_hot_i[13];
  assign data_masked[1772] = data_i[1772] & sel_one_hot_i[13];
  assign data_masked[1771] = data_i[1771] & sel_one_hot_i[13];
  assign data_masked[1770] = data_i[1770] & sel_one_hot_i[13];
  assign data_masked[1769] = data_i[1769] & sel_one_hot_i[13];
  assign data_masked[1768] = data_i[1768] & sel_one_hot_i[13];
  assign data_masked[1767] = data_i[1767] & sel_one_hot_i[13];
  assign data_masked[1766] = data_i[1766] & sel_one_hot_i[13];
  assign data_masked[1765] = data_i[1765] & sel_one_hot_i[13];
  assign data_masked[1764] = data_i[1764] & sel_one_hot_i[13];
  assign data_masked[1763] = data_i[1763] & sel_one_hot_i[13];
  assign data_masked[1762] = data_i[1762] & sel_one_hot_i[13];
  assign data_masked[1761] = data_i[1761] & sel_one_hot_i[13];
  assign data_masked[1760] = data_i[1760] & sel_one_hot_i[13];
  assign data_masked[1759] = data_i[1759] & sel_one_hot_i[13];
  assign data_masked[1758] = data_i[1758] & sel_one_hot_i[13];
  assign data_masked[1757] = data_i[1757] & sel_one_hot_i[13];
  assign data_masked[1756] = data_i[1756] & sel_one_hot_i[13];
  assign data_masked[1755] = data_i[1755] & sel_one_hot_i[13];
  assign data_masked[1754] = data_i[1754] & sel_one_hot_i[13];
  assign data_masked[1753] = data_i[1753] & sel_one_hot_i[13];
  assign data_masked[1752] = data_i[1752] & sel_one_hot_i[13];
  assign data_masked[1751] = data_i[1751] & sel_one_hot_i[13];
  assign data_masked[1750] = data_i[1750] & sel_one_hot_i[13];
  assign data_masked[1749] = data_i[1749] & sel_one_hot_i[13];
  assign data_masked[1748] = data_i[1748] & sel_one_hot_i[13];
  assign data_masked[1747] = data_i[1747] & sel_one_hot_i[13];
  assign data_masked[1746] = data_i[1746] & sel_one_hot_i[13];
  assign data_masked[1745] = data_i[1745] & sel_one_hot_i[13];
  assign data_masked[1744] = data_i[1744] & sel_one_hot_i[13];
  assign data_masked[1743] = data_i[1743] & sel_one_hot_i[13];
  assign data_masked[1742] = data_i[1742] & sel_one_hot_i[13];
  assign data_masked[1741] = data_i[1741] & sel_one_hot_i[13];
  assign data_masked[1740] = data_i[1740] & sel_one_hot_i[13];
  assign data_masked[1739] = data_i[1739] & sel_one_hot_i[13];
  assign data_masked[1738] = data_i[1738] & sel_one_hot_i[13];
  assign data_masked[1737] = data_i[1737] & sel_one_hot_i[13];
  assign data_masked[1736] = data_i[1736] & sel_one_hot_i[13];
  assign data_masked[1735] = data_i[1735] & sel_one_hot_i[13];
  assign data_masked[1734] = data_i[1734] & sel_one_hot_i[13];
  assign data_masked[1733] = data_i[1733] & sel_one_hot_i[13];
  assign data_masked[1732] = data_i[1732] & sel_one_hot_i[13];
  assign data_masked[1731] = data_i[1731] & sel_one_hot_i[13];
  assign data_masked[1730] = data_i[1730] & sel_one_hot_i[13];
  assign data_masked[1729] = data_i[1729] & sel_one_hot_i[13];
  assign data_masked[1728] = data_i[1728] & sel_one_hot_i[13];
  assign data_masked[1727] = data_i[1727] & sel_one_hot_i[13];
  assign data_masked[1726] = data_i[1726] & sel_one_hot_i[13];
  assign data_masked[1725] = data_i[1725] & sel_one_hot_i[13];
  assign data_masked[1724] = data_i[1724] & sel_one_hot_i[13];
  assign data_masked[1723] = data_i[1723] & sel_one_hot_i[13];
  assign data_masked[1722] = data_i[1722] & sel_one_hot_i[13];
  assign data_masked[1721] = data_i[1721] & sel_one_hot_i[13];
  assign data_masked[1720] = data_i[1720] & sel_one_hot_i[13];
  assign data_masked[1719] = data_i[1719] & sel_one_hot_i[13];
  assign data_masked[1718] = data_i[1718] & sel_one_hot_i[13];
  assign data_masked[1717] = data_i[1717] & sel_one_hot_i[13];
  assign data_masked[1716] = data_i[1716] & sel_one_hot_i[13];
  assign data_masked[1715] = data_i[1715] & sel_one_hot_i[13];
  assign data_masked[1714] = data_i[1714] & sel_one_hot_i[13];
  assign data_masked[1713] = data_i[1713] & sel_one_hot_i[13];
  assign data_masked[1712] = data_i[1712] & sel_one_hot_i[13];
  assign data_masked[1711] = data_i[1711] & sel_one_hot_i[13];
  assign data_masked[1710] = data_i[1710] & sel_one_hot_i[13];
  assign data_masked[1709] = data_i[1709] & sel_one_hot_i[13];
  assign data_masked[1708] = data_i[1708] & sel_one_hot_i[13];
  assign data_masked[1707] = data_i[1707] & sel_one_hot_i[13];
  assign data_masked[1706] = data_i[1706] & sel_one_hot_i[13];
  assign data_masked[1705] = data_i[1705] & sel_one_hot_i[13];
  assign data_masked[1704] = data_i[1704] & sel_one_hot_i[13];
  assign data_masked[1703] = data_i[1703] & sel_one_hot_i[13];
  assign data_masked[1702] = data_i[1702] & sel_one_hot_i[13];
  assign data_masked[1701] = data_i[1701] & sel_one_hot_i[13];
  assign data_masked[1700] = data_i[1700] & sel_one_hot_i[13];
  assign data_masked[1699] = data_i[1699] & sel_one_hot_i[13];
  assign data_masked[1698] = data_i[1698] & sel_one_hot_i[13];
  assign data_masked[1697] = data_i[1697] & sel_one_hot_i[13];
  assign data_masked[1696] = data_i[1696] & sel_one_hot_i[13];
  assign data_masked[1695] = data_i[1695] & sel_one_hot_i[13];
  assign data_masked[1694] = data_i[1694] & sel_one_hot_i[13];
  assign data_masked[1693] = data_i[1693] & sel_one_hot_i[13];
  assign data_masked[1692] = data_i[1692] & sel_one_hot_i[13];
  assign data_masked[1691] = data_i[1691] & sel_one_hot_i[13];
  assign data_masked[1690] = data_i[1690] & sel_one_hot_i[13];
  assign data_masked[1689] = data_i[1689] & sel_one_hot_i[13];
  assign data_masked[1688] = data_i[1688] & sel_one_hot_i[13];
  assign data_masked[1687] = data_i[1687] & sel_one_hot_i[13];
  assign data_masked[1686] = data_i[1686] & sel_one_hot_i[13];
  assign data_masked[1685] = data_i[1685] & sel_one_hot_i[13];
  assign data_masked[1684] = data_i[1684] & sel_one_hot_i[13];
  assign data_masked[1683] = data_i[1683] & sel_one_hot_i[13];
  assign data_masked[1682] = data_i[1682] & sel_one_hot_i[13];
  assign data_masked[1681] = data_i[1681] & sel_one_hot_i[13];
  assign data_masked[1680] = data_i[1680] & sel_one_hot_i[13];
  assign data_masked[1679] = data_i[1679] & sel_one_hot_i[13];
  assign data_masked[1678] = data_i[1678] & sel_one_hot_i[13];
  assign data_masked[1677] = data_i[1677] & sel_one_hot_i[13];
  assign data_masked[1676] = data_i[1676] & sel_one_hot_i[13];
  assign data_masked[1675] = data_i[1675] & sel_one_hot_i[13];
  assign data_masked[1674] = data_i[1674] & sel_one_hot_i[13];
  assign data_masked[1673] = data_i[1673] & sel_one_hot_i[13];
  assign data_masked[1672] = data_i[1672] & sel_one_hot_i[13];
  assign data_masked[1671] = data_i[1671] & sel_one_hot_i[13];
  assign data_masked[1670] = data_i[1670] & sel_one_hot_i[13];
  assign data_masked[1669] = data_i[1669] & sel_one_hot_i[13];
  assign data_masked[1668] = data_i[1668] & sel_one_hot_i[13];
  assign data_masked[1667] = data_i[1667] & sel_one_hot_i[13];
  assign data_masked[1666] = data_i[1666] & sel_one_hot_i[13];
  assign data_masked[1665] = data_i[1665] & sel_one_hot_i[13];
  assign data_masked[1664] = data_i[1664] & sel_one_hot_i[13];
  assign data_masked[1919] = data_i[1919] & sel_one_hot_i[14];
  assign data_masked[1918] = data_i[1918] & sel_one_hot_i[14];
  assign data_masked[1917] = data_i[1917] & sel_one_hot_i[14];
  assign data_masked[1916] = data_i[1916] & sel_one_hot_i[14];
  assign data_masked[1915] = data_i[1915] & sel_one_hot_i[14];
  assign data_masked[1914] = data_i[1914] & sel_one_hot_i[14];
  assign data_masked[1913] = data_i[1913] & sel_one_hot_i[14];
  assign data_masked[1912] = data_i[1912] & sel_one_hot_i[14];
  assign data_masked[1911] = data_i[1911] & sel_one_hot_i[14];
  assign data_masked[1910] = data_i[1910] & sel_one_hot_i[14];
  assign data_masked[1909] = data_i[1909] & sel_one_hot_i[14];
  assign data_masked[1908] = data_i[1908] & sel_one_hot_i[14];
  assign data_masked[1907] = data_i[1907] & sel_one_hot_i[14];
  assign data_masked[1906] = data_i[1906] & sel_one_hot_i[14];
  assign data_masked[1905] = data_i[1905] & sel_one_hot_i[14];
  assign data_masked[1904] = data_i[1904] & sel_one_hot_i[14];
  assign data_masked[1903] = data_i[1903] & sel_one_hot_i[14];
  assign data_masked[1902] = data_i[1902] & sel_one_hot_i[14];
  assign data_masked[1901] = data_i[1901] & sel_one_hot_i[14];
  assign data_masked[1900] = data_i[1900] & sel_one_hot_i[14];
  assign data_masked[1899] = data_i[1899] & sel_one_hot_i[14];
  assign data_masked[1898] = data_i[1898] & sel_one_hot_i[14];
  assign data_masked[1897] = data_i[1897] & sel_one_hot_i[14];
  assign data_masked[1896] = data_i[1896] & sel_one_hot_i[14];
  assign data_masked[1895] = data_i[1895] & sel_one_hot_i[14];
  assign data_masked[1894] = data_i[1894] & sel_one_hot_i[14];
  assign data_masked[1893] = data_i[1893] & sel_one_hot_i[14];
  assign data_masked[1892] = data_i[1892] & sel_one_hot_i[14];
  assign data_masked[1891] = data_i[1891] & sel_one_hot_i[14];
  assign data_masked[1890] = data_i[1890] & sel_one_hot_i[14];
  assign data_masked[1889] = data_i[1889] & sel_one_hot_i[14];
  assign data_masked[1888] = data_i[1888] & sel_one_hot_i[14];
  assign data_masked[1887] = data_i[1887] & sel_one_hot_i[14];
  assign data_masked[1886] = data_i[1886] & sel_one_hot_i[14];
  assign data_masked[1885] = data_i[1885] & sel_one_hot_i[14];
  assign data_masked[1884] = data_i[1884] & sel_one_hot_i[14];
  assign data_masked[1883] = data_i[1883] & sel_one_hot_i[14];
  assign data_masked[1882] = data_i[1882] & sel_one_hot_i[14];
  assign data_masked[1881] = data_i[1881] & sel_one_hot_i[14];
  assign data_masked[1880] = data_i[1880] & sel_one_hot_i[14];
  assign data_masked[1879] = data_i[1879] & sel_one_hot_i[14];
  assign data_masked[1878] = data_i[1878] & sel_one_hot_i[14];
  assign data_masked[1877] = data_i[1877] & sel_one_hot_i[14];
  assign data_masked[1876] = data_i[1876] & sel_one_hot_i[14];
  assign data_masked[1875] = data_i[1875] & sel_one_hot_i[14];
  assign data_masked[1874] = data_i[1874] & sel_one_hot_i[14];
  assign data_masked[1873] = data_i[1873] & sel_one_hot_i[14];
  assign data_masked[1872] = data_i[1872] & sel_one_hot_i[14];
  assign data_masked[1871] = data_i[1871] & sel_one_hot_i[14];
  assign data_masked[1870] = data_i[1870] & sel_one_hot_i[14];
  assign data_masked[1869] = data_i[1869] & sel_one_hot_i[14];
  assign data_masked[1868] = data_i[1868] & sel_one_hot_i[14];
  assign data_masked[1867] = data_i[1867] & sel_one_hot_i[14];
  assign data_masked[1866] = data_i[1866] & sel_one_hot_i[14];
  assign data_masked[1865] = data_i[1865] & sel_one_hot_i[14];
  assign data_masked[1864] = data_i[1864] & sel_one_hot_i[14];
  assign data_masked[1863] = data_i[1863] & sel_one_hot_i[14];
  assign data_masked[1862] = data_i[1862] & sel_one_hot_i[14];
  assign data_masked[1861] = data_i[1861] & sel_one_hot_i[14];
  assign data_masked[1860] = data_i[1860] & sel_one_hot_i[14];
  assign data_masked[1859] = data_i[1859] & sel_one_hot_i[14];
  assign data_masked[1858] = data_i[1858] & sel_one_hot_i[14];
  assign data_masked[1857] = data_i[1857] & sel_one_hot_i[14];
  assign data_masked[1856] = data_i[1856] & sel_one_hot_i[14];
  assign data_masked[1855] = data_i[1855] & sel_one_hot_i[14];
  assign data_masked[1854] = data_i[1854] & sel_one_hot_i[14];
  assign data_masked[1853] = data_i[1853] & sel_one_hot_i[14];
  assign data_masked[1852] = data_i[1852] & sel_one_hot_i[14];
  assign data_masked[1851] = data_i[1851] & sel_one_hot_i[14];
  assign data_masked[1850] = data_i[1850] & sel_one_hot_i[14];
  assign data_masked[1849] = data_i[1849] & sel_one_hot_i[14];
  assign data_masked[1848] = data_i[1848] & sel_one_hot_i[14];
  assign data_masked[1847] = data_i[1847] & sel_one_hot_i[14];
  assign data_masked[1846] = data_i[1846] & sel_one_hot_i[14];
  assign data_masked[1845] = data_i[1845] & sel_one_hot_i[14];
  assign data_masked[1844] = data_i[1844] & sel_one_hot_i[14];
  assign data_masked[1843] = data_i[1843] & sel_one_hot_i[14];
  assign data_masked[1842] = data_i[1842] & sel_one_hot_i[14];
  assign data_masked[1841] = data_i[1841] & sel_one_hot_i[14];
  assign data_masked[1840] = data_i[1840] & sel_one_hot_i[14];
  assign data_masked[1839] = data_i[1839] & sel_one_hot_i[14];
  assign data_masked[1838] = data_i[1838] & sel_one_hot_i[14];
  assign data_masked[1837] = data_i[1837] & sel_one_hot_i[14];
  assign data_masked[1836] = data_i[1836] & sel_one_hot_i[14];
  assign data_masked[1835] = data_i[1835] & sel_one_hot_i[14];
  assign data_masked[1834] = data_i[1834] & sel_one_hot_i[14];
  assign data_masked[1833] = data_i[1833] & sel_one_hot_i[14];
  assign data_masked[1832] = data_i[1832] & sel_one_hot_i[14];
  assign data_masked[1831] = data_i[1831] & sel_one_hot_i[14];
  assign data_masked[1830] = data_i[1830] & sel_one_hot_i[14];
  assign data_masked[1829] = data_i[1829] & sel_one_hot_i[14];
  assign data_masked[1828] = data_i[1828] & sel_one_hot_i[14];
  assign data_masked[1827] = data_i[1827] & sel_one_hot_i[14];
  assign data_masked[1826] = data_i[1826] & sel_one_hot_i[14];
  assign data_masked[1825] = data_i[1825] & sel_one_hot_i[14];
  assign data_masked[1824] = data_i[1824] & sel_one_hot_i[14];
  assign data_masked[1823] = data_i[1823] & sel_one_hot_i[14];
  assign data_masked[1822] = data_i[1822] & sel_one_hot_i[14];
  assign data_masked[1821] = data_i[1821] & sel_one_hot_i[14];
  assign data_masked[1820] = data_i[1820] & sel_one_hot_i[14];
  assign data_masked[1819] = data_i[1819] & sel_one_hot_i[14];
  assign data_masked[1818] = data_i[1818] & sel_one_hot_i[14];
  assign data_masked[1817] = data_i[1817] & sel_one_hot_i[14];
  assign data_masked[1816] = data_i[1816] & sel_one_hot_i[14];
  assign data_masked[1815] = data_i[1815] & sel_one_hot_i[14];
  assign data_masked[1814] = data_i[1814] & sel_one_hot_i[14];
  assign data_masked[1813] = data_i[1813] & sel_one_hot_i[14];
  assign data_masked[1812] = data_i[1812] & sel_one_hot_i[14];
  assign data_masked[1811] = data_i[1811] & sel_one_hot_i[14];
  assign data_masked[1810] = data_i[1810] & sel_one_hot_i[14];
  assign data_masked[1809] = data_i[1809] & sel_one_hot_i[14];
  assign data_masked[1808] = data_i[1808] & sel_one_hot_i[14];
  assign data_masked[1807] = data_i[1807] & sel_one_hot_i[14];
  assign data_masked[1806] = data_i[1806] & sel_one_hot_i[14];
  assign data_masked[1805] = data_i[1805] & sel_one_hot_i[14];
  assign data_masked[1804] = data_i[1804] & sel_one_hot_i[14];
  assign data_masked[1803] = data_i[1803] & sel_one_hot_i[14];
  assign data_masked[1802] = data_i[1802] & sel_one_hot_i[14];
  assign data_masked[1801] = data_i[1801] & sel_one_hot_i[14];
  assign data_masked[1800] = data_i[1800] & sel_one_hot_i[14];
  assign data_masked[1799] = data_i[1799] & sel_one_hot_i[14];
  assign data_masked[1798] = data_i[1798] & sel_one_hot_i[14];
  assign data_masked[1797] = data_i[1797] & sel_one_hot_i[14];
  assign data_masked[1796] = data_i[1796] & sel_one_hot_i[14];
  assign data_masked[1795] = data_i[1795] & sel_one_hot_i[14];
  assign data_masked[1794] = data_i[1794] & sel_one_hot_i[14];
  assign data_masked[1793] = data_i[1793] & sel_one_hot_i[14];
  assign data_masked[1792] = data_i[1792] & sel_one_hot_i[14];
  assign data_masked[2047] = data_i[2047] & sel_one_hot_i[15];
  assign data_masked[2046] = data_i[2046] & sel_one_hot_i[15];
  assign data_masked[2045] = data_i[2045] & sel_one_hot_i[15];
  assign data_masked[2044] = data_i[2044] & sel_one_hot_i[15];
  assign data_masked[2043] = data_i[2043] & sel_one_hot_i[15];
  assign data_masked[2042] = data_i[2042] & sel_one_hot_i[15];
  assign data_masked[2041] = data_i[2041] & sel_one_hot_i[15];
  assign data_masked[2040] = data_i[2040] & sel_one_hot_i[15];
  assign data_masked[2039] = data_i[2039] & sel_one_hot_i[15];
  assign data_masked[2038] = data_i[2038] & sel_one_hot_i[15];
  assign data_masked[2037] = data_i[2037] & sel_one_hot_i[15];
  assign data_masked[2036] = data_i[2036] & sel_one_hot_i[15];
  assign data_masked[2035] = data_i[2035] & sel_one_hot_i[15];
  assign data_masked[2034] = data_i[2034] & sel_one_hot_i[15];
  assign data_masked[2033] = data_i[2033] & sel_one_hot_i[15];
  assign data_masked[2032] = data_i[2032] & sel_one_hot_i[15];
  assign data_masked[2031] = data_i[2031] & sel_one_hot_i[15];
  assign data_masked[2030] = data_i[2030] & sel_one_hot_i[15];
  assign data_masked[2029] = data_i[2029] & sel_one_hot_i[15];
  assign data_masked[2028] = data_i[2028] & sel_one_hot_i[15];
  assign data_masked[2027] = data_i[2027] & sel_one_hot_i[15];
  assign data_masked[2026] = data_i[2026] & sel_one_hot_i[15];
  assign data_masked[2025] = data_i[2025] & sel_one_hot_i[15];
  assign data_masked[2024] = data_i[2024] & sel_one_hot_i[15];
  assign data_masked[2023] = data_i[2023] & sel_one_hot_i[15];
  assign data_masked[2022] = data_i[2022] & sel_one_hot_i[15];
  assign data_masked[2021] = data_i[2021] & sel_one_hot_i[15];
  assign data_masked[2020] = data_i[2020] & sel_one_hot_i[15];
  assign data_masked[2019] = data_i[2019] & sel_one_hot_i[15];
  assign data_masked[2018] = data_i[2018] & sel_one_hot_i[15];
  assign data_masked[2017] = data_i[2017] & sel_one_hot_i[15];
  assign data_masked[2016] = data_i[2016] & sel_one_hot_i[15];
  assign data_masked[2015] = data_i[2015] & sel_one_hot_i[15];
  assign data_masked[2014] = data_i[2014] & sel_one_hot_i[15];
  assign data_masked[2013] = data_i[2013] & sel_one_hot_i[15];
  assign data_masked[2012] = data_i[2012] & sel_one_hot_i[15];
  assign data_masked[2011] = data_i[2011] & sel_one_hot_i[15];
  assign data_masked[2010] = data_i[2010] & sel_one_hot_i[15];
  assign data_masked[2009] = data_i[2009] & sel_one_hot_i[15];
  assign data_masked[2008] = data_i[2008] & sel_one_hot_i[15];
  assign data_masked[2007] = data_i[2007] & sel_one_hot_i[15];
  assign data_masked[2006] = data_i[2006] & sel_one_hot_i[15];
  assign data_masked[2005] = data_i[2005] & sel_one_hot_i[15];
  assign data_masked[2004] = data_i[2004] & sel_one_hot_i[15];
  assign data_masked[2003] = data_i[2003] & sel_one_hot_i[15];
  assign data_masked[2002] = data_i[2002] & sel_one_hot_i[15];
  assign data_masked[2001] = data_i[2001] & sel_one_hot_i[15];
  assign data_masked[2000] = data_i[2000] & sel_one_hot_i[15];
  assign data_masked[1999] = data_i[1999] & sel_one_hot_i[15];
  assign data_masked[1998] = data_i[1998] & sel_one_hot_i[15];
  assign data_masked[1997] = data_i[1997] & sel_one_hot_i[15];
  assign data_masked[1996] = data_i[1996] & sel_one_hot_i[15];
  assign data_masked[1995] = data_i[1995] & sel_one_hot_i[15];
  assign data_masked[1994] = data_i[1994] & sel_one_hot_i[15];
  assign data_masked[1993] = data_i[1993] & sel_one_hot_i[15];
  assign data_masked[1992] = data_i[1992] & sel_one_hot_i[15];
  assign data_masked[1991] = data_i[1991] & sel_one_hot_i[15];
  assign data_masked[1990] = data_i[1990] & sel_one_hot_i[15];
  assign data_masked[1989] = data_i[1989] & sel_one_hot_i[15];
  assign data_masked[1988] = data_i[1988] & sel_one_hot_i[15];
  assign data_masked[1987] = data_i[1987] & sel_one_hot_i[15];
  assign data_masked[1986] = data_i[1986] & sel_one_hot_i[15];
  assign data_masked[1985] = data_i[1985] & sel_one_hot_i[15];
  assign data_masked[1984] = data_i[1984] & sel_one_hot_i[15];
  assign data_masked[1983] = data_i[1983] & sel_one_hot_i[15];
  assign data_masked[1982] = data_i[1982] & sel_one_hot_i[15];
  assign data_masked[1981] = data_i[1981] & sel_one_hot_i[15];
  assign data_masked[1980] = data_i[1980] & sel_one_hot_i[15];
  assign data_masked[1979] = data_i[1979] & sel_one_hot_i[15];
  assign data_masked[1978] = data_i[1978] & sel_one_hot_i[15];
  assign data_masked[1977] = data_i[1977] & sel_one_hot_i[15];
  assign data_masked[1976] = data_i[1976] & sel_one_hot_i[15];
  assign data_masked[1975] = data_i[1975] & sel_one_hot_i[15];
  assign data_masked[1974] = data_i[1974] & sel_one_hot_i[15];
  assign data_masked[1973] = data_i[1973] & sel_one_hot_i[15];
  assign data_masked[1972] = data_i[1972] & sel_one_hot_i[15];
  assign data_masked[1971] = data_i[1971] & sel_one_hot_i[15];
  assign data_masked[1970] = data_i[1970] & sel_one_hot_i[15];
  assign data_masked[1969] = data_i[1969] & sel_one_hot_i[15];
  assign data_masked[1968] = data_i[1968] & sel_one_hot_i[15];
  assign data_masked[1967] = data_i[1967] & sel_one_hot_i[15];
  assign data_masked[1966] = data_i[1966] & sel_one_hot_i[15];
  assign data_masked[1965] = data_i[1965] & sel_one_hot_i[15];
  assign data_masked[1964] = data_i[1964] & sel_one_hot_i[15];
  assign data_masked[1963] = data_i[1963] & sel_one_hot_i[15];
  assign data_masked[1962] = data_i[1962] & sel_one_hot_i[15];
  assign data_masked[1961] = data_i[1961] & sel_one_hot_i[15];
  assign data_masked[1960] = data_i[1960] & sel_one_hot_i[15];
  assign data_masked[1959] = data_i[1959] & sel_one_hot_i[15];
  assign data_masked[1958] = data_i[1958] & sel_one_hot_i[15];
  assign data_masked[1957] = data_i[1957] & sel_one_hot_i[15];
  assign data_masked[1956] = data_i[1956] & sel_one_hot_i[15];
  assign data_masked[1955] = data_i[1955] & sel_one_hot_i[15];
  assign data_masked[1954] = data_i[1954] & sel_one_hot_i[15];
  assign data_masked[1953] = data_i[1953] & sel_one_hot_i[15];
  assign data_masked[1952] = data_i[1952] & sel_one_hot_i[15];
  assign data_masked[1951] = data_i[1951] & sel_one_hot_i[15];
  assign data_masked[1950] = data_i[1950] & sel_one_hot_i[15];
  assign data_masked[1949] = data_i[1949] & sel_one_hot_i[15];
  assign data_masked[1948] = data_i[1948] & sel_one_hot_i[15];
  assign data_masked[1947] = data_i[1947] & sel_one_hot_i[15];
  assign data_masked[1946] = data_i[1946] & sel_one_hot_i[15];
  assign data_masked[1945] = data_i[1945] & sel_one_hot_i[15];
  assign data_masked[1944] = data_i[1944] & sel_one_hot_i[15];
  assign data_masked[1943] = data_i[1943] & sel_one_hot_i[15];
  assign data_masked[1942] = data_i[1942] & sel_one_hot_i[15];
  assign data_masked[1941] = data_i[1941] & sel_one_hot_i[15];
  assign data_masked[1940] = data_i[1940] & sel_one_hot_i[15];
  assign data_masked[1939] = data_i[1939] & sel_one_hot_i[15];
  assign data_masked[1938] = data_i[1938] & sel_one_hot_i[15];
  assign data_masked[1937] = data_i[1937] & sel_one_hot_i[15];
  assign data_masked[1936] = data_i[1936] & sel_one_hot_i[15];
  assign data_masked[1935] = data_i[1935] & sel_one_hot_i[15];
  assign data_masked[1934] = data_i[1934] & sel_one_hot_i[15];
  assign data_masked[1933] = data_i[1933] & sel_one_hot_i[15];
  assign data_masked[1932] = data_i[1932] & sel_one_hot_i[15];
  assign data_masked[1931] = data_i[1931] & sel_one_hot_i[15];
  assign data_masked[1930] = data_i[1930] & sel_one_hot_i[15];
  assign data_masked[1929] = data_i[1929] & sel_one_hot_i[15];
  assign data_masked[1928] = data_i[1928] & sel_one_hot_i[15];
  assign data_masked[1927] = data_i[1927] & sel_one_hot_i[15];
  assign data_masked[1926] = data_i[1926] & sel_one_hot_i[15];
  assign data_masked[1925] = data_i[1925] & sel_one_hot_i[15];
  assign data_masked[1924] = data_i[1924] & sel_one_hot_i[15];
  assign data_masked[1923] = data_i[1923] & sel_one_hot_i[15];
  assign data_masked[1922] = data_i[1922] & sel_one_hot_i[15];
  assign data_masked[1921] = data_i[1921] & sel_one_hot_i[15];
  assign data_masked[1920] = data_i[1920] & sel_one_hot_i[15];
  assign data_masked[2175] = data_i[2175] & sel_one_hot_i[16];
  assign data_masked[2174] = data_i[2174] & sel_one_hot_i[16];
  assign data_masked[2173] = data_i[2173] & sel_one_hot_i[16];
  assign data_masked[2172] = data_i[2172] & sel_one_hot_i[16];
  assign data_masked[2171] = data_i[2171] & sel_one_hot_i[16];
  assign data_masked[2170] = data_i[2170] & sel_one_hot_i[16];
  assign data_masked[2169] = data_i[2169] & sel_one_hot_i[16];
  assign data_masked[2168] = data_i[2168] & sel_one_hot_i[16];
  assign data_masked[2167] = data_i[2167] & sel_one_hot_i[16];
  assign data_masked[2166] = data_i[2166] & sel_one_hot_i[16];
  assign data_masked[2165] = data_i[2165] & sel_one_hot_i[16];
  assign data_masked[2164] = data_i[2164] & sel_one_hot_i[16];
  assign data_masked[2163] = data_i[2163] & sel_one_hot_i[16];
  assign data_masked[2162] = data_i[2162] & sel_one_hot_i[16];
  assign data_masked[2161] = data_i[2161] & sel_one_hot_i[16];
  assign data_masked[2160] = data_i[2160] & sel_one_hot_i[16];
  assign data_masked[2159] = data_i[2159] & sel_one_hot_i[16];
  assign data_masked[2158] = data_i[2158] & sel_one_hot_i[16];
  assign data_masked[2157] = data_i[2157] & sel_one_hot_i[16];
  assign data_masked[2156] = data_i[2156] & sel_one_hot_i[16];
  assign data_masked[2155] = data_i[2155] & sel_one_hot_i[16];
  assign data_masked[2154] = data_i[2154] & sel_one_hot_i[16];
  assign data_masked[2153] = data_i[2153] & sel_one_hot_i[16];
  assign data_masked[2152] = data_i[2152] & sel_one_hot_i[16];
  assign data_masked[2151] = data_i[2151] & sel_one_hot_i[16];
  assign data_masked[2150] = data_i[2150] & sel_one_hot_i[16];
  assign data_masked[2149] = data_i[2149] & sel_one_hot_i[16];
  assign data_masked[2148] = data_i[2148] & sel_one_hot_i[16];
  assign data_masked[2147] = data_i[2147] & sel_one_hot_i[16];
  assign data_masked[2146] = data_i[2146] & sel_one_hot_i[16];
  assign data_masked[2145] = data_i[2145] & sel_one_hot_i[16];
  assign data_masked[2144] = data_i[2144] & sel_one_hot_i[16];
  assign data_masked[2143] = data_i[2143] & sel_one_hot_i[16];
  assign data_masked[2142] = data_i[2142] & sel_one_hot_i[16];
  assign data_masked[2141] = data_i[2141] & sel_one_hot_i[16];
  assign data_masked[2140] = data_i[2140] & sel_one_hot_i[16];
  assign data_masked[2139] = data_i[2139] & sel_one_hot_i[16];
  assign data_masked[2138] = data_i[2138] & sel_one_hot_i[16];
  assign data_masked[2137] = data_i[2137] & sel_one_hot_i[16];
  assign data_masked[2136] = data_i[2136] & sel_one_hot_i[16];
  assign data_masked[2135] = data_i[2135] & sel_one_hot_i[16];
  assign data_masked[2134] = data_i[2134] & sel_one_hot_i[16];
  assign data_masked[2133] = data_i[2133] & sel_one_hot_i[16];
  assign data_masked[2132] = data_i[2132] & sel_one_hot_i[16];
  assign data_masked[2131] = data_i[2131] & sel_one_hot_i[16];
  assign data_masked[2130] = data_i[2130] & sel_one_hot_i[16];
  assign data_masked[2129] = data_i[2129] & sel_one_hot_i[16];
  assign data_masked[2128] = data_i[2128] & sel_one_hot_i[16];
  assign data_masked[2127] = data_i[2127] & sel_one_hot_i[16];
  assign data_masked[2126] = data_i[2126] & sel_one_hot_i[16];
  assign data_masked[2125] = data_i[2125] & sel_one_hot_i[16];
  assign data_masked[2124] = data_i[2124] & sel_one_hot_i[16];
  assign data_masked[2123] = data_i[2123] & sel_one_hot_i[16];
  assign data_masked[2122] = data_i[2122] & sel_one_hot_i[16];
  assign data_masked[2121] = data_i[2121] & sel_one_hot_i[16];
  assign data_masked[2120] = data_i[2120] & sel_one_hot_i[16];
  assign data_masked[2119] = data_i[2119] & sel_one_hot_i[16];
  assign data_masked[2118] = data_i[2118] & sel_one_hot_i[16];
  assign data_masked[2117] = data_i[2117] & sel_one_hot_i[16];
  assign data_masked[2116] = data_i[2116] & sel_one_hot_i[16];
  assign data_masked[2115] = data_i[2115] & sel_one_hot_i[16];
  assign data_masked[2114] = data_i[2114] & sel_one_hot_i[16];
  assign data_masked[2113] = data_i[2113] & sel_one_hot_i[16];
  assign data_masked[2112] = data_i[2112] & sel_one_hot_i[16];
  assign data_masked[2111] = data_i[2111] & sel_one_hot_i[16];
  assign data_masked[2110] = data_i[2110] & sel_one_hot_i[16];
  assign data_masked[2109] = data_i[2109] & sel_one_hot_i[16];
  assign data_masked[2108] = data_i[2108] & sel_one_hot_i[16];
  assign data_masked[2107] = data_i[2107] & sel_one_hot_i[16];
  assign data_masked[2106] = data_i[2106] & sel_one_hot_i[16];
  assign data_masked[2105] = data_i[2105] & sel_one_hot_i[16];
  assign data_masked[2104] = data_i[2104] & sel_one_hot_i[16];
  assign data_masked[2103] = data_i[2103] & sel_one_hot_i[16];
  assign data_masked[2102] = data_i[2102] & sel_one_hot_i[16];
  assign data_masked[2101] = data_i[2101] & sel_one_hot_i[16];
  assign data_masked[2100] = data_i[2100] & sel_one_hot_i[16];
  assign data_masked[2099] = data_i[2099] & sel_one_hot_i[16];
  assign data_masked[2098] = data_i[2098] & sel_one_hot_i[16];
  assign data_masked[2097] = data_i[2097] & sel_one_hot_i[16];
  assign data_masked[2096] = data_i[2096] & sel_one_hot_i[16];
  assign data_masked[2095] = data_i[2095] & sel_one_hot_i[16];
  assign data_masked[2094] = data_i[2094] & sel_one_hot_i[16];
  assign data_masked[2093] = data_i[2093] & sel_one_hot_i[16];
  assign data_masked[2092] = data_i[2092] & sel_one_hot_i[16];
  assign data_masked[2091] = data_i[2091] & sel_one_hot_i[16];
  assign data_masked[2090] = data_i[2090] & sel_one_hot_i[16];
  assign data_masked[2089] = data_i[2089] & sel_one_hot_i[16];
  assign data_masked[2088] = data_i[2088] & sel_one_hot_i[16];
  assign data_masked[2087] = data_i[2087] & sel_one_hot_i[16];
  assign data_masked[2086] = data_i[2086] & sel_one_hot_i[16];
  assign data_masked[2085] = data_i[2085] & sel_one_hot_i[16];
  assign data_masked[2084] = data_i[2084] & sel_one_hot_i[16];
  assign data_masked[2083] = data_i[2083] & sel_one_hot_i[16];
  assign data_masked[2082] = data_i[2082] & sel_one_hot_i[16];
  assign data_masked[2081] = data_i[2081] & sel_one_hot_i[16];
  assign data_masked[2080] = data_i[2080] & sel_one_hot_i[16];
  assign data_masked[2079] = data_i[2079] & sel_one_hot_i[16];
  assign data_masked[2078] = data_i[2078] & sel_one_hot_i[16];
  assign data_masked[2077] = data_i[2077] & sel_one_hot_i[16];
  assign data_masked[2076] = data_i[2076] & sel_one_hot_i[16];
  assign data_masked[2075] = data_i[2075] & sel_one_hot_i[16];
  assign data_masked[2074] = data_i[2074] & sel_one_hot_i[16];
  assign data_masked[2073] = data_i[2073] & sel_one_hot_i[16];
  assign data_masked[2072] = data_i[2072] & sel_one_hot_i[16];
  assign data_masked[2071] = data_i[2071] & sel_one_hot_i[16];
  assign data_masked[2070] = data_i[2070] & sel_one_hot_i[16];
  assign data_masked[2069] = data_i[2069] & sel_one_hot_i[16];
  assign data_masked[2068] = data_i[2068] & sel_one_hot_i[16];
  assign data_masked[2067] = data_i[2067] & sel_one_hot_i[16];
  assign data_masked[2066] = data_i[2066] & sel_one_hot_i[16];
  assign data_masked[2065] = data_i[2065] & sel_one_hot_i[16];
  assign data_masked[2064] = data_i[2064] & sel_one_hot_i[16];
  assign data_masked[2063] = data_i[2063] & sel_one_hot_i[16];
  assign data_masked[2062] = data_i[2062] & sel_one_hot_i[16];
  assign data_masked[2061] = data_i[2061] & sel_one_hot_i[16];
  assign data_masked[2060] = data_i[2060] & sel_one_hot_i[16];
  assign data_masked[2059] = data_i[2059] & sel_one_hot_i[16];
  assign data_masked[2058] = data_i[2058] & sel_one_hot_i[16];
  assign data_masked[2057] = data_i[2057] & sel_one_hot_i[16];
  assign data_masked[2056] = data_i[2056] & sel_one_hot_i[16];
  assign data_masked[2055] = data_i[2055] & sel_one_hot_i[16];
  assign data_masked[2054] = data_i[2054] & sel_one_hot_i[16];
  assign data_masked[2053] = data_i[2053] & sel_one_hot_i[16];
  assign data_masked[2052] = data_i[2052] & sel_one_hot_i[16];
  assign data_masked[2051] = data_i[2051] & sel_one_hot_i[16];
  assign data_masked[2050] = data_i[2050] & sel_one_hot_i[16];
  assign data_masked[2049] = data_i[2049] & sel_one_hot_i[16];
  assign data_masked[2048] = data_i[2048] & sel_one_hot_i[16];
  assign data_masked[2303] = data_i[2303] & sel_one_hot_i[17];
  assign data_masked[2302] = data_i[2302] & sel_one_hot_i[17];
  assign data_masked[2301] = data_i[2301] & sel_one_hot_i[17];
  assign data_masked[2300] = data_i[2300] & sel_one_hot_i[17];
  assign data_masked[2299] = data_i[2299] & sel_one_hot_i[17];
  assign data_masked[2298] = data_i[2298] & sel_one_hot_i[17];
  assign data_masked[2297] = data_i[2297] & sel_one_hot_i[17];
  assign data_masked[2296] = data_i[2296] & sel_one_hot_i[17];
  assign data_masked[2295] = data_i[2295] & sel_one_hot_i[17];
  assign data_masked[2294] = data_i[2294] & sel_one_hot_i[17];
  assign data_masked[2293] = data_i[2293] & sel_one_hot_i[17];
  assign data_masked[2292] = data_i[2292] & sel_one_hot_i[17];
  assign data_masked[2291] = data_i[2291] & sel_one_hot_i[17];
  assign data_masked[2290] = data_i[2290] & sel_one_hot_i[17];
  assign data_masked[2289] = data_i[2289] & sel_one_hot_i[17];
  assign data_masked[2288] = data_i[2288] & sel_one_hot_i[17];
  assign data_masked[2287] = data_i[2287] & sel_one_hot_i[17];
  assign data_masked[2286] = data_i[2286] & sel_one_hot_i[17];
  assign data_masked[2285] = data_i[2285] & sel_one_hot_i[17];
  assign data_masked[2284] = data_i[2284] & sel_one_hot_i[17];
  assign data_masked[2283] = data_i[2283] & sel_one_hot_i[17];
  assign data_masked[2282] = data_i[2282] & sel_one_hot_i[17];
  assign data_masked[2281] = data_i[2281] & sel_one_hot_i[17];
  assign data_masked[2280] = data_i[2280] & sel_one_hot_i[17];
  assign data_masked[2279] = data_i[2279] & sel_one_hot_i[17];
  assign data_masked[2278] = data_i[2278] & sel_one_hot_i[17];
  assign data_masked[2277] = data_i[2277] & sel_one_hot_i[17];
  assign data_masked[2276] = data_i[2276] & sel_one_hot_i[17];
  assign data_masked[2275] = data_i[2275] & sel_one_hot_i[17];
  assign data_masked[2274] = data_i[2274] & sel_one_hot_i[17];
  assign data_masked[2273] = data_i[2273] & sel_one_hot_i[17];
  assign data_masked[2272] = data_i[2272] & sel_one_hot_i[17];
  assign data_masked[2271] = data_i[2271] & sel_one_hot_i[17];
  assign data_masked[2270] = data_i[2270] & sel_one_hot_i[17];
  assign data_masked[2269] = data_i[2269] & sel_one_hot_i[17];
  assign data_masked[2268] = data_i[2268] & sel_one_hot_i[17];
  assign data_masked[2267] = data_i[2267] & sel_one_hot_i[17];
  assign data_masked[2266] = data_i[2266] & sel_one_hot_i[17];
  assign data_masked[2265] = data_i[2265] & sel_one_hot_i[17];
  assign data_masked[2264] = data_i[2264] & sel_one_hot_i[17];
  assign data_masked[2263] = data_i[2263] & sel_one_hot_i[17];
  assign data_masked[2262] = data_i[2262] & sel_one_hot_i[17];
  assign data_masked[2261] = data_i[2261] & sel_one_hot_i[17];
  assign data_masked[2260] = data_i[2260] & sel_one_hot_i[17];
  assign data_masked[2259] = data_i[2259] & sel_one_hot_i[17];
  assign data_masked[2258] = data_i[2258] & sel_one_hot_i[17];
  assign data_masked[2257] = data_i[2257] & sel_one_hot_i[17];
  assign data_masked[2256] = data_i[2256] & sel_one_hot_i[17];
  assign data_masked[2255] = data_i[2255] & sel_one_hot_i[17];
  assign data_masked[2254] = data_i[2254] & sel_one_hot_i[17];
  assign data_masked[2253] = data_i[2253] & sel_one_hot_i[17];
  assign data_masked[2252] = data_i[2252] & sel_one_hot_i[17];
  assign data_masked[2251] = data_i[2251] & sel_one_hot_i[17];
  assign data_masked[2250] = data_i[2250] & sel_one_hot_i[17];
  assign data_masked[2249] = data_i[2249] & sel_one_hot_i[17];
  assign data_masked[2248] = data_i[2248] & sel_one_hot_i[17];
  assign data_masked[2247] = data_i[2247] & sel_one_hot_i[17];
  assign data_masked[2246] = data_i[2246] & sel_one_hot_i[17];
  assign data_masked[2245] = data_i[2245] & sel_one_hot_i[17];
  assign data_masked[2244] = data_i[2244] & sel_one_hot_i[17];
  assign data_masked[2243] = data_i[2243] & sel_one_hot_i[17];
  assign data_masked[2242] = data_i[2242] & sel_one_hot_i[17];
  assign data_masked[2241] = data_i[2241] & sel_one_hot_i[17];
  assign data_masked[2240] = data_i[2240] & sel_one_hot_i[17];
  assign data_masked[2239] = data_i[2239] & sel_one_hot_i[17];
  assign data_masked[2238] = data_i[2238] & sel_one_hot_i[17];
  assign data_masked[2237] = data_i[2237] & sel_one_hot_i[17];
  assign data_masked[2236] = data_i[2236] & sel_one_hot_i[17];
  assign data_masked[2235] = data_i[2235] & sel_one_hot_i[17];
  assign data_masked[2234] = data_i[2234] & sel_one_hot_i[17];
  assign data_masked[2233] = data_i[2233] & sel_one_hot_i[17];
  assign data_masked[2232] = data_i[2232] & sel_one_hot_i[17];
  assign data_masked[2231] = data_i[2231] & sel_one_hot_i[17];
  assign data_masked[2230] = data_i[2230] & sel_one_hot_i[17];
  assign data_masked[2229] = data_i[2229] & sel_one_hot_i[17];
  assign data_masked[2228] = data_i[2228] & sel_one_hot_i[17];
  assign data_masked[2227] = data_i[2227] & sel_one_hot_i[17];
  assign data_masked[2226] = data_i[2226] & sel_one_hot_i[17];
  assign data_masked[2225] = data_i[2225] & sel_one_hot_i[17];
  assign data_masked[2224] = data_i[2224] & sel_one_hot_i[17];
  assign data_masked[2223] = data_i[2223] & sel_one_hot_i[17];
  assign data_masked[2222] = data_i[2222] & sel_one_hot_i[17];
  assign data_masked[2221] = data_i[2221] & sel_one_hot_i[17];
  assign data_masked[2220] = data_i[2220] & sel_one_hot_i[17];
  assign data_masked[2219] = data_i[2219] & sel_one_hot_i[17];
  assign data_masked[2218] = data_i[2218] & sel_one_hot_i[17];
  assign data_masked[2217] = data_i[2217] & sel_one_hot_i[17];
  assign data_masked[2216] = data_i[2216] & sel_one_hot_i[17];
  assign data_masked[2215] = data_i[2215] & sel_one_hot_i[17];
  assign data_masked[2214] = data_i[2214] & sel_one_hot_i[17];
  assign data_masked[2213] = data_i[2213] & sel_one_hot_i[17];
  assign data_masked[2212] = data_i[2212] & sel_one_hot_i[17];
  assign data_masked[2211] = data_i[2211] & sel_one_hot_i[17];
  assign data_masked[2210] = data_i[2210] & sel_one_hot_i[17];
  assign data_masked[2209] = data_i[2209] & sel_one_hot_i[17];
  assign data_masked[2208] = data_i[2208] & sel_one_hot_i[17];
  assign data_masked[2207] = data_i[2207] & sel_one_hot_i[17];
  assign data_masked[2206] = data_i[2206] & sel_one_hot_i[17];
  assign data_masked[2205] = data_i[2205] & sel_one_hot_i[17];
  assign data_masked[2204] = data_i[2204] & sel_one_hot_i[17];
  assign data_masked[2203] = data_i[2203] & sel_one_hot_i[17];
  assign data_masked[2202] = data_i[2202] & sel_one_hot_i[17];
  assign data_masked[2201] = data_i[2201] & sel_one_hot_i[17];
  assign data_masked[2200] = data_i[2200] & sel_one_hot_i[17];
  assign data_masked[2199] = data_i[2199] & sel_one_hot_i[17];
  assign data_masked[2198] = data_i[2198] & sel_one_hot_i[17];
  assign data_masked[2197] = data_i[2197] & sel_one_hot_i[17];
  assign data_masked[2196] = data_i[2196] & sel_one_hot_i[17];
  assign data_masked[2195] = data_i[2195] & sel_one_hot_i[17];
  assign data_masked[2194] = data_i[2194] & sel_one_hot_i[17];
  assign data_masked[2193] = data_i[2193] & sel_one_hot_i[17];
  assign data_masked[2192] = data_i[2192] & sel_one_hot_i[17];
  assign data_masked[2191] = data_i[2191] & sel_one_hot_i[17];
  assign data_masked[2190] = data_i[2190] & sel_one_hot_i[17];
  assign data_masked[2189] = data_i[2189] & sel_one_hot_i[17];
  assign data_masked[2188] = data_i[2188] & sel_one_hot_i[17];
  assign data_masked[2187] = data_i[2187] & sel_one_hot_i[17];
  assign data_masked[2186] = data_i[2186] & sel_one_hot_i[17];
  assign data_masked[2185] = data_i[2185] & sel_one_hot_i[17];
  assign data_masked[2184] = data_i[2184] & sel_one_hot_i[17];
  assign data_masked[2183] = data_i[2183] & sel_one_hot_i[17];
  assign data_masked[2182] = data_i[2182] & sel_one_hot_i[17];
  assign data_masked[2181] = data_i[2181] & sel_one_hot_i[17];
  assign data_masked[2180] = data_i[2180] & sel_one_hot_i[17];
  assign data_masked[2179] = data_i[2179] & sel_one_hot_i[17];
  assign data_masked[2178] = data_i[2178] & sel_one_hot_i[17];
  assign data_masked[2177] = data_i[2177] & sel_one_hot_i[17];
  assign data_masked[2176] = data_i[2176] & sel_one_hot_i[17];
  assign data_masked[2431] = data_i[2431] & sel_one_hot_i[18];
  assign data_masked[2430] = data_i[2430] & sel_one_hot_i[18];
  assign data_masked[2429] = data_i[2429] & sel_one_hot_i[18];
  assign data_masked[2428] = data_i[2428] & sel_one_hot_i[18];
  assign data_masked[2427] = data_i[2427] & sel_one_hot_i[18];
  assign data_masked[2426] = data_i[2426] & sel_one_hot_i[18];
  assign data_masked[2425] = data_i[2425] & sel_one_hot_i[18];
  assign data_masked[2424] = data_i[2424] & sel_one_hot_i[18];
  assign data_masked[2423] = data_i[2423] & sel_one_hot_i[18];
  assign data_masked[2422] = data_i[2422] & sel_one_hot_i[18];
  assign data_masked[2421] = data_i[2421] & sel_one_hot_i[18];
  assign data_masked[2420] = data_i[2420] & sel_one_hot_i[18];
  assign data_masked[2419] = data_i[2419] & sel_one_hot_i[18];
  assign data_masked[2418] = data_i[2418] & sel_one_hot_i[18];
  assign data_masked[2417] = data_i[2417] & sel_one_hot_i[18];
  assign data_masked[2416] = data_i[2416] & sel_one_hot_i[18];
  assign data_masked[2415] = data_i[2415] & sel_one_hot_i[18];
  assign data_masked[2414] = data_i[2414] & sel_one_hot_i[18];
  assign data_masked[2413] = data_i[2413] & sel_one_hot_i[18];
  assign data_masked[2412] = data_i[2412] & sel_one_hot_i[18];
  assign data_masked[2411] = data_i[2411] & sel_one_hot_i[18];
  assign data_masked[2410] = data_i[2410] & sel_one_hot_i[18];
  assign data_masked[2409] = data_i[2409] & sel_one_hot_i[18];
  assign data_masked[2408] = data_i[2408] & sel_one_hot_i[18];
  assign data_masked[2407] = data_i[2407] & sel_one_hot_i[18];
  assign data_masked[2406] = data_i[2406] & sel_one_hot_i[18];
  assign data_masked[2405] = data_i[2405] & sel_one_hot_i[18];
  assign data_masked[2404] = data_i[2404] & sel_one_hot_i[18];
  assign data_masked[2403] = data_i[2403] & sel_one_hot_i[18];
  assign data_masked[2402] = data_i[2402] & sel_one_hot_i[18];
  assign data_masked[2401] = data_i[2401] & sel_one_hot_i[18];
  assign data_masked[2400] = data_i[2400] & sel_one_hot_i[18];
  assign data_masked[2399] = data_i[2399] & sel_one_hot_i[18];
  assign data_masked[2398] = data_i[2398] & sel_one_hot_i[18];
  assign data_masked[2397] = data_i[2397] & sel_one_hot_i[18];
  assign data_masked[2396] = data_i[2396] & sel_one_hot_i[18];
  assign data_masked[2395] = data_i[2395] & sel_one_hot_i[18];
  assign data_masked[2394] = data_i[2394] & sel_one_hot_i[18];
  assign data_masked[2393] = data_i[2393] & sel_one_hot_i[18];
  assign data_masked[2392] = data_i[2392] & sel_one_hot_i[18];
  assign data_masked[2391] = data_i[2391] & sel_one_hot_i[18];
  assign data_masked[2390] = data_i[2390] & sel_one_hot_i[18];
  assign data_masked[2389] = data_i[2389] & sel_one_hot_i[18];
  assign data_masked[2388] = data_i[2388] & sel_one_hot_i[18];
  assign data_masked[2387] = data_i[2387] & sel_one_hot_i[18];
  assign data_masked[2386] = data_i[2386] & sel_one_hot_i[18];
  assign data_masked[2385] = data_i[2385] & sel_one_hot_i[18];
  assign data_masked[2384] = data_i[2384] & sel_one_hot_i[18];
  assign data_masked[2383] = data_i[2383] & sel_one_hot_i[18];
  assign data_masked[2382] = data_i[2382] & sel_one_hot_i[18];
  assign data_masked[2381] = data_i[2381] & sel_one_hot_i[18];
  assign data_masked[2380] = data_i[2380] & sel_one_hot_i[18];
  assign data_masked[2379] = data_i[2379] & sel_one_hot_i[18];
  assign data_masked[2378] = data_i[2378] & sel_one_hot_i[18];
  assign data_masked[2377] = data_i[2377] & sel_one_hot_i[18];
  assign data_masked[2376] = data_i[2376] & sel_one_hot_i[18];
  assign data_masked[2375] = data_i[2375] & sel_one_hot_i[18];
  assign data_masked[2374] = data_i[2374] & sel_one_hot_i[18];
  assign data_masked[2373] = data_i[2373] & sel_one_hot_i[18];
  assign data_masked[2372] = data_i[2372] & sel_one_hot_i[18];
  assign data_masked[2371] = data_i[2371] & sel_one_hot_i[18];
  assign data_masked[2370] = data_i[2370] & sel_one_hot_i[18];
  assign data_masked[2369] = data_i[2369] & sel_one_hot_i[18];
  assign data_masked[2368] = data_i[2368] & sel_one_hot_i[18];
  assign data_masked[2367] = data_i[2367] & sel_one_hot_i[18];
  assign data_masked[2366] = data_i[2366] & sel_one_hot_i[18];
  assign data_masked[2365] = data_i[2365] & sel_one_hot_i[18];
  assign data_masked[2364] = data_i[2364] & sel_one_hot_i[18];
  assign data_masked[2363] = data_i[2363] & sel_one_hot_i[18];
  assign data_masked[2362] = data_i[2362] & sel_one_hot_i[18];
  assign data_masked[2361] = data_i[2361] & sel_one_hot_i[18];
  assign data_masked[2360] = data_i[2360] & sel_one_hot_i[18];
  assign data_masked[2359] = data_i[2359] & sel_one_hot_i[18];
  assign data_masked[2358] = data_i[2358] & sel_one_hot_i[18];
  assign data_masked[2357] = data_i[2357] & sel_one_hot_i[18];
  assign data_masked[2356] = data_i[2356] & sel_one_hot_i[18];
  assign data_masked[2355] = data_i[2355] & sel_one_hot_i[18];
  assign data_masked[2354] = data_i[2354] & sel_one_hot_i[18];
  assign data_masked[2353] = data_i[2353] & sel_one_hot_i[18];
  assign data_masked[2352] = data_i[2352] & sel_one_hot_i[18];
  assign data_masked[2351] = data_i[2351] & sel_one_hot_i[18];
  assign data_masked[2350] = data_i[2350] & sel_one_hot_i[18];
  assign data_masked[2349] = data_i[2349] & sel_one_hot_i[18];
  assign data_masked[2348] = data_i[2348] & sel_one_hot_i[18];
  assign data_masked[2347] = data_i[2347] & sel_one_hot_i[18];
  assign data_masked[2346] = data_i[2346] & sel_one_hot_i[18];
  assign data_masked[2345] = data_i[2345] & sel_one_hot_i[18];
  assign data_masked[2344] = data_i[2344] & sel_one_hot_i[18];
  assign data_masked[2343] = data_i[2343] & sel_one_hot_i[18];
  assign data_masked[2342] = data_i[2342] & sel_one_hot_i[18];
  assign data_masked[2341] = data_i[2341] & sel_one_hot_i[18];
  assign data_masked[2340] = data_i[2340] & sel_one_hot_i[18];
  assign data_masked[2339] = data_i[2339] & sel_one_hot_i[18];
  assign data_masked[2338] = data_i[2338] & sel_one_hot_i[18];
  assign data_masked[2337] = data_i[2337] & sel_one_hot_i[18];
  assign data_masked[2336] = data_i[2336] & sel_one_hot_i[18];
  assign data_masked[2335] = data_i[2335] & sel_one_hot_i[18];
  assign data_masked[2334] = data_i[2334] & sel_one_hot_i[18];
  assign data_masked[2333] = data_i[2333] & sel_one_hot_i[18];
  assign data_masked[2332] = data_i[2332] & sel_one_hot_i[18];
  assign data_masked[2331] = data_i[2331] & sel_one_hot_i[18];
  assign data_masked[2330] = data_i[2330] & sel_one_hot_i[18];
  assign data_masked[2329] = data_i[2329] & sel_one_hot_i[18];
  assign data_masked[2328] = data_i[2328] & sel_one_hot_i[18];
  assign data_masked[2327] = data_i[2327] & sel_one_hot_i[18];
  assign data_masked[2326] = data_i[2326] & sel_one_hot_i[18];
  assign data_masked[2325] = data_i[2325] & sel_one_hot_i[18];
  assign data_masked[2324] = data_i[2324] & sel_one_hot_i[18];
  assign data_masked[2323] = data_i[2323] & sel_one_hot_i[18];
  assign data_masked[2322] = data_i[2322] & sel_one_hot_i[18];
  assign data_masked[2321] = data_i[2321] & sel_one_hot_i[18];
  assign data_masked[2320] = data_i[2320] & sel_one_hot_i[18];
  assign data_masked[2319] = data_i[2319] & sel_one_hot_i[18];
  assign data_masked[2318] = data_i[2318] & sel_one_hot_i[18];
  assign data_masked[2317] = data_i[2317] & sel_one_hot_i[18];
  assign data_masked[2316] = data_i[2316] & sel_one_hot_i[18];
  assign data_masked[2315] = data_i[2315] & sel_one_hot_i[18];
  assign data_masked[2314] = data_i[2314] & sel_one_hot_i[18];
  assign data_masked[2313] = data_i[2313] & sel_one_hot_i[18];
  assign data_masked[2312] = data_i[2312] & sel_one_hot_i[18];
  assign data_masked[2311] = data_i[2311] & sel_one_hot_i[18];
  assign data_masked[2310] = data_i[2310] & sel_one_hot_i[18];
  assign data_masked[2309] = data_i[2309] & sel_one_hot_i[18];
  assign data_masked[2308] = data_i[2308] & sel_one_hot_i[18];
  assign data_masked[2307] = data_i[2307] & sel_one_hot_i[18];
  assign data_masked[2306] = data_i[2306] & sel_one_hot_i[18];
  assign data_masked[2305] = data_i[2305] & sel_one_hot_i[18];
  assign data_masked[2304] = data_i[2304] & sel_one_hot_i[18];
  assign data_masked[2559] = data_i[2559] & sel_one_hot_i[19];
  assign data_masked[2558] = data_i[2558] & sel_one_hot_i[19];
  assign data_masked[2557] = data_i[2557] & sel_one_hot_i[19];
  assign data_masked[2556] = data_i[2556] & sel_one_hot_i[19];
  assign data_masked[2555] = data_i[2555] & sel_one_hot_i[19];
  assign data_masked[2554] = data_i[2554] & sel_one_hot_i[19];
  assign data_masked[2553] = data_i[2553] & sel_one_hot_i[19];
  assign data_masked[2552] = data_i[2552] & sel_one_hot_i[19];
  assign data_masked[2551] = data_i[2551] & sel_one_hot_i[19];
  assign data_masked[2550] = data_i[2550] & sel_one_hot_i[19];
  assign data_masked[2549] = data_i[2549] & sel_one_hot_i[19];
  assign data_masked[2548] = data_i[2548] & sel_one_hot_i[19];
  assign data_masked[2547] = data_i[2547] & sel_one_hot_i[19];
  assign data_masked[2546] = data_i[2546] & sel_one_hot_i[19];
  assign data_masked[2545] = data_i[2545] & sel_one_hot_i[19];
  assign data_masked[2544] = data_i[2544] & sel_one_hot_i[19];
  assign data_masked[2543] = data_i[2543] & sel_one_hot_i[19];
  assign data_masked[2542] = data_i[2542] & sel_one_hot_i[19];
  assign data_masked[2541] = data_i[2541] & sel_one_hot_i[19];
  assign data_masked[2540] = data_i[2540] & sel_one_hot_i[19];
  assign data_masked[2539] = data_i[2539] & sel_one_hot_i[19];
  assign data_masked[2538] = data_i[2538] & sel_one_hot_i[19];
  assign data_masked[2537] = data_i[2537] & sel_one_hot_i[19];
  assign data_masked[2536] = data_i[2536] & sel_one_hot_i[19];
  assign data_masked[2535] = data_i[2535] & sel_one_hot_i[19];
  assign data_masked[2534] = data_i[2534] & sel_one_hot_i[19];
  assign data_masked[2533] = data_i[2533] & sel_one_hot_i[19];
  assign data_masked[2532] = data_i[2532] & sel_one_hot_i[19];
  assign data_masked[2531] = data_i[2531] & sel_one_hot_i[19];
  assign data_masked[2530] = data_i[2530] & sel_one_hot_i[19];
  assign data_masked[2529] = data_i[2529] & sel_one_hot_i[19];
  assign data_masked[2528] = data_i[2528] & sel_one_hot_i[19];
  assign data_masked[2527] = data_i[2527] & sel_one_hot_i[19];
  assign data_masked[2526] = data_i[2526] & sel_one_hot_i[19];
  assign data_masked[2525] = data_i[2525] & sel_one_hot_i[19];
  assign data_masked[2524] = data_i[2524] & sel_one_hot_i[19];
  assign data_masked[2523] = data_i[2523] & sel_one_hot_i[19];
  assign data_masked[2522] = data_i[2522] & sel_one_hot_i[19];
  assign data_masked[2521] = data_i[2521] & sel_one_hot_i[19];
  assign data_masked[2520] = data_i[2520] & sel_one_hot_i[19];
  assign data_masked[2519] = data_i[2519] & sel_one_hot_i[19];
  assign data_masked[2518] = data_i[2518] & sel_one_hot_i[19];
  assign data_masked[2517] = data_i[2517] & sel_one_hot_i[19];
  assign data_masked[2516] = data_i[2516] & sel_one_hot_i[19];
  assign data_masked[2515] = data_i[2515] & sel_one_hot_i[19];
  assign data_masked[2514] = data_i[2514] & sel_one_hot_i[19];
  assign data_masked[2513] = data_i[2513] & sel_one_hot_i[19];
  assign data_masked[2512] = data_i[2512] & sel_one_hot_i[19];
  assign data_masked[2511] = data_i[2511] & sel_one_hot_i[19];
  assign data_masked[2510] = data_i[2510] & sel_one_hot_i[19];
  assign data_masked[2509] = data_i[2509] & sel_one_hot_i[19];
  assign data_masked[2508] = data_i[2508] & sel_one_hot_i[19];
  assign data_masked[2507] = data_i[2507] & sel_one_hot_i[19];
  assign data_masked[2506] = data_i[2506] & sel_one_hot_i[19];
  assign data_masked[2505] = data_i[2505] & sel_one_hot_i[19];
  assign data_masked[2504] = data_i[2504] & sel_one_hot_i[19];
  assign data_masked[2503] = data_i[2503] & sel_one_hot_i[19];
  assign data_masked[2502] = data_i[2502] & sel_one_hot_i[19];
  assign data_masked[2501] = data_i[2501] & sel_one_hot_i[19];
  assign data_masked[2500] = data_i[2500] & sel_one_hot_i[19];
  assign data_masked[2499] = data_i[2499] & sel_one_hot_i[19];
  assign data_masked[2498] = data_i[2498] & sel_one_hot_i[19];
  assign data_masked[2497] = data_i[2497] & sel_one_hot_i[19];
  assign data_masked[2496] = data_i[2496] & sel_one_hot_i[19];
  assign data_masked[2495] = data_i[2495] & sel_one_hot_i[19];
  assign data_masked[2494] = data_i[2494] & sel_one_hot_i[19];
  assign data_masked[2493] = data_i[2493] & sel_one_hot_i[19];
  assign data_masked[2492] = data_i[2492] & sel_one_hot_i[19];
  assign data_masked[2491] = data_i[2491] & sel_one_hot_i[19];
  assign data_masked[2490] = data_i[2490] & sel_one_hot_i[19];
  assign data_masked[2489] = data_i[2489] & sel_one_hot_i[19];
  assign data_masked[2488] = data_i[2488] & sel_one_hot_i[19];
  assign data_masked[2487] = data_i[2487] & sel_one_hot_i[19];
  assign data_masked[2486] = data_i[2486] & sel_one_hot_i[19];
  assign data_masked[2485] = data_i[2485] & sel_one_hot_i[19];
  assign data_masked[2484] = data_i[2484] & sel_one_hot_i[19];
  assign data_masked[2483] = data_i[2483] & sel_one_hot_i[19];
  assign data_masked[2482] = data_i[2482] & sel_one_hot_i[19];
  assign data_masked[2481] = data_i[2481] & sel_one_hot_i[19];
  assign data_masked[2480] = data_i[2480] & sel_one_hot_i[19];
  assign data_masked[2479] = data_i[2479] & sel_one_hot_i[19];
  assign data_masked[2478] = data_i[2478] & sel_one_hot_i[19];
  assign data_masked[2477] = data_i[2477] & sel_one_hot_i[19];
  assign data_masked[2476] = data_i[2476] & sel_one_hot_i[19];
  assign data_masked[2475] = data_i[2475] & sel_one_hot_i[19];
  assign data_masked[2474] = data_i[2474] & sel_one_hot_i[19];
  assign data_masked[2473] = data_i[2473] & sel_one_hot_i[19];
  assign data_masked[2472] = data_i[2472] & sel_one_hot_i[19];
  assign data_masked[2471] = data_i[2471] & sel_one_hot_i[19];
  assign data_masked[2470] = data_i[2470] & sel_one_hot_i[19];
  assign data_masked[2469] = data_i[2469] & sel_one_hot_i[19];
  assign data_masked[2468] = data_i[2468] & sel_one_hot_i[19];
  assign data_masked[2467] = data_i[2467] & sel_one_hot_i[19];
  assign data_masked[2466] = data_i[2466] & sel_one_hot_i[19];
  assign data_masked[2465] = data_i[2465] & sel_one_hot_i[19];
  assign data_masked[2464] = data_i[2464] & sel_one_hot_i[19];
  assign data_masked[2463] = data_i[2463] & sel_one_hot_i[19];
  assign data_masked[2462] = data_i[2462] & sel_one_hot_i[19];
  assign data_masked[2461] = data_i[2461] & sel_one_hot_i[19];
  assign data_masked[2460] = data_i[2460] & sel_one_hot_i[19];
  assign data_masked[2459] = data_i[2459] & sel_one_hot_i[19];
  assign data_masked[2458] = data_i[2458] & sel_one_hot_i[19];
  assign data_masked[2457] = data_i[2457] & sel_one_hot_i[19];
  assign data_masked[2456] = data_i[2456] & sel_one_hot_i[19];
  assign data_masked[2455] = data_i[2455] & sel_one_hot_i[19];
  assign data_masked[2454] = data_i[2454] & sel_one_hot_i[19];
  assign data_masked[2453] = data_i[2453] & sel_one_hot_i[19];
  assign data_masked[2452] = data_i[2452] & sel_one_hot_i[19];
  assign data_masked[2451] = data_i[2451] & sel_one_hot_i[19];
  assign data_masked[2450] = data_i[2450] & sel_one_hot_i[19];
  assign data_masked[2449] = data_i[2449] & sel_one_hot_i[19];
  assign data_masked[2448] = data_i[2448] & sel_one_hot_i[19];
  assign data_masked[2447] = data_i[2447] & sel_one_hot_i[19];
  assign data_masked[2446] = data_i[2446] & sel_one_hot_i[19];
  assign data_masked[2445] = data_i[2445] & sel_one_hot_i[19];
  assign data_masked[2444] = data_i[2444] & sel_one_hot_i[19];
  assign data_masked[2443] = data_i[2443] & sel_one_hot_i[19];
  assign data_masked[2442] = data_i[2442] & sel_one_hot_i[19];
  assign data_masked[2441] = data_i[2441] & sel_one_hot_i[19];
  assign data_masked[2440] = data_i[2440] & sel_one_hot_i[19];
  assign data_masked[2439] = data_i[2439] & sel_one_hot_i[19];
  assign data_masked[2438] = data_i[2438] & sel_one_hot_i[19];
  assign data_masked[2437] = data_i[2437] & sel_one_hot_i[19];
  assign data_masked[2436] = data_i[2436] & sel_one_hot_i[19];
  assign data_masked[2435] = data_i[2435] & sel_one_hot_i[19];
  assign data_masked[2434] = data_i[2434] & sel_one_hot_i[19];
  assign data_masked[2433] = data_i[2433] & sel_one_hot_i[19];
  assign data_masked[2432] = data_i[2432] & sel_one_hot_i[19];
  assign data_masked[2687] = data_i[2687] & sel_one_hot_i[20];
  assign data_masked[2686] = data_i[2686] & sel_one_hot_i[20];
  assign data_masked[2685] = data_i[2685] & sel_one_hot_i[20];
  assign data_masked[2684] = data_i[2684] & sel_one_hot_i[20];
  assign data_masked[2683] = data_i[2683] & sel_one_hot_i[20];
  assign data_masked[2682] = data_i[2682] & sel_one_hot_i[20];
  assign data_masked[2681] = data_i[2681] & sel_one_hot_i[20];
  assign data_masked[2680] = data_i[2680] & sel_one_hot_i[20];
  assign data_masked[2679] = data_i[2679] & sel_one_hot_i[20];
  assign data_masked[2678] = data_i[2678] & sel_one_hot_i[20];
  assign data_masked[2677] = data_i[2677] & sel_one_hot_i[20];
  assign data_masked[2676] = data_i[2676] & sel_one_hot_i[20];
  assign data_masked[2675] = data_i[2675] & sel_one_hot_i[20];
  assign data_masked[2674] = data_i[2674] & sel_one_hot_i[20];
  assign data_masked[2673] = data_i[2673] & sel_one_hot_i[20];
  assign data_masked[2672] = data_i[2672] & sel_one_hot_i[20];
  assign data_masked[2671] = data_i[2671] & sel_one_hot_i[20];
  assign data_masked[2670] = data_i[2670] & sel_one_hot_i[20];
  assign data_masked[2669] = data_i[2669] & sel_one_hot_i[20];
  assign data_masked[2668] = data_i[2668] & sel_one_hot_i[20];
  assign data_masked[2667] = data_i[2667] & sel_one_hot_i[20];
  assign data_masked[2666] = data_i[2666] & sel_one_hot_i[20];
  assign data_masked[2665] = data_i[2665] & sel_one_hot_i[20];
  assign data_masked[2664] = data_i[2664] & sel_one_hot_i[20];
  assign data_masked[2663] = data_i[2663] & sel_one_hot_i[20];
  assign data_masked[2662] = data_i[2662] & sel_one_hot_i[20];
  assign data_masked[2661] = data_i[2661] & sel_one_hot_i[20];
  assign data_masked[2660] = data_i[2660] & sel_one_hot_i[20];
  assign data_masked[2659] = data_i[2659] & sel_one_hot_i[20];
  assign data_masked[2658] = data_i[2658] & sel_one_hot_i[20];
  assign data_masked[2657] = data_i[2657] & sel_one_hot_i[20];
  assign data_masked[2656] = data_i[2656] & sel_one_hot_i[20];
  assign data_masked[2655] = data_i[2655] & sel_one_hot_i[20];
  assign data_masked[2654] = data_i[2654] & sel_one_hot_i[20];
  assign data_masked[2653] = data_i[2653] & sel_one_hot_i[20];
  assign data_masked[2652] = data_i[2652] & sel_one_hot_i[20];
  assign data_masked[2651] = data_i[2651] & sel_one_hot_i[20];
  assign data_masked[2650] = data_i[2650] & sel_one_hot_i[20];
  assign data_masked[2649] = data_i[2649] & sel_one_hot_i[20];
  assign data_masked[2648] = data_i[2648] & sel_one_hot_i[20];
  assign data_masked[2647] = data_i[2647] & sel_one_hot_i[20];
  assign data_masked[2646] = data_i[2646] & sel_one_hot_i[20];
  assign data_masked[2645] = data_i[2645] & sel_one_hot_i[20];
  assign data_masked[2644] = data_i[2644] & sel_one_hot_i[20];
  assign data_masked[2643] = data_i[2643] & sel_one_hot_i[20];
  assign data_masked[2642] = data_i[2642] & sel_one_hot_i[20];
  assign data_masked[2641] = data_i[2641] & sel_one_hot_i[20];
  assign data_masked[2640] = data_i[2640] & sel_one_hot_i[20];
  assign data_masked[2639] = data_i[2639] & sel_one_hot_i[20];
  assign data_masked[2638] = data_i[2638] & sel_one_hot_i[20];
  assign data_masked[2637] = data_i[2637] & sel_one_hot_i[20];
  assign data_masked[2636] = data_i[2636] & sel_one_hot_i[20];
  assign data_masked[2635] = data_i[2635] & sel_one_hot_i[20];
  assign data_masked[2634] = data_i[2634] & sel_one_hot_i[20];
  assign data_masked[2633] = data_i[2633] & sel_one_hot_i[20];
  assign data_masked[2632] = data_i[2632] & sel_one_hot_i[20];
  assign data_masked[2631] = data_i[2631] & sel_one_hot_i[20];
  assign data_masked[2630] = data_i[2630] & sel_one_hot_i[20];
  assign data_masked[2629] = data_i[2629] & sel_one_hot_i[20];
  assign data_masked[2628] = data_i[2628] & sel_one_hot_i[20];
  assign data_masked[2627] = data_i[2627] & sel_one_hot_i[20];
  assign data_masked[2626] = data_i[2626] & sel_one_hot_i[20];
  assign data_masked[2625] = data_i[2625] & sel_one_hot_i[20];
  assign data_masked[2624] = data_i[2624] & sel_one_hot_i[20];
  assign data_masked[2623] = data_i[2623] & sel_one_hot_i[20];
  assign data_masked[2622] = data_i[2622] & sel_one_hot_i[20];
  assign data_masked[2621] = data_i[2621] & sel_one_hot_i[20];
  assign data_masked[2620] = data_i[2620] & sel_one_hot_i[20];
  assign data_masked[2619] = data_i[2619] & sel_one_hot_i[20];
  assign data_masked[2618] = data_i[2618] & sel_one_hot_i[20];
  assign data_masked[2617] = data_i[2617] & sel_one_hot_i[20];
  assign data_masked[2616] = data_i[2616] & sel_one_hot_i[20];
  assign data_masked[2615] = data_i[2615] & sel_one_hot_i[20];
  assign data_masked[2614] = data_i[2614] & sel_one_hot_i[20];
  assign data_masked[2613] = data_i[2613] & sel_one_hot_i[20];
  assign data_masked[2612] = data_i[2612] & sel_one_hot_i[20];
  assign data_masked[2611] = data_i[2611] & sel_one_hot_i[20];
  assign data_masked[2610] = data_i[2610] & sel_one_hot_i[20];
  assign data_masked[2609] = data_i[2609] & sel_one_hot_i[20];
  assign data_masked[2608] = data_i[2608] & sel_one_hot_i[20];
  assign data_masked[2607] = data_i[2607] & sel_one_hot_i[20];
  assign data_masked[2606] = data_i[2606] & sel_one_hot_i[20];
  assign data_masked[2605] = data_i[2605] & sel_one_hot_i[20];
  assign data_masked[2604] = data_i[2604] & sel_one_hot_i[20];
  assign data_masked[2603] = data_i[2603] & sel_one_hot_i[20];
  assign data_masked[2602] = data_i[2602] & sel_one_hot_i[20];
  assign data_masked[2601] = data_i[2601] & sel_one_hot_i[20];
  assign data_masked[2600] = data_i[2600] & sel_one_hot_i[20];
  assign data_masked[2599] = data_i[2599] & sel_one_hot_i[20];
  assign data_masked[2598] = data_i[2598] & sel_one_hot_i[20];
  assign data_masked[2597] = data_i[2597] & sel_one_hot_i[20];
  assign data_masked[2596] = data_i[2596] & sel_one_hot_i[20];
  assign data_masked[2595] = data_i[2595] & sel_one_hot_i[20];
  assign data_masked[2594] = data_i[2594] & sel_one_hot_i[20];
  assign data_masked[2593] = data_i[2593] & sel_one_hot_i[20];
  assign data_masked[2592] = data_i[2592] & sel_one_hot_i[20];
  assign data_masked[2591] = data_i[2591] & sel_one_hot_i[20];
  assign data_masked[2590] = data_i[2590] & sel_one_hot_i[20];
  assign data_masked[2589] = data_i[2589] & sel_one_hot_i[20];
  assign data_masked[2588] = data_i[2588] & sel_one_hot_i[20];
  assign data_masked[2587] = data_i[2587] & sel_one_hot_i[20];
  assign data_masked[2586] = data_i[2586] & sel_one_hot_i[20];
  assign data_masked[2585] = data_i[2585] & sel_one_hot_i[20];
  assign data_masked[2584] = data_i[2584] & sel_one_hot_i[20];
  assign data_masked[2583] = data_i[2583] & sel_one_hot_i[20];
  assign data_masked[2582] = data_i[2582] & sel_one_hot_i[20];
  assign data_masked[2581] = data_i[2581] & sel_one_hot_i[20];
  assign data_masked[2580] = data_i[2580] & sel_one_hot_i[20];
  assign data_masked[2579] = data_i[2579] & sel_one_hot_i[20];
  assign data_masked[2578] = data_i[2578] & sel_one_hot_i[20];
  assign data_masked[2577] = data_i[2577] & sel_one_hot_i[20];
  assign data_masked[2576] = data_i[2576] & sel_one_hot_i[20];
  assign data_masked[2575] = data_i[2575] & sel_one_hot_i[20];
  assign data_masked[2574] = data_i[2574] & sel_one_hot_i[20];
  assign data_masked[2573] = data_i[2573] & sel_one_hot_i[20];
  assign data_masked[2572] = data_i[2572] & sel_one_hot_i[20];
  assign data_masked[2571] = data_i[2571] & sel_one_hot_i[20];
  assign data_masked[2570] = data_i[2570] & sel_one_hot_i[20];
  assign data_masked[2569] = data_i[2569] & sel_one_hot_i[20];
  assign data_masked[2568] = data_i[2568] & sel_one_hot_i[20];
  assign data_masked[2567] = data_i[2567] & sel_one_hot_i[20];
  assign data_masked[2566] = data_i[2566] & sel_one_hot_i[20];
  assign data_masked[2565] = data_i[2565] & sel_one_hot_i[20];
  assign data_masked[2564] = data_i[2564] & sel_one_hot_i[20];
  assign data_masked[2563] = data_i[2563] & sel_one_hot_i[20];
  assign data_masked[2562] = data_i[2562] & sel_one_hot_i[20];
  assign data_masked[2561] = data_i[2561] & sel_one_hot_i[20];
  assign data_masked[2560] = data_i[2560] & sel_one_hot_i[20];
  assign data_masked[2815] = data_i[2815] & sel_one_hot_i[21];
  assign data_masked[2814] = data_i[2814] & sel_one_hot_i[21];
  assign data_masked[2813] = data_i[2813] & sel_one_hot_i[21];
  assign data_masked[2812] = data_i[2812] & sel_one_hot_i[21];
  assign data_masked[2811] = data_i[2811] & sel_one_hot_i[21];
  assign data_masked[2810] = data_i[2810] & sel_one_hot_i[21];
  assign data_masked[2809] = data_i[2809] & sel_one_hot_i[21];
  assign data_masked[2808] = data_i[2808] & sel_one_hot_i[21];
  assign data_masked[2807] = data_i[2807] & sel_one_hot_i[21];
  assign data_masked[2806] = data_i[2806] & sel_one_hot_i[21];
  assign data_masked[2805] = data_i[2805] & sel_one_hot_i[21];
  assign data_masked[2804] = data_i[2804] & sel_one_hot_i[21];
  assign data_masked[2803] = data_i[2803] & sel_one_hot_i[21];
  assign data_masked[2802] = data_i[2802] & sel_one_hot_i[21];
  assign data_masked[2801] = data_i[2801] & sel_one_hot_i[21];
  assign data_masked[2800] = data_i[2800] & sel_one_hot_i[21];
  assign data_masked[2799] = data_i[2799] & sel_one_hot_i[21];
  assign data_masked[2798] = data_i[2798] & sel_one_hot_i[21];
  assign data_masked[2797] = data_i[2797] & sel_one_hot_i[21];
  assign data_masked[2796] = data_i[2796] & sel_one_hot_i[21];
  assign data_masked[2795] = data_i[2795] & sel_one_hot_i[21];
  assign data_masked[2794] = data_i[2794] & sel_one_hot_i[21];
  assign data_masked[2793] = data_i[2793] & sel_one_hot_i[21];
  assign data_masked[2792] = data_i[2792] & sel_one_hot_i[21];
  assign data_masked[2791] = data_i[2791] & sel_one_hot_i[21];
  assign data_masked[2790] = data_i[2790] & sel_one_hot_i[21];
  assign data_masked[2789] = data_i[2789] & sel_one_hot_i[21];
  assign data_masked[2788] = data_i[2788] & sel_one_hot_i[21];
  assign data_masked[2787] = data_i[2787] & sel_one_hot_i[21];
  assign data_masked[2786] = data_i[2786] & sel_one_hot_i[21];
  assign data_masked[2785] = data_i[2785] & sel_one_hot_i[21];
  assign data_masked[2784] = data_i[2784] & sel_one_hot_i[21];
  assign data_masked[2783] = data_i[2783] & sel_one_hot_i[21];
  assign data_masked[2782] = data_i[2782] & sel_one_hot_i[21];
  assign data_masked[2781] = data_i[2781] & sel_one_hot_i[21];
  assign data_masked[2780] = data_i[2780] & sel_one_hot_i[21];
  assign data_masked[2779] = data_i[2779] & sel_one_hot_i[21];
  assign data_masked[2778] = data_i[2778] & sel_one_hot_i[21];
  assign data_masked[2777] = data_i[2777] & sel_one_hot_i[21];
  assign data_masked[2776] = data_i[2776] & sel_one_hot_i[21];
  assign data_masked[2775] = data_i[2775] & sel_one_hot_i[21];
  assign data_masked[2774] = data_i[2774] & sel_one_hot_i[21];
  assign data_masked[2773] = data_i[2773] & sel_one_hot_i[21];
  assign data_masked[2772] = data_i[2772] & sel_one_hot_i[21];
  assign data_masked[2771] = data_i[2771] & sel_one_hot_i[21];
  assign data_masked[2770] = data_i[2770] & sel_one_hot_i[21];
  assign data_masked[2769] = data_i[2769] & sel_one_hot_i[21];
  assign data_masked[2768] = data_i[2768] & sel_one_hot_i[21];
  assign data_masked[2767] = data_i[2767] & sel_one_hot_i[21];
  assign data_masked[2766] = data_i[2766] & sel_one_hot_i[21];
  assign data_masked[2765] = data_i[2765] & sel_one_hot_i[21];
  assign data_masked[2764] = data_i[2764] & sel_one_hot_i[21];
  assign data_masked[2763] = data_i[2763] & sel_one_hot_i[21];
  assign data_masked[2762] = data_i[2762] & sel_one_hot_i[21];
  assign data_masked[2761] = data_i[2761] & sel_one_hot_i[21];
  assign data_masked[2760] = data_i[2760] & sel_one_hot_i[21];
  assign data_masked[2759] = data_i[2759] & sel_one_hot_i[21];
  assign data_masked[2758] = data_i[2758] & sel_one_hot_i[21];
  assign data_masked[2757] = data_i[2757] & sel_one_hot_i[21];
  assign data_masked[2756] = data_i[2756] & sel_one_hot_i[21];
  assign data_masked[2755] = data_i[2755] & sel_one_hot_i[21];
  assign data_masked[2754] = data_i[2754] & sel_one_hot_i[21];
  assign data_masked[2753] = data_i[2753] & sel_one_hot_i[21];
  assign data_masked[2752] = data_i[2752] & sel_one_hot_i[21];
  assign data_masked[2751] = data_i[2751] & sel_one_hot_i[21];
  assign data_masked[2750] = data_i[2750] & sel_one_hot_i[21];
  assign data_masked[2749] = data_i[2749] & sel_one_hot_i[21];
  assign data_masked[2748] = data_i[2748] & sel_one_hot_i[21];
  assign data_masked[2747] = data_i[2747] & sel_one_hot_i[21];
  assign data_masked[2746] = data_i[2746] & sel_one_hot_i[21];
  assign data_masked[2745] = data_i[2745] & sel_one_hot_i[21];
  assign data_masked[2744] = data_i[2744] & sel_one_hot_i[21];
  assign data_masked[2743] = data_i[2743] & sel_one_hot_i[21];
  assign data_masked[2742] = data_i[2742] & sel_one_hot_i[21];
  assign data_masked[2741] = data_i[2741] & sel_one_hot_i[21];
  assign data_masked[2740] = data_i[2740] & sel_one_hot_i[21];
  assign data_masked[2739] = data_i[2739] & sel_one_hot_i[21];
  assign data_masked[2738] = data_i[2738] & sel_one_hot_i[21];
  assign data_masked[2737] = data_i[2737] & sel_one_hot_i[21];
  assign data_masked[2736] = data_i[2736] & sel_one_hot_i[21];
  assign data_masked[2735] = data_i[2735] & sel_one_hot_i[21];
  assign data_masked[2734] = data_i[2734] & sel_one_hot_i[21];
  assign data_masked[2733] = data_i[2733] & sel_one_hot_i[21];
  assign data_masked[2732] = data_i[2732] & sel_one_hot_i[21];
  assign data_masked[2731] = data_i[2731] & sel_one_hot_i[21];
  assign data_masked[2730] = data_i[2730] & sel_one_hot_i[21];
  assign data_masked[2729] = data_i[2729] & sel_one_hot_i[21];
  assign data_masked[2728] = data_i[2728] & sel_one_hot_i[21];
  assign data_masked[2727] = data_i[2727] & sel_one_hot_i[21];
  assign data_masked[2726] = data_i[2726] & sel_one_hot_i[21];
  assign data_masked[2725] = data_i[2725] & sel_one_hot_i[21];
  assign data_masked[2724] = data_i[2724] & sel_one_hot_i[21];
  assign data_masked[2723] = data_i[2723] & sel_one_hot_i[21];
  assign data_masked[2722] = data_i[2722] & sel_one_hot_i[21];
  assign data_masked[2721] = data_i[2721] & sel_one_hot_i[21];
  assign data_masked[2720] = data_i[2720] & sel_one_hot_i[21];
  assign data_masked[2719] = data_i[2719] & sel_one_hot_i[21];
  assign data_masked[2718] = data_i[2718] & sel_one_hot_i[21];
  assign data_masked[2717] = data_i[2717] & sel_one_hot_i[21];
  assign data_masked[2716] = data_i[2716] & sel_one_hot_i[21];
  assign data_masked[2715] = data_i[2715] & sel_one_hot_i[21];
  assign data_masked[2714] = data_i[2714] & sel_one_hot_i[21];
  assign data_masked[2713] = data_i[2713] & sel_one_hot_i[21];
  assign data_masked[2712] = data_i[2712] & sel_one_hot_i[21];
  assign data_masked[2711] = data_i[2711] & sel_one_hot_i[21];
  assign data_masked[2710] = data_i[2710] & sel_one_hot_i[21];
  assign data_masked[2709] = data_i[2709] & sel_one_hot_i[21];
  assign data_masked[2708] = data_i[2708] & sel_one_hot_i[21];
  assign data_masked[2707] = data_i[2707] & sel_one_hot_i[21];
  assign data_masked[2706] = data_i[2706] & sel_one_hot_i[21];
  assign data_masked[2705] = data_i[2705] & sel_one_hot_i[21];
  assign data_masked[2704] = data_i[2704] & sel_one_hot_i[21];
  assign data_masked[2703] = data_i[2703] & sel_one_hot_i[21];
  assign data_masked[2702] = data_i[2702] & sel_one_hot_i[21];
  assign data_masked[2701] = data_i[2701] & sel_one_hot_i[21];
  assign data_masked[2700] = data_i[2700] & sel_one_hot_i[21];
  assign data_masked[2699] = data_i[2699] & sel_one_hot_i[21];
  assign data_masked[2698] = data_i[2698] & sel_one_hot_i[21];
  assign data_masked[2697] = data_i[2697] & sel_one_hot_i[21];
  assign data_masked[2696] = data_i[2696] & sel_one_hot_i[21];
  assign data_masked[2695] = data_i[2695] & sel_one_hot_i[21];
  assign data_masked[2694] = data_i[2694] & sel_one_hot_i[21];
  assign data_masked[2693] = data_i[2693] & sel_one_hot_i[21];
  assign data_masked[2692] = data_i[2692] & sel_one_hot_i[21];
  assign data_masked[2691] = data_i[2691] & sel_one_hot_i[21];
  assign data_masked[2690] = data_i[2690] & sel_one_hot_i[21];
  assign data_masked[2689] = data_i[2689] & sel_one_hot_i[21];
  assign data_masked[2688] = data_i[2688] & sel_one_hot_i[21];
  assign data_masked[2943] = data_i[2943] & sel_one_hot_i[22];
  assign data_masked[2942] = data_i[2942] & sel_one_hot_i[22];
  assign data_masked[2941] = data_i[2941] & sel_one_hot_i[22];
  assign data_masked[2940] = data_i[2940] & sel_one_hot_i[22];
  assign data_masked[2939] = data_i[2939] & sel_one_hot_i[22];
  assign data_masked[2938] = data_i[2938] & sel_one_hot_i[22];
  assign data_masked[2937] = data_i[2937] & sel_one_hot_i[22];
  assign data_masked[2936] = data_i[2936] & sel_one_hot_i[22];
  assign data_masked[2935] = data_i[2935] & sel_one_hot_i[22];
  assign data_masked[2934] = data_i[2934] & sel_one_hot_i[22];
  assign data_masked[2933] = data_i[2933] & sel_one_hot_i[22];
  assign data_masked[2932] = data_i[2932] & sel_one_hot_i[22];
  assign data_masked[2931] = data_i[2931] & sel_one_hot_i[22];
  assign data_masked[2930] = data_i[2930] & sel_one_hot_i[22];
  assign data_masked[2929] = data_i[2929] & sel_one_hot_i[22];
  assign data_masked[2928] = data_i[2928] & sel_one_hot_i[22];
  assign data_masked[2927] = data_i[2927] & sel_one_hot_i[22];
  assign data_masked[2926] = data_i[2926] & sel_one_hot_i[22];
  assign data_masked[2925] = data_i[2925] & sel_one_hot_i[22];
  assign data_masked[2924] = data_i[2924] & sel_one_hot_i[22];
  assign data_masked[2923] = data_i[2923] & sel_one_hot_i[22];
  assign data_masked[2922] = data_i[2922] & sel_one_hot_i[22];
  assign data_masked[2921] = data_i[2921] & sel_one_hot_i[22];
  assign data_masked[2920] = data_i[2920] & sel_one_hot_i[22];
  assign data_masked[2919] = data_i[2919] & sel_one_hot_i[22];
  assign data_masked[2918] = data_i[2918] & sel_one_hot_i[22];
  assign data_masked[2917] = data_i[2917] & sel_one_hot_i[22];
  assign data_masked[2916] = data_i[2916] & sel_one_hot_i[22];
  assign data_masked[2915] = data_i[2915] & sel_one_hot_i[22];
  assign data_masked[2914] = data_i[2914] & sel_one_hot_i[22];
  assign data_masked[2913] = data_i[2913] & sel_one_hot_i[22];
  assign data_masked[2912] = data_i[2912] & sel_one_hot_i[22];
  assign data_masked[2911] = data_i[2911] & sel_one_hot_i[22];
  assign data_masked[2910] = data_i[2910] & sel_one_hot_i[22];
  assign data_masked[2909] = data_i[2909] & sel_one_hot_i[22];
  assign data_masked[2908] = data_i[2908] & sel_one_hot_i[22];
  assign data_masked[2907] = data_i[2907] & sel_one_hot_i[22];
  assign data_masked[2906] = data_i[2906] & sel_one_hot_i[22];
  assign data_masked[2905] = data_i[2905] & sel_one_hot_i[22];
  assign data_masked[2904] = data_i[2904] & sel_one_hot_i[22];
  assign data_masked[2903] = data_i[2903] & sel_one_hot_i[22];
  assign data_masked[2902] = data_i[2902] & sel_one_hot_i[22];
  assign data_masked[2901] = data_i[2901] & sel_one_hot_i[22];
  assign data_masked[2900] = data_i[2900] & sel_one_hot_i[22];
  assign data_masked[2899] = data_i[2899] & sel_one_hot_i[22];
  assign data_masked[2898] = data_i[2898] & sel_one_hot_i[22];
  assign data_masked[2897] = data_i[2897] & sel_one_hot_i[22];
  assign data_masked[2896] = data_i[2896] & sel_one_hot_i[22];
  assign data_masked[2895] = data_i[2895] & sel_one_hot_i[22];
  assign data_masked[2894] = data_i[2894] & sel_one_hot_i[22];
  assign data_masked[2893] = data_i[2893] & sel_one_hot_i[22];
  assign data_masked[2892] = data_i[2892] & sel_one_hot_i[22];
  assign data_masked[2891] = data_i[2891] & sel_one_hot_i[22];
  assign data_masked[2890] = data_i[2890] & sel_one_hot_i[22];
  assign data_masked[2889] = data_i[2889] & sel_one_hot_i[22];
  assign data_masked[2888] = data_i[2888] & sel_one_hot_i[22];
  assign data_masked[2887] = data_i[2887] & sel_one_hot_i[22];
  assign data_masked[2886] = data_i[2886] & sel_one_hot_i[22];
  assign data_masked[2885] = data_i[2885] & sel_one_hot_i[22];
  assign data_masked[2884] = data_i[2884] & sel_one_hot_i[22];
  assign data_masked[2883] = data_i[2883] & sel_one_hot_i[22];
  assign data_masked[2882] = data_i[2882] & sel_one_hot_i[22];
  assign data_masked[2881] = data_i[2881] & sel_one_hot_i[22];
  assign data_masked[2880] = data_i[2880] & sel_one_hot_i[22];
  assign data_masked[2879] = data_i[2879] & sel_one_hot_i[22];
  assign data_masked[2878] = data_i[2878] & sel_one_hot_i[22];
  assign data_masked[2877] = data_i[2877] & sel_one_hot_i[22];
  assign data_masked[2876] = data_i[2876] & sel_one_hot_i[22];
  assign data_masked[2875] = data_i[2875] & sel_one_hot_i[22];
  assign data_masked[2874] = data_i[2874] & sel_one_hot_i[22];
  assign data_masked[2873] = data_i[2873] & sel_one_hot_i[22];
  assign data_masked[2872] = data_i[2872] & sel_one_hot_i[22];
  assign data_masked[2871] = data_i[2871] & sel_one_hot_i[22];
  assign data_masked[2870] = data_i[2870] & sel_one_hot_i[22];
  assign data_masked[2869] = data_i[2869] & sel_one_hot_i[22];
  assign data_masked[2868] = data_i[2868] & sel_one_hot_i[22];
  assign data_masked[2867] = data_i[2867] & sel_one_hot_i[22];
  assign data_masked[2866] = data_i[2866] & sel_one_hot_i[22];
  assign data_masked[2865] = data_i[2865] & sel_one_hot_i[22];
  assign data_masked[2864] = data_i[2864] & sel_one_hot_i[22];
  assign data_masked[2863] = data_i[2863] & sel_one_hot_i[22];
  assign data_masked[2862] = data_i[2862] & sel_one_hot_i[22];
  assign data_masked[2861] = data_i[2861] & sel_one_hot_i[22];
  assign data_masked[2860] = data_i[2860] & sel_one_hot_i[22];
  assign data_masked[2859] = data_i[2859] & sel_one_hot_i[22];
  assign data_masked[2858] = data_i[2858] & sel_one_hot_i[22];
  assign data_masked[2857] = data_i[2857] & sel_one_hot_i[22];
  assign data_masked[2856] = data_i[2856] & sel_one_hot_i[22];
  assign data_masked[2855] = data_i[2855] & sel_one_hot_i[22];
  assign data_masked[2854] = data_i[2854] & sel_one_hot_i[22];
  assign data_masked[2853] = data_i[2853] & sel_one_hot_i[22];
  assign data_masked[2852] = data_i[2852] & sel_one_hot_i[22];
  assign data_masked[2851] = data_i[2851] & sel_one_hot_i[22];
  assign data_masked[2850] = data_i[2850] & sel_one_hot_i[22];
  assign data_masked[2849] = data_i[2849] & sel_one_hot_i[22];
  assign data_masked[2848] = data_i[2848] & sel_one_hot_i[22];
  assign data_masked[2847] = data_i[2847] & sel_one_hot_i[22];
  assign data_masked[2846] = data_i[2846] & sel_one_hot_i[22];
  assign data_masked[2845] = data_i[2845] & sel_one_hot_i[22];
  assign data_masked[2844] = data_i[2844] & sel_one_hot_i[22];
  assign data_masked[2843] = data_i[2843] & sel_one_hot_i[22];
  assign data_masked[2842] = data_i[2842] & sel_one_hot_i[22];
  assign data_masked[2841] = data_i[2841] & sel_one_hot_i[22];
  assign data_masked[2840] = data_i[2840] & sel_one_hot_i[22];
  assign data_masked[2839] = data_i[2839] & sel_one_hot_i[22];
  assign data_masked[2838] = data_i[2838] & sel_one_hot_i[22];
  assign data_masked[2837] = data_i[2837] & sel_one_hot_i[22];
  assign data_masked[2836] = data_i[2836] & sel_one_hot_i[22];
  assign data_masked[2835] = data_i[2835] & sel_one_hot_i[22];
  assign data_masked[2834] = data_i[2834] & sel_one_hot_i[22];
  assign data_masked[2833] = data_i[2833] & sel_one_hot_i[22];
  assign data_masked[2832] = data_i[2832] & sel_one_hot_i[22];
  assign data_masked[2831] = data_i[2831] & sel_one_hot_i[22];
  assign data_masked[2830] = data_i[2830] & sel_one_hot_i[22];
  assign data_masked[2829] = data_i[2829] & sel_one_hot_i[22];
  assign data_masked[2828] = data_i[2828] & sel_one_hot_i[22];
  assign data_masked[2827] = data_i[2827] & sel_one_hot_i[22];
  assign data_masked[2826] = data_i[2826] & sel_one_hot_i[22];
  assign data_masked[2825] = data_i[2825] & sel_one_hot_i[22];
  assign data_masked[2824] = data_i[2824] & sel_one_hot_i[22];
  assign data_masked[2823] = data_i[2823] & sel_one_hot_i[22];
  assign data_masked[2822] = data_i[2822] & sel_one_hot_i[22];
  assign data_masked[2821] = data_i[2821] & sel_one_hot_i[22];
  assign data_masked[2820] = data_i[2820] & sel_one_hot_i[22];
  assign data_masked[2819] = data_i[2819] & sel_one_hot_i[22];
  assign data_masked[2818] = data_i[2818] & sel_one_hot_i[22];
  assign data_masked[2817] = data_i[2817] & sel_one_hot_i[22];
  assign data_masked[2816] = data_i[2816] & sel_one_hot_i[22];
  assign data_masked[3071] = data_i[3071] & sel_one_hot_i[23];
  assign data_masked[3070] = data_i[3070] & sel_one_hot_i[23];
  assign data_masked[3069] = data_i[3069] & sel_one_hot_i[23];
  assign data_masked[3068] = data_i[3068] & sel_one_hot_i[23];
  assign data_masked[3067] = data_i[3067] & sel_one_hot_i[23];
  assign data_masked[3066] = data_i[3066] & sel_one_hot_i[23];
  assign data_masked[3065] = data_i[3065] & sel_one_hot_i[23];
  assign data_masked[3064] = data_i[3064] & sel_one_hot_i[23];
  assign data_masked[3063] = data_i[3063] & sel_one_hot_i[23];
  assign data_masked[3062] = data_i[3062] & sel_one_hot_i[23];
  assign data_masked[3061] = data_i[3061] & sel_one_hot_i[23];
  assign data_masked[3060] = data_i[3060] & sel_one_hot_i[23];
  assign data_masked[3059] = data_i[3059] & sel_one_hot_i[23];
  assign data_masked[3058] = data_i[3058] & sel_one_hot_i[23];
  assign data_masked[3057] = data_i[3057] & sel_one_hot_i[23];
  assign data_masked[3056] = data_i[3056] & sel_one_hot_i[23];
  assign data_masked[3055] = data_i[3055] & sel_one_hot_i[23];
  assign data_masked[3054] = data_i[3054] & sel_one_hot_i[23];
  assign data_masked[3053] = data_i[3053] & sel_one_hot_i[23];
  assign data_masked[3052] = data_i[3052] & sel_one_hot_i[23];
  assign data_masked[3051] = data_i[3051] & sel_one_hot_i[23];
  assign data_masked[3050] = data_i[3050] & sel_one_hot_i[23];
  assign data_masked[3049] = data_i[3049] & sel_one_hot_i[23];
  assign data_masked[3048] = data_i[3048] & sel_one_hot_i[23];
  assign data_masked[3047] = data_i[3047] & sel_one_hot_i[23];
  assign data_masked[3046] = data_i[3046] & sel_one_hot_i[23];
  assign data_masked[3045] = data_i[3045] & sel_one_hot_i[23];
  assign data_masked[3044] = data_i[3044] & sel_one_hot_i[23];
  assign data_masked[3043] = data_i[3043] & sel_one_hot_i[23];
  assign data_masked[3042] = data_i[3042] & sel_one_hot_i[23];
  assign data_masked[3041] = data_i[3041] & sel_one_hot_i[23];
  assign data_masked[3040] = data_i[3040] & sel_one_hot_i[23];
  assign data_masked[3039] = data_i[3039] & sel_one_hot_i[23];
  assign data_masked[3038] = data_i[3038] & sel_one_hot_i[23];
  assign data_masked[3037] = data_i[3037] & sel_one_hot_i[23];
  assign data_masked[3036] = data_i[3036] & sel_one_hot_i[23];
  assign data_masked[3035] = data_i[3035] & sel_one_hot_i[23];
  assign data_masked[3034] = data_i[3034] & sel_one_hot_i[23];
  assign data_masked[3033] = data_i[3033] & sel_one_hot_i[23];
  assign data_masked[3032] = data_i[3032] & sel_one_hot_i[23];
  assign data_masked[3031] = data_i[3031] & sel_one_hot_i[23];
  assign data_masked[3030] = data_i[3030] & sel_one_hot_i[23];
  assign data_masked[3029] = data_i[3029] & sel_one_hot_i[23];
  assign data_masked[3028] = data_i[3028] & sel_one_hot_i[23];
  assign data_masked[3027] = data_i[3027] & sel_one_hot_i[23];
  assign data_masked[3026] = data_i[3026] & sel_one_hot_i[23];
  assign data_masked[3025] = data_i[3025] & sel_one_hot_i[23];
  assign data_masked[3024] = data_i[3024] & sel_one_hot_i[23];
  assign data_masked[3023] = data_i[3023] & sel_one_hot_i[23];
  assign data_masked[3022] = data_i[3022] & sel_one_hot_i[23];
  assign data_masked[3021] = data_i[3021] & sel_one_hot_i[23];
  assign data_masked[3020] = data_i[3020] & sel_one_hot_i[23];
  assign data_masked[3019] = data_i[3019] & sel_one_hot_i[23];
  assign data_masked[3018] = data_i[3018] & sel_one_hot_i[23];
  assign data_masked[3017] = data_i[3017] & sel_one_hot_i[23];
  assign data_masked[3016] = data_i[3016] & sel_one_hot_i[23];
  assign data_masked[3015] = data_i[3015] & sel_one_hot_i[23];
  assign data_masked[3014] = data_i[3014] & sel_one_hot_i[23];
  assign data_masked[3013] = data_i[3013] & sel_one_hot_i[23];
  assign data_masked[3012] = data_i[3012] & sel_one_hot_i[23];
  assign data_masked[3011] = data_i[3011] & sel_one_hot_i[23];
  assign data_masked[3010] = data_i[3010] & sel_one_hot_i[23];
  assign data_masked[3009] = data_i[3009] & sel_one_hot_i[23];
  assign data_masked[3008] = data_i[3008] & sel_one_hot_i[23];
  assign data_masked[3007] = data_i[3007] & sel_one_hot_i[23];
  assign data_masked[3006] = data_i[3006] & sel_one_hot_i[23];
  assign data_masked[3005] = data_i[3005] & sel_one_hot_i[23];
  assign data_masked[3004] = data_i[3004] & sel_one_hot_i[23];
  assign data_masked[3003] = data_i[3003] & sel_one_hot_i[23];
  assign data_masked[3002] = data_i[3002] & sel_one_hot_i[23];
  assign data_masked[3001] = data_i[3001] & sel_one_hot_i[23];
  assign data_masked[3000] = data_i[3000] & sel_one_hot_i[23];
  assign data_masked[2999] = data_i[2999] & sel_one_hot_i[23];
  assign data_masked[2998] = data_i[2998] & sel_one_hot_i[23];
  assign data_masked[2997] = data_i[2997] & sel_one_hot_i[23];
  assign data_masked[2996] = data_i[2996] & sel_one_hot_i[23];
  assign data_masked[2995] = data_i[2995] & sel_one_hot_i[23];
  assign data_masked[2994] = data_i[2994] & sel_one_hot_i[23];
  assign data_masked[2993] = data_i[2993] & sel_one_hot_i[23];
  assign data_masked[2992] = data_i[2992] & sel_one_hot_i[23];
  assign data_masked[2991] = data_i[2991] & sel_one_hot_i[23];
  assign data_masked[2990] = data_i[2990] & sel_one_hot_i[23];
  assign data_masked[2989] = data_i[2989] & sel_one_hot_i[23];
  assign data_masked[2988] = data_i[2988] & sel_one_hot_i[23];
  assign data_masked[2987] = data_i[2987] & sel_one_hot_i[23];
  assign data_masked[2986] = data_i[2986] & sel_one_hot_i[23];
  assign data_masked[2985] = data_i[2985] & sel_one_hot_i[23];
  assign data_masked[2984] = data_i[2984] & sel_one_hot_i[23];
  assign data_masked[2983] = data_i[2983] & sel_one_hot_i[23];
  assign data_masked[2982] = data_i[2982] & sel_one_hot_i[23];
  assign data_masked[2981] = data_i[2981] & sel_one_hot_i[23];
  assign data_masked[2980] = data_i[2980] & sel_one_hot_i[23];
  assign data_masked[2979] = data_i[2979] & sel_one_hot_i[23];
  assign data_masked[2978] = data_i[2978] & sel_one_hot_i[23];
  assign data_masked[2977] = data_i[2977] & sel_one_hot_i[23];
  assign data_masked[2976] = data_i[2976] & sel_one_hot_i[23];
  assign data_masked[2975] = data_i[2975] & sel_one_hot_i[23];
  assign data_masked[2974] = data_i[2974] & sel_one_hot_i[23];
  assign data_masked[2973] = data_i[2973] & sel_one_hot_i[23];
  assign data_masked[2972] = data_i[2972] & sel_one_hot_i[23];
  assign data_masked[2971] = data_i[2971] & sel_one_hot_i[23];
  assign data_masked[2970] = data_i[2970] & sel_one_hot_i[23];
  assign data_masked[2969] = data_i[2969] & sel_one_hot_i[23];
  assign data_masked[2968] = data_i[2968] & sel_one_hot_i[23];
  assign data_masked[2967] = data_i[2967] & sel_one_hot_i[23];
  assign data_masked[2966] = data_i[2966] & sel_one_hot_i[23];
  assign data_masked[2965] = data_i[2965] & sel_one_hot_i[23];
  assign data_masked[2964] = data_i[2964] & sel_one_hot_i[23];
  assign data_masked[2963] = data_i[2963] & sel_one_hot_i[23];
  assign data_masked[2962] = data_i[2962] & sel_one_hot_i[23];
  assign data_masked[2961] = data_i[2961] & sel_one_hot_i[23];
  assign data_masked[2960] = data_i[2960] & sel_one_hot_i[23];
  assign data_masked[2959] = data_i[2959] & sel_one_hot_i[23];
  assign data_masked[2958] = data_i[2958] & sel_one_hot_i[23];
  assign data_masked[2957] = data_i[2957] & sel_one_hot_i[23];
  assign data_masked[2956] = data_i[2956] & sel_one_hot_i[23];
  assign data_masked[2955] = data_i[2955] & sel_one_hot_i[23];
  assign data_masked[2954] = data_i[2954] & sel_one_hot_i[23];
  assign data_masked[2953] = data_i[2953] & sel_one_hot_i[23];
  assign data_masked[2952] = data_i[2952] & sel_one_hot_i[23];
  assign data_masked[2951] = data_i[2951] & sel_one_hot_i[23];
  assign data_masked[2950] = data_i[2950] & sel_one_hot_i[23];
  assign data_masked[2949] = data_i[2949] & sel_one_hot_i[23];
  assign data_masked[2948] = data_i[2948] & sel_one_hot_i[23];
  assign data_masked[2947] = data_i[2947] & sel_one_hot_i[23];
  assign data_masked[2946] = data_i[2946] & sel_one_hot_i[23];
  assign data_masked[2945] = data_i[2945] & sel_one_hot_i[23];
  assign data_masked[2944] = data_i[2944] & sel_one_hot_i[23];
  assign data_masked[3199] = data_i[3199] & sel_one_hot_i[24];
  assign data_masked[3198] = data_i[3198] & sel_one_hot_i[24];
  assign data_masked[3197] = data_i[3197] & sel_one_hot_i[24];
  assign data_masked[3196] = data_i[3196] & sel_one_hot_i[24];
  assign data_masked[3195] = data_i[3195] & sel_one_hot_i[24];
  assign data_masked[3194] = data_i[3194] & sel_one_hot_i[24];
  assign data_masked[3193] = data_i[3193] & sel_one_hot_i[24];
  assign data_masked[3192] = data_i[3192] & sel_one_hot_i[24];
  assign data_masked[3191] = data_i[3191] & sel_one_hot_i[24];
  assign data_masked[3190] = data_i[3190] & sel_one_hot_i[24];
  assign data_masked[3189] = data_i[3189] & sel_one_hot_i[24];
  assign data_masked[3188] = data_i[3188] & sel_one_hot_i[24];
  assign data_masked[3187] = data_i[3187] & sel_one_hot_i[24];
  assign data_masked[3186] = data_i[3186] & sel_one_hot_i[24];
  assign data_masked[3185] = data_i[3185] & sel_one_hot_i[24];
  assign data_masked[3184] = data_i[3184] & sel_one_hot_i[24];
  assign data_masked[3183] = data_i[3183] & sel_one_hot_i[24];
  assign data_masked[3182] = data_i[3182] & sel_one_hot_i[24];
  assign data_masked[3181] = data_i[3181] & sel_one_hot_i[24];
  assign data_masked[3180] = data_i[3180] & sel_one_hot_i[24];
  assign data_masked[3179] = data_i[3179] & sel_one_hot_i[24];
  assign data_masked[3178] = data_i[3178] & sel_one_hot_i[24];
  assign data_masked[3177] = data_i[3177] & sel_one_hot_i[24];
  assign data_masked[3176] = data_i[3176] & sel_one_hot_i[24];
  assign data_masked[3175] = data_i[3175] & sel_one_hot_i[24];
  assign data_masked[3174] = data_i[3174] & sel_one_hot_i[24];
  assign data_masked[3173] = data_i[3173] & sel_one_hot_i[24];
  assign data_masked[3172] = data_i[3172] & sel_one_hot_i[24];
  assign data_masked[3171] = data_i[3171] & sel_one_hot_i[24];
  assign data_masked[3170] = data_i[3170] & sel_one_hot_i[24];
  assign data_masked[3169] = data_i[3169] & sel_one_hot_i[24];
  assign data_masked[3168] = data_i[3168] & sel_one_hot_i[24];
  assign data_masked[3167] = data_i[3167] & sel_one_hot_i[24];
  assign data_masked[3166] = data_i[3166] & sel_one_hot_i[24];
  assign data_masked[3165] = data_i[3165] & sel_one_hot_i[24];
  assign data_masked[3164] = data_i[3164] & sel_one_hot_i[24];
  assign data_masked[3163] = data_i[3163] & sel_one_hot_i[24];
  assign data_masked[3162] = data_i[3162] & sel_one_hot_i[24];
  assign data_masked[3161] = data_i[3161] & sel_one_hot_i[24];
  assign data_masked[3160] = data_i[3160] & sel_one_hot_i[24];
  assign data_masked[3159] = data_i[3159] & sel_one_hot_i[24];
  assign data_masked[3158] = data_i[3158] & sel_one_hot_i[24];
  assign data_masked[3157] = data_i[3157] & sel_one_hot_i[24];
  assign data_masked[3156] = data_i[3156] & sel_one_hot_i[24];
  assign data_masked[3155] = data_i[3155] & sel_one_hot_i[24];
  assign data_masked[3154] = data_i[3154] & sel_one_hot_i[24];
  assign data_masked[3153] = data_i[3153] & sel_one_hot_i[24];
  assign data_masked[3152] = data_i[3152] & sel_one_hot_i[24];
  assign data_masked[3151] = data_i[3151] & sel_one_hot_i[24];
  assign data_masked[3150] = data_i[3150] & sel_one_hot_i[24];
  assign data_masked[3149] = data_i[3149] & sel_one_hot_i[24];
  assign data_masked[3148] = data_i[3148] & sel_one_hot_i[24];
  assign data_masked[3147] = data_i[3147] & sel_one_hot_i[24];
  assign data_masked[3146] = data_i[3146] & sel_one_hot_i[24];
  assign data_masked[3145] = data_i[3145] & sel_one_hot_i[24];
  assign data_masked[3144] = data_i[3144] & sel_one_hot_i[24];
  assign data_masked[3143] = data_i[3143] & sel_one_hot_i[24];
  assign data_masked[3142] = data_i[3142] & sel_one_hot_i[24];
  assign data_masked[3141] = data_i[3141] & sel_one_hot_i[24];
  assign data_masked[3140] = data_i[3140] & sel_one_hot_i[24];
  assign data_masked[3139] = data_i[3139] & sel_one_hot_i[24];
  assign data_masked[3138] = data_i[3138] & sel_one_hot_i[24];
  assign data_masked[3137] = data_i[3137] & sel_one_hot_i[24];
  assign data_masked[3136] = data_i[3136] & sel_one_hot_i[24];
  assign data_masked[3135] = data_i[3135] & sel_one_hot_i[24];
  assign data_masked[3134] = data_i[3134] & sel_one_hot_i[24];
  assign data_masked[3133] = data_i[3133] & sel_one_hot_i[24];
  assign data_masked[3132] = data_i[3132] & sel_one_hot_i[24];
  assign data_masked[3131] = data_i[3131] & sel_one_hot_i[24];
  assign data_masked[3130] = data_i[3130] & sel_one_hot_i[24];
  assign data_masked[3129] = data_i[3129] & sel_one_hot_i[24];
  assign data_masked[3128] = data_i[3128] & sel_one_hot_i[24];
  assign data_masked[3127] = data_i[3127] & sel_one_hot_i[24];
  assign data_masked[3126] = data_i[3126] & sel_one_hot_i[24];
  assign data_masked[3125] = data_i[3125] & sel_one_hot_i[24];
  assign data_masked[3124] = data_i[3124] & sel_one_hot_i[24];
  assign data_masked[3123] = data_i[3123] & sel_one_hot_i[24];
  assign data_masked[3122] = data_i[3122] & sel_one_hot_i[24];
  assign data_masked[3121] = data_i[3121] & sel_one_hot_i[24];
  assign data_masked[3120] = data_i[3120] & sel_one_hot_i[24];
  assign data_masked[3119] = data_i[3119] & sel_one_hot_i[24];
  assign data_masked[3118] = data_i[3118] & sel_one_hot_i[24];
  assign data_masked[3117] = data_i[3117] & sel_one_hot_i[24];
  assign data_masked[3116] = data_i[3116] & sel_one_hot_i[24];
  assign data_masked[3115] = data_i[3115] & sel_one_hot_i[24];
  assign data_masked[3114] = data_i[3114] & sel_one_hot_i[24];
  assign data_masked[3113] = data_i[3113] & sel_one_hot_i[24];
  assign data_masked[3112] = data_i[3112] & sel_one_hot_i[24];
  assign data_masked[3111] = data_i[3111] & sel_one_hot_i[24];
  assign data_masked[3110] = data_i[3110] & sel_one_hot_i[24];
  assign data_masked[3109] = data_i[3109] & sel_one_hot_i[24];
  assign data_masked[3108] = data_i[3108] & sel_one_hot_i[24];
  assign data_masked[3107] = data_i[3107] & sel_one_hot_i[24];
  assign data_masked[3106] = data_i[3106] & sel_one_hot_i[24];
  assign data_masked[3105] = data_i[3105] & sel_one_hot_i[24];
  assign data_masked[3104] = data_i[3104] & sel_one_hot_i[24];
  assign data_masked[3103] = data_i[3103] & sel_one_hot_i[24];
  assign data_masked[3102] = data_i[3102] & sel_one_hot_i[24];
  assign data_masked[3101] = data_i[3101] & sel_one_hot_i[24];
  assign data_masked[3100] = data_i[3100] & sel_one_hot_i[24];
  assign data_masked[3099] = data_i[3099] & sel_one_hot_i[24];
  assign data_masked[3098] = data_i[3098] & sel_one_hot_i[24];
  assign data_masked[3097] = data_i[3097] & sel_one_hot_i[24];
  assign data_masked[3096] = data_i[3096] & sel_one_hot_i[24];
  assign data_masked[3095] = data_i[3095] & sel_one_hot_i[24];
  assign data_masked[3094] = data_i[3094] & sel_one_hot_i[24];
  assign data_masked[3093] = data_i[3093] & sel_one_hot_i[24];
  assign data_masked[3092] = data_i[3092] & sel_one_hot_i[24];
  assign data_masked[3091] = data_i[3091] & sel_one_hot_i[24];
  assign data_masked[3090] = data_i[3090] & sel_one_hot_i[24];
  assign data_masked[3089] = data_i[3089] & sel_one_hot_i[24];
  assign data_masked[3088] = data_i[3088] & sel_one_hot_i[24];
  assign data_masked[3087] = data_i[3087] & sel_one_hot_i[24];
  assign data_masked[3086] = data_i[3086] & sel_one_hot_i[24];
  assign data_masked[3085] = data_i[3085] & sel_one_hot_i[24];
  assign data_masked[3084] = data_i[3084] & sel_one_hot_i[24];
  assign data_masked[3083] = data_i[3083] & sel_one_hot_i[24];
  assign data_masked[3082] = data_i[3082] & sel_one_hot_i[24];
  assign data_masked[3081] = data_i[3081] & sel_one_hot_i[24];
  assign data_masked[3080] = data_i[3080] & sel_one_hot_i[24];
  assign data_masked[3079] = data_i[3079] & sel_one_hot_i[24];
  assign data_masked[3078] = data_i[3078] & sel_one_hot_i[24];
  assign data_masked[3077] = data_i[3077] & sel_one_hot_i[24];
  assign data_masked[3076] = data_i[3076] & sel_one_hot_i[24];
  assign data_masked[3075] = data_i[3075] & sel_one_hot_i[24];
  assign data_masked[3074] = data_i[3074] & sel_one_hot_i[24];
  assign data_masked[3073] = data_i[3073] & sel_one_hot_i[24];
  assign data_masked[3072] = data_i[3072] & sel_one_hot_i[24];
  assign data_masked[3327] = data_i[3327] & sel_one_hot_i[25];
  assign data_masked[3326] = data_i[3326] & sel_one_hot_i[25];
  assign data_masked[3325] = data_i[3325] & sel_one_hot_i[25];
  assign data_masked[3324] = data_i[3324] & sel_one_hot_i[25];
  assign data_masked[3323] = data_i[3323] & sel_one_hot_i[25];
  assign data_masked[3322] = data_i[3322] & sel_one_hot_i[25];
  assign data_masked[3321] = data_i[3321] & sel_one_hot_i[25];
  assign data_masked[3320] = data_i[3320] & sel_one_hot_i[25];
  assign data_masked[3319] = data_i[3319] & sel_one_hot_i[25];
  assign data_masked[3318] = data_i[3318] & sel_one_hot_i[25];
  assign data_masked[3317] = data_i[3317] & sel_one_hot_i[25];
  assign data_masked[3316] = data_i[3316] & sel_one_hot_i[25];
  assign data_masked[3315] = data_i[3315] & sel_one_hot_i[25];
  assign data_masked[3314] = data_i[3314] & sel_one_hot_i[25];
  assign data_masked[3313] = data_i[3313] & sel_one_hot_i[25];
  assign data_masked[3312] = data_i[3312] & sel_one_hot_i[25];
  assign data_masked[3311] = data_i[3311] & sel_one_hot_i[25];
  assign data_masked[3310] = data_i[3310] & sel_one_hot_i[25];
  assign data_masked[3309] = data_i[3309] & sel_one_hot_i[25];
  assign data_masked[3308] = data_i[3308] & sel_one_hot_i[25];
  assign data_masked[3307] = data_i[3307] & sel_one_hot_i[25];
  assign data_masked[3306] = data_i[3306] & sel_one_hot_i[25];
  assign data_masked[3305] = data_i[3305] & sel_one_hot_i[25];
  assign data_masked[3304] = data_i[3304] & sel_one_hot_i[25];
  assign data_masked[3303] = data_i[3303] & sel_one_hot_i[25];
  assign data_masked[3302] = data_i[3302] & sel_one_hot_i[25];
  assign data_masked[3301] = data_i[3301] & sel_one_hot_i[25];
  assign data_masked[3300] = data_i[3300] & sel_one_hot_i[25];
  assign data_masked[3299] = data_i[3299] & sel_one_hot_i[25];
  assign data_masked[3298] = data_i[3298] & sel_one_hot_i[25];
  assign data_masked[3297] = data_i[3297] & sel_one_hot_i[25];
  assign data_masked[3296] = data_i[3296] & sel_one_hot_i[25];
  assign data_masked[3295] = data_i[3295] & sel_one_hot_i[25];
  assign data_masked[3294] = data_i[3294] & sel_one_hot_i[25];
  assign data_masked[3293] = data_i[3293] & sel_one_hot_i[25];
  assign data_masked[3292] = data_i[3292] & sel_one_hot_i[25];
  assign data_masked[3291] = data_i[3291] & sel_one_hot_i[25];
  assign data_masked[3290] = data_i[3290] & sel_one_hot_i[25];
  assign data_masked[3289] = data_i[3289] & sel_one_hot_i[25];
  assign data_masked[3288] = data_i[3288] & sel_one_hot_i[25];
  assign data_masked[3287] = data_i[3287] & sel_one_hot_i[25];
  assign data_masked[3286] = data_i[3286] & sel_one_hot_i[25];
  assign data_masked[3285] = data_i[3285] & sel_one_hot_i[25];
  assign data_masked[3284] = data_i[3284] & sel_one_hot_i[25];
  assign data_masked[3283] = data_i[3283] & sel_one_hot_i[25];
  assign data_masked[3282] = data_i[3282] & sel_one_hot_i[25];
  assign data_masked[3281] = data_i[3281] & sel_one_hot_i[25];
  assign data_masked[3280] = data_i[3280] & sel_one_hot_i[25];
  assign data_masked[3279] = data_i[3279] & sel_one_hot_i[25];
  assign data_masked[3278] = data_i[3278] & sel_one_hot_i[25];
  assign data_masked[3277] = data_i[3277] & sel_one_hot_i[25];
  assign data_masked[3276] = data_i[3276] & sel_one_hot_i[25];
  assign data_masked[3275] = data_i[3275] & sel_one_hot_i[25];
  assign data_masked[3274] = data_i[3274] & sel_one_hot_i[25];
  assign data_masked[3273] = data_i[3273] & sel_one_hot_i[25];
  assign data_masked[3272] = data_i[3272] & sel_one_hot_i[25];
  assign data_masked[3271] = data_i[3271] & sel_one_hot_i[25];
  assign data_masked[3270] = data_i[3270] & sel_one_hot_i[25];
  assign data_masked[3269] = data_i[3269] & sel_one_hot_i[25];
  assign data_masked[3268] = data_i[3268] & sel_one_hot_i[25];
  assign data_masked[3267] = data_i[3267] & sel_one_hot_i[25];
  assign data_masked[3266] = data_i[3266] & sel_one_hot_i[25];
  assign data_masked[3265] = data_i[3265] & sel_one_hot_i[25];
  assign data_masked[3264] = data_i[3264] & sel_one_hot_i[25];
  assign data_masked[3263] = data_i[3263] & sel_one_hot_i[25];
  assign data_masked[3262] = data_i[3262] & sel_one_hot_i[25];
  assign data_masked[3261] = data_i[3261] & sel_one_hot_i[25];
  assign data_masked[3260] = data_i[3260] & sel_one_hot_i[25];
  assign data_masked[3259] = data_i[3259] & sel_one_hot_i[25];
  assign data_masked[3258] = data_i[3258] & sel_one_hot_i[25];
  assign data_masked[3257] = data_i[3257] & sel_one_hot_i[25];
  assign data_masked[3256] = data_i[3256] & sel_one_hot_i[25];
  assign data_masked[3255] = data_i[3255] & sel_one_hot_i[25];
  assign data_masked[3254] = data_i[3254] & sel_one_hot_i[25];
  assign data_masked[3253] = data_i[3253] & sel_one_hot_i[25];
  assign data_masked[3252] = data_i[3252] & sel_one_hot_i[25];
  assign data_masked[3251] = data_i[3251] & sel_one_hot_i[25];
  assign data_masked[3250] = data_i[3250] & sel_one_hot_i[25];
  assign data_masked[3249] = data_i[3249] & sel_one_hot_i[25];
  assign data_masked[3248] = data_i[3248] & sel_one_hot_i[25];
  assign data_masked[3247] = data_i[3247] & sel_one_hot_i[25];
  assign data_masked[3246] = data_i[3246] & sel_one_hot_i[25];
  assign data_masked[3245] = data_i[3245] & sel_one_hot_i[25];
  assign data_masked[3244] = data_i[3244] & sel_one_hot_i[25];
  assign data_masked[3243] = data_i[3243] & sel_one_hot_i[25];
  assign data_masked[3242] = data_i[3242] & sel_one_hot_i[25];
  assign data_masked[3241] = data_i[3241] & sel_one_hot_i[25];
  assign data_masked[3240] = data_i[3240] & sel_one_hot_i[25];
  assign data_masked[3239] = data_i[3239] & sel_one_hot_i[25];
  assign data_masked[3238] = data_i[3238] & sel_one_hot_i[25];
  assign data_masked[3237] = data_i[3237] & sel_one_hot_i[25];
  assign data_masked[3236] = data_i[3236] & sel_one_hot_i[25];
  assign data_masked[3235] = data_i[3235] & sel_one_hot_i[25];
  assign data_masked[3234] = data_i[3234] & sel_one_hot_i[25];
  assign data_masked[3233] = data_i[3233] & sel_one_hot_i[25];
  assign data_masked[3232] = data_i[3232] & sel_one_hot_i[25];
  assign data_masked[3231] = data_i[3231] & sel_one_hot_i[25];
  assign data_masked[3230] = data_i[3230] & sel_one_hot_i[25];
  assign data_masked[3229] = data_i[3229] & sel_one_hot_i[25];
  assign data_masked[3228] = data_i[3228] & sel_one_hot_i[25];
  assign data_masked[3227] = data_i[3227] & sel_one_hot_i[25];
  assign data_masked[3226] = data_i[3226] & sel_one_hot_i[25];
  assign data_masked[3225] = data_i[3225] & sel_one_hot_i[25];
  assign data_masked[3224] = data_i[3224] & sel_one_hot_i[25];
  assign data_masked[3223] = data_i[3223] & sel_one_hot_i[25];
  assign data_masked[3222] = data_i[3222] & sel_one_hot_i[25];
  assign data_masked[3221] = data_i[3221] & sel_one_hot_i[25];
  assign data_masked[3220] = data_i[3220] & sel_one_hot_i[25];
  assign data_masked[3219] = data_i[3219] & sel_one_hot_i[25];
  assign data_masked[3218] = data_i[3218] & sel_one_hot_i[25];
  assign data_masked[3217] = data_i[3217] & sel_one_hot_i[25];
  assign data_masked[3216] = data_i[3216] & sel_one_hot_i[25];
  assign data_masked[3215] = data_i[3215] & sel_one_hot_i[25];
  assign data_masked[3214] = data_i[3214] & sel_one_hot_i[25];
  assign data_masked[3213] = data_i[3213] & sel_one_hot_i[25];
  assign data_masked[3212] = data_i[3212] & sel_one_hot_i[25];
  assign data_masked[3211] = data_i[3211] & sel_one_hot_i[25];
  assign data_masked[3210] = data_i[3210] & sel_one_hot_i[25];
  assign data_masked[3209] = data_i[3209] & sel_one_hot_i[25];
  assign data_masked[3208] = data_i[3208] & sel_one_hot_i[25];
  assign data_masked[3207] = data_i[3207] & sel_one_hot_i[25];
  assign data_masked[3206] = data_i[3206] & sel_one_hot_i[25];
  assign data_masked[3205] = data_i[3205] & sel_one_hot_i[25];
  assign data_masked[3204] = data_i[3204] & sel_one_hot_i[25];
  assign data_masked[3203] = data_i[3203] & sel_one_hot_i[25];
  assign data_masked[3202] = data_i[3202] & sel_one_hot_i[25];
  assign data_masked[3201] = data_i[3201] & sel_one_hot_i[25];
  assign data_masked[3200] = data_i[3200] & sel_one_hot_i[25];
  assign data_masked[3455] = data_i[3455] & sel_one_hot_i[26];
  assign data_masked[3454] = data_i[3454] & sel_one_hot_i[26];
  assign data_masked[3453] = data_i[3453] & sel_one_hot_i[26];
  assign data_masked[3452] = data_i[3452] & sel_one_hot_i[26];
  assign data_masked[3451] = data_i[3451] & sel_one_hot_i[26];
  assign data_masked[3450] = data_i[3450] & sel_one_hot_i[26];
  assign data_masked[3449] = data_i[3449] & sel_one_hot_i[26];
  assign data_masked[3448] = data_i[3448] & sel_one_hot_i[26];
  assign data_masked[3447] = data_i[3447] & sel_one_hot_i[26];
  assign data_masked[3446] = data_i[3446] & sel_one_hot_i[26];
  assign data_masked[3445] = data_i[3445] & sel_one_hot_i[26];
  assign data_masked[3444] = data_i[3444] & sel_one_hot_i[26];
  assign data_masked[3443] = data_i[3443] & sel_one_hot_i[26];
  assign data_masked[3442] = data_i[3442] & sel_one_hot_i[26];
  assign data_masked[3441] = data_i[3441] & sel_one_hot_i[26];
  assign data_masked[3440] = data_i[3440] & sel_one_hot_i[26];
  assign data_masked[3439] = data_i[3439] & sel_one_hot_i[26];
  assign data_masked[3438] = data_i[3438] & sel_one_hot_i[26];
  assign data_masked[3437] = data_i[3437] & sel_one_hot_i[26];
  assign data_masked[3436] = data_i[3436] & sel_one_hot_i[26];
  assign data_masked[3435] = data_i[3435] & sel_one_hot_i[26];
  assign data_masked[3434] = data_i[3434] & sel_one_hot_i[26];
  assign data_masked[3433] = data_i[3433] & sel_one_hot_i[26];
  assign data_masked[3432] = data_i[3432] & sel_one_hot_i[26];
  assign data_masked[3431] = data_i[3431] & sel_one_hot_i[26];
  assign data_masked[3430] = data_i[3430] & sel_one_hot_i[26];
  assign data_masked[3429] = data_i[3429] & sel_one_hot_i[26];
  assign data_masked[3428] = data_i[3428] & sel_one_hot_i[26];
  assign data_masked[3427] = data_i[3427] & sel_one_hot_i[26];
  assign data_masked[3426] = data_i[3426] & sel_one_hot_i[26];
  assign data_masked[3425] = data_i[3425] & sel_one_hot_i[26];
  assign data_masked[3424] = data_i[3424] & sel_one_hot_i[26];
  assign data_masked[3423] = data_i[3423] & sel_one_hot_i[26];
  assign data_masked[3422] = data_i[3422] & sel_one_hot_i[26];
  assign data_masked[3421] = data_i[3421] & sel_one_hot_i[26];
  assign data_masked[3420] = data_i[3420] & sel_one_hot_i[26];
  assign data_masked[3419] = data_i[3419] & sel_one_hot_i[26];
  assign data_masked[3418] = data_i[3418] & sel_one_hot_i[26];
  assign data_masked[3417] = data_i[3417] & sel_one_hot_i[26];
  assign data_masked[3416] = data_i[3416] & sel_one_hot_i[26];
  assign data_masked[3415] = data_i[3415] & sel_one_hot_i[26];
  assign data_masked[3414] = data_i[3414] & sel_one_hot_i[26];
  assign data_masked[3413] = data_i[3413] & sel_one_hot_i[26];
  assign data_masked[3412] = data_i[3412] & sel_one_hot_i[26];
  assign data_masked[3411] = data_i[3411] & sel_one_hot_i[26];
  assign data_masked[3410] = data_i[3410] & sel_one_hot_i[26];
  assign data_masked[3409] = data_i[3409] & sel_one_hot_i[26];
  assign data_masked[3408] = data_i[3408] & sel_one_hot_i[26];
  assign data_masked[3407] = data_i[3407] & sel_one_hot_i[26];
  assign data_masked[3406] = data_i[3406] & sel_one_hot_i[26];
  assign data_masked[3405] = data_i[3405] & sel_one_hot_i[26];
  assign data_masked[3404] = data_i[3404] & sel_one_hot_i[26];
  assign data_masked[3403] = data_i[3403] & sel_one_hot_i[26];
  assign data_masked[3402] = data_i[3402] & sel_one_hot_i[26];
  assign data_masked[3401] = data_i[3401] & sel_one_hot_i[26];
  assign data_masked[3400] = data_i[3400] & sel_one_hot_i[26];
  assign data_masked[3399] = data_i[3399] & sel_one_hot_i[26];
  assign data_masked[3398] = data_i[3398] & sel_one_hot_i[26];
  assign data_masked[3397] = data_i[3397] & sel_one_hot_i[26];
  assign data_masked[3396] = data_i[3396] & sel_one_hot_i[26];
  assign data_masked[3395] = data_i[3395] & sel_one_hot_i[26];
  assign data_masked[3394] = data_i[3394] & sel_one_hot_i[26];
  assign data_masked[3393] = data_i[3393] & sel_one_hot_i[26];
  assign data_masked[3392] = data_i[3392] & sel_one_hot_i[26];
  assign data_masked[3391] = data_i[3391] & sel_one_hot_i[26];
  assign data_masked[3390] = data_i[3390] & sel_one_hot_i[26];
  assign data_masked[3389] = data_i[3389] & sel_one_hot_i[26];
  assign data_masked[3388] = data_i[3388] & sel_one_hot_i[26];
  assign data_masked[3387] = data_i[3387] & sel_one_hot_i[26];
  assign data_masked[3386] = data_i[3386] & sel_one_hot_i[26];
  assign data_masked[3385] = data_i[3385] & sel_one_hot_i[26];
  assign data_masked[3384] = data_i[3384] & sel_one_hot_i[26];
  assign data_masked[3383] = data_i[3383] & sel_one_hot_i[26];
  assign data_masked[3382] = data_i[3382] & sel_one_hot_i[26];
  assign data_masked[3381] = data_i[3381] & sel_one_hot_i[26];
  assign data_masked[3380] = data_i[3380] & sel_one_hot_i[26];
  assign data_masked[3379] = data_i[3379] & sel_one_hot_i[26];
  assign data_masked[3378] = data_i[3378] & sel_one_hot_i[26];
  assign data_masked[3377] = data_i[3377] & sel_one_hot_i[26];
  assign data_masked[3376] = data_i[3376] & sel_one_hot_i[26];
  assign data_masked[3375] = data_i[3375] & sel_one_hot_i[26];
  assign data_masked[3374] = data_i[3374] & sel_one_hot_i[26];
  assign data_masked[3373] = data_i[3373] & sel_one_hot_i[26];
  assign data_masked[3372] = data_i[3372] & sel_one_hot_i[26];
  assign data_masked[3371] = data_i[3371] & sel_one_hot_i[26];
  assign data_masked[3370] = data_i[3370] & sel_one_hot_i[26];
  assign data_masked[3369] = data_i[3369] & sel_one_hot_i[26];
  assign data_masked[3368] = data_i[3368] & sel_one_hot_i[26];
  assign data_masked[3367] = data_i[3367] & sel_one_hot_i[26];
  assign data_masked[3366] = data_i[3366] & sel_one_hot_i[26];
  assign data_masked[3365] = data_i[3365] & sel_one_hot_i[26];
  assign data_masked[3364] = data_i[3364] & sel_one_hot_i[26];
  assign data_masked[3363] = data_i[3363] & sel_one_hot_i[26];
  assign data_masked[3362] = data_i[3362] & sel_one_hot_i[26];
  assign data_masked[3361] = data_i[3361] & sel_one_hot_i[26];
  assign data_masked[3360] = data_i[3360] & sel_one_hot_i[26];
  assign data_masked[3359] = data_i[3359] & sel_one_hot_i[26];
  assign data_masked[3358] = data_i[3358] & sel_one_hot_i[26];
  assign data_masked[3357] = data_i[3357] & sel_one_hot_i[26];
  assign data_masked[3356] = data_i[3356] & sel_one_hot_i[26];
  assign data_masked[3355] = data_i[3355] & sel_one_hot_i[26];
  assign data_masked[3354] = data_i[3354] & sel_one_hot_i[26];
  assign data_masked[3353] = data_i[3353] & sel_one_hot_i[26];
  assign data_masked[3352] = data_i[3352] & sel_one_hot_i[26];
  assign data_masked[3351] = data_i[3351] & sel_one_hot_i[26];
  assign data_masked[3350] = data_i[3350] & sel_one_hot_i[26];
  assign data_masked[3349] = data_i[3349] & sel_one_hot_i[26];
  assign data_masked[3348] = data_i[3348] & sel_one_hot_i[26];
  assign data_masked[3347] = data_i[3347] & sel_one_hot_i[26];
  assign data_masked[3346] = data_i[3346] & sel_one_hot_i[26];
  assign data_masked[3345] = data_i[3345] & sel_one_hot_i[26];
  assign data_masked[3344] = data_i[3344] & sel_one_hot_i[26];
  assign data_masked[3343] = data_i[3343] & sel_one_hot_i[26];
  assign data_masked[3342] = data_i[3342] & sel_one_hot_i[26];
  assign data_masked[3341] = data_i[3341] & sel_one_hot_i[26];
  assign data_masked[3340] = data_i[3340] & sel_one_hot_i[26];
  assign data_masked[3339] = data_i[3339] & sel_one_hot_i[26];
  assign data_masked[3338] = data_i[3338] & sel_one_hot_i[26];
  assign data_masked[3337] = data_i[3337] & sel_one_hot_i[26];
  assign data_masked[3336] = data_i[3336] & sel_one_hot_i[26];
  assign data_masked[3335] = data_i[3335] & sel_one_hot_i[26];
  assign data_masked[3334] = data_i[3334] & sel_one_hot_i[26];
  assign data_masked[3333] = data_i[3333] & sel_one_hot_i[26];
  assign data_masked[3332] = data_i[3332] & sel_one_hot_i[26];
  assign data_masked[3331] = data_i[3331] & sel_one_hot_i[26];
  assign data_masked[3330] = data_i[3330] & sel_one_hot_i[26];
  assign data_masked[3329] = data_i[3329] & sel_one_hot_i[26];
  assign data_masked[3328] = data_i[3328] & sel_one_hot_i[26];
  assign data_masked[3583] = data_i[3583] & sel_one_hot_i[27];
  assign data_masked[3582] = data_i[3582] & sel_one_hot_i[27];
  assign data_masked[3581] = data_i[3581] & sel_one_hot_i[27];
  assign data_masked[3580] = data_i[3580] & sel_one_hot_i[27];
  assign data_masked[3579] = data_i[3579] & sel_one_hot_i[27];
  assign data_masked[3578] = data_i[3578] & sel_one_hot_i[27];
  assign data_masked[3577] = data_i[3577] & sel_one_hot_i[27];
  assign data_masked[3576] = data_i[3576] & sel_one_hot_i[27];
  assign data_masked[3575] = data_i[3575] & sel_one_hot_i[27];
  assign data_masked[3574] = data_i[3574] & sel_one_hot_i[27];
  assign data_masked[3573] = data_i[3573] & sel_one_hot_i[27];
  assign data_masked[3572] = data_i[3572] & sel_one_hot_i[27];
  assign data_masked[3571] = data_i[3571] & sel_one_hot_i[27];
  assign data_masked[3570] = data_i[3570] & sel_one_hot_i[27];
  assign data_masked[3569] = data_i[3569] & sel_one_hot_i[27];
  assign data_masked[3568] = data_i[3568] & sel_one_hot_i[27];
  assign data_masked[3567] = data_i[3567] & sel_one_hot_i[27];
  assign data_masked[3566] = data_i[3566] & sel_one_hot_i[27];
  assign data_masked[3565] = data_i[3565] & sel_one_hot_i[27];
  assign data_masked[3564] = data_i[3564] & sel_one_hot_i[27];
  assign data_masked[3563] = data_i[3563] & sel_one_hot_i[27];
  assign data_masked[3562] = data_i[3562] & sel_one_hot_i[27];
  assign data_masked[3561] = data_i[3561] & sel_one_hot_i[27];
  assign data_masked[3560] = data_i[3560] & sel_one_hot_i[27];
  assign data_masked[3559] = data_i[3559] & sel_one_hot_i[27];
  assign data_masked[3558] = data_i[3558] & sel_one_hot_i[27];
  assign data_masked[3557] = data_i[3557] & sel_one_hot_i[27];
  assign data_masked[3556] = data_i[3556] & sel_one_hot_i[27];
  assign data_masked[3555] = data_i[3555] & sel_one_hot_i[27];
  assign data_masked[3554] = data_i[3554] & sel_one_hot_i[27];
  assign data_masked[3553] = data_i[3553] & sel_one_hot_i[27];
  assign data_masked[3552] = data_i[3552] & sel_one_hot_i[27];
  assign data_masked[3551] = data_i[3551] & sel_one_hot_i[27];
  assign data_masked[3550] = data_i[3550] & sel_one_hot_i[27];
  assign data_masked[3549] = data_i[3549] & sel_one_hot_i[27];
  assign data_masked[3548] = data_i[3548] & sel_one_hot_i[27];
  assign data_masked[3547] = data_i[3547] & sel_one_hot_i[27];
  assign data_masked[3546] = data_i[3546] & sel_one_hot_i[27];
  assign data_masked[3545] = data_i[3545] & sel_one_hot_i[27];
  assign data_masked[3544] = data_i[3544] & sel_one_hot_i[27];
  assign data_masked[3543] = data_i[3543] & sel_one_hot_i[27];
  assign data_masked[3542] = data_i[3542] & sel_one_hot_i[27];
  assign data_masked[3541] = data_i[3541] & sel_one_hot_i[27];
  assign data_masked[3540] = data_i[3540] & sel_one_hot_i[27];
  assign data_masked[3539] = data_i[3539] & sel_one_hot_i[27];
  assign data_masked[3538] = data_i[3538] & sel_one_hot_i[27];
  assign data_masked[3537] = data_i[3537] & sel_one_hot_i[27];
  assign data_masked[3536] = data_i[3536] & sel_one_hot_i[27];
  assign data_masked[3535] = data_i[3535] & sel_one_hot_i[27];
  assign data_masked[3534] = data_i[3534] & sel_one_hot_i[27];
  assign data_masked[3533] = data_i[3533] & sel_one_hot_i[27];
  assign data_masked[3532] = data_i[3532] & sel_one_hot_i[27];
  assign data_masked[3531] = data_i[3531] & sel_one_hot_i[27];
  assign data_masked[3530] = data_i[3530] & sel_one_hot_i[27];
  assign data_masked[3529] = data_i[3529] & sel_one_hot_i[27];
  assign data_masked[3528] = data_i[3528] & sel_one_hot_i[27];
  assign data_masked[3527] = data_i[3527] & sel_one_hot_i[27];
  assign data_masked[3526] = data_i[3526] & sel_one_hot_i[27];
  assign data_masked[3525] = data_i[3525] & sel_one_hot_i[27];
  assign data_masked[3524] = data_i[3524] & sel_one_hot_i[27];
  assign data_masked[3523] = data_i[3523] & sel_one_hot_i[27];
  assign data_masked[3522] = data_i[3522] & sel_one_hot_i[27];
  assign data_masked[3521] = data_i[3521] & sel_one_hot_i[27];
  assign data_masked[3520] = data_i[3520] & sel_one_hot_i[27];
  assign data_masked[3519] = data_i[3519] & sel_one_hot_i[27];
  assign data_masked[3518] = data_i[3518] & sel_one_hot_i[27];
  assign data_masked[3517] = data_i[3517] & sel_one_hot_i[27];
  assign data_masked[3516] = data_i[3516] & sel_one_hot_i[27];
  assign data_masked[3515] = data_i[3515] & sel_one_hot_i[27];
  assign data_masked[3514] = data_i[3514] & sel_one_hot_i[27];
  assign data_masked[3513] = data_i[3513] & sel_one_hot_i[27];
  assign data_masked[3512] = data_i[3512] & sel_one_hot_i[27];
  assign data_masked[3511] = data_i[3511] & sel_one_hot_i[27];
  assign data_masked[3510] = data_i[3510] & sel_one_hot_i[27];
  assign data_masked[3509] = data_i[3509] & sel_one_hot_i[27];
  assign data_masked[3508] = data_i[3508] & sel_one_hot_i[27];
  assign data_masked[3507] = data_i[3507] & sel_one_hot_i[27];
  assign data_masked[3506] = data_i[3506] & sel_one_hot_i[27];
  assign data_masked[3505] = data_i[3505] & sel_one_hot_i[27];
  assign data_masked[3504] = data_i[3504] & sel_one_hot_i[27];
  assign data_masked[3503] = data_i[3503] & sel_one_hot_i[27];
  assign data_masked[3502] = data_i[3502] & sel_one_hot_i[27];
  assign data_masked[3501] = data_i[3501] & sel_one_hot_i[27];
  assign data_masked[3500] = data_i[3500] & sel_one_hot_i[27];
  assign data_masked[3499] = data_i[3499] & sel_one_hot_i[27];
  assign data_masked[3498] = data_i[3498] & sel_one_hot_i[27];
  assign data_masked[3497] = data_i[3497] & sel_one_hot_i[27];
  assign data_masked[3496] = data_i[3496] & sel_one_hot_i[27];
  assign data_masked[3495] = data_i[3495] & sel_one_hot_i[27];
  assign data_masked[3494] = data_i[3494] & sel_one_hot_i[27];
  assign data_masked[3493] = data_i[3493] & sel_one_hot_i[27];
  assign data_masked[3492] = data_i[3492] & sel_one_hot_i[27];
  assign data_masked[3491] = data_i[3491] & sel_one_hot_i[27];
  assign data_masked[3490] = data_i[3490] & sel_one_hot_i[27];
  assign data_masked[3489] = data_i[3489] & sel_one_hot_i[27];
  assign data_masked[3488] = data_i[3488] & sel_one_hot_i[27];
  assign data_masked[3487] = data_i[3487] & sel_one_hot_i[27];
  assign data_masked[3486] = data_i[3486] & sel_one_hot_i[27];
  assign data_masked[3485] = data_i[3485] & sel_one_hot_i[27];
  assign data_masked[3484] = data_i[3484] & sel_one_hot_i[27];
  assign data_masked[3483] = data_i[3483] & sel_one_hot_i[27];
  assign data_masked[3482] = data_i[3482] & sel_one_hot_i[27];
  assign data_masked[3481] = data_i[3481] & sel_one_hot_i[27];
  assign data_masked[3480] = data_i[3480] & sel_one_hot_i[27];
  assign data_masked[3479] = data_i[3479] & sel_one_hot_i[27];
  assign data_masked[3478] = data_i[3478] & sel_one_hot_i[27];
  assign data_masked[3477] = data_i[3477] & sel_one_hot_i[27];
  assign data_masked[3476] = data_i[3476] & sel_one_hot_i[27];
  assign data_masked[3475] = data_i[3475] & sel_one_hot_i[27];
  assign data_masked[3474] = data_i[3474] & sel_one_hot_i[27];
  assign data_masked[3473] = data_i[3473] & sel_one_hot_i[27];
  assign data_masked[3472] = data_i[3472] & sel_one_hot_i[27];
  assign data_masked[3471] = data_i[3471] & sel_one_hot_i[27];
  assign data_masked[3470] = data_i[3470] & sel_one_hot_i[27];
  assign data_masked[3469] = data_i[3469] & sel_one_hot_i[27];
  assign data_masked[3468] = data_i[3468] & sel_one_hot_i[27];
  assign data_masked[3467] = data_i[3467] & sel_one_hot_i[27];
  assign data_masked[3466] = data_i[3466] & sel_one_hot_i[27];
  assign data_masked[3465] = data_i[3465] & sel_one_hot_i[27];
  assign data_masked[3464] = data_i[3464] & sel_one_hot_i[27];
  assign data_masked[3463] = data_i[3463] & sel_one_hot_i[27];
  assign data_masked[3462] = data_i[3462] & sel_one_hot_i[27];
  assign data_masked[3461] = data_i[3461] & sel_one_hot_i[27];
  assign data_masked[3460] = data_i[3460] & sel_one_hot_i[27];
  assign data_masked[3459] = data_i[3459] & sel_one_hot_i[27];
  assign data_masked[3458] = data_i[3458] & sel_one_hot_i[27];
  assign data_masked[3457] = data_i[3457] & sel_one_hot_i[27];
  assign data_masked[3456] = data_i[3456] & sel_one_hot_i[27];
  assign data_masked[3711] = data_i[3711] & sel_one_hot_i[28];
  assign data_masked[3710] = data_i[3710] & sel_one_hot_i[28];
  assign data_masked[3709] = data_i[3709] & sel_one_hot_i[28];
  assign data_masked[3708] = data_i[3708] & sel_one_hot_i[28];
  assign data_masked[3707] = data_i[3707] & sel_one_hot_i[28];
  assign data_masked[3706] = data_i[3706] & sel_one_hot_i[28];
  assign data_masked[3705] = data_i[3705] & sel_one_hot_i[28];
  assign data_masked[3704] = data_i[3704] & sel_one_hot_i[28];
  assign data_masked[3703] = data_i[3703] & sel_one_hot_i[28];
  assign data_masked[3702] = data_i[3702] & sel_one_hot_i[28];
  assign data_masked[3701] = data_i[3701] & sel_one_hot_i[28];
  assign data_masked[3700] = data_i[3700] & sel_one_hot_i[28];
  assign data_masked[3699] = data_i[3699] & sel_one_hot_i[28];
  assign data_masked[3698] = data_i[3698] & sel_one_hot_i[28];
  assign data_masked[3697] = data_i[3697] & sel_one_hot_i[28];
  assign data_masked[3696] = data_i[3696] & sel_one_hot_i[28];
  assign data_masked[3695] = data_i[3695] & sel_one_hot_i[28];
  assign data_masked[3694] = data_i[3694] & sel_one_hot_i[28];
  assign data_masked[3693] = data_i[3693] & sel_one_hot_i[28];
  assign data_masked[3692] = data_i[3692] & sel_one_hot_i[28];
  assign data_masked[3691] = data_i[3691] & sel_one_hot_i[28];
  assign data_masked[3690] = data_i[3690] & sel_one_hot_i[28];
  assign data_masked[3689] = data_i[3689] & sel_one_hot_i[28];
  assign data_masked[3688] = data_i[3688] & sel_one_hot_i[28];
  assign data_masked[3687] = data_i[3687] & sel_one_hot_i[28];
  assign data_masked[3686] = data_i[3686] & sel_one_hot_i[28];
  assign data_masked[3685] = data_i[3685] & sel_one_hot_i[28];
  assign data_masked[3684] = data_i[3684] & sel_one_hot_i[28];
  assign data_masked[3683] = data_i[3683] & sel_one_hot_i[28];
  assign data_masked[3682] = data_i[3682] & sel_one_hot_i[28];
  assign data_masked[3681] = data_i[3681] & sel_one_hot_i[28];
  assign data_masked[3680] = data_i[3680] & sel_one_hot_i[28];
  assign data_masked[3679] = data_i[3679] & sel_one_hot_i[28];
  assign data_masked[3678] = data_i[3678] & sel_one_hot_i[28];
  assign data_masked[3677] = data_i[3677] & sel_one_hot_i[28];
  assign data_masked[3676] = data_i[3676] & sel_one_hot_i[28];
  assign data_masked[3675] = data_i[3675] & sel_one_hot_i[28];
  assign data_masked[3674] = data_i[3674] & sel_one_hot_i[28];
  assign data_masked[3673] = data_i[3673] & sel_one_hot_i[28];
  assign data_masked[3672] = data_i[3672] & sel_one_hot_i[28];
  assign data_masked[3671] = data_i[3671] & sel_one_hot_i[28];
  assign data_masked[3670] = data_i[3670] & sel_one_hot_i[28];
  assign data_masked[3669] = data_i[3669] & sel_one_hot_i[28];
  assign data_masked[3668] = data_i[3668] & sel_one_hot_i[28];
  assign data_masked[3667] = data_i[3667] & sel_one_hot_i[28];
  assign data_masked[3666] = data_i[3666] & sel_one_hot_i[28];
  assign data_masked[3665] = data_i[3665] & sel_one_hot_i[28];
  assign data_masked[3664] = data_i[3664] & sel_one_hot_i[28];
  assign data_masked[3663] = data_i[3663] & sel_one_hot_i[28];
  assign data_masked[3662] = data_i[3662] & sel_one_hot_i[28];
  assign data_masked[3661] = data_i[3661] & sel_one_hot_i[28];
  assign data_masked[3660] = data_i[3660] & sel_one_hot_i[28];
  assign data_masked[3659] = data_i[3659] & sel_one_hot_i[28];
  assign data_masked[3658] = data_i[3658] & sel_one_hot_i[28];
  assign data_masked[3657] = data_i[3657] & sel_one_hot_i[28];
  assign data_masked[3656] = data_i[3656] & sel_one_hot_i[28];
  assign data_masked[3655] = data_i[3655] & sel_one_hot_i[28];
  assign data_masked[3654] = data_i[3654] & sel_one_hot_i[28];
  assign data_masked[3653] = data_i[3653] & sel_one_hot_i[28];
  assign data_masked[3652] = data_i[3652] & sel_one_hot_i[28];
  assign data_masked[3651] = data_i[3651] & sel_one_hot_i[28];
  assign data_masked[3650] = data_i[3650] & sel_one_hot_i[28];
  assign data_masked[3649] = data_i[3649] & sel_one_hot_i[28];
  assign data_masked[3648] = data_i[3648] & sel_one_hot_i[28];
  assign data_masked[3647] = data_i[3647] & sel_one_hot_i[28];
  assign data_masked[3646] = data_i[3646] & sel_one_hot_i[28];
  assign data_masked[3645] = data_i[3645] & sel_one_hot_i[28];
  assign data_masked[3644] = data_i[3644] & sel_one_hot_i[28];
  assign data_masked[3643] = data_i[3643] & sel_one_hot_i[28];
  assign data_masked[3642] = data_i[3642] & sel_one_hot_i[28];
  assign data_masked[3641] = data_i[3641] & sel_one_hot_i[28];
  assign data_masked[3640] = data_i[3640] & sel_one_hot_i[28];
  assign data_masked[3639] = data_i[3639] & sel_one_hot_i[28];
  assign data_masked[3638] = data_i[3638] & sel_one_hot_i[28];
  assign data_masked[3637] = data_i[3637] & sel_one_hot_i[28];
  assign data_masked[3636] = data_i[3636] & sel_one_hot_i[28];
  assign data_masked[3635] = data_i[3635] & sel_one_hot_i[28];
  assign data_masked[3634] = data_i[3634] & sel_one_hot_i[28];
  assign data_masked[3633] = data_i[3633] & sel_one_hot_i[28];
  assign data_masked[3632] = data_i[3632] & sel_one_hot_i[28];
  assign data_masked[3631] = data_i[3631] & sel_one_hot_i[28];
  assign data_masked[3630] = data_i[3630] & sel_one_hot_i[28];
  assign data_masked[3629] = data_i[3629] & sel_one_hot_i[28];
  assign data_masked[3628] = data_i[3628] & sel_one_hot_i[28];
  assign data_masked[3627] = data_i[3627] & sel_one_hot_i[28];
  assign data_masked[3626] = data_i[3626] & sel_one_hot_i[28];
  assign data_masked[3625] = data_i[3625] & sel_one_hot_i[28];
  assign data_masked[3624] = data_i[3624] & sel_one_hot_i[28];
  assign data_masked[3623] = data_i[3623] & sel_one_hot_i[28];
  assign data_masked[3622] = data_i[3622] & sel_one_hot_i[28];
  assign data_masked[3621] = data_i[3621] & sel_one_hot_i[28];
  assign data_masked[3620] = data_i[3620] & sel_one_hot_i[28];
  assign data_masked[3619] = data_i[3619] & sel_one_hot_i[28];
  assign data_masked[3618] = data_i[3618] & sel_one_hot_i[28];
  assign data_masked[3617] = data_i[3617] & sel_one_hot_i[28];
  assign data_masked[3616] = data_i[3616] & sel_one_hot_i[28];
  assign data_masked[3615] = data_i[3615] & sel_one_hot_i[28];
  assign data_masked[3614] = data_i[3614] & sel_one_hot_i[28];
  assign data_masked[3613] = data_i[3613] & sel_one_hot_i[28];
  assign data_masked[3612] = data_i[3612] & sel_one_hot_i[28];
  assign data_masked[3611] = data_i[3611] & sel_one_hot_i[28];
  assign data_masked[3610] = data_i[3610] & sel_one_hot_i[28];
  assign data_masked[3609] = data_i[3609] & sel_one_hot_i[28];
  assign data_masked[3608] = data_i[3608] & sel_one_hot_i[28];
  assign data_masked[3607] = data_i[3607] & sel_one_hot_i[28];
  assign data_masked[3606] = data_i[3606] & sel_one_hot_i[28];
  assign data_masked[3605] = data_i[3605] & sel_one_hot_i[28];
  assign data_masked[3604] = data_i[3604] & sel_one_hot_i[28];
  assign data_masked[3603] = data_i[3603] & sel_one_hot_i[28];
  assign data_masked[3602] = data_i[3602] & sel_one_hot_i[28];
  assign data_masked[3601] = data_i[3601] & sel_one_hot_i[28];
  assign data_masked[3600] = data_i[3600] & sel_one_hot_i[28];
  assign data_masked[3599] = data_i[3599] & sel_one_hot_i[28];
  assign data_masked[3598] = data_i[3598] & sel_one_hot_i[28];
  assign data_masked[3597] = data_i[3597] & sel_one_hot_i[28];
  assign data_masked[3596] = data_i[3596] & sel_one_hot_i[28];
  assign data_masked[3595] = data_i[3595] & sel_one_hot_i[28];
  assign data_masked[3594] = data_i[3594] & sel_one_hot_i[28];
  assign data_masked[3593] = data_i[3593] & sel_one_hot_i[28];
  assign data_masked[3592] = data_i[3592] & sel_one_hot_i[28];
  assign data_masked[3591] = data_i[3591] & sel_one_hot_i[28];
  assign data_masked[3590] = data_i[3590] & sel_one_hot_i[28];
  assign data_masked[3589] = data_i[3589] & sel_one_hot_i[28];
  assign data_masked[3588] = data_i[3588] & sel_one_hot_i[28];
  assign data_masked[3587] = data_i[3587] & sel_one_hot_i[28];
  assign data_masked[3586] = data_i[3586] & sel_one_hot_i[28];
  assign data_masked[3585] = data_i[3585] & sel_one_hot_i[28];
  assign data_masked[3584] = data_i[3584] & sel_one_hot_i[28];
  assign data_masked[3839] = data_i[3839] & sel_one_hot_i[29];
  assign data_masked[3838] = data_i[3838] & sel_one_hot_i[29];
  assign data_masked[3837] = data_i[3837] & sel_one_hot_i[29];
  assign data_masked[3836] = data_i[3836] & sel_one_hot_i[29];
  assign data_masked[3835] = data_i[3835] & sel_one_hot_i[29];
  assign data_masked[3834] = data_i[3834] & sel_one_hot_i[29];
  assign data_masked[3833] = data_i[3833] & sel_one_hot_i[29];
  assign data_masked[3832] = data_i[3832] & sel_one_hot_i[29];
  assign data_masked[3831] = data_i[3831] & sel_one_hot_i[29];
  assign data_masked[3830] = data_i[3830] & sel_one_hot_i[29];
  assign data_masked[3829] = data_i[3829] & sel_one_hot_i[29];
  assign data_masked[3828] = data_i[3828] & sel_one_hot_i[29];
  assign data_masked[3827] = data_i[3827] & sel_one_hot_i[29];
  assign data_masked[3826] = data_i[3826] & sel_one_hot_i[29];
  assign data_masked[3825] = data_i[3825] & sel_one_hot_i[29];
  assign data_masked[3824] = data_i[3824] & sel_one_hot_i[29];
  assign data_masked[3823] = data_i[3823] & sel_one_hot_i[29];
  assign data_masked[3822] = data_i[3822] & sel_one_hot_i[29];
  assign data_masked[3821] = data_i[3821] & sel_one_hot_i[29];
  assign data_masked[3820] = data_i[3820] & sel_one_hot_i[29];
  assign data_masked[3819] = data_i[3819] & sel_one_hot_i[29];
  assign data_masked[3818] = data_i[3818] & sel_one_hot_i[29];
  assign data_masked[3817] = data_i[3817] & sel_one_hot_i[29];
  assign data_masked[3816] = data_i[3816] & sel_one_hot_i[29];
  assign data_masked[3815] = data_i[3815] & sel_one_hot_i[29];
  assign data_masked[3814] = data_i[3814] & sel_one_hot_i[29];
  assign data_masked[3813] = data_i[3813] & sel_one_hot_i[29];
  assign data_masked[3812] = data_i[3812] & sel_one_hot_i[29];
  assign data_masked[3811] = data_i[3811] & sel_one_hot_i[29];
  assign data_masked[3810] = data_i[3810] & sel_one_hot_i[29];
  assign data_masked[3809] = data_i[3809] & sel_one_hot_i[29];
  assign data_masked[3808] = data_i[3808] & sel_one_hot_i[29];
  assign data_masked[3807] = data_i[3807] & sel_one_hot_i[29];
  assign data_masked[3806] = data_i[3806] & sel_one_hot_i[29];
  assign data_masked[3805] = data_i[3805] & sel_one_hot_i[29];
  assign data_masked[3804] = data_i[3804] & sel_one_hot_i[29];
  assign data_masked[3803] = data_i[3803] & sel_one_hot_i[29];
  assign data_masked[3802] = data_i[3802] & sel_one_hot_i[29];
  assign data_masked[3801] = data_i[3801] & sel_one_hot_i[29];
  assign data_masked[3800] = data_i[3800] & sel_one_hot_i[29];
  assign data_masked[3799] = data_i[3799] & sel_one_hot_i[29];
  assign data_masked[3798] = data_i[3798] & sel_one_hot_i[29];
  assign data_masked[3797] = data_i[3797] & sel_one_hot_i[29];
  assign data_masked[3796] = data_i[3796] & sel_one_hot_i[29];
  assign data_masked[3795] = data_i[3795] & sel_one_hot_i[29];
  assign data_masked[3794] = data_i[3794] & sel_one_hot_i[29];
  assign data_masked[3793] = data_i[3793] & sel_one_hot_i[29];
  assign data_masked[3792] = data_i[3792] & sel_one_hot_i[29];
  assign data_masked[3791] = data_i[3791] & sel_one_hot_i[29];
  assign data_masked[3790] = data_i[3790] & sel_one_hot_i[29];
  assign data_masked[3789] = data_i[3789] & sel_one_hot_i[29];
  assign data_masked[3788] = data_i[3788] & sel_one_hot_i[29];
  assign data_masked[3787] = data_i[3787] & sel_one_hot_i[29];
  assign data_masked[3786] = data_i[3786] & sel_one_hot_i[29];
  assign data_masked[3785] = data_i[3785] & sel_one_hot_i[29];
  assign data_masked[3784] = data_i[3784] & sel_one_hot_i[29];
  assign data_masked[3783] = data_i[3783] & sel_one_hot_i[29];
  assign data_masked[3782] = data_i[3782] & sel_one_hot_i[29];
  assign data_masked[3781] = data_i[3781] & sel_one_hot_i[29];
  assign data_masked[3780] = data_i[3780] & sel_one_hot_i[29];
  assign data_masked[3779] = data_i[3779] & sel_one_hot_i[29];
  assign data_masked[3778] = data_i[3778] & sel_one_hot_i[29];
  assign data_masked[3777] = data_i[3777] & sel_one_hot_i[29];
  assign data_masked[3776] = data_i[3776] & sel_one_hot_i[29];
  assign data_masked[3775] = data_i[3775] & sel_one_hot_i[29];
  assign data_masked[3774] = data_i[3774] & sel_one_hot_i[29];
  assign data_masked[3773] = data_i[3773] & sel_one_hot_i[29];
  assign data_masked[3772] = data_i[3772] & sel_one_hot_i[29];
  assign data_masked[3771] = data_i[3771] & sel_one_hot_i[29];
  assign data_masked[3770] = data_i[3770] & sel_one_hot_i[29];
  assign data_masked[3769] = data_i[3769] & sel_one_hot_i[29];
  assign data_masked[3768] = data_i[3768] & sel_one_hot_i[29];
  assign data_masked[3767] = data_i[3767] & sel_one_hot_i[29];
  assign data_masked[3766] = data_i[3766] & sel_one_hot_i[29];
  assign data_masked[3765] = data_i[3765] & sel_one_hot_i[29];
  assign data_masked[3764] = data_i[3764] & sel_one_hot_i[29];
  assign data_masked[3763] = data_i[3763] & sel_one_hot_i[29];
  assign data_masked[3762] = data_i[3762] & sel_one_hot_i[29];
  assign data_masked[3761] = data_i[3761] & sel_one_hot_i[29];
  assign data_masked[3760] = data_i[3760] & sel_one_hot_i[29];
  assign data_masked[3759] = data_i[3759] & sel_one_hot_i[29];
  assign data_masked[3758] = data_i[3758] & sel_one_hot_i[29];
  assign data_masked[3757] = data_i[3757] & sel_one_hot_i[29];
  assign data_masked[3756] = data_i[3756] & sel_one_hot_i[29];
  assign data_masked[3755] = data_i[3755] & sel_one_hot_i[29];
  assign data_masked[3754] = data_i[3754] & sel_one_hot_i[29];
  assign data_masked[3753] = data_i[3753] & sel_one_hot_i[29];
  assign data_masked[3752] = data_i[3752] & sel_one_hot_i[29];
  assign data_masked[3751] = data_i[3751] & sel_one_hot_i[29];
  assign data_masked[3750] = data_i[3750] & sel_one_hot_i[29];
  assign data_masked[3749] = data_i[3749] & sel_one_hot_i[29];
  assign data_masked[3748] = data_i[3748] & sel_one_hot_i[29];
  assign data_masked[3747] = data_i[3747] & sel_one_hot_i[29];
  assign data_masked[3746] = data_i[3746] & sel_one_hot_i[29];
  assign data_masked[3745] = data_i[3745] & sel_one_hot_i[29];
  assign data_masked[3744] = data_i[3744] & sel_one_hot_i[29];
  assign data_masked[3743] = data_i[3743] & sel_one_hot_i[29];
  assign data_masked[3742] = data_i[3742] & sel_one_hot_i[29];
  assign data_masked[3741] = data_i[3741] & sel_one_hot_i[29];
  assign data_masked[3740] = data_i[3740] & sel_one_hot_i[29];
  assign data_masked[3739] = data_i[3739] & sel_one_hot_i[29];
  assign data_masked[3738] = data_i[3738] & sel_one_hot_i[29];
  assign data_masked[3737] = data_i[3737] & sel_one_hot_i[29];
  assign data_masked[3736] = data_i[3736] & sel_one_hot_i[29];
  assign data_masked[3735] = data_i[3735] & sel_one_hot_i[29];
  assign data_masked[3734] = data_i[3734] & sel_one_hot_i[29];
  assign data_masked[3733] = data_i[3733] & sel_one_hot_i[29];
  assign data_masked[3732] = data_i[3732] & sel_one_hot_i[29];
  assign data_masked[3731] = data_i[3731] & sel_one_hot_i[29];
  assign data_masked[3730] = data_i[3730] & sel_one_hot_i[29];
  assign data_masked[3729] = data_i[3729] & sel_one_hot_i[29];
  assign data_masked[3728] = data_i[3728] & sel_one_hot_i[29];
  assign data_masked[3727] = data_i[3727] & sel_one_hot_i[29];
  assign data_masked[3726] = data_i[3726] & sel_one_hot_i[29];
  assign data_masked[3725] = data_i[3725] & sel_one_hot_i[29];
  assign data_masked[3724] = data_i[3724] & sel_one_hot_i[29];
  assign data_masked[3723] = data_i[3723] & sel_one_hot_i[29];
  assign data_masked[3722] = data_i[3722] & sel_one_hot_i[29];
  assign data_masked[3721] = data_i[3721] & sel_one_hot_i[29];
  assign data_masked[3720] = data_i[3720] & sel_one_hot_i[29];
  assign data_masked[3719] = data_i[3719] & sel_one_hot_i[29];
  assign data_masked[3718] = data_i[3718] & sel_one_hot_i[29];
  assign data_masked[3717] = data_i[3717] & sel_one_hot_i[29];
  assign data_masked[3716] = data_i[3716] & sel_one_hot_i[29];
  assign data_masked[3715] = data_i[3715] & sel_one_hot_i[29];
  assign data_masked[3714] = data_i[3714] & sel_one_hot_i[29];
  assign data_masked[3713] = data_i[3713] & sel_one_hot_i[29];
  assign data_masked[3712] = data_i[3712] & sel_one_hot_i[29];
  assign data_masked[3967] = data_i[3967] & sel_one_hot_i[30];
  assign data_masked[3966] = data_i[3966] & sel_one_hot_i[30];
  assign data_masked[3965] = data_i[3965] & sel_one_hot_i[30];
  assign data_masked[3964] = data_i[3964] & sel_one_hot_i[30];
  assign data_masked[3963] = data_i[3963] & sel_one_hot_i[30];
  assign data_masked[3962] = data_i[3962] & sel_one_hot_i[30];
  assign data_masked[3961] = data_i[3961] & sel_one_hot_i[30];
  assign data_masked[3960] = data_i[3960] & sel_one_hot_i[30];
  assign data_masked[3959] = data_i[3959] & sel_one_hot_i[30];
  assign data_masked[3958] = data_i[3958] & sel_one_hot_i[30];
  assign data_masked[3957] = data_i[3957] & sel_one_hot_i[30];
  assign data_masked[3956] = data_i[3956] & sel_one_hot_i[30];
  assign data_masked[3955] = data_i[3955] & sel_one_hot_i[30];
  assign data_masked[3954] = data_i[3954] & sel_one_hot_i[30];
  assign data_masked[3953] = data_i[3953] & sel_one_hot_i[30];
  assign data_masked[3952] = data_i[3952] & sel_one_hot_i[30];
  assign data_masked[3951] = data_i[3951] & sel_one_hot_i[30];
  assign data_masked[3950] = data_i[3950] & sel_one_hot_i[30];
  assign data_masked[3949] = data_i[3949] & sel_one_hot_i[30];
  assign data_masked[3948] = data_i[3948] & sel_one_hot_i[30];
  assign data_masked[3947] = data_i[3947] & sel_one_hot_i[30];
  assign data_masked[3946] = data_i[3946] & sel_one_hot_i[30];
  assign data_masked[3945] = data_i[3945] & sel_one_hot_i[30];
  assign data_masked[3944] = data_i[3944] & sel_one_hot_i[30];
  assign data_masked[3943] = data_i[3943] & sel_one_hot_i[30];
  assign data_masked[3942] = data_i[3942] & sel_one_hot_i[30];
  assign data_masked[3941] = data_i[3941] & sel_one_hot_i[30];
  assign data_masked[3940] = data_i[3940] & sel_one_hot_i[30];
  assign data_masked[3939] = data_i[3939] & sel_one_hot_i[30];
  assign data_masked[3938] = data_i[3938] & sel_one_hot_i[30];
  assign data_masked[3937] = data_i[3937] & sel_one_hot_i[30];
  assign data_masked[3936] = data_i[3936] & sel_one_hot_i[30];
  assign data_masked[3935] = data_i[3935] & sel_one_hot_i[30];
  assign data_masked[3934] = data_i[3934] & sel_one_hot_i[30];
  assign data_masked[3933] = data_i[3933] & sel_one_hot_i[30];
  assign data_masked[3932] = data_i[3932] & sel_one_hot_i[30];
  assign data_masked[3931] = data_i[3931] & sel_one_hot_i[30];
  assign data_masked[3930] = data_i[3930] & sel_one_hot_i[30];
  assign data_masked[3929] = data_i[3929] & sel_one_hot_i[30];
  assign data_masked[3928] = data_i[3928] & sel_one_hot_i[30];
  assign data_masked[3927] = data_i[3927] & sel_one_hot_i[30];
  assign data_masked[3926] = data_i[3926] & sel_one_hot_i[30];
  assign data_masked[3925] = data_i[3925] & sel_one_hot_i[30];
  assign data_masked[3924] = data_i[3924] & sel_one_hot_i[30];
  assign data_masked[3923] = data_i[3923] & sel_one_hot_i[30];
  assign data_masked[3922] = data_i[3922] & sel_one_hot_i[30];
  assign data_masked[3921] = data_i[3921] & sel_one_hot_i[30];
  assign data_masked[3920] = data_i[3920] & sel_one_hot_i[30];
  assign data_masked[3919] = data_i[3919] & sel_one_hot_i[30];
  assign data_masked[3918] = data_i[3918] & sel_one_hot_i[30];
  assign data_masked[3917] = data_i[3917] & sel_one_hot_i[30];
  assign data_masked[3916] = data_i[3916] & sel_one_hot_i[30];
  assign data_masked[3915] = data_i[3915] & sel_one_hot_i[30];
  assign data_masked[3914] = data_i[3914] & sel_one_hot_i[30];
  assign data_masked[3913] = data_i[3913] & sel_one_hot_i[30];
  assign data_masked[3912] = data_i[3912] & sel_one_hot_i[30];
  assign data_masked[3911] = data_i[3911] & sel_one_hot_i[30];
  assign data_masked[3910] = data_i[3910] & sel_one_hot_i[30];
  assign data_masked[3909] = data_i[3909] & sel_one_hot_i[30];
  assign data_masked[3908] = data_i[3908] & sel_one_hot_i[30];
  assign data_masked[3907] = data_i[3907] & sel_one_hot_i[30];
  assign data_masked[3906] = data_i[3906] & sel_one_hot_i[30];
  assign data_masked[3905] = data_i[3905] & sel_one_hot_i[30];
  assign data_masked[3904] = data_i[3904] & sel_one_hot_i[30];
  assign data_masked[3903] = data_i[3903] & sel_one_hot_i[30];
  assign data_masked[3902] = data_i[3902] & sel_one_hot_i[30];
  assign data_masked[3901] = data_i[3901] & sel_one_hot_i[30];
  assign data_masked[3900] = data_i[3900] & sel_one_hot_i[30];
  assign data_masked[3899] = data_i[3899] & sel_one_hot_i[30];
  assign data_masked[3898] = data_i[3898] & sel_one_hot_i[30];
  assign data_masked[3897] = data_i[3897] & sel_one_hot_i[30];
  assign data_masked[3896] = data_i[3896] & sel_one_hot_i[30];
  assign data_masked[3895] = data_i[3895] & sel_one_hot_i[30];
  assign data_masked[3894] = data_i[3894] & sel_one_hot_i[30];
  assign data_masked[3893] = data_i[3893] & sel_one_hot_i[30];
  assign data_masked[3892] = data_i[3892] & sel_one_hot_i[30];
  assign data_masked[3891] = data_i[3891] & sel_one_hot_i[30];
  assign data_masked[3890] = data_i[3890] & sel_one_hot_i[30];
  assign data_masked[3889] = data_i[3889] & sel_one_hot_i[30];
  assign data_masked[3888] = data_i[3888] & sel_one_hot_i[30];
  assign data_masked[3887] = data_i[3887] & sel_one_hot_i[30];
  assign data_masked[3886] = data_i[3886] & sel_one_hot_i[30];
  assign data_masked[3885] = data_i[3885] & sel_one_hot_i[30];
  assign data_masked[3884] = data_i[3884] & sel_one_hot_i[30];
  assign data_masked[3883] = data_i[3883] & sel_one_hot_i[30];
  assign data_masked[3882] = data_i[3882] & sel_one_hot_i[30];
  assign data_masked[3881] = data_i[3881] & sel_one_hot_i[30];
  assign data_masked[3880] = data_i[3880] & sel_one_hot_i[30];
  assign data_masked[3879] = data_i[3879] & sel_one_hot_i[30];
  assign data_masked[3878] = data_i[3878] & sel_one_hot_i[30];
  assign data_masked[3877] = data_i[3877] & sel_one_hot_i[30];
  assign data_masked[3876] = data_i[3876] & sel_one_hot_i[30];
  assign data_masked[3875] = data_i[3875] & sel_one_hot_i[30];
  assign data_masked[3874] = data_i[3874] & sel_one_hot_i[30];
  assign data_masked[3873] = data_i[3873] & sel_one_hot_i[30];
  assign data_masked[3872] = data_i[3872] & sel_one_hot_i[30];
  assign data_masked[3871] = data_i[3871] & sel_one_hot_i[30];
  assign data_masked[3870] = data_i[3870] & sel_one_hot_i[30];
  assign data_masked[3869] = data_i[3869] & sel_one_hot_i[30];
  assign data_masked[3868] = data_i[3868] & sel_one_hot_i[30];
  assign data_masked[3867] = data_i[3867] & sel_one_hot_i[30];
  assign data_masked[3866] = data_i[3866] & sel_one_hot_i[30];
  assign data_masked[3865] = data_i[3865] & sel_one_hot_i[30];
  assign data_masked[3864] = data_i[3864] & sel_one_hot_i[30];
  assign data_masked[3863] = data_i[3863] & sel_one_hot_i[30];
  assign data_masked[3862] = data_i[3862] & sel_one_hot_i[30];
  assign data_masked[3861] = data_i[3861] & sel_one_hot_i[30];
  assign data_masked[3860] = data_i[3860] & sel_one_hot_i[30];
  assign data_masked[3859] = data_i[3859] & sel_one_hot_i[30];
  assign data_masked[3858] = data_i[3858] & sel_one_hot_i[30];
  assign data_masked[3857] = data_i[3857] & sel_one_hot_i[30];
  assign data_masked[3856] = data_i[3856] & sel_one_hot_i[30];
  assign data_masked[3855] = data_i[3855] & sel_one_hot_i[30];
  assign data_masked[3854] = data_i[3854] & sel_one_hot_i[30];
  assign data_masked[3853] = data_i[3853] & sel_one_hot_i[30];
  assign data_masked[3852] = data_i[3852] & sel_one_hot_i[30];
  assign data_masked[3851] = data_i[3851] & sel_one_hot_i[30];
  assign data_masked[3850] = data_i[3850] & sel_one_hot_i[30];
  assign data_masked[3849] = data_i[3849] & sel_one_hot_i[30];
  assign data_masked[3848] = data_i[3848] & sel_one_hot_i[30];
  assign data_masked[3847] = data_i[3847] & sel_one_hot_i[30];
  assign data_masked[3846] = data_i[3846] & sel_one_hot_i[30];
  assign data_masked[3845] = data_i[3845] & sel_one_hot_i[30];
  assign data_masked[3844] = data_i[3844] & sel_one_hot_i[30];
  assign data_masked[3843] = data_i[3843] & sel_one_hot_i[30];
  assign data_masked[3842] = data_i[3842] & sel_one_hot_i[30];
  assign data_masked[3841] = data_i[3841] & sel_one_hot_i[30];
  assign data_masked[3840] = data_i[3840] & sel_one_hot_i[30];
  assign data_masked[4095] = data_i[4095] & sel_one_hot_i[31];
  assign data_masked[4094] = data_i[4094] & sel_one_hot_i[31];
  assign data_masked[4093] = data_i[4093] & sel_one_hot_i[31];
  assign data_masked[4092] = data_i[4092] & sel_one_hot_i[31];
  assign data_masked[4091] = data_i[4091] & sel_one_hot_i[31];
  assign data_masked[4090] = data_i[4090] & sel_one_hot_i[31];
  assign data_masked[4089] = data_i[4089] & sel_one_hot_i[31];
  assign data_masked[4088] = data_i[4088] & sel_one_hot_i[31];
  assign data_masked[4087] = data_i[4087] & sel_one_hot_i[31];
  assign data_masked[4086] = data_i[4086] & sel_one_hot_i[31];
  assign data_masked[4085] = data_i[4085] & sel_one_hot_i[31];
  assign data_masked[4084] = data_i[4084] & sel_one_hot_i[31];
  assign data_masked[4083] = data_i[4083] & sel_one_hot_i[31];
  assign data_masked[4082] = data_i[4082] & sel_one_hot_i[31];
  assign data_masked[4081] = data_i[4081] & sel_one_hot_i[31];
  assign data_masked[4080] = data_i[4080] & sel_one_hot_i[31];
  assign data_masked[4079] = data_i[4079] & sel_one_hot_i[31];
  assign data_masked[4078] = data_i[4078] & sel_one_hot_i[31];
  assign data_masked[4077] = data_i[4077] & sel_one_hot_i[31];
  assign data_masked[4076] = data_i[4076] & sel_one_hot_i[31];
  assign data_masked[4075] = data_i[4075] & sel_one_hot_i[31];
  assign data_masked[4074] = data_i[4074] & sel_one_hot_i[31];
  assign data_masked[4073] = data_i[4073] & sel_one_hot_i[31];
  assign data_masked[4072] = data_i[4072] & sel_one_hot_i[31];
  assign data_masked[4071] = data_i[4071] & sel_one_hot_i[31];
  assign data_masked[4070] = data_i[4070] & sel_one_hot_i[31];
  assign data_masked[4069] = data_i[4069] & sel_one_hot_i[31];
  assign data_masked[4068] = data_i[4068] & sel_one_hot_i[31];
  assign data_masked[4067] = data_i[4067] & sel_one_hot_i[31];
  assign data_masked[4066] = data_i[4066] & sel_one_hot_i[31];
  assign data_masked[4065] = data_i[4065] & sel_one_hot_i[31];
  assign data_masked[4064] = data_i[4064] & sel_one_hot_i[31];
  assign data_masked[4063] = data_i[4063] & sel_one_hot_i[31];
  assign data_masked[4062] = data_i[4062] & sel_one_hot_i[31];
  assign data_masked[4061] = data_i[4061] & sel_one_hot_i[31];
  assign data_masked[4060] = data_i[4060] & sel_one_hot_i[31];
  assign data_masked[4059] = data_i[4059] & sel_one_hot_i[31];
  assign data_masked[4058] = data_i[4058] & sel_one_hot_i[31];
  assign data_masked[4057] = data_i[4057] & sel_one_hot_i[31];
  assign data_masked[4056] = data_i[4056] & sel_one_hot_i[31];
  assign data_masked[4055] = data_i[4055] & sel_one_hot_i[31];
  assign data_masked[4054] = data_i[4054] & sel_one_hot_i[31];
  assign data_masked[4053] = data_i[4053] & sel_one_hot_i[31];
  assign data_masked[4052] = data_i[4052] & sel_one_hot_i[31];
  assign data_masked[4051] = data_i[4051] & sel_one_hot_i[31];
  assign data_masked[4050] = data_i[4050] & sel_one_hot_i[31];
  assign data_masked[4049] = data_i[4049] & sel_one_hot_i[31];
  assign data_masked[4048] = data_i[4048] & sel_one_hot_i[31];
  assign data_masked[4047] = data_i[4047] & sel_one_hot_i[31];
  assign data_masked[4046] = data_i[4046] & sel_one_hot_i[31];
  assign data_masked[4045] = data_i[4045] & sel_one_hot_i[31];
  assign data_masked[4044] = data_i[4044] & sel_one_hot_i[31];
  assign data_masked[4043] = data_i[4043] & sel_one_hot_i[31];
  assign data_masked[4042] = data_i[4042] & sel_one_hot_i[31];
  assign data_masked[4041] = data_i[4041] & sel_one_hot_i[31];
  assign data_masked[4040] = data_i[4040] & sel_one_hot_i[31];
  assign data_masked[4039] = data_i[4039] & sel_one_hot_i[31];
  assign data_masked[4038] = data_i[4038] & sel_one_hot_i[31];
  assign data_masked[4037] = data_i[4037] & sel_one_hot_i[31];
  assign data_masked[4036] = data_i[4036] & sel_one_hot_i[31];
  assign data_masked[4035] = data_i[4035] & sel_one_hot_i[31];
  assign data_masked[4034] = data_i[4034] & sel_one_hot_i[31];
  assign data_masked[4033] = data_i[4033] & sel_one_hot_i[31];
  assign data_masked[4032] = data_i[4032] & sel_one_hot_i[31];
  assign data_masked[4031] = data_i[4031] & sel_one_hot_i[31];
  assign data_masked[4030] = data_i[4030] & sel_one_hot_i[31];
  assign data_masked[4029] = data_i[4029] & sel_one_hot_i[31];
  assign data_masked[4028] = data_i[4028] & sel_one_hot_i[31];
  assign data_masked[4027] = data_i[4027] & sel_one_hot_i[31];
  assign data_masked[4026] = data_i[4026] & sel_one_hot_i[31];
  assign data_masked[4025] = data_i[4025] & sel_one_hot_i[31];
  assign data_masked[4024] = data_i[4024] & sel_one_hot_i[31];
  assign data_masked[4023] = data_i[4023] & sel_one_hot_i[31];
  assign data_masked[4022] = data_i[4022] & sel_one_hot_i[31];
  assign data_masked[4021] = data_i[4021] & sel_one_hot_i[31];
  assign data_masked[4020] = data_i[4020] & sel_one_hot_i[31];
  assign data_masked[4019] = data_i[4019] & sel_one_hot_i[31];
  assign data_masked[4018] = data_i[4018] & sel_one_hot_i[31];
  assign data_masked[4017] = data_i[4017] & sel_one_hot_i[31];
  assign data_masked[4016] = data_i[4016] & sel_one_hot_i[31];
  assign data_masked[4015] = data_i[4015] & sel_one_hot_i[31];
  assign data_masked[4014] = data_i[4014] & sel_one_hot_i[31];
  assign data_masked[4013] = data_i[4013] & sel_one_hot_i[31];
  assign data_masked[4012] = data_i[4012] & sel_one_hot_i[31];
  assign data_masked[4011] = data_i[4011] & sel_one_hot_i[31];
  assign data_masked[4010] = data_i[4010] & sel_one_hot_i[31];
  assign data_masked[4009] = data_i[4009] & sel_one_hot_i[31];
  assign data_masked[4008] = data_i[4008] & sel_one_hot_i[31];
  assign data_masked[4007] = data_i[4007] & sel_one_hot_i[31];
  assign data_masked[4006] = data_i[4006] & sel_one_hot_i[31];
  assign data_masked[4005] = data_i[4005] & sel_one_hot_i[31];
  assign data_masked[4004] = data_i[4004] & sel_one_hot_i[31];
  assign data_masked[4003] = data_i[4003] & sel_one_hot_i[31];
  assign data_masked[4002] = data_i[4002] & sel_one_hot_i[31];
  assign data_masked[4001] = data_i[4001] & sel_one_hot_i[31];
  assign data_masked[4000] = data_i[4000] & sel_one_hot_i[31];
  assign data_masked[3999] = data_i[3999] & sel_one_hot_i[31];
  assign data_masked[3998] = data_i[3998] & sel_one_hot_i[31];
  assign data_masked[3997] = data_i[3997] & sel_one_hot_i[31];
  assign data_masked[3996] = data_i[3996] & sel_one_hot_i[31];
  assign data_masked[3995] = data_i[3995] & sel_one_hot_i[31];
  assign data_masked[3994] = data_i[3994] & sel_one_hot_i[31];
  assign data_masked[3993] = data_i[3993] & sel_one_hot_i[31];
  assign data_masked[3992] = data_i[3992] & sel_one_hot_i[31];
  assign data_masked[3991] = data_i[3991] & sel_one_hot_i[31];
  assign data_masked[3990] = data_i[3990] & sel_one_hot_i[31];
  assign data_masked[3989] = data_i[3989] & sel_one_hot_i[31];
  assign data_masked[3988] = data_i[3988] & sel_one_hot_i[31];
  assign data_masked[3987] = data_i[3987] & sel_one_hot_i[31];
  assign data_masked[3986] = data_i[3986] & sel_one_hot_i[31];
  assign data_masked[3985] = data_i[3985] & sel_one_hot_i[31];
  assign data_masked[3984] = data_i[3984] & sel_one_hot_i[31];
  assign data_masked[3983] = data_i[3983] & sel_one_hot_i[31];
  assign data_masked[3982] = data_i[3982] & sel_one_hot_i[31];
  assign data_masked[3981] = data_i[3981] & sel_one_hot_i[31];
  assign data_masked[3980] = data_i[3980] & sel_one_hot_i[31];
  assign data_masked[3979] = data_i[3979] & sel_one_hot_i[31];
  assign data_masked[3978] = data_i[3978] & sel_one_hot_i[31];
  assign data_masked[3977] = data_i[3977] & sel_one_hot_i[31];
  assign data_masked[3976] = data_i[3976] & sel_one_hot_i[31];
  assign data_masked[3975] = data_i[3975] & sel_one_hot_i[31];
  assign data_masked[3974] = data_i[3974] & sel_one_hot_i[31];
  assign data_masked[3973] = data_i[3973] & sel_one_hot_i[31];
  assign data_masked[3972] = data_i[3972] & sel_one_hot_i[31];
  assign data_masked[3971] = data_i[3971] & sel_one_hot_i[31];
  assign data_masked[3970] = data_i[3970] & sel_one_hot_i[31];
  assign data_masked[3969] = data_i[3969] & sel_one_hot_i[31];
  assign data_masked[3968] = data_i[3968] & sel_one_hot_i[31];
  assign data_masked[4223] = data_i[4223] & sel_one_hot_i[32];
  assign data_masked[4222] = data_i[4222] & sel_one_hot_i[32];
  assign data_masked[4221] = data_i[4221] & sel_one_hot_i[32];
  assign data_masked[4220] = data_i[4220] & sel_one_hot_i[32];
  assign data_masked[4219] = data_i[4219] & sel_one_hot_i[32];
  assign data_masked[4218] = data_i[4218] & sel_one_hot_i[32];
  assign data_masked[4217] = data_i[4217] & sel_one_hot_i[32];
  assign data_masked[4216] = data_i[4216] & sel_one_hot_i[32];
  assign data_masked[4215] = data_i[4215] & sel_one_hot_i[32];
  assign data_masked[4214] = data_i[4214] & sel_one_hot_i[32];
  assign data_masked[4213] = data_i[4213] & sel_one_hot_i[32];
  assign data_masked[4212] = data_i[4212] & sel_one_hot_i[32];
  assign data_masked[4211] = data_i[4211] & sel_one_hot_i[32];
  assign data_masked[4210] = data_i[4210] & sel_one_hot_i[32];
  assign data_masked[4209] = data_i[4209] & sel_one_hot_i[32];
  assign data_masked[4208] = data_i[4208] & sel_one_hot_i[32];
  assign data_masked[4207] = data_i[4207] & sel_one_hot_i[32];
  assign data_masked[4206] = data_i[4206] & sel_one_hot_i[32];
  assign data_masked[4205] = data_i[4205] & sel_one_hot_i[32];
  assign data_masked[4204] = data_i[4204] & sel_one_hot_i[32];
  assign data_masked[4203] = data_i[4203] & sel_one_hot_i[32];
  assign data_masked[4202] = data_i[4202] & sel_one_hot_i[32];
  assign data_masked[4201] = data_i[4201] & sel_one_hot_i[32];
  assign data_masked[4200] = data_i[4200] & sel_one_hot_i[32];
  assign data_masked[4199] = data_i[4199] & sel_one_hot_i[32];
  assign data_masked[4198] = data_i[4198] & sel_one_hot_i[32];
  assign data_masked[4197] = data_i[4197] & sel_one_hot_i[32];
  assign data_masked[4196] = data_i[4196] & sel_one_hot_i[32];
  assign data_masked[4195] = data_i[4195] & sel_one_hot_i[32];
  assign data_masked[4194] = data_i[4194] & sel_one_hot_i[32];
  assign data_masked[4193] = data_i[4193] & sel_one_hot_i[32];
  assign data_masked[4192] = data_i[4192] & sel_one_hot_i[32];
  assign data_masked[4191] = data_i[4191] & sel_one_hot_i[32];
  assign data_masked[4190] = data_i[4190] & sel_one_hot_i[32];
  assign data_masked[4189] = data_i[4189] & sel_one_hot_i[32];
  assign data_masked[4188] = data_i[4188] & sel_one_hot_i[32];
  assign data_masked[4187] = data_i[4187] & sel_one_hot_i[32];
  assign data_masked[4186] = data_i[4186] & sel_one_hot_i[32];
  assign data_masked[4185] = data_i[4185] & sel_one_hot_i[32];
  assign data_masked[4184] = data_i[4184] & sel_one_hot_i[32];
  assign data_masked[4183] = data_i[4183] & sel_one_hot_i[32];
  assign data_masked[4182] = data_i[4182] & sel_one_hot_i[32];
  assign data_masked[4181] = data_i[4181] & sel_one_hot_i[32];
  assign data_masked[4180] = data_i[4180] & sel_one_hot_i[32];
  assign data_masked[4179] = data_i[4179] & sel_one_hot_i[32];
  assign data_masked[4178] = data_i[4178] & sel_one_hot_i[32];
  assign data_masked[4177] = data_i[4177] & sel_one_hot_i[32];
  assign data_masked[4176] = data_i[4176] & sel_one_hot_i[32];
  assign data_masked[4175] = data_i[4175] & sel_one_hot_i[32];
  assign data_masked[4174] = data_i[4174] & sel_one_hot_i[32];
  assign data_masked[4173] = data_i[4173] & sel_one_hot_i[32];
  assign data_masked[4172] = data_i[4172] & sel_one_hot_i[32];
  assign data_masked[4171] = data_i[4171] & sel_one_hot_i[32];
  assign data_masked[4170] = data_i[4170] & sel_one_hot_i[32];
  assign data_masked[4169] = data_i[4169] & sel_one_hot_i[32];
  assign data_masked[4168] = data_i[4168] & sel_one_hot_i[32];
  assign data_masked[4167] = data_i[4167] & sel_one_hot_i[32];
  assign data_masked[4166] = data_i[4166] & sel_one_hot_i[32];
  assign data_masked[4165] = data_i[4165] & sel_one_hot_i[32];
  assign data_masked[4164] = data_i[4164] & sel_one_hot_i[32];
  assign data_masked[4163] = data_i[4163] & sel_one_hot_i[32];
  assign data_masked[4162] = data_i[4162] & sel_one_hot_i[32];
  assign data_masked[4161] = data_i[4161] & sel_one_hot_i[32];
  assign data_masked[4160] = data_i[4160] & sel_one_hot_i[32];
  assign data_masked[4159] = data_i[4159] & sel_one_hot_i[32];
  assign data_masked[4158] = data_i[4158] & sel_one_hot_i[32];
  assign data_masked[4157] = data_i[4157] & sel_one_hot_i[32];
  assign data_masked[4156] = data_i[4156] & sel_one_hot_i[32];
  assign data_masked[4155] = data_i[4155] & sel_one_hot_i[32];
  assign data_masked[4154] = data_i[4154] & sel_one_hot_i[32];
  assign data_masked[4153] = data_i[4153] & sel_one_hot_i[32];
  assign data_masked[4152] = data_i[4152] & sel_one_hot_i[32];
  assign data_masked[4151] = data_i[4151] & sel_one_hot_i[32];
  assign data_masked[4150] = data_i[4150] & sel_one_hot_i[32];
  assign data_masked[4149] = data_i[4149] & sel_one_hot_i[32];
  assign data_masked[4148] = data_i[4148] & sel_one_hot_i[32];
  assign data_masked[4147] = data_i[4147] & sel_one_hot_i[32];
  assign data_masked[4146] = data_i[4146] & sel_one_hot_i[32];
  assign data_masked[4145] = data_i[4145] & sel_one_hot_i[32];
  assign data_masked[4144] = data_i[4144] & sel_one_hot_i[32];
  assign data_masked[4143] = data_i[4143] & sel_one_hot_i[32];
  assign data_masked[4142] = data_i[4142] & sel_one_hot_i[32];
  assign data_masked[4141] = data_i[4141] & sel_one_hot_i[32];
  assign data_masked[4140] = data_i[4140] & sel_one_hot_i[32];
  assign data_masked[4139] = data_i[4139] & sel_one_hot_i[32];
  assign data_masked[4138] = data_i[4138] & sel_one_hot_i[32];
  assign data_masked[4137] = data_i[4137] & sel_one_hot_i[32];
  assign data_masked[4136] = data_i[4136] & sel_one_hot_i[32];
  assign data_masked[4135] = data_i[4135] & sel_one_hot_i[32];
  assign data_masked[4134] = data_i[4134] & sel_one_hot_i[32];
  assign data_masked[4133] = data_i[4133] & sel_one_hot_i[32];
  assign data_masked[4132] = data_i[4132] & sel_one_hot_i[32];
  assign data_masked[4131] = data_i[4131] & sel_one_hot_i[32];
  assign data_masked[4130] = data_i[4130] & sel_one_hot_i[32];
  assign data_masked[4129] = data_i[4129] & sel_one_hot_i[32];
  assign data_masked[4128] = data_i[4128] & sel_one_hot_i[32];
  assign data_masked[4127] = data_i[4127] & sel_one_hot_i[32];
  assign data_masked[4126] = data_i[4126] & sel_one_hot_i[32];
  assign data_masked[4125] = data_i[4125] & sel_one_hot_i[32];
  assign data_masked[4124] = data_i[4124] & sel_one_hot_i[32];
  assign data_masked[4123] = data_i[4123] & sel_one_hot_i[32];
  assign data_masked[4122] = data_i[4122] & sel_one_hot_i[32];
  assign data_masked[4121] = data_i[4121] & sel_one_hot_i[32];
  assign data_masked[4120] = data_i[4120] & sel_one_hot_i[32];
  assign data_masked[4119] = data_i[4119] & sel_one_hot_i[32];
  assign data_masked[4118] = data_i[4118] & sel_one_hot_i[32];
  assign data_masked[4117] = data_i[4117] & sel_one_hot_i[32];
  assign data_masked[4116] = data_i[4116] & sel_one_hot_i[32];
  assign data_masked[4115] = data_i[4115] & sel_one_hot_i[32];
  assign data_masked[4114] = data_i[4114] & sel_one_hot_i[32];
  assign data_masked[4113] = data_i[4113] & sel_one_hot_i[32];
  assign data_masked[4112] = data_i[4112] & sel_one_hot_i[32];
  assign data_masked[4111] = data_i[4111] & sel_one_hot_i[32];
  assign data_masked[4110] = data_i[4110] & sel_one_hot_i[32];
  assign data_masked[4109] = data_i[4109] & sel_one_hot_i[32];
  assign data_masked[4108] = data_i[4108] & sel_one_hot_i[32];
  assign data_masked[4107] = data_i[4107] & sel_one_hot_i[32];
  assign data_masked[4106] = data_i[4106] & sel_one_hot_i[32];
  assign data_masked[4105] = data_i[4105] & sel_one_hot_i[32];
  assign data_masked[4104] = data_i[4104] & sel_one_hot_i[32];
  assign data_masked[4103] = data_i[4103] & sel_one_hot_i[32];
  assign data_masked[4102] = data_i[4102] & sel_one_hot_i[32];
  assign data_masked[4101] = data_i[4101] & sel_one_hot_i[32];
  assign data_masked[4100] = data_i[4100] & sel_one_hot_i[32];
  assign data_masked[4099] = data_i[4099] & sel_one_hot_i[32];
  assign data_masked[4098] = data_i[4098] & sel_one_hot_i[32];
  assign data_masked[4097] = data_i[4097] & sel_one_hot_i[32];
  assign data_masked[4096] = data_i[4096] & sel_one_hot_i[32];
  assign data_masked[4351] = data_i[4351] & sel_one_hot_i[33];
  assign data_masked[4350] = data_i[4350] & sel_one_hot_i[33];
  assign data_masked[4349] = data_i[4349] & sel_one_hot_i[33];
  assign data_masked[4348] = data_i[4348] & sel_one_hot_i[33];
  assign data_masked[4347] = data_i[4347] & sel_one_hot_i[33];
  assign data_masked[4346] = data_i[4346] & sel_one_hot_i[33];
  assign data_masked[4345] = data_i[4345] & sel_one_hot_i[33];
  assign data_masked[4344] = data_i[4344] & sel_one_hot_i[33];
  assign data_masked[4343] = data_i[4343] & sel_one_hot_i[33];
  assign data_masked[4342] = data_i[4342] & sel_one_hot_i[33];
  assign data_masked[4341] = data_i[4341] & sel_one_hot_i[33];
  assign data_masked[4340] = data_i[4340] & sel_one_hot_i[33];
  assign data_masked[4339] = data_i[4339] & sel_one_hot_i[33];
  assign data_masked[4338] = data_i[4338] & sel_one_hot_i[33];
  assign data_masked[4337] = data_i[4337] & sel_one_hot_i[33];
  assign data_masked[4336] = data_i[4336] & sel_one_hot_i[33];
  assign data_masked[4335] = data_i[4335] & sel_one_hot_i[33];
  assign data_masked[4334] = data_i[4334] & sel_one_hot_i[33];
  assign data_masked[4333] = data_i[4333] & sel_one_hot_i[33];
  assign data_masked[4332] = data_i[4332] & sel_one_hot_i[33];
  assign data_masked[4331] = data_i[4331] & sel_one_hot_i[33];
  assign data_masked[4330] = data_i[4330] & sel_one_hot_i[33];
  assign data_masked[4329] = data_i[4329] & sel_one_hot_i[33];
  assign data_masked[4328] = data_i[4328] & sel_one_hot_i[33];
  assign data_masked[4327] = data_i[4327] & sel_one_hot_i[33];
  assign data_masked[4326] = data_i[4326] & sel_one_hot_i[33];
  assign data_masked[4325] = data_i[4325] & sel_one_hot_i[33];
  assign data_masked[4324] = data_i[4324] & sel_one_hot_i[33];
  assign data_masked[4323] = data_i[4323] & sel_one_hot_i[33];
  assign data_masked[4322] = data_i[4322] & sel_one_hot_i[33];
  assign data_masked[4321] = data_i[4321] & sel_one_hot_i[33];
  assign data_masked[4320] = data_i[4320] & sel_one_hot_i[33];
  assign data_masked[4319] = data_i[4319] & sel_one_hot_i[33];
  assign data_masked[4318] = data_i[4318] & sel_one_hot_i[33];
  assign data_masked[4317] = data_i[4317] & sel_one_hot_i[33];
  assign data_masked[4316] = data_i[4316] & sel_one_hot_i[33];
  assign data_masked[4315] = data_i[4315] & sel_one_hot_i[33];
  assign data_masked[4314] = data_i[4314] & sel_one_hot_i[33];
  assign data_masked[4313] = data_i[4313] & sel_one_hot_i[33];
  assign data_masked[4312] = data_i[4312] & sel_one_hot_i[33];
  assign data_masked[4311] = data_i[4311] & sel_one_hot_i[33];
  assign data_masked[4310] = data_i[4310] & sel_one_hot_i[33];
  assign data_masked[4309] = data_i[4309] & sel_one_hot_i[33];
  assign data_masked[4308] = data_i[4308] & sel_one_hot_i[33];
  assign data_masked[4307] = data_i[4307] & sel_one_hot_i[33];
  assign data_masked[4306] = data_i[4306] & sel_one_hot_i[33];
  assign data_masked[4305] = data_i[4305] & sel_one_hot_i[33];
  assign data_masked[4304] = data_i[4304] & sel_one_hot_i[33];
  assign data_masked[4303] = data_i[4303] & sel_one_hot_i[33];
  assign data_masked[4302] = data_i[4302] & sel_one_hot_i[33];
  assign data_masked[4301] = data_i[4301] & sel_one_hot_i[33];
  assign data_masked[4300] = data_i[4300] & sel_one_hot_i[33];
  assign data_masked[4299] = data_i[4299] & sel_one_hot_i[33];
  assign data_masked[4298] = data_i[4298] & sel_one_hot_i[33];
  assign data_masked[4297] = data_i[4297] & sel_one_hot_i[33];
  assign data_masked[4296] = data_i[4296] & sel_one_hot_i[33];
  assign data_masked[4295] = data_i[4295] & sel_one_hot_i[33];
  assign data_masked[4294] = data_i[4294] & sel_one_hot_i[33];
  assign data_masked[4293] = data_i[4293] & sel_one_hot_i[33];
  assign data_masked[4292] = data_i[4292] & sel_one_hot_i[33];
  assign data_masked[4291] = data_i[4291] & sel_one_hot_i[33];
  assign data_masked[4290] = data_i[4290] & sel_one_hot_i[33];
  assign data_masked[4289] = data_i[4289] & sel_one_hot_i[33];
  assign data_masked[4288] = data_i[4288] & sel_one_hot_i[33];
  assign data_masked[4287] = data_i[4287] & sel_one_hot_i[33];
  assign data_masked[4286] = data_i[4286] & sel_one_hot_i[33];
  assign data_masked[4285] = data_i[4285] & sel_one_hot_i[33];
  assign data_masked[4284] = data_i[4284] & sel_one_hot_i[33];
  assign data_masked[4283] = data_i[4283] & sel_one_hot_i[33];
  assign data_masked[4282] = data_i[4282] & sel_one_hot_i[33];
  assign data_masked[4281] = data_i[4281] & sel_one_hot_i[33];
  assign data_masked[4280] = data_i[4280] & sel_one_hot_i[33];
  assign data_masked[4279] = data_i[4279] & sel_one_hot_i[33];
  assign data_masked[4278] = data_i[4278] & sel_one_hot_i[33];
  assign data_masked[4277] = data_i[4277] & sel_one_hot_i[33];
  assign data_masked[4276] = data_i[4276] & sel_one_hot_i[33];
  assign data_masked[4275] = data_i[4275] & sel_one_hot_i[33];
  assign data_masked[4274] = data_i[4274] & sel_one_hot_i[33];
  assign data_masked[4273] = data_i[4273] & sel_one_hot_i[33];
  assign data_masked[4272] = data_i[4272] & sel_one_hot_i[33];
  assign data_masked[4271] = data_i[4271] & sel_one_hot_i[33];
  assign data_masked[4270] = data_i[4270] & sel_one_hot_i[33];
  assign data_masked[4269] = data_i[4269] & sel_one_hot_i[33];
  assign data_masked[4268] = data_i[4268] & sel_one_hot_i[33];
  assign data_masked[4267] = data_i[4267] & sel_one_hot_i[33];
  assign data_masked[4266] = data_i[4266] & sel_one_hot_i[33];
  assign data_masked[4265] = data_i[4265] & sel_one_hot_i[33];
  assign data_masked[4264] = data_i[4264] & sel_one_hot_i[33];
  assign data_masked[4263] = data_i[4263] & sel_one_hot_i[33];
  assign data_masked[4262] = data_i[4262] & sel_one_hot_i[33];
  assign data_masked[4261] = data_i[4261] & sel_one_hot_i[33];
  assign data_masked[4260] = data_i[4260] & sel_one_hot_i[33];
  assign data_masked[4259] = data_i[4259] & sel_one_hot_i[33];
  assign data_masked[4258] = data_i[4258] & sel_one_hot_i[33];
  assign data_masked[4257] = data_i[4257] & sel_one_hot_i[33];
  assign data_masked[4256] = data_i[4256] & sel_one_hot_i[33];
  assign data_masked[4255] = data_i[4255] & sel_one_hot_i[33];
  assign data_masked[4254] = data_i[4254] & sel_one_hot_i[33];
  assign data_masked[4253] = data_i[4253] & sel_one_hot_i[33];
  assign data_masked[4252] = data_i[4252] & sel_one_hot_i[33];
  assign data_masked[4251] = data_i[4251] & sel_one_hot_i[33];
  assign data_masked[4250] = data_i[4250] & sel_one_hot_i[33];
  assign data_masked[4249] = data_i[4249] & sel_one_hot_i[33];
  assign data_masked[4248] = data_i[4248] & sel_one_hot_i[33];
  assign data_masked[4247] = data_i[4247] & sel_one_hot_i[33];
  assign data_masked[4246] = data_i[4246] & sel_one_hot_i[33];
  assign data_masked[4245] = data_i[4245] & sel_one_hot_i[33];
  assign data_masked[4244] = data_i[4244] & sel_one_hot_i[33];
  assign data_masked[4243] = data_i[4243] & sel_one_hot_i[33];
  assign data_masked[4242] = data_i[4242] & sel_one_hot_i[33];
  assign data_masked[4241] = data_i[4241] & sel_one_hot_i[33];
  assign data_masked[4240] = data_i[4240] & sel_one_hot_i[33];
  assign data_masked[4239] = data_i[4239] & sel_one_hot_i[33];
  assign data_masked[4238] = data_i[4238] & sel_one_hot_i[33];
  assign data_masked[4237] = data_i[4237] & sel_one_hot_i[33];
  assign data_masked[4236] = data_i[4236] & sel_one_hot_i[33];
  assign data_masked[4235] = data_i[4235] & sel_one_hot_i[33];
  assign data_masked[4234] = data_i[4234] & sel_one_hot_i[33];
  assign data_masked[4233] = data_i[4233] & sel_one_hot_i[33];
  assign data_masked[4232] = data_i[4232] & sel_one_hot_i[33];
  assign data_masked[4231] = data_i[4231] & sel_one_hot_i[33];
  assign data_masked[4230] = data_i[4230] & sel_one_hot_i[33];
  assign data_masked[4229] = data_i[4229] & sel_one_hot_i[33];
  assign data_masked[4228] = data_i[4228] & sel_one_hot_i[33];
  assign data_masked[4227] = data_i[4227] & sel_one_hot_i[33];
  assign data_masked[4226] = data_i[4226] & sel_one_hot_i[33];
  assign data_masked[4225] = data_i[4225] & sel_one_hot_i[33];
  assign data_masked[4224] = data_i[4224] & sel_one_hot_i[33];
  assign data_masked[4479] = data_i[4479] & sel_one_hot_i[34];
  assign data_masked[4478] = data_i[4478] & sel_one_hot_i[34];
  assign data_masked[4477] = data_i[4477] & sel_one_hot_i[34];
  assign data_masked[4476] = data_i[4476] & sel_one_hot_i[34];
  assign data_masked[4475] = data_i[4475] & sel_one_hot_i[34];
  assign data_masked[4474] = data_i[4474] & sel_one_hot_i[34];
  assign data_masked[4473] = data_i[4473] & sel_one_hot_i[34];
  assign data_masked[4472] = data_i[4472] & sel_one_hot_i[34];
  assign data_masked[4471] = data_i[4471] & sel_one_hot_i[34];
  assign data_masked[4470] = data_i[4470] & sel_one_hot_i[34];
  assign data_masked[4469] = data_i[4469] & sel_one_hot_i[34];
  assign data_masked[4468] = data_i[4468] & sel_one_hot_i[34];
  assign data_masked[4467] = data_i[4467] & sel_one_hot_i[34];
  assign data_masked[4466] = data_i[4466] & sel_one_hot_i[34];
  assign data_masked[4465] = data_i[4465] & sel_one_hot_i[34];
  assign data_masked[4464] = data_i[4464] & sel_one_hot_i[34];
  assign data_masked[4463] = data_i[4463] & sel_one_hot_i[34];
  assign data_masked[4462] = data_i[4462] & sel_one_hot_i[34];
  assign data_masked[4461] = data_i[4461] & sel_one_hot_i[34];
  assign data_masked[4460] = data_i[4460] & sel_one_hot_i[34];
  assign data_masked[4459] = data_i[4459] & sel_one_hot_i[34];
  assign data_masked[4458] = data_i[4458] & sel_one_hot_i[34];
  assign data_masked[4457] = data_i[4457] & sel_one_hot_i[34];
  assign data_masked[4456] = data_i[4456] & sel_one_hot_i[34];
  assign data_masked[4455] = data_i[4455] & sel_one_hot_i[34];
  assign data_masked[4454] = data_i[4454] & sel_one_hot_i[34];
  assign data_masked[4453] = data_i[4453] & sel_one_hot_i[34];
  assign data_masked[4452] = data_i[4452] & sel_one_hot_i[34];
  assign data_masked[4451] = data_i[4451] & sel_one_hot_i[34];
  assign data_masked[4450] = data_i[4450] & sel_one_hot_i[34];
  assign data_masked[4449] = data_i[4449] & sel_one_hot_i[34];
  assign data_masked[4448] = data_i[4448] & sel_one_hot_i[34];
  assign data_masked[4447] = data_i[4447] & sel_one_hot_i[34];
  assign data_masked[4446] = data_i[4446] & sel_one_hot_i[34];
  assign data_masked[4445] = data_i[4445] & sel_one_hot_i[34];
  assign data_masked[4444] = data_i[4444] & sel_one_hot_i[34];
  assign data_masked[4443] = data_i[4443] & sel_one_hot_i[34];
  assign data_masked[4442] = data_i[4442] & sel_one_hot_i[34];
  assign data_masked[4441] = data_i[4441] & sel_one_hot_i[34];
  assign data_masked[4440] = data_i[4440] & sel_one_hot_i[34];
  assign data_masked[4439] = data_i[4439] & sel_one_hot_i[34];
  assign data_masked[4438] = data_i[4438] & sel_one_hot_i[34];
  assign data_masked[4437] = data_i[4437] & sel_one_hot_i[34];
  assign data_masked[4436] = data_i[4436] & sel_one_hot_i[34];
  assign data_masked[4435] = data_i[4435] & sel_one_hot_i[34];
  assign data_masked[4434] = data_i[4434] & sel_one_hot_i[34];
  assign data_masked[4433] = data_i[4433] & sel_one_hot_i[34];
  assign data_masked[4432] = data_i[4432] & sel_one_hot_i[34];
  assign data_masked[4431] = data_i[4431] & sel_one_hot_i[34];
  assign data_masked[4430] = data_i[4430] & sel_one_hot_i[34];
  assign data_masked[4429] = data_i[4429] & sel_one_hot_i[34];
  assign data_masked[4428] = data_i[4428] & sel_one_hot_i[34];
  assign data_masked[4427] = data_i[4427] & sel_one_hot_i[34];
  assign data_masked[4426] = data_i[4426] & sel_one_hot_i[34];
  assign data_masked[4425] = data_i[4425] & sel_one_hot_i[34];
  assign data_masked[4424] = data_i[4424] & sel_one_hot_i[34];
  assign data_masked[4423] = data_i[4423] & sel_one_hot_i[34];
  assign data_masked[4422] = data_i[4422] & sel_one_hot_i[34];
  assign data_masked[4421] = data_i[4421] & sel_one_hot_i[34];
  assign data_masked[4420] = data_i[4420] & sel_one_hot_i[34];
  assign data_masked[4419] = data_i[4419] & sel_one_hot_i[34];
  assign data_masked[4418] = data_i[4418] & sel_one_hot_i[34];
  assign data_masked[4417] = data_i[4417] & sel_one_hot_i[34];
  assign data_masked[4416] = data_i[4416] & sel_one_hot_i[34];
  assign data_masked[4415] = data_i[4415] & sel_one_hot_i[34];
  assign data_masked[4414] = data_i[4414] & sel_one_hot_i[34];
  assign data_masked[4413] = data_i[4413] & sel_one_hot_i[34];
  assign data_masked[4412] = data_i[4412] & sel_one_hot_i[34];
  assign data_masked[4411] = data_i[4411] & sel_one_hot_i[34];
  assign data_masked[4410] = data_i[4410] & sel_one_hot_i[34];
  assign data_masked[4409] = data_i[4409] & sel_one_hot_i[34];
  assign data_masked[4408] = data_i[4408] & sel_one_hot_i[34];
  assign data_masked[4407] = data_i[4407] & sel_one_hot_i[34];
  assign data_masked[4406] = data_i[4406] & sel_one_hot_i[34];
  assign data_masked[4405] = data_i[4405] & sel_one_hot_i[34];
  assign data_masked[4404] = data_i[4404] & sel_one_hot_i[34];
  assign data_masked[4403] = data_i[4403] & sel_one_hot_i[34];
  assign data_masked[4402] = data_i[4402] & sel_one_hot_i[34];
  assign data_masked[4401] = data_i[4401] & sel_one_hot_i[34];
  assign data_masked[4400] = data_i[4400] & sel_one_hot_i[34];
  assign data_masked[4399] = data_i[4399] & sel_one_hot_i[34];
  assign data_masked[4398] = data_i[4398] & sel_one_hot_i[34];
  assign data_masked[4397] = data_i[4397] & sel_one_hot_i[34];
  assign data_masked[4396] = data_i[4396] & sel_one_hot_i[34];
  assign data_masked[4395] = data_i[4395] & sel_one_hot_i[34];
  assign data_masked[4394] = data_i[4394] & sel_one_hot_i[34];
  assign data_masked[4393] = data_i[4393] & sel_one_hot_i[34];
  assign data_masked[4392] = data_i[4392] & sel_one_hot_i[34];
  assign data_masked[4391] = data_i[4391] & sel_one_hot_i[34];
  assign data_masked[4390] = data_i[4390] & sel_one_hot_i[34];
  assign data_masked[4389] = data_i[4389] & sel_one_hot_i[34];
  assign data_masked[4388] = data_i[4388] & sel_one_hot_i[34];
  assign data_masked[4387] = data_i[4387] & sel_one_hot_i[34];
  assign data_masked[4386] = data_i[4386] & sel_one_hot_i[34];
  assign data_masked[4385] = data_i[4385] & sel_one_hot_i[34];
  assign data_masked[4384] = data_i[4384] & sel_one_hot_i[34];
  assign data_masked[4383] = data_i[4383] & sel_one_hot_i[34];
  assign data_masked[4382] = data_i[4382] & sel_one_hot_i[34];
  assign data_masked[4381] = data_i[4381] & sel_one_hot_i[34];
  assign data_masked[4380] = data_i[4380] & sel_one_hot_i[34];
  assign data_masked[4379] = data_i[4379] & sel_one_hot_i[34];
  assign data_masked[4378] = data_i[4378] & sel_one_hot_i[34];
  assign data_masked[4377] = data_i[4377] & sel_one_hot_i[34];
  assign data_masked[4376] = data_i[4376] & sel_one_hot_i[34];
  assign data_masked[4375] = data_i[4375] & sel_one_hot_i[34];
  assign data_masked[4374] = data_i[4374] & sel_one_hot_i[34];
  assign data_masked[4373] = data_i[4373] & sel_one_hot_i[34];
  assign data_masked[4372] = data_i[4372] & sel_one_hot_i[34];
  assign data_masked[4371] = data_i[4371] & sel_one_hot_i[34];
  assign data_masked[4370] = data_i[4370] & sel_one_hot_i[34];
  assign data_masked[4369] = data_i[4369] & sel_one_hot_i[34];
  assign data_masked[4368] = data_i[4368] & sel_one_hot_i[34];
  assign data_masked[4367] = data_i[4367] & sel_one_hot_i[34];
  assign data_masked[4366] = data_i[4366] & sel_one_hot_i[34];
  assign data_masked[4365] = data_i[4365] & sel_one_hot_i[34];
  assign data_masked[4364] = data_i[4364] & sel_one_hot_i[34];
  assign data_masked[4363] = data_i[4363] & sel_one_hot_i[34];
  assign data_masked[4362] = data_i[4362] & sel_one_hot_i[34];
  assign data_masked[4361] = data_i[4361] & sel_one_hot_i[34];
  assign data_masked[4360] = data_i[4360] & sel_one_hot_i[34];
  assign data_masked[4359] = data_i[4359] & sel_one_hot_i[34];
  assign data_masked[4358] = data_i[4358] & sel_one_hot_i[34];
  assign data_masked[4357] = data_i[4357] & sel_one_hot_i[34];
  assign data_masked[4356] = data_i[4356] & sel_one_hot_i[34];
  assign data_masked[4355] = data_i[4355] & sel_one_hot_i[34];
  assign data_masked[4354] = data_i[4354] & sel_one_hot_i[34];
  assign data_masked[4353] = data_i[4353] & sel_one_hot_i[34];
  assign data_masked[4352] = data_i[4352] & sel_one_hot_i[34];
  assign data_masked[4607] = data_i[4607] & sel_one_hot_i[35];
  assign data_masked[4606] = data_i[4606] & sel_one_hot_i[35];
  assign data_masked[4605] = data_i[4605] & sel_one_hot_i[35];
  assign data_masked[4604] = data_i[4604] & sel_one_hot_i[35];
  assign data_masked[4603] = data_i[4603] & sel_one_hot_i[35];
  assign data_masked[4602] = data_i[4602] & sel_one_hot_i[35];
  assign data_masked[4601] = data_i[4601] & sel_one_hot_i[35];
  assign data_masked[4600] = data_i[4600] & sel_one_hot_i[35];
  assign data_masked[4599] = data_i[4599] & sel_one_hot_i[35];
  assign data_masked[4598] = data_i[4598] & sel_one_hot_i[35];
  assign data_masked[4597] = data_i[4597] & sel_one_hot_i[35];
  assign data_masked[4596] = data_i[4596] & sel_one_hot_i[35];
  assign data_masked[4595] = data_i[4595] & sel_one_hot_i[35];
  assign data_masked[4594] = data_i[4594] & sel_one_hot_i[35];
  assign data_masked[4593] = data_i[4593] & sel_one_hot_i[35];
  assign data_masked[4592] = data_i[4592] & sel_one_hot_i[35];
  assign data_masked[4591] = data_i[4591] & sel_one_hot_i[35];
  assign data_masked[4590] = data_i[4590] & sel_one_hot_i[35];
  assign data_masked[4589] = data_i[4589] & sel_one_hot_i[35];
  assign data_masked[4588] = data_i[4588] & sel_one_hot_i[35];
  assign data_masked[4587] = data_i[4587] & sel_one_hot_i[35];
  assign data_masked[4586] = data_i[4586] & sel_one_hot_i[35];
  assign data_masked[4585] = data_i[4585] & sel_one_hot_i[35];
  assign data_masked[4584] = data_i[4584] & sel_one_hot_i[35];
  assign data_masked[4583] = data_i[4583] & sel_one_hot_i[35];
  assign data_masked[4582] = data_i[4582] & sel_one_hot_i[35];
  assign data_masked[4581] = data_i[4581] & sel_one_hot_i[35];
  assign data_masked[4580] = data_i[4580] & sel_one_hot_i[35];
  assign data_masked[4579] = data_i[4579] & sel_one_hot_i[35];
  assign data_masked[4578] = data_i[4578] & sel_one_hot_i[35];
  assign data_masked[4577] = data_i[4577] & sel_one_hot_i[35];
  assign data_masked[4576] = data_i[4576] & sel_one_hot_i[35];
  assign data_masked[4575] = data_i[4575] & sel_one_hot_i[35];
  assign data_masked[4574] = data_i[4574] & sel_one_hot_i[35];
  assign data_masked[4573] = data_i[4573] & sel_one_hot_i[35];
  assign data_masked[4572] = data_i[4572] & sel_one_hot_i[35];
  assign data_masked[4571] = data_i[4571] & sel_one_hot_i[35];
  assign data_masked[4570] = data_i[4570] & sel_one_hot_i[35];
  assign data_masked[4569] = data_i[4569] & sel_one_hot_i[35];
  assign data_masked[4568] = data_i[4568] & sel_one_hot_i[35];
  assign data_masked[4567] = data_i[4567] & sel_one_hot_i[35];
  assign data_masked[4566] = data_i[4566] & sel_one_hot_i[35];
  assign data_masked[4565] = data_i[4565] & sel_one_hot_i[35];
  assign data_masked[4564] = data_i[4564] & sel_one_hot_i[35];
  assign data_masked[4563] = data_i[4563] & sel_one_hot_i[35];
  assign data_masked[4562] = data_i[4562] & sel_one_hot_i[35];
  assign data_masked[4561] = data_i[4561] & sel_one_hot_i[35];
  assign data_masked[4560] = data_i[4560] & sel_one_hot_i[35];
  assign data_masked[4559] = data_i[4559] & sel_one_hot_i[35];
  assign data_masked[4558] = data_i[4558] & sel_one_hot_i[35];
  assign data_masked[4557] = data_i[4557] & sel_one_hot_i[35];
  assign data_masked[4556] = data_i[4556] & sel_one_hot_i[35];
  assign data_masked[4555] = data_i[4555] & sel_one_hot_i[35];
  assign data_masked[4554] = data_i[4554] & sel_one_hot_i[35];
  assign data_masked[4553] = data_i[4553] & sel_one_hot_i[35];
  assign data_masked[4552] = data_i[4552] & sel_one_hot_i[35];
  assign data_masked[4551] = data_i[4551] & sel_one_hot_i[35];
  assign data_masked[4550] = data_i[4550] & sel_one_hot_i[35];
  assign data_masked[4549] = data_i[4549] & sel_one_hot_i[35];
  assign data_masked[4548] = data_i[4548] & sel_one_hot_i[35];
  assign data_masked[4547] = data_i[4547] & sel_one_hot_i[35];
  assign data_masked[4546] = data_i[4546] & sel_one_hot_i[35];
  assign data_masked[4545] = data_i[4545] & sel_one_hot_i[35];
  assign data_masked[4544] = data_i[4544] & sel_one_hot_i[35];
  assign data_masked[4543] = data_i[4543] & sel_one_hot_i[35];
  assign data_masked[4542] = data_i[4542] & sel_one_hot_i[35];
  assign data_masked[4541] = data_i[4541] & sel_one_hot_i[35];
  assign data_masked[4540] = data_i[4540] & sel_one_hot_i[35];
  assign data_masked[4539] = data_i[4539] & sel_one_hot_i[35];
  assign data_masked[4538] = data_i[4538] & sel_one_hot_i[35];
  assign data_masked[4537] = data_i[4537] & sel_one_hot_i[35];
  assign data_masked[4536] = data_i[4536] & sel_one_hot_i[35];
  assign data_masked[4535] = data_i[4535] & sel_one_hot_i[35];
  assign data_masked[4534] = data_i[4534] & sel_one_hot_i[35];
  assign data_masked[4533] = data_i[4533] & sel_one_hot_i[35];
  assign data_masked[4532] = data_i[4532] & sel_one_hot_i[35];
  assign data_masked[4531] = data_i[4531] & sel_one_hot_i[35];
  assign data_masked[4530] = data_i[4530] & sel_one_hot_i[35];
  assign data_masked[4529] = data_i[4529] & sel_one_hot_i[35];
  assign data_masked[4528] = data_i[4528] & sel_one_hot_i[35];
  assign data_masked[4527] = data_i[4527] & sel_one_hot_i[35];
  assign data_masked[4526] = data_i[4526] & sel_one_hot_i[35];
  assign data_masked[4525] = data_i[4525] & sel_one_hot_i[35];
  assign data_masked[4524] = data_i[4524] & sel_one_hot_i[35];
  assign data_masked[4523] = data_i[4523] & sel_one_hot_i[35];
  assign data_masked[4522] = data_i[4522] & sel_one_hot_i[35];
  assign data_masked[4521] = data_i[4521] & sel_one_hot_i[35];
  assign data_masked[4520] = data_i[4520] & sel_one_hot_i[35];
  assign data_masked[4519] = data_i[4519] & sel_one_hot_i[35];
  assign data_masked[4518] = data_i[4518] & sel_one_hot_i[35];
  assign data_masked[4517] = data_i[4517] & sel_one_hot_i[35];
  assign data_masked[4516] = data_i[4516] & sel_one_hot_i[35];
  assign data_masked[4515] = data_i[4515] & sel_one_hot_i[35];
  assign data_masked[4514] = data_i[4514] & sel_one_hot_i[35];
  assign data_masked[4513] = data_i[4513] & sel_one_hot_i[35];
  assign data_masked[4512] = data_i[4512] & sel_one_hot_i[35];
  assign data_masked[4511] = data_i[4511] & sel_one_hot_i[35];
  assign data_masked[4510] = data_i[4510] & sel_one_hot_i[35];
  assign data_masked[4509] = data_i[4509] & sel_one_hot_i[35];
  assign data_masked[4508] = data_i[4508] & sel_one_hot_i[35];
  assign data_masked[4507] = data_i[4507] & sel_one_hot_i[35];
  assign data_masked[4506] = data_i[4506] & sel_one_hot_i[35];
  assign data_masked[4505] = data_i[4505] & sel_one_hot_i[35];
  assign data_masked[4504] = data_i[4504] & sel_one_hot_i[35];
  assign data_masked[4503] = data_i[4503] & sel_one_hot_i[35];
  assign data_masked[4502] = data_i[4502] & sel_one_hot_i[35];
  assign data_masked[4501] = data_i[4501] & sel_one_hot_i[35];
  assign data_masked[4500] = data_i[4500] & sel_one_hot_i[35];
  assign data_masked[4499] = data_i[4499] & sel_one_hot_i[35];
  assign data_masked[4498] = data_i[4498] & sel_one_hot_i[35];
  assign data_masked[4497] = data_i[4497] & sel_one_hot_i[35];
  assign data_masked[4496] = data_i[4496] & sel_one_hot_i[35];
  assign data_masked[4495] = data_i[4495] & sel_one_hot_i[35];
  assign data_masked[4494] = data_i[4494] & sel_one_hot_i[35];
  assign data_masked[4493] = data_i[4493] & sel_one_hot_i[35];
  assign data_masked[4492] = data_i[4492] & sel_one_hot_i[35];
  assign data_masked[4491] = data_i[4491] & sel_one_hot_i[35];
  assign data_masked[4490] = data_i[4490] & sel_one_hot_i[35];
  assign data_masked[4489] = data_i[4489] & sel_one_hot_i[35];
  assign data_masked[4488] = data_i[4488] & sel_one_hot_i[35];
  assign data_masked[4487] = data_i[4487] & sel_one_hot_i[35];
  assign data_masked[4486] = data_i[4486] & sel_one_hot_i[35];
  assign data_masked[4485] = data_i[4485] & sel_one_hot_i[35];
  assign data_masked[4484] = data_i[4484] & sel_one_hot_i[35];
  assign data_masked[4483] = data_i[4483] & sel_one_hot_i[35];
  assign data_masked[4482] = data_i[4482] & sel_one_hot_i[35];
  assign data_masked[4481] = data_i[4481] & sel_one_hot_i[35];
  assign data_masked[4480] = data_i[4480] & sel_one_hot_i[35];
  assign data_masked[4735] = data_i[4735] & sel_one_hot_i[36];
  assign data_masked[4734] = data_i[4734] & sel_one_hot_i[36];
  assign data_masked[4733] = data_i[4733] & sel_one_hot_i[36];
  assign data_masked[4732] = data_i[4732] & sel_one_hot_i[36];
  assign data_masked[4731] = data_i[4731] & sel_one_hot_i[36];
  assign data_masked[4730] = data_i[4730] & sel_one_hot_i[36];
  assign data_masked[4729] = data_i[4729] & sel_one_hot_i[36];
  assign data_masked[4728] = data_i[4728] & sel_one_hot_i[36];
  assign data_masked[4727] = data_i[4727] & sel_one_hot_i[36];
  assign data_masked[4726] = data_i[4726] & sel_one_hot_i[36];
  assign data_masked[4725] = data_i[4725] & sel_one_hot_i[36];
  assign data_masked[4724] = data_i[4724] & sel_one_hot_i[36];
  assign data_masked[4723] = data_i[4723] & sel_one_hot_i[36];
  assign data_masked[4722] = data_i[4722] & sel_one_hot_i[36];
  assign data_masked[4721] = data_i[4721] & sel_one_hot_i[36];
  assign data_masked[4720] = data_i[4720] & sel_one_hot_i[36];
  assign data_masked[4719] = data_i[4719] & sel_one_hot_i[36];
  assign data_masked[4718] = data_i[4718] & sel_one_hot_i[36];
  assign data_masked[4717] = data_i[4717] & sel_one_hot_i[36];
  assign data_masked[4716] = data_i[4716] & sel_one_hot_i[36];
  assign data_masked[4715] = data_i[4715] & sel_one_hot_i[36];
  assign data_masked[4714] = data_i[4714] & sel_one_hot_i[36];
  assign data_masked[4713] = data_i[4713] & sel_one_hot_i[36];
  assign data_masked[4712] = data_i[4712] & sel_one_hot_i[36];
  assign data_masked[4711] = data_i[4711] & sel_one_hot_i[36];
  assign data_masked[4710] = data_i[4710] & sel_one_hot_i[36];
  assign data_masked[4709] = data_i[4709] & sel_one_hot_i[36];
  assign data_masked[4708] = data_i[4708] & sel_one_hot_i[36];
  assign data_masked[4707] = data_i[4707] & sel_one_hot_i[36];
  assign data_masked[4706] = data_i[4706] & sel_one_hot_i[36];
  assign data_masked[4705] = data_i[4705] & sel_one_hot_i[36];
  assign data_masked[4704] = data_i[4704] & sel_one_hot_i[36];
  assign data_masked[4703] = data_i[4703] & sel_one_hot_i[36];
  assign data_masked[4702] = data_i[4702] & sel_one_hot_i[36];
  assign data_masked[4701] = data_i[4701] & sel_one_hot_i[36];
  assign data_masked[4700] = data_i[4700] & sel_one_hot_i[36];
  assign data_masked[4699] = data_i[4699] & sel_one_hot_i[36];
  assign data_masked[4698] = data_i[4698] & sel_one_hot_i[36];
  assign data_masked[4697] = data_i[4697] & sel_one_hot_i[36];
  assign data_masked[4696] = data_i[4696] & sel_one_hot_i[36];
  assign data_masked[4695] = data_i[4695] & sel_one_hot_i[36];
  assign data_masked[4694] = data_i[4694] & sel_one_hot_i[36];
  assign data_masked[4693] = data_i[4693] & sel_one_hot_i[36];
  assign data_masked[4692] = data_i[4692] & sel_one_hot_i[36];
  assign data_masked[4691] = data_i[4691] & sel_one_hot_i[36];
  assign data_masked[4690] = data_i[4690] & sel_one_hot_i[36];
  assign data_masked[4689] = data_i[4689] & sel_one_hot_i[36];
  assign data_masked[4688] = data_i[4688] & sel_one_hot_i[36];
  assign data_masked[4687] = data_i[4687] & sel_one_hot_i[36];
  assign data_masked[4686] = data_i[4686] & sel_one_hot_i[36];
  assign data_masked[4685] = data_i[4685] & sel_one_hot_i[36];
  assign data_masked[4684] = data_i[4684] & sel_one_hot_i[36];
  assign data_masked[4683] = data_i[4683] & sel_one_hot_i[36];
  assign data_masked[4682] = data_i[4682] & sel_one_hot_i[36];
  assign data_masked[4681] = data_i[4681] & sel_one_hot_i[36];
  assign data_masked[4680] = data_i[4680] & sel_one_hot_i[36];
  assign data_masked[4679] = data_i[4679] & sel_one_hot_i[36];
  assign data_masked[4678] = data_i[4678] & sel_one_hot_i[36];
  assign data_masked[4677] = data_i[4677] & sel_one_hot_i[36];
  assign data_masked[4676] = data_i[4676] & sel_one_hot_i[36];
  assign data_masked[4675] = data_i[4675] & sel_one_hot_i[36];
  assign data_masked[4674] = data_i[4674] & sel_one_hot_i[36];
  assign data_masked[4673] = data_i[4673] & sel_one_hot_i[36];
  assign data_masked[4672] = data_i[4672] & sel_one_hot_i[36];
  assign data_masked[4671] = data_i[4671] & sel_one_hot_i[36];
  assign data_masked[4670] = data_i[4670] & sel_one_hot_i[36];
  assign data_masked[4669] = data_i[4669] & sel_one_hot_i[36];
  assign data_masked[4668] = data_i[4668] & sel_one_hot_i[36];
  assign data_masked[4667] = data_i[4667] & sel_one_hot_i[36];
  assign data_masked[4666] = data_i[4666] & sel_one_hot_i[36];
  assign data_masked[4665] = data_i[4665] & sel_one_hot_i[36];
  assign data_masked[4664] = data_i[4664] & sel_one_hot_i[36];
  assign data_masked[4663] = data_i[4663] & sel_one_hot_i[36];
  assign data_masked[4662] = data_i[4662] & sel_one_hot_i[36];
  assign data_masked[4661] = data_i[4661] & sel_one_hot_i[36];
  assign data_masked[4660] = data_i[4660] & sel_one_hot_i[36];
  assign data_masked[4659] = data_i[4659] & sel_one_hot_i[36];
  assign data_masked[4658] = data_i[4658] & sel_one_hot_i[36];
  assign data_masked[4657] = data_i[4657] & sel_one_hot_i[36];
  assign data_masked[4656] = data_i[4656] & sel_one_hot_i[36];
  assign data_masked[4655] = data_i[4655] & sel_one_hot_i[36];
  assign data_masked[4654] = data_i[4654] & sel_one_hot_i[36];
  assign data_masked[4653] = data_i[4653] & sel_one_hot_i[36];
  assign data_masked[4652] = data_i[4652] & sel_one_hot_i[36];
  assign data_masked[4651] = data_i[4651] & sel_one_hot_i[36];
  assign data_masked[4650] = data_i[4650] & sel_one_hot_i[36];
  assign data_masked[4649] = data_i[4649] & sel_one_hot_i[36];
  assign data_masked[4648] = data_i[4648] & sel_one_hot_i[36];
  assign data_masked[4647] = data_i[4647] & sel_one_hot_i[36];
  assign data_masked[4646] = data_i[4646] & sel_one_hot_i[36];
  assign data_masked[4645] = data_i[4645] & sel_one_hot_i[36];
  assign data_masked[4644] = data_i[4644] & sel_one_hot_i[36];
  assign data_masked[4643] = data_i[4643] & sel_one_hot_i[36];
  assign data_masked[4642] = data_i[4642] & sel_one_hot_i[36];
  assign data_masked[4641] = data_i[4641] & sel_one_hot_i[36];
  assign data_masked[4640] = data_i[4640] & sel_one_hot_i[36];
  assign data_masked[4639] = data_i[4639] & sel_one_hot_i[36];
  assign data_masked[4638] = data_i[4638] & sel_one_hot_i[36];
  assign data_masked[4637] = data_i[4637] & sel_one_hot_i[36];
  assign data_masked[4636] = data_i[4636] & sel_one_hot_i[36];
  assign data_masked[4635] = data_i[4635] & sel_one_hot_i[36];
  assign data_masked[4634] = data_i[4634] & sel_one_hot_i[36];
  assign data_masked[4633] = data_i[4633] & sel_one_hot_i[36];
  assign data_masked[4632] = data_i[4632] & sel_one_hot_i[36];
  assign data_masked[4631] = data_i[4631] & sel_one_hot_i[36];
  assign data_masked[4630] = data_i[4630] & sel_one_hot_i[36];
  assign data_masked[4629] = data_i[4629] & sel_one_hot_i[36];
  assign data_masked[4628] = data_i[4628] & sel_one_hot_i[36];
  assign data_masked[4627] = data_i[4627] & sel_one_hot_i[36];
  assign data_masked[4626] = data_i[4626] & sel_one_hot_i[36];
  assign data_masked[4625] = data_i[4625] & sel_one_hot_i[36];
  assign data_masked[4624] = data_i[4624] & sel_one_hot_i[36];
  assign data_masked[4623] = data_i[4623] & sel_one_hot_i[36];
  assign data_masked[4622] = data_i[4622] & sel_one_hot_i[36];
  assign data_masked[4621] = data_i[4621] & sel_one_hot_i[36];
  assign data_masked[4620] = data_i[4620] & sel_one_hot_i[36];
  assign data_masked[4619] = data_i[4619] & sel_one_hot_i[36];
  assign data_masked[4618] = data_i[4618] & sel_one_hot_i[36];
  assign data_masked[4617] = data_i[4617] & sel_one_hot_i[36];
  assign data_masked[4616] = data_i[4616] & sel_one_hot_i[36];
  assign data_masked[4615] = data_i[4615] & sel_one_hot_i[36];
  assign data_masked[4614] = data_i[4614] & sel_one_hot_i[36];
  assign data_masked[4613] = data_i[4613] & sel_one_hot_i[36];
  assign data_masked[4612] = data_i[4612] & sel_one_hot_i[36];
  assign data_masked[4611] = data_i[4611] & sel_one_hot_i[36];
  assign data_masked[4610] = data_i[4610] & sel_one_hot_i[36];
  assign data_masked[4609] = data_i[4609] & sel_one_hot_i[36];
  assign data_masked[4608] = data_i[4608] & sel_one_hot_i[36];
  assign data_masked[4863] = data_i[4863] & sel_one_hot_i[37];
  assign data_masked[4862] = data_i[4862] & sel_one_hot_i[37];
  assign data_masked[4861] = data_i[4861] & sel_one_hot_i[37];
  assign data_masked[4860] = data_i[4860] & sel_one_hot_i[37];
  assign data_masked[4859] = data_i[4859] & sel_one_hot_i[37];
  assign data_masked[4858] = data_i[4858] & sel_one_hot_i[37];
  assign data_masked[4857] = data_i[4857] & sel_one_hot_i[37];
  assign data_masked[4856] = data_i[4856] & sel_one_hot_i[37];
  assign data_masked[4855] = data_i[4855] & sel_one_hot_i[37];
  assign data_masked[4854] = data_i[4854] & sel_one_hot_i[37];
  assign data_masked[4853] = data_i[4853] & sel_one_hot_i[37];
  assign data_masked[4852] = data_i[4852] & sel_one_hot_i[37];
  assign data_masked[4851] = data_i[4851] & sel_one_hot_i[37];
  assign data_masked[4850] = data_i[4850] & sel_one_hot_i[37];
  assign data_masked[4849] = data_i[4849] & sel_one_hot_i[37];
  assign data_masked[4848] = data_i[4848] & sel_one_hot_i[37];
  assign data_masked[4847] = data_i[4847] & sel_one_hot_i[37];
  assign data_masked[4846] = data_i[4846] & sel_one_hot_i[37];
  assign data_masked[4845] = data_i[4845] & sel_one_hot_i[37];
  assign data_masked[4844] = data_i[4844] & sel_one_hot_i[37];
  assign data_masked[4843] = data_i[4843] & sel_one_hot_i[37];
  assign data_masked[4842] = data_i[4842] & sel_one_hot_i[37];
  assign data_masked[4841] = data_i[4841] & sel_one_hot_i[37];
  assign data_masked[4840] = data_i[4840] & sel_one_hot_i[37];
  assign data_masked[4839] = data_i[4839] & sel_one_hot_i[37];
  assign data_masked[4838] = data_i[4838] & sel_one_hot_i[37];
  assign data_masked[4837] = data_i[4837] & sel_one_hot_i[37];
  assign data_masked[4836] = data_i[4836] & sel_one_hot_i[37];
  assign data_masked[4835] = data_i[4835] & sel_one_hot_i[37];
  assign data_masked[4834] = data_i[4834] & sel_one_hot_i[37];
  assign data_masked[4833] = data_i[4833] & sel_one_hot_i[37];
  assign data_masked[4832] = data_i[4832] & sel_one_hot_i[37];
  assign data_masked[4831] = data_i[4831] & sel_one_hot_i[37];
  assign data_masked[4830] = data_i[4830] & sel_one_hot_i[37];
  assign data_masked[4829] = data_i[4829] & sel_one_hot_i[37];
  assign data_masked[4828] = data_i[4828] & sel_one_hot_i[37];
  assign data_masked[4827] = data_i[4827] & sel_one_hot_i[37];
  assign data_masked[4826] = data_i[4826] & sel_one_hot_i[37];
  assign data_masked[4825] = data_i[4825] & sel_one_hot_i[37];
  assign data_masked[4824] = data_i[4824] & sel_one_hot_i[37];
  assign data_masked[4823] = data_i[4823] & sel_one_hot_i[37];
  assign data_masked[4822] = data_i[4822] & sel_one_hot_i[37];
  assign data_masked[4821] = data_i[4821] & sel_one_hot_i[37];
  assign data_masked[4820] = data_i[4820] & sel_one_hot_i[37];
  assign data_masked[4819] = data_i[4819] & sel_one_hot_i[37];
  assign data_masked[4818] = data_i[4818] & sel_one_hot_i[37];
  assign data_masked[4817] = data_i[4817] & sel_one_hot_i[37];
  assign data_masked[4816] = data_i[4816] & sel_one_hot_i[37];
  assign data_masked[4815] = data_i[4815] & sel_one_hot_i[37];
  assign data_masked[4814] = data_i[4814] & sel_one_hot_i[37];
  assign data_masked[4813] = data_i[4813] & sel_one_hot_i[37];
  assign data_masked[4812] = data_i[4812] & sel_one_hot_i[37];
  assign data_masked[4811] = data_i[4811] & sel_one_hot_i[37];
  assign data_masked[4810] = data_i[4810] & sel_one_hot_i[37];
  assign data_masked[4809] = data_i[4809] & sel_one_hot_i[37];
  assign data_masked[4808] = data_i[4808] & sel_one_hot_i[37];
  assign data_masked[4807] = data_i[4807] & sel_one_hot_i[37];
  assign data_masked[4806] = data_i[4806] & sel_one_hot_i[37];
  assign data_masked[4805] = data_i[4805] & sel_one_hot_i[37];
  assign data_masked[4804] = data_i[4804] & sel_one_hot_i[37];
  assign data_masked[4803] = data_i[4803] & sel_one_hot_i[37];
  assign data_masked[4802] = data_i[4802] & sel_one_hot_i[37];
  assign data_masked[4801] = data_i[4801] & sel_one_hot_i[37];
  assign data_masked[4800] = data_i[4800] & sel_one_hot_i[37];
  assign data_masked[4799] = data_i[4799] & sel_one_hot_i[37];
  assign data_masked[4798] = data_i[4798] & sel_one_hot_i[37];
  assign data_masked[4797] = data_i[4797] & sel_one_hot_i[37];
  assign data_masked[4796] = data_i[4796] & sel_one_hot_i[37];
  assign data_masked[4795] = data_i[4795] & sel_one_hot_i[37];
  assign data_masked[4794] = data_i[4794] & sel_one_hot_i[37];
  assign data_masked[4793] = data_i[4793] & sel_one_hot_i[37];
  assign data_masked[4792] = data_i[4792] & sel_one_hot_i[37];
  assign data_masked[4791] = data_i[4791] & sel_one_hot_i[37];
  assign data_masked[4790] = data_i[4790] & sel_one_hot_i[37];
  assign data_masked[4789] = data_i[4789] & sel_one_hot_i[37];
  assign data_masked[4788] = data_i[4788] & sel_one_hot_i[37];
  assign data_masked[4787] = data_i[4787] & sel_one_hot_i[37];
  assign data_masked[4786] = data_i[4786] & sel_one_hot_i[37];
  assign data_masked[4785] = data_i[4785] & sel_one_hot_i[37];
  assign data_masked[4784] = data_i[4784] & sel_one_hot_i[37];
  assign data_masked[4783] = data_i[4783] & sel_one_hot_i[37];
  assign data_masked[4782] = data_i[4782] & sel_one_hot_i[37];
  assign data_masked[4781] = data_i[4781] & sel_one_hot_i[37];
  assign data_masked[4780] = data_i[4780] & sel_one_hot_i[37];
  assign data_masked[4779] = data_i[4779] & sel_one_hot_i[37];
  assign data_masked[4778] = data_i[4778] & sel_one_hot_i[37];
  assign data_masked[4777] = data_i[4777] & sel_one_hot_i[37];
  assign data_masked[4776] = data_i[4776] & sel_one_hot_i[37];
  assign data_masked[4775] = data_i[4775] & sel_one_hot_i[37];
  assign data_masked[4774] = data_i[4774] & sel_one_hot_i[37];
  assign data_masked[4773] = data_i[4773] & sel_one_hot_i[37];
  assign data_masked[4772] = data_i[4772] & sel_one_hot_i[37];
  assign data_masked[4771] = data_i[4771] & sel_one_hot_i[37];
  assign data_masked[4770] = data_i[4770] & sel_one_hot_i[37];
  assign data_masked[4769] = data_i[4769] & sel_one_hot_i[37];
  assign data_masked[4768] = data_i[4768] & sel_one_hot_i[37];
  assign data_masked[4767] = data_i[4767] & sel_one_hot_i[37];
  assign data_masked[4766] = data_i[4766] & sel_one_hot_i[37];
  assign data_masked[4765] = data_i[4765] & sel_one_hot_i[37];
  assign data_masked[4764] = data_i[4764] & sel_one_hot_i[37];
  assign data_masked[4763] = data_i[4763] & sel_one_hot_i[37];
  assign data_masked[4762] = data_i[4762] & sel_one_hot_i[37];
  assign data_masked[4761] = data_i[4761] & sel_one_hot_i[37];
  assign data_masked[4760] = data_i[4760] & sel_one_hot_i[37];
  assign data_masked[4759] = data_i[4759] & sel_one_hot_i[37];
  assign data_masked[4758] = data_i[4758] & sel_one_hot_i[37];
  assign data_masked[4757] = data_i[4757] & sel_one_hot_i[37];
  assign data_masked[4756] = data_i[4756] & sel_one_hot_i[37];
  assign data_masked[4755] = data_i[4755] & sel_one_hot_i[37];
  assign data_masked[4754] = data_i[4754] & sel_one_hot_i[37];
  assign data_masked[4753] = data_i[4753] & sel_one_hot_i[37];
  assign data_masked[4752] = data_i[4752] & sel_one_hot_i[37];
  assign data_masked[4751] = data_i[4751] & sel_one_hot_i[37];
  assign data_masked[4750] = data_i[4750] & sel_one_hot_i[37];
  assign data_masked[4749] = data_i[4749] & sel_one_hot_i[37];
  assign data_masked[4748] = data_i[4748] & sel_one_hot_i[37];
  assign data_masked[4747] = data_i[4747] & sel_one_hot_i[37];
  assign data_masked[4746] = data_i[4746] & sel_one_hot_i[37];
  assign data_masked[4745] = data_i[4745] & sel_one_hot_i[37];
  assign data_masked[4744] = data_i[4744] & sel_one_hot_i[37];
  assign data_masked[4743] = data_i[4743] & sel_one_hot_i[37];
  assign data_masked[4742] = data_i[4742] & sel_one_hot_i[37];
  assign data_masked[4741] = data_i[4741] & sel_one_hot_i[37];
  assign data_masked[4740] = data_i[4740] & sel_one_hot_i[37];
  assign data_masked[4739] = data_i[4739] & sel_one_hot_i[37];
  assign data_masked[4738] = data_i[4738] & sel_one_hot_i[37];
  assign data_masked[4737] = data_i[4737] & sel_one_hot_i[37];
  assign data_masked[4736] = data_i[4736] & sel_one_hot_i[37];
  assign data_masked[4991] = data_i[4991] & sel_one_hot_i[38];
  assign data_masked[4990] = data_i[4990] & sel_one_hot_i[38];
  assign data_masked[4989] = data_i[4989] & sel_one_hot_i[38];
  assign data_masked[4988] = data_i[4988] & sel_one_hot_i[38];
  assign data_masked[4987] = data_i[4987] & sel_one_hot_i[38];
  assign data_masked[4986] = data_i[4986] & sel_one_hot_i[38];
  assign data_masked[4985] = data_i[4985] & sel_one_hot_i[38];
  assign data_masked[4984] = data_i[4984] & sel_one_hot_i[38];
  assign data_masked[4983] = data_i[4983] & sel_one_hot_i[38];
  assign data_masked[4982] = data_i[4982] & sel_one_hot_i[38];
  assign data_masked[4981] = data_i[4981] & sel_one_hot_i[38];
  assign data_masked[4980] = data_i[4980] & sel_one_hot_i[38];
  assign data_masked[4979] = data_i[4979] & sel_one_hot_i[38];
  assign data_masked[4978] = data_i[4978] & sel_one_hot_i[38];
  assign data_masked[4977] = data_i[4977] & sel_one_hot_i[38];
  assign data_masked[4976] = data_i[4976] & sel_one_hot_i[38];
  assign data_masked[4975] = data_i[4975] & sel_one_hot_i[38];
  assign data_masked[4974] = data_i[4974] & sel_one_hot_i[38];
  assign data_masked[4973] = data_i[4973] & sel_one_hot_i[38];
  assign data_masked[4972] = data_i[4972] & sel_one_hot_i[38];
  assign data_masked[4971] = data_i[4971] & sel_one_hot_i[38];
  assign data_masked[4970] = data_i[4970] & sel_one_hot_i[38];
  assign data_masked[4969] = data_i[4969] & sel_one_hot_i[38];
  assign data_masked[4968] = data_i[4968] & sel_one_hot_i[38];
  assign data_masked[4967] = data_i[4967] & sel_one_hot_i[38];
  assign data_masked[4966] = data_i[4966] & sel_one_hot_i[38];
  assign data_masked[4965] = data_i[4965] & sel_one_hot_i[38];
  assign data_masked[4964] = data_i[4964] & sel_one_hot_i[38];
  assign data_masked[4963] = data_i[4963] & sel_one_hot_i[38];
  assign data_masked[4962] = data_i[4962] & sel_one_hot_i[38];
  assign data_masked[4961] = data_i[4961] & sel_one_hot_i[38];
  assign data_masked[4960] = data_i[4960] & sel_one_hot_i[38];
  assign data_masked[4959] = data_i[4959] & sel_one_hot_i[38];
  assign data_masked[4958] = data_i[4958] & sel_one_hot_i[38];
  assign data_masked[4957] = data_i[4957] & sel_one_hot_i[38];
  assign data_masked[4956] = data_i[4956] & sel_one_hot_i[38];
  assign data_masked[4955] = data_i[4955] & sel_one_hot_i[38];
  assign data_masked[4954] = data_i[4954] & sel_one_hot_i[38];
  assign data_masked[4953] = data_i[4953] & sel_one_hot_i[38];
  assign data_masked[4952] = data_i[4952] & sel_one_hot_i[38];
  assign data_masked[4951] = data_i[4951] & sel_one_hot_i[38];
  assign data_masked[4950] = data_i[4950] & sel_one_hot_i[38];
  assign data_masked[4949] = data_i[4949] & sel_one_hot_i[38];
  assign data_masked[4948] = data_i[4948] & sel_one_hot_i[38];
  assign data_masked[4947] = data_i[4947] & sel_one_hot_i[38];
  assign data_masked[4946] = data_i[4946] & sel_one_hot_i[38];
  assign data_masked[4945] = data_i[4945] & sel_one_hot_i[38];
  assign data_masked[4944] = data_i[4944] & sel_one_hot_i[38];
  assign data_masked[4943] = data_i[4943] & sel_one_hot_i[38];
  assign data_masked[4942] = data_i[4942] & sel_one_hot_i[38];
  assign data_masked[4941] = data_i[4941] & sel_one_hot_i[38];
  assign data_masked[4940] = data_i[4940] & sel_one_hot_i[38];
  assign data_masked[4939] = data_i[4939] & sel_one_hot_i[38];
  assign data_masked[4938] = data_i[4938] & sel_one_hot_i[38];
  assign data_masked[4937] = data_i[4937] & sel_one_hot_i[38];
  assign data_masked[4936] = data_i[4936] & sel_one_hot_i[38];
  assign data_masked[4935] = data_i[4935] & sel_one_hot_i[38];
  assign data_masked[4934] = data_i[4934] & sel_one_hot_i[38];
  assign data_masked[4933] = data_i[4933] & sel_one_hot_i[38];
  assign data_masked[4932] = data_i[4932] & sel_one_hot_i[38];
  assign data_masked[4931] = data_i[4931] & sel_one_hot_i[38];
  assign data_masked[4930] = data_i[4930] & sel_one_hot_i[38];
  assign data_masked[4929] = data_i[4929] & sel_one_hot_i[38];
  assign data_masked[4928] = data_i[4928] & sel_one_hot_i[38];
  assign data_masked[4927] = data_i[4927] & sel_one_hot_i[38];
  assign data_masked[4926] = data_i[4926] & sel_one_hot_i[38];
  assign data_masked[4925] = data_i[4925] & sel_one_hot_i[38];
  assign data_masked[4924] = data_i[4924] & sel_one_hot_i[38];
  assign data_masked[4923] = data_i[4923] & sel_one_hot_i[38];
  assign data_masked[4922] = data_i[4922] & sel_one_hot_i[38];
  assign data_masked[4921] = data_i[4921] & sel_one_hot_i[38];
  assign data_masked[4920] = data_i[4920] & sel_one_hot_i[38];
  assign data_masked[4919] = data_i[4919] & sel_one_hot_i[38];
  assign data_masked[4918] = data_i[4918] & sel_one_hot_i[38];
  assign data_masked[4917] = data_i[4917] & sel_one_hot_i[38];
  assign data_masked[4916] = data_i[4916] & sel_one_hot_i[38];
  assign data_masked[4915] = data_i[4915] & sel_one_hot_i[38];
  assign data_masked[4914] = data_i[4914] & sel_one_hot_i[38];
  assign data_masked[4913] = data_i[4913] & sel_one_hot_i[38];
  assign data_masked[4912] = data_i[4912] & sel_one_hot_i[38];
  assign data_masked[4911] = data_i[4911] & sel_one_hot_i[38];
  assign data_masked[4910] = data_i[4910] & sel_one_hot_i[38];
  assign data_masked[4909] = data_i[4909] & sel_one_hot_i[38];
  assign data_masked[4908] = data_i[4908] & sel_one_hot_i[38];
  assign data_masked[4907] = data_i[4907] & sel_one_hot_i[38];
  assign data_masked[4906] = data_i[4906] & sel_one_hot_i[38];
  assign data_masked[4905] = data_i[4905] & sel_one_hot_i[38];
  assign data_masked[4904] = data_i[4904] & sel_one_hot_i[38];
  assign data_masked[4903] = data_i[4903] & sel_one_hot_i[38];
  assign data_masked[4902] = data_i[4902] & sel_one_hot_i[38];
  assign data_masked[4901] = data_i[4901] & sel_one_hot_i[38];
  assign data_masked[4900] = data_i[4900] & sel_one_hot_i[38];
  assign data_masked[4899] = data_i[4899] & sel_one_hot_i[38];
  assign data_masked[4898] = data_i[4898] & sel_one_hot_i[38];
  assign data_masked[4897] = data_i[4897] & sel_one_hot_i[38];
  assign data_masked[4896] = data_i[4896] & sel_one_hot_i[38];
  assign data_masked[4895] = data_i[4895] & sel_one_hot_i[38];
  assign data_masked[4894] = data_i[4894] & sel_one_hot_i[38];
  assign data_masked[4893] = data_i[4893] & sel_one_hot_i[38];
  assign data_masked[4892] = data_i[4892] & sel_one_hot_i[38];
  assign data_masked[4891] = data_i[4891] & sel_one_hot_i[38];
  assign data_masked[4890] = data_i[4890] & sel_one_hot_i[38];
  assign data_masked[4889] = data_i[4889] & sel_one_hot_i[38];
  assign data_masked[4888] = data_i[4888] & sel_one_hot_i[38];
  assign data_masked[4887] = data_i[4887] & sel_one_hot_i[38];
  assign data_masked[4886] = data_i[4886] & sel_one_hot_i[38];
  assign data_masked[4885] = data_i[4885] & sel_one_hot_i[38];
  assign data_masked[4884] = data_i[4884] & sel_one_hot_i[38];
  assign data_masked[4883] = data_i[4883] & sel_one_hot_i[38];
  assign data_masked[4882] = data_i[4882] & sel_one_hot_i[38];
  assign data_masked[4881] = data_i[4881] & sel_one_hot_i[38];
  assign data_masked[4880] = data_i[4880] & sel_one_hot_i[38];
  assign data_masked[4879] = data_i[4879] & sel_one_hot_i[38];
  assign data_masked[4878] = data_i[4878] & sel_one_hot_i[38];
  assign data_masked[4877] = data_i[4877] & sel_one_hot_i[38];
  assign data_masked[4876] = data_i[4876] & sel_one_hot_i[38];
  assign data_masked[4875] = data_i[4875] & sel_one_hot_i[38];
  assign data_masked[4874] = data_i[4874] & sel_one_hot_i[38];
  assign data_masked[4873] = data_i[4873] & sel_one_hot_i[38];
  assign data_masked[4872] = data_i[4872] & sel_one_hot_i[38];
  assign data_masked[4871] = data_i[4871] & sel_one_hot_i[38];
  assign data_masked[4870] = data_i[4870] & sel_one_hot_i[38];
  assign data_masked[4869] = data_i[4869] & sel_one_hot_i[38];
  assign data_masked[4868] = data_i[4868] & sel_one_hot_i[38];
  assign data_masked[4867] = data_i[4867] & sel_one_hot_i[38];
  assign data_masked[4866] = data_i[4866] & sel_one_hot_i[38];
  assign data_masked[4865] = data_i[4865] & sel_one_hot_i[38];
  assign data_masked[4864] = data_i[4864] & sel_one_hot_i[38];
  assign data_masked[5119] = data_i[5119] & sel_one_hot_i[39];
  assign data_masked[5118] = data_i[5118] & sel_one_hot_i[39];
  assign data_masked[5117] = data_i[5117] & sel_one_hot_i[39];
  assign data_masked[5116] = data_i[5116] & sel_one_hot_i[39];
  assign data_masked[5115] = data_i[5115] & sel_one_hot_i[39];
  assign data_masked[5114] = data_i[5114] & sel_one_hot_i[39];
  assign data_masked[5113] = data_i[5113] & sel_one_hot_i[39];
  assign data_masked[5112] = data_i[5112] & sel_one_hot_i[39];
  assign data_masked[5111] = data_i[5111] & sel_one_hot_i[39];
  assign data_masked[5110] = data_i[5110] & sel_one_hot_i[39];
  assign data_masked[5109] = data_i[5109] & sel_one_hot_i[39];
  assign data_masked[5108] = data_i[5108] & sel_one_hot_i[39];
  assign data_masked[5107] = data_i[5107] & sel_one_hot_i[39];
  assign data_masked[5106] = data_i[5106] & sel_one_hot_i[39];
  assign data_masked[5105] = data_i[5105] & sel_one_hot_i[39];
  assign data_masked[5104] = data_i[5104] & sel_one_hot_i[39];
  assign data_masked[5103] = data_i[5103] & sel_one_hot_i[39];
  assign data_masked[5102] = data_i[5102] & sel_one_hot_i[39];
  assign data_masked[5101] = data_i[5101] & sel_one_hot_i[39];
  assign data_masked[5100] = data_i[5100] & sel_one_hot_i[39];
  assign data_masked[5099] = data_i[5099] & sel_one_hot_i[39];
  assign data_masked[5098] = data_i[5098] & sel_one_hot_i[39];
  assign data_masked[5097] = data_i[5097] & sel_one_hot_i[39];
  assign data_masked[5096] = data_i[5096] & sel_one_hot_i[39];
  assign data_masked[5095] = data_i[5095] & sel_one_hot_i[39];
  assign data_masked[5094] = data_i[5094] & sel_one_hot_i[39];
  assign data_masked[5093] = data_i[5093] & sel_one_hot_i[39];
  assign data_masked[5092] = data_i[5092] & sel_one_hot_i[39];
  assign data_masked[5091] = data_i[5091] & sel_one_hot_i[39];
  assign data_masked[5090] = data_i[5090] & sel_one_hot_i[39];
  assign data_masked[5089] = data_i[5089] & sel_one_hot_i[39];
  assign data_masked[5088] = data_i[5088] & sel_one_hot_i[39];
  assign data_masked[5087] = data_i[5087] & sel_one_hot_i[39];
  assign data_masked[5086] = data_i[5086] & sel_one_hot_i[39];
  assign data_masked[5085] = data_i[5085] & sel_one_hot_i[39];
  assign data_masked[5084] = data_i[5084] & sel_one_hot_i[39];
  assign data_masked[5083] = data_i[5083] & sel_one_hot_i[39];
  assign data_masked[5082] = data_i[5082] & sel_one_hot_i[39];
  assign data_masked[5081] = data_i[5081] & sel_one_hot_i[39];
  assign data_masked[5080] = data_i[5080] & sel_one_hot_i[39];
  assign data_masked[5079] = data_i[5079] & sel_one_hot_i[39];
  assign data_masked[5078] = data_i[5078] & sel_one_hot_i[39];
  assign data_masked[5077] = data_i[5077] & sel_one_hot_i[39];
  assign data_masked[5076] = data_i[5076] & sel_one_hot_i[39];
  assign data_masked[5075] = data_i[5075] & sel_one_hot_i[39];
  assign data_masked[5074] = data_i[5074] & sel_one_hot_i[39];
  assign data_masked[5073] = data_i[5073] & sel_one_hot_i[39];
  assign data_masked[5072] = data_i[5072] & sel_one_hot_i[39];
  assign data_masked[5071] = data_i[5071] & sel_one_hot_i[39];
  assign data_masked[5070] = data_i[5070] & sel_one_hot_i[39];
  assign data_masked[5069] = data_i[5069] & sel_one_hot_i[39];
  assign data_masked[5068] = data_i[5068] & sel_one_hot_i[39];
  assign data_masked[5067] = data_i[5067] & sel_one_hot_i[39];
  assign data_masked[5066] = data_i[5066] & sel_one_hot_i[39];
  assign data_masked[5065] = data_i[5065] & sel_one_hot_i[39];
  assign data_masked[5064] = data_i[5064] & sel_one_hot_i[39];
  assign data_masked[5063] = data_i[5063] & sel_one_hot_i[39];
  assign data_masked[5062] = data_i[5062] & sel_one_hot_i[39];
  assign data_masked[5061] = data_i[5061] & sel_one_hot_i[39];
  assign data_masked[5060] = data_i[5060] & sel_one_hot_i[39];
  assign data_masked[5059] = data_i[5059] & sel_one_hot_i[39];
  assign data_masked[5058] = data_i[5058] & sel_one_hot_i[39];
  assign data_masked[5057] = data_i[5057] & sel_one_hot_i[39];
  assign data_masked[5056] = data_i[5056] & sel_one_hot_i[39];
  assign data_masked[5055] = data_i[5055] & sel_one_hot_i[39];
  assign data_masked[5054] = data_i[5054] & sel_one_hot_i[39];
  assign data_masked[5053] = data_i[5053] & sel_one_hot_i[39];
  assign data_masked[5052] = data_i[5052] & sel_one_hot_i[39];
  assign data_masked[5051] = data_i[5051] & sel_one_hot_i[39];
  assign data_masked[5050] = data_i[5050] & sel_one_hot_i[39];
  assign data_masked[5049] = data_i[5049] & sel_one_hot_i[39];
  assign data_masked[5048] = data_i[5048] & sel_one_hot_i[39];
  assign data_masked[5047] = data_i[5047] & sel_one_hot_i[39];
  assign data_masked[5046] = data_i[5046] & sel_one_hot_i[39];
  assign data_masked[5045] = data_i[5045] & sel_one_hot_i[39];
  assign data_masked[5044] = data_i[5044] & sel_one_hot_i[39];
  assign data_masked[5043] = data_i[5043] & sel_one_hot_i[39];
  assign data_masked[5042] = data_i[5042] & sel_one_hot_i[39];
  assign data_masked[5041] = data_i[5041] & sel_one_hot_i[39];
  assign data_masked[5040] = data_i[5040] & sel_one_hot_i[39];
  assign data_masked[5039] = data_i[5039] & sel_one_hot_i[39];
  assign data_masked[5038] = data_i[5038] & sel_one_hot_i[39];
  assign data_masked[5037] = data_i[5037] & sel_one_hot_i[39];
  assign data_masked[5036] = data_i[5036] & sel_one_hot_i[39];
  assign data_masked[5035] = data_i[5035] & sel_one_hot_i[39];
  assign data_masked[5034] = data_i[5034] & sel_one_hot_i[39];
  assign data_masked[5033] = data_i[5033] & sel_one_hot_i[39];
  assign data_masked[5032] = data_i[5032] & sel_one_hot_i[39];
  assign data_masked[5031] = data_i[5031] & sel_one_hot_i[39];
  assign data_masked[5030] = data_i[5030] & sel_one_hot_i[39];
  assign data_masked[5029] = data_i[5029] & sel_one_hot_i[39];
  assign data_masked[5028] = data_i[5028] & sel_one_hot_i[39];
  assign data_masked[5027] = data_i[5027] & sel_one_hot_i[39];
  assign data_masked[5026] = data_i[5026] & sel_one_hot_i[39];
  assign data_masked[5025] = data_i[5025] & sel_one_hot_i[39];
  assign data_masked[5024] = data_i[5024] & sel_one_hot_i[39];
  assign data_masked[5023] = data_i[5023] & sel_one_hot_i[39];
  assign data_masked[5022] = data_i[5022] & sel_one_hot_i[39];
  assign data_masked[5021] = data_i[5021] & sel_one_hot_i[39];
  assign data_masked[5020] = data_i[5020] & sel_one_hot_i[39];
  assign data_masked[5019] = data_i[5019] & sel_one_hot_i[39];
  assign data_masked[5018] = data_i[5018] & sel_one_hot_i[39];
  assign data_masked[5017] = data_i[5017] & sel_one_hot_i[39];
  assign data_masked[5016] = data_i[5016] & sel_one_hot_i[39];
  assign data_masked[5015] = data_i[5015] & sel_one_hot_i[39];
  assign data_masked[5014] = data_i[5014] & sel_one_hot_i[39];
  assign data_masked[5013] = data_i[5013] & sel_one_hot_i[39];
  assign data_masked[5012] = data_i[5012] & sel_one_hot_i[39];
  assign data_masked[5011] = data_i[5011] & sel_one_hot_i[39];
  assign data_masked[5010] = data_i[5010] & sel_one_hot_i[39];
  assign data_masked[5009] = data_i[5009] & sel_one_hot_i[39];
  assign data_masked[5008] = data_i[5008] & sel_one_hot_i[39];
  assign data_masked[5007] = data_i[5007] & sel_one_hot_i[39];
  assign data_masked[5006] = data_i[5006] & sel_one_hot_i[39];
  assign data_masked[5005] = data_i[5005] & sel_one_hot_i[39];
  assign data_masked[5004] = data_i[5004] & sel_one_hot_i[39];
  assign data_masked[5003] = data_i[5003] & sel_one_hot_i[39];
  assign data_masked[5002] = data_i[5002] & sel_one_hot_i[39];
  assign data_masked[5001] = data_i[5001] & sel_one_hot_i[39];
  assign data_masked[5000] = data_i[5000] & sel_one_hot_i[39];
  assign data_masked[4999] = data_i[4999] & sel_one_hot_i[39];
  assign data_masked[4998] = data_i[4998] & sel_one_hot_i[39];
  assign data_masked[4997] = data_i[4997] & sel_one_hot_i[39];
  assign data_masked[4996] = data_i[4996] & sel_one_hot_i[39];
  assign data_masked[4995] = data_i[4995] & sel_one_hot_i[39];
  assign data_masked[4994] = data_i[4994] & sel_one_hot_i[39];
  assign data_masked[4993] = data_i[4993] & sel_one_hot_i[39];
  assign data_masked[4992] = data_i[4992] & sel_one_hot_i[39];
  assign data_masked[5247] = data_i[5247] & sel_one_hot_i[40];
  assign data_masked[5246] = data_i[5246] & sel_one_hot_i[40];
  assign data_masked[5245] = data_i[5245] & sel_one_hot_i[40];
  assign data_masked[5244] = data_i[5244] & sel_one_hot_i[40];
  assign data_masked[5243] = data_i[5243] & sel_one_hot_i[40];
  assign data_masked[5242] = data_i[5242] & sel_one_hot_i[40];
  assign data_masked[5241] = data_i[5241] & sel_one_hot_i[40];
  assign data_masked[5240] = data_i[5240] & sel_one_hot_i[40];
  assign data_masked[5239] = data_i[5239] & sel_one_hot_i[40];
  assign data_masked[5238] = data_i[5238] & sel_one_hot_i[40];
  assign data_masked[5237] = data_i[5237] & sel_one_hot_i[40];
  assign data_masked[5236] = data_i[5236] & sel_one_hot_i[40];
  assign data_masked[5235] = data_i[5235] & sel_one_hot_i[40];
  assign data_masked[5234] = data_i[5234] & sel_one_hot_i[40];
  assign data_masked[5233] = data_i[5233] & sel_one_hot_i[40];
  assign data_masked[5232] = data_i[5232] & sel_one_hot_i[40];
  assign data_masked[5231] = data_i[5231] & sel_one_hot_i[40];
  assign data_masked[5230] = data_i[5230] & sel_one_hot_i[40];
  assign data_masked[5229] = data_i[5229] & sel_one_hot_i[40];
  assign data_masked[5228] = data_i[5228] & sel_one_hot_i[40];
  assign data_masked[5227] = data_i[5227] & sel_one_hot_i[40];
  assign data_masked[5226] = data_i[5226] & sel_one_hot_i[40];
  assign data_masked[5225] = data_i[5225] & sel_one_hot_i[40];
  assign data_masked[5224] = data_i[5224] & sel_one_hot_i[40];
  assign data_masked[5223] = data_i[5223] & sel_one_hot_i[40];
  assign data_masked[5222] = data_i[5222] & sel_one_hot_i[40];
  assign data_masked[5221] = data_i[5221] & sel_one_hot_i[40];
  assign data_masked[5220] = data_i[5220] & sel_one_hot_i[40];
  assign data_masked[5219] = data_i[5219] & sel_one_hot_i[40];
  assign data_masked[5218] = data_i[5218] & sel_one_hot_i[40];
  assign data_masked[5217] = data_i[5217] & sel_one_hot_i[40];
  assign data_masked[5216] = data_i[5216] & sel_one_hot_i[40];
  assign data_masked[5215] = data_i[5215] & sel_one_hot_i[40];
  assign data_masked[5214] = data_i[5214] & sel_one_hot_i[40];
  assign data_masked[5213] = data_i[5213] & sel_one_hot_i[40];
  assign data_masked[5212] = data_i[5212] & sel_one_hot_i[40];
  assign data_masked[5211] = data_i[5211] & sel_one_hot_i[40];
  assign data_masked[5210] = data_i[5210] & sel_one_hot_i[40];
  assign data_masked[5209] = data_i[5209] & sel_one_hot_i[40];
  assign data_masked[5208] = data_i[5208] & sel_one_hot_i[40];
  assign data_masked[5207] = data_i[5207] & sel_one_hot_i[40];
  assign data_masked[5206] = data_i[5206] & sel_one_hot_i[40];
  assign data_masked[5205] = data_i[5205] & sel_one_hot_i[40];
  assign data_masked[5204] = data_i[5204] & sel_one_hot_i[40];
  assign data_masked[5203] = data_i[5203] & sel_one_hot_i[40];
  assign data_masked[5202] = data_i[5202] & sel_one_hot_i[40];
  assign data_masked[5201] = data_i[5201] & sel_one_hot_i[40];
  assign data_masked[5200] = data_i[5200] & sel_one_hot_i[40];
  assign data_masked[5199] = data_i[5199] & sel_one_hot_i[40];
  assign data_masked[5198] = data_i[5198] & sel_one_hot_i[40];
  assign data_masked[5197] = data_i[5197] & sel_one_hot_i[40];
  assign data_masked[5196] = data_i[5196] & sel_one_hot_i[40];
  assign data_masked[5195] = data_i[5195] & sel_one_hot_i[40];
  assign data_masked[5194] = data_i[5194] & sel_one_hot_i[40];
  assign data_masked[5193] = data_i[5193] & sel_one_hot_i[40];
  assign data_masked[5192] = data_i[5192] & sel_one_hot_i[40];
  assign data_masked[5191] = data_i[5191] & sel_one_hot_i[40];
  assign data_masked[5190] = data_i[5190] & sel_one_hot_i[40];
  assign data_masked[5189] = data_i[5189] & sel_one_hot_i[40];
  assign data_masked[5188] = data_i[5188] & sel_one_hot_i[40];
  assign data_masked[5187] = data_i[5187] & sel_one_hot_i[40];
  assign data_masked[5186] = data_i[5186] & sel_one_hot_i[40];
  assign data_masked[5185] = data_i[5185] & sel_one_hot_i[40];
  assign data_masked[5184] = data_i[5184] & sel_one_hot_i[40];
  assign data_masked[5183] = data_i[5183] & sel_one_hot_i[40];
  assign data_masked[5182] = data_i[5182] & sel_one_hot_i[40];
  assign data_masked[5181] = data_i[5181] & sel_one_hot_i[40];
  assign data_masked[5180] = data_i[5180] & sel_one_hot_i[40];
  assign data_masked[5179] = data_i[5179] & sel_one_hot_i[40];
  assign data_masked[5178] = data_i[5178] & sel_one_hot_i[40];
  assign data_masked[5177] = data_i[5177] & sel_one_hot_i[40];
  assign data_masked[5176] = data_i[5176] & sel_one_hot_i[40];
  assign data_masked[5175] = data_i[5175] & sel_one_hot_i[40];
  assign data_masked[5174] = data_i[5174] & sel_one_hot_i[40];
  assign data_masked[5173] = data_i[5173] & sel_one_hot_i[40];
  assign data_masked[5172] = data_i[5172] & sel_one_hot_i[40];
  assign data_masked[5171] = data_i[5171] & sel_one_hot_i[40];
  assign data_masked[5170] = data_i[5170] & sel_one_hot_i[40];
  assign data_masked[5169] = data_i[5169] & sel_one_hot_i[40];
  assign data_masked[5168] = data_i[5168] & sel_one_hot_i[40];
  assign data_masked[5167] = data_i[5167] & sel_one_hot_i[40];
  assign data_masked[5166] = data_i[5166] & sel_one_hot_i[40];
  assign data_masked[5165] = data_i[5165] & sel_one_hot_i[40];
  assign data_masked[5164] = data_i[5164] & sel_one_hot_i[40];
  assign data_masked[5163] = data_i[5163] & sel_one_hot_i[40];
  assign data_masked[5162] = data_i[5162] & sel_one_hot_i[40];
  assign data_masked[5161] = data_i[5161] & sel_one_hot_i[40];
  assign data_masked[5160] = data_i[5160] & sel_one_hot_i[40];
  assign data_masked[5159] = data_i[5159] & sel_one_hot_i[40];
  assign data_masked[5158] = data_i[5158] & sel_one_hot_i[40];
  assign data_masked[5157] = data_i[5157] & sel_one_hot_i[40];
  assign data_masked[5156] = data_i[5156] & sel_one_hot_i[40];
  assign data_masked[5155] = data_i[5155] & sel_one_hot_i[40];
  assign data_masked[5154] = data_i[5154] & sel_one_hot_i[40];
  assign data_masked[5153] = data_i[5153] & sel_one_hot_i[40];
  assign data_masked[5152] = data_i[5152] & sel_one_hot_i[40];
  assign data_masked[5151] = data_i[5151] & sel_one_hot_i[40];
  assign data_masked[5150] = data_i[5150] & sel_one_hot_i[40];
  assign data_masked[5149] = data_i[5149] & sel_one_hot_i[40];
  assign data_masked[5148] = data_i[5148] & sel_one_hot_i[40];
  assign data_masked[5147] = data_i[5147] & sel_one_hot_i[40];
  assign data_masked[5146] = data_i[5146] & sel_one_hot_i[40];
  assign data_masked[5145] = data_i[5145] & sel_one_hot_i[40];
  assign data_masked[5144] = data_i[5144] & sel_one_hot_i[40];
  assign data_masked[5143] = data_i[5143] & sel_one_hot_i[40];
  assign data_masked[5142] = data_i[5142] & sel_one_hot_i[40];
  assign data_masked[5141] = data_i[5141] & sel_one_hot_i[40];
  assign data_masked[5140] = data_i[5140] & sel_one_hot_i[40];
  assign data_masked[5139] = data_i[5139] & sel_one_hot_i[40];
  assign data_masked[5138] = data_i[5138] & sel_one_hot_i[40];
  assign data_masked[5137] = data_i[5137] & sel_one_hot_i[40];
  assign data_masked[5136] = data_i[5136] & sel_one_hot_i[40];
  assign data_masked[5135] = data_i[5135] & sel_one_hot_i[40];
  assign data_masked[5134] = data_i[5134] & sel_one_hot_i[40];
  assign data_masked[5133] = data_i[5133] & sel_one_hot_i[40];
  assign data_masked[5132] = data_i[5132] & sel_one_hot_i[40];
  assign data_masked[5131] = data_i[5131] & sel_one_hot_i[40];
  assign data_masked[5130] = data_i[5130] & sel_one_hot_i[40];
  assign data_masked[5129] = data_i[5129] & sel_one_hot_i[40];
  assign data_masked[5128] = data_i[5128] & sel_one_hot_i[40];
  assign data_masked[5127] = data_i[5127] & sel_one_hot_i[40];
  assign data_masked[5126] = data_i[5126] & sel_one_hot_i[40];
  assign data_masked[5125] = data_i[5125] & sel_one_hot_i[40];
  assign data_masked[5124] = data_i[5124] & sel_one_hot_i[40];
  assign data_masked[5123] = data_i[5123] & sel_one_hot_i[40];
  assign data_masked[5122] = data_i[5122] & sel_one_hot_i[40];
  assign data_masked[5121] = data_i[5121] & sel_one_hot_i[40];
  assign data_masked[5120] = data_i[5120] & sel_one_hot_i[40];
  assign data_masked[5375] = data_i[5375] & sel_one_hot_i[41];
  assign data_masked[5374] = data_i[5374] & sel_one_hot_i[41];
  assign data_masked[5373] = data_i[5373] & sel_one_hot_i[41];
  assign data_masked[5372] = data_i[5372] & sel_one_hot_i[41];
  assign data_masked[5371] = data_i[5371] & sel_one_hot_i[41];
  assign data_masked[5370] = data_i[5370] & sel_one_hot_i[41];
  assign data_masked[5369] = data_i[5369] & sel_one_hot_i[41];
  assign data_masked[5368] = data_i[5368] & sel_one_hot_i[41];
  assign data_masked[5367] = data_i[5367] & sel_one_hot_i[41];
  assign data_masked[5366] = data_i[5366] & sel_one_hot_i[41];
  assign data_masked[5365] = data_i[5365] & sel_one_hot_i[41];
  assign data_masked[5364] = data_i[5364] & sel_one_hot_i[41];
  assign data_masked[5363] = data_i[5363] & sel_one_hot_i[41];
  assign data_masked[5362] = data_i[5362] & sel_one_hot_i[41];
  assign data_masked[5361] = data_i[5361] & sel_one_hot_i[41];
  assign data_masked[5360] = data_i[5360] & sel_one_hot_i[41];
  assign data_masked[5359] = data_i[5359] & sel_one_hot_i[41];
  assign data_masked[5358] = data_i[5358] & sel_one_hot_i[41];
  assign data_masked[5357] = data_i[5357] & sel_one_hot_i[41];
  assign data_masked[5356] = data_i[5356] & sel_one_hot_i[41];
  assign data_masked[5355] = data_i[5355] & sel_one_hot_i[41];
  assign data_masked[5354] = data_i[5354] & sel_one_hot_i[41];
  assign data_masked[5353] = data_i[5353] & sel_one_hot_i[41];
  assign data_masked[5352] = data_i[5352] & sel_one_hot_i[41];
  assign data_masked[5351] = data_i[5351] & sel_one_hot_i[41];
  assign data_masked[5350] = data_i[5350] & sel_one_hot_i[41];
  assign data_masked[5349] = data_i[5349] & sel_one_hot_i[41];
  assign data_masked[5348] = data_i[5348] & sel_one_hot_i[41];
  assign data_masked[5347] = data_i[5347] & sel_one_hot_i[41];
  assign data_masked[5346] = data_i[5346] & sel_one_hot_i[41];
  assign data_masked[5345] = data_i[5345] & sel_one_hot_i[41];
  assign data_masked[5344] = data_i[5344] & sel_one_hot_i[41];
  assign data_masked[5343] = data_i[5343] & sel_one_hot_i[41];
  assign data_masked[5342] = data_i[5342] & sel_one_hot_i[41];
  assign data_masked[5341] = data_i[5341] & sel_one_hot_i[41];
  assign data_masked[5340] = data_i[5340] & sel_one_hot_i[41];
  assign data_masked[5339] = data_i[5339] & sel_one_hot_i[41];
  assign data_masked[5338] = data_i[5338] & sel_one_hot_i[41];
  assign data_masked[5337] = data_i[5337] & sel_one_hot_i[41];
  assign data_masked[5336] = data_i[5336] & sel_one_hot_i[41];
  assign data_masked[5335] = data_i[5335] & sel_one_hot_i[41];
  assign data_masked[5334] = data_i[5334] & sel_one_hot_i[41];
  assign data_masked[5333] = data_i[5333] & sel_one_hot_i[41];
  assign data_masked[5332] = data_i[5332] & sel_one_hot_i[41];
  assign data_masked[5331] = data_i[5331] & sel_one_hot_i[41];
  assign data_masked[5330] = data_i[5330] & sel_one_hot_i[41];
  assign data_masked[5329] = data_i[5329] & sel_one_hot_i[41];
  assign data_masked[5328] = data_i[5328] & sel_one_hot_i[41];
  assign data_masked[5327] = data_i[5327] & sel_one_hot_i[41];
  assign data_masked[5326] = data_i[5326] & sel_one_hot_i[41];
  assign data_masked[5325] = data_i[5325] & sel_one_hot_i[41];
  assign data_masked[5324] = data_i[5324] & sel_one_hot_i[41];
  assign data_masked[5323] = data_i[5323] & sel_one_hot_i[41];
  assign data_masked[5322] = data_i[5322] & sel_one_hot_i[41];
  assign data_masked[5321] = data_i[5321] & sel_one_hot_i[41];
  assign data_masked[5320] = data_i[5320] & sel_one_hot_i[41];
  assign data_masked[5319] = data_i[5319] & sel_one_hot_i[41];
  assign data_masked[5318] = data_i[5318] & sel_one_hot_i[41];
  assign data_masked[5317] = data_i[5317] & sel_one_hot_i[41];
  assign data_masked[5316] = data_i[5316] & sel_one_hot_i[41];
  assign data_masked[5315] = data_i[5315] & sel_one_hot_i[41];
  assign data_masked[5314] = data_i[5314] & sel_one_hot_i[41];
  assign data_masked[5313] = data_i[5313] & sel_one_hot_i[41];
  assign data_masked[5312] = data_i[5312] & sel_one_hot_i[41];
  assign data_masked[5311] = data_i[5311] & sel_one_hot_i[41];
  assign data_masked[5310] = data_i[5310] & sel_one_hot_i[41];
  assign data_masked[5309] = data_i[5309] & sel_one_hot_i[41];
  assign data_masked[5308] = data_i[5308] & sel_one_hot_i[41];
  assign data_masked[5307] = data_i[5307] & sel_one_hot_i[41];
  assign data_masked[5306] = data_i[5306] & sel_one_hot_i[41];
  assign data_masked[5305] = data_i[5305] & sel_one_hot_i[41];
  assign data_masked[5304] = data_i[5304] & sel_one_hot_i[41];
  assign data_masked[5303] = data_i[5303] & sel_one_hot_i[41];
  assign data_masked[5302] = data_i[5302] & sel_one_hot_i[41];
  assign data_masked[5301] = data_i[5301] & sel_one_hot_i[41];
  assign data_masked[5300] = data_i[5300] & sel_one_hot_i[41];
  assign data_masked[5299] = data_i[5299] & sel_one_hot_i[41];
  assign data_masked[5298] = data_i[5298] & sel_one_hot_i[41];
  assign data_masked[5297] = data_i[5297] & sel_one_hot_i[41];
  assign data_masked[5296] = data_i[5296] & sel_one_hot_i[41];
  assign data_masked[5295] = data_i[5295] & sel_one_hot_i[41];
  assign data_masked[5294] = data_i[5294] & sel_one_hot_i[41];
  assign data_masked[5293] = data_i[5293] & sel_one_hot_i[41];
  assign data_masked[5292] = data_i[5292] & sel_one_hot_i[41];
  assign data_masked[5291] = data_i[5291] & sel_one_hot_i[41];
  assign data_masked[5290] = data_i[5290] & sel_one_hot_i[41];
  assign data_masked[5289] = data_i[5289] & sel_one_hot_i[41];
  assign data_masked[5288] = data_i[5288] & sel_one_hot_i[41];
  assign data_masked[5287] = data_i[5287] & sel_one_hot_i[41];
  assign data_masked[5286] = data_i[5286] & sel_one_hot_i[41];
  assign data_masked[5285] = data_i[5285] & sel_one_hot_i[41];
  assign data_masked[5284] = data_i[5284] & sel_one_hot_i[41];
  assign data_masked[5283] = data_i[5283] & sel_one_hot_i[41];
  assign data_masked[5282] = data_i[5282] & sel_one_hot_i[41];
  assign data_masked[5281] = data_i[5281] & sel_one_hot_i[41];
  assign data_masked[5280] = data_i[5280] & sel_one_hot_i[41];
  assign data_masked[5279] = data_i[5279] & sel_one_hot_i[41];
  assign data_masked[5278] = data_i[5278] & sel_one_hot_i[41];
  assign data_masked[5277] = data_i[5277] & sel_one_hot_i[41];
  assign data_masked[5276] = data_i[5276] & sel_one_hot_i[41];
  assign data_masked[5275] = data_i[5275] & sel_one_hot_i[41];
  assign data_masked[5274] = data_i[5274] & sel_one_hot_i[41];
  assign data_masked[5273] = data_i[5273] & sel_one_hot_i[41];
  assign data_masked[5272] = data_i[5272] & sel_one_hot_i[41];
  assign data_masked[5271] = data_i[5271] & sel_one_hot_i[41];
  assign data_masked[5270] = data_i[5270] & sel_one_hot_i[41];
  assign data_masked[5269] = data_i[5269] & sel_one_hot_i[41];
  assign data_masked[5268] = data_i[5268] & sel_one_hot_i[41];
  assign data_masked[5267] = data_i[5267] & sel_one_hot_i[41];
  assign data_masked[5266] = data_i[5266] & sel_one_hot_i[41];
  assign data_masked[5265] = data_i[5265] & sel_one_hot_i[41];
  assign data_masked[5264] = data_i[5264] & sel_one_hot_i[41];
  assign data_masked[5263] = data_i[5263] & sel_one_hot_i[41];
  assign data_masked[5262] = data_i[5262] & sel_one_hot_i[41];
  assign data_masked[5261] = data_i[5261] & sel_one_hot_i[41];
  assign data_masked[5260] = data_i[5260] & sel_one_hot_i[41];
  assign data_masked[5259] = data_i[5259] & sel_one_hot_i[41];
  assign data_masked[5258] = data_i[5258] & sel_one_hot_i[41];
  assign data_masked[5257] = data_i[5257] & sel_one_hot_i[41];
  assign data_masked[5256] = data_i[5256] & sel_one_hot_i[41];
  assign data_masked[5255] = data_i[5255] & sel_one_hot_i[41];
  assign data_masked[5254] = data_i[5254] & sel_one_hot_i[41];
  assign data_masked[5253] = data_i[5253] & sel_one_hot_i[41];
  assign data_masked[5252] = data_i[5252] & sel_one_hot_i[41];
  assign data_masked[5251] = data_i[5251] & sel_one_hot_i[41];
  assign data_masked[5250] = data_i[5250] & sel_one_hot_i[41];
  assign data_masked[5249] = data_i[5249] & sel_one_hot_i[41];
  assign data_masked[5248] = data_i[5248] & sel_one_hot_i[41];
  assign data_masked[5503] = data_i[5503] & sel_one_hot_i[42];
  assign data_masked[5502] = data_i[5502] & sel_one_hot_i[42];
  assign data_masked[5501] = data_i[5501] & sel_one_hot_i[42];
  assign data_masked[5500] = data_i[5500] & sel_one_hot_i[42];
  assign data_masked[5499] = data_i[5499] & sel_one_hot_i[42];
  assign data_masked[5498] = data_i[5498] & sel_one_hot_i[42];
  assign data_masked[5497] = data_i[5497] & sel_one_hot_i[42];
  assign data_masked[5496] = data_i[5496] & sel_one_hot_i[42];
  assign data_masked[5495] = data_i[5495] & sel_one_hot_i[42];
  assign data_masked[5494] = data_i[5494] & sel_one_hot_i[42];
  assign data_masked[5493] = data_i[5493] & sel_one_hot_i[42];
  assign data_masked[5492] = data_i[5492] & sel_one_hot_i[42];
  assign data_masked[5491] = data_i[5491] & sel_one_hot_i[42];
  assign data_masked[5490] = data_i[5490] & sel_one_hot_i[42];
  assign data_masked[5489] = data_i[5489] & sel_one_hot_i[42];
  assign data_masked[5488] = data_i[5488] & sel_one_hot_i[42];
  assign data_masked[5487] = data_i[5487] & sel_one_hot_i[42];
  assign data_masked[5486] = data_i[5486] & sel_one_hot_i[42];
  assign data_masked[5485] = data_i[5485] & sel_one_hot_i[42];
  assign data_masked[5484] = data_i[5484] & sel_one_hot_i[42];
  assign data_masked[5483] = data_i[5483] & sel_one_hot_i[42];
  assign data_masked[5482] = data_i[5482] & sel_one_hot_i[42];
  assign data_masked[5481] = data_i[5481] & sel_one_hot_i[42];
  assign data_masked[5480] = data_i[5480] & sel_one_hot_i[42];
  assign data_masked[5479] = data_i[5479] & sel_one_hot_i[42];
  assign data_masked[5478] = data_i[5478] & sel_one_hot_i[42];
  assign data_masked[5477] = data_i[5477] & sel_one_hot_i[42];
  assign data_masked[5476] = data_i[5476] & sel_one_hot_i[42];
  assign data_masked[5475] = data_i[5475] & sel_one_hot_i[42];
  assign data_masked[5474] = data_i[5474] & sel_one_hot_i[42];
  assign data_masked[5473] = data_i[5473] & sel_one_hot_i[42];
  assign data_masked[5472] = data_i[5472] & sel_one_hot_i[42];
  assign data_masked[5471] = data_i[5471] & sel_one_hot_i[42];
  assign data_masked[5470] = data_i[5470] & sel_one_hot_i[42];
  assign data_masked[5469] = data_i[5469] & sel_one_hot_i[42];
  assign data_masked[5468] = data_i[5468] & sel_one_hot_i[42];
  assign data_masked[5467] = data_i[5467] & sel_one_hot_i[42];
  assign data_masked[5466] = data_i[5466] & sel_one_hot_i[42];
  assign data_masked[5465] = data_i[5465] & sel_one_hot_i[42];
  assign data_masked[5464] = data_i[5464] & sel_one_hot_i[42];
  assign data_masked[5463] = data_i[5463] & sel_one_hot_i[42];
  assign data_masked[5462] = data_i[5462] & sel_one_hot_i[42];
  assign data_masked[5461] = data_i[5461] & sel_one_hot_i[42];
  assign data_masked[5460] = data_i[5460] & sel_one_hot_i[42];
  assign data_masked[5459] = data_i[5459] & sel_one_hot_i[42];
  assign data_masked[5458] = data_i[5458] & sel_one_hot_i[42];
  assign data_masked[5457] = data_i[5457] & sel_one_hot_i[42];
  assign data_masked[5456] = data_i[5456] & sel_one_hot_i[42];
  assign data_masked[5455] = data_i[5455] & sel_one_hot_i[42];
  assign data_masked[5454] = data_i[5454] & sel_one_hot_i[42];
  assign data_masked[5453] = data_i[5453] & sel_one_hot_i[42];
  assign data_masked[5452] = data_i[5452] & sel_one_hot_i[42];
  assign data_masked[5451] = data_i[5451] & sel_one_hot_i[42];
  assign data_masked[5450] = data_i[5450] & sel_one_hot_i[42];
  assign data_masked[5449] = data_i[5449] & sel_one_hot_i[42];
  assign data_masked[5448] = data_i[5448] & sel_one_hot_i[42];
  assign data_masked[5447] = data_i[5447] & sel_one_hot_i[42];
  assign data_masked[5446] = data_i[5446] & sel_one_hot_i[42];
  assign data_masked[5445] = data_i[5445] & sel_one_hot_i[42];
  assign data_masked[5444] = data_i[5444] & sel_one_hot_i[42];
  assign data_masked[5443] = data_i[5443] & sel_one_hot_i[42];
  assign data_masked[5442] = data_i[5442] & sel_one_hot_i[42];
  assign data_masked[5441] = data_i[5441] & sel_one_hot_i[42];
  assign data_masked[5440] = data_i[5440] & sel_one_hot_i[42];
  assign data_masked[5439] = data_i[5439] & sel_one_hot_i[42];
  assign data_masked[5438] = data_i[5438] & sel_one_hot_i[42];
  assign data_masked[5437] = data_i[5437] & sel_one_hot_i[42];
  assign data_masked[5436] = data_i[5436] & sel_one_hot_i[42];
  assign data_masked[5435] = data_i[5435] & sel_one_hot_i[42];
  assign data_masked[5434] = data_i[5434] & sel_one_hot_i[42];
  assign data_masked[5433] = data_i[5433] & sel_one_hot_i[42];
  assign data_masked[5432] = data_i[5432] & sel_one_hot_i[42];
  assign data_masked[5431] = data_i[5431] & sel_one_hot_i[42];
  assign data_masked[5430] = data_i[5430] & sel_one_hot_i[42];
  assign data_masked[5429] = data_i[5429] & sel_one_hot_i[42];
  assign data_masked[5428] = data_i[5428] & sel_one_hot_i[42];
  assign data_masked[5427] = data_i[5427] & sel_one_hot_i[42];
  assign data_masked[5426] = data_i[5426] & sel_one_hot_i[42];
  assign data_masked[5425] = data_i[5425] & sel_one_hot_i[42];
  assign data_masked[5424] = data_i[5424] & sel_one_hot_i[42];
  assign data_masked[5423] = data_i[5423] & sel_one_hot_i[42];
  assign data_masked[5422] = data_i[5422] & sel_one_hot_i[42];
  assign data_masked[5421] = data_i[5421] & sel_one_hot_i[42];
  assign data_masked[5420] = data_i[5420] & sel_one_hot_i[42];
  assign data_masked[5419] = data_i[5419] & sel_one_hot_i[42];
  assign data_masked[5418] = data_i[5418] & sel_one_hot_i[42];
  assign data_masked[5417] = data_i[5417] & sel_one_hot_i[42];
  assign data_masked[5416] = data_i[5416] & sel_one_hot_i[42];
  assign data_masked[5415] = data_i[5415] & sel_one_hot_i[42];
  assign data_masked[5414] = data_i[5414] & sel_one_hot_i[42];
  assign data_masked[5413] = data_i[5413] & sel_one_hot_i[42];
  assign data_masked[5412] = data_i[5412] & sel_one_hot_i[42];
  assign data_masked[5411] = data_i[5411] & sel_one_hot_i[42];
  assign data_masked[5410] = data_i[5410] & sel_one_hot_i[42];
  assign data_masked[5409] = data_i[5409] & sel_one_hot_i[42];
  assign data_masked[5408] = data_i[5408] & sel_one_hot_i[42];
  assign data_masked[5407] = data_i[5407] & sel_one_hot_i[42];
  assign data_masked[5406] = data_i[5406] & sel_one_hot_i[42];
  assign data_masked[5405] = data_i[5405] & sel_one_hot_i[42];
  assign data_masked[5404] = data_i[5404] & sel_one_hot_i[42];
  assign data_masked[5403] = data_i[5403] & sel_one_hot_i[42];
  assign data_masked[5402] = data_i[5402] & sel_one_hot_i[42];
  assign data_masked[5401] = data_i[5401] & sel_one_hot_i[42];
  assign data_masked[5400] = data_i[5400] & sel_one_hot_i[42];
  assign data_masked[5399] = data_i[5399] & sel_one_hot_i[42];
  assign data_masked[5398] = data_i[5398] & sel_one_hot_i[42];
  assign data_masked[5397] = data_i[5397] & sel_one_hot_i[42];
  assign data_masked[5396] = data_i[5396] & sel_one_hot_i[42];
  assign data_masked[5395] = data_i[5395] & sel_one_hot_i[42];
  assign data_masked[5394] = data_i[5394] & sel_one_hot_i[42];
  assign data_masked[5393] = data_i[5393] & sel_one_hot_i[42];
  assign data_masked[5392] = data_i[5392] & sel_one_hot_i[42];
  assign data_masked[5391] = data_i[5391] & sel_one_hot_i[42];
  assign data_masked[5390] = data_i[5390] & sel_one_hot_i[42];
  assign data_masked[5389] = data_i[5389] & sel_one_hot_i[42];
  assign data_masked[5388] = data_i[5388] & sel_one_hot_i[42];
  assign data_masked[5387] = data_i[5387] & sel_one_hot_i[42];
  assign data_masked[5386] = data_i[5386] & sel_one_hot_i[42];
  assign data_masked[5385] = data_i[5385] & sel_one_hot_i[42];
  assign data_masked[5384] = data_i[5384] & sel_one_hot_i[42];
  assign data_masked[5383] = data_i[5383] & sel_one_hot_i[42];
  assign data_masked[5382] = data_i[5382] & sel_one_hot_i[42];
  assign data_masked[5381] = data_i[5381] & sel_one_hot_i[42];
  assign data_masked[5380] = data_i[5380] & sel_one_hot_i[42];
  assign data_masked[5379] = data_i[5379] & sel_one_hot_i[42];
  assign data_masked[5378] = data_i[5378] & sel_one_hot_i[42];
  assign data_masked[5377] = data_i[5377] & sel_one_hot_i[42];
  assign data_masked[5376] = data_i[5376] & sel_one_hot_i[42];
  assign data_masked[5631] = data_i[5631] & sel_one_hot_i[43];
  assign data_masked[5630] = data_i[5630] & sel_one_hot_i[43];
  assign data_masked[5629] = data_i[5629] & sel_one_hot_i[43];
  assign data_masked[5628] = data_i[5628] & sel_one_hot_i[43];
  assign data_masked[5627] = data_i[5627] & sel_one_hot_i[43];
  assign data_masked[5626] = data_i[5626] & sel_one_hot_i[43];
  assign data_masked[5625] = data_i[5625] & sel_one_hot_i[43];
  assign data_masked[5624] = data_i[5624] & sel_one_hot_i[43];
  assign data_masked[5623] = data_i[5623] & sel_one_hot_i[43];
  assign data_masked[5622] = data_i[5622] & sel_one_hot_i[43];
  assign data_masked[5621] = data_i[5621] & sel_one_hot_i[43];
  assign data_masked[5620] = data_i[5620] & sel_one_hot_i[43];
  assign data_masked[5619] = data_i[5619] & sel_one_hot_i[43];
  assign data_masked[5618] = data_i[5618] & sel_one_hot_i[43];
  assign data_masked[5617] = data_i[5617] & sel_one_hot_i[43];
  assign data_masked[5616] = data_i[5616] & sel_one_hot_i[43];
  assign data_masked[5615] = data_i[5615] & sel_one_hot_i[43];
  assign data_masked[5614] = data_i[5614] & sel_one_hot_i[43];
  assign data_masked[5613] = data_i[5613] & sel_one_hot_i[43];
  assign data_masked[5612] = data_i[5612] & sel_one_hot_i[43];
  assign data_masked[5611] = data_i[5611] & sel_one_hot_i[43];
  assign data_masked[5610] = data_i[5610] & sel_one_hot_i[43];
  assign data_masked[5609] = data_i[5609] & sel_one_hot_i[43];
  assign data_masked[5608] = data_i[5608] & sel_one_hot_i[43];
  assign data_masked[5607] = data_i[5607] & sel_one_hot_i[43];
  assign data_masked[5606] = data_i[5606] & sel_one_hot_i[43];
  assign data_masked[5605] = data_i[5605] & sel_one_hot_i[43];
  assign data_masked[5604] = data_i[5604] & sel_one_hot_i[43];
  assign data_masked[5603] = data_i[5603] & sel_one_hot_i[43];
  assign data_masked[5602] = data_i[5602] & sel_one_hot_i[43];
  assign data_masked[5601] = data_i[5601] & sel_one_hot_i[43];
  assign data_masked[5600] = data_i[5600] & sel_one_hot_i[43];
  assign data_masked[5599] = data_i[5599] & sel_one_hot_i[43];
  assign data_masked[5598] = data_i[5598] & sel_one_hot_i[43];
  assign data_masked[5597] = data_i[5597] & sel_one_hot_i[43];
  assign data_masked[5596] = data_i[5596] & sel_one_hot_i[43];
  assign data_masked[5595] = data_i[5595] & sel_one_hot_i[43];
  assign data_masked[5594] = data_i[5594] & sel_one_hot_i[43];
  assign data_masked[5593] = data_i[5593] & sel_one_hot_i[43];
  assign data_masked[5592] = data_i[5592] & sel_one_hot_i[43];
  assign data_masked[5591] = data_i[5591] & sel_one_hot_i[43];
  assign data_masked[5590] = data_i[5590] & sel_one_hot_i[43];
  assign data_masked[5589] = data_i[5589] & sel_one_hot_i[43];
  assign data_masked[5588] = data_i[5588] & sel_one_hot_i[43];
  assign data_masked[5587] = data_i[5587] & sel_one_hot_i[43];
  assign data_masked[5586] = data_i[5586] & sel_one_hot_i[43];
  assign data_masked[5585] = data_i[5585] & sel_one_hot_i[43];
  assign data_masked[5584] = data_i[5584] & sel_one_hot_i[43];
  assign data_masked[5583] = data_i[5583] & sel_one_hot_i[43];
  assign data_masked[5582] = data_i[5582] & sel_one_hot_i[43];
  assign data_masked[5581] = data_i[5581] & sel_one_hot_i[43];
  assign data_masked[5580] = data_i[5580] & sel_one_hot_i[43];
  assign data_masked[5579] = data_i[5579] & sel_one_hot_i[43];
  assign data_masked[5578] = data_i[5578] & sel_one_hot_i[43];
  assign data_masked[5577] = data_i[5577] & sel_one_hot_i[43];
  assign data_masked[5576] = data_i[5576] & sel_one_hot_i[43];
  assign data_masked[5575] = data_i[5575] & sel_one_hot_i[43];
  assign data_masked[5574] = data_i[5574] & sel_one_hot_i[43];
  assign data_masked[5573] = data_i[5573] & sel_one_hot_i[43];
  assign data_masked[5572] = data_i[5572] & sel_one_hot_i[43];
  assign data_masked[5571] = data_i[5571] & sel_one_hot_i[43];
  assign data_masked[5570] = data_i[5570] & sel_one_hot_i[43];
  assign data_masked[5569] = data_i[5569] & sel_one_hot_i[43];
  assign data_masked[5568] = data_i[5568] & sel_one_hot_i[43];
  assign data_masked[5567] = data_i[5567] & sel_one_hot_i[43];
  assign data_masked[5566] = data_i[5566] & sel_one_hot_i[43];
  assign data_masked[5565] = data_i[5565] & sel_one_hot_i[43];
  assign data_masked[5564] = data_i[5564] & sel_one_hot_i[43];
  assign data_masked[5563] = data_i[5563] & sel_one_hot_i[43];
  assign data_masked[5562] = data_i[5562] & sel_one_hot_i[43];
  assign data_masked[5561] = data_i[5561] & sel_one_hot_i[43];
  assign data_masked[5560] = data_i[5560] & sel_one_hot_i[43];
  assign data_masked[5559] = data_i[5559] & sel_one_hot_i[43];
  assign data_masked[5558] = data_i[5558] & sel_one_hot_i[43];
  assign data_masked[5557] = data_i[5557] & sel_one_hot_i[43];
  assign data_masked[5556] = data_i[5556] & sel_one_hot_i[43];
  assign data_masked[5555] = data_i[5555] & sel_one_hot_i[43];
  assign data_masked[5554] = data_i[5554] & sel_one_hot_i[43];
  assign data_masked[5553] = data_i[5553] & sel_one_hot_i[43];
  assign data_masked[5552] = data_i[5552] & sel_one_hot_i[43];
  assign data_masked[5551] = data_i[5551] & sel_one_hot_i[43];
  assign data_masked[5550] = data_i[5550] & sel_one_hot_i[43];
  assign data_masked[5549] = data_i[5549] & sel_one_hot_i[43];
  assign data_masked[5548] = data_i[5548] & sel_one_hot_i[43];
  assign data_masked[5547] = data_i[5547] & sel_one_hot_i[43];
  assign data_masked[5546] = data_i[5546] & sel_one_hot_i[43];
  assign data_masked[5545] = data_i[5545] & sel_one_hot_i[43];
  assign data_masked[5544] = data_i[5544] & sel_one_hot_i[43];
  assign data_masked[5543] = data_i[5543] & sel_one_hot_i[43];
  assign data_masked[5542] = data_i[5542] & sel_one_hot_i[43];
  assign data_masked[5541] = data_i[5541] & sel_one_hot_i[43];
  assign data_masked[5540] = data_i[5540] & sel_one_hot_i[43];
  assign data_masked[5539] = data_i[5539] & sel_one_hot_i[43];
  assign data_masked[5538] = data_i[5538] & sel_one_hot_i[43];
  assign data_masked[5537] = data_i[5537] & sel_one_hot_i[43];
  assign data_masked[5536] = data_i[5536] & sel_one_hot_i[43];
  assign data_masked[5535] = data_i[5535] & sel_one_hot_i[43];
  assign data_masked[5534] = data_i[5534] & sel_one_hot_i[43];
  assign data_masked[5533] = data_i[5533] & sel_one_hot_i[43];
  assign data_masked[5532] = data_i[5532] & sel_one_hot_i[43];
  assign data_masked[5531] = data_i[5531] & sel_one_hot_i[43];
  assign data_masked[5530] = data_i[5530] & sel_one_hot_i[43];
  assign data_masked[5529] = data_i[5529] & sel_one_hot_i[43];
  assign data_masked[5528] = data_i[5528] & sel_one_hot_i[43];
  assign data_masked[5527] = data_i[5527] & sel_one_hot_i[43];
  assign data_masked[5526] = data_i[5526] & sel_one_hot_i[43];
  assign data_masked[5525] = data_i[5525] & sel_one_hot_i[43];
  assign data_masked[5524] = data_i[5524] & sel_one_hot_i[43];
  assign data_masked[5523] = data_i[5523] & sel_one_hot_i[43];
  assign data_masked[5522] = data_i[5522] & sel_one_hot_i[43];
  assign data_masked[5521] = data_i[5521] & sel_one_hot_i[43];
  assign data_masked[5520] = data_i[5520] & sel_one_hot_i[43];
  assign data_masked[5519] = data_i[5519] & sel_one_hot_i[43];
  assign data_masked[5518] = data_i[5518] & sel_one_hot_i[43];
  assign data_masked[5517] = data_i[5517] & sel_one_hot_i[43];
  assign data_masked[5516] = data_i[5516] & sel_one_hot_i[43];
  assign data_masked[5515] = data_i[5515] & sel_one_hot_i[43];
  assign data_masked[5514] = data_i[5514] & sel_one_hot_i[43];
  assign data_masked[5513] = data_i[5513] & sel_one_hot_i[43];
  assign data_masked[5512] = data_i[5512] & sel_one_hot_i[43];
  assign data_masked[5511] = data_i[5511] & sel_one_hot_i[43];
  assign data_masked[5510] = data_i[5510] & sel_one_hot_i[43];
  assign data_masked[5509] = data_i[5509] & sel_one_hot_i[43];
  assign data_masked[5508] = data_i[5508] & sel_one_hot_i[43];
  assign data_masked[5507] = data_i[5507] & sel_one_hot_i[43];
  assign data_masked[5506] = data_i[5506] & sel_one_hot_i[43];
  assign data_masked[5505] = data_i[5505] & sel_one_hot_i[43];
  assign data_masked[5504] = data_i[5504] & sel_one_hot_i[43];
  assign data_masked[5759] = data_i[5759] & sel_one_hot_i[44];
  assign data_masked[5758] = data_i[5758] & sel_one_hot_i[44];
  assign data_masked[5757] = data_i[5757] & sel_one_hot_i[44];
  assign data_masked[5756] = data_i[5756] & sel_one_hot_i[44];
  assign data_masked[5755] = data_i[5755] & sel_one_hot_i[44];
  assign data_masked[5754] = data_i[5754] & sel_one_hot_i[44];
  assign data_masked[5753] = data_i[5753] & sel_one_hot_i[44];
  assign data_masked[5752] = data_i[5752] & sel_one_hot_i[44];
  assign data_masked[5751] = data_i[5751] & sel_one_hot_i[44];
  assign data_masked[5750] = data_i[5750] & sel_one_hot_i[44];
  assign data_masked[5749] = data_i[5749] & sel_one_hot_i[44];
  assign data_masked[5748] = data_i[5748] & sel_one_hot_i[44];
  assign data_masked[5747] = data_i[5747] & sel_one_hot_i[44];
  assign data_masked[5746] = data_i[5746] & sel_one_hot_i[44];
  assign data_masked[5745] = data_i[5745] & sel_one_hot_i[44];
  assign data_masked[5744] = data_i[5744] & sel_one_hot_i[44];
  assign data_masked[5743] = data_i[5743] & sel_one_hot_i[44];
  assign data_masked[5742] = data_i[5742] & sel_one_hot_i[44];
  assign data_masked[5741] = data_i[5741] & sel_one_hot_i[44];
  assign data_masked[5740] = data_i[5740] & sel_one_hot_i[44];
  assign data_masked[5739] = data_i[5739] & sel_one_hot_i[44];
  assign data_masked[5738] = data_i[5738] & sel_one_hot_i[44];
  assign data_masked[5737] = data_i[5737] & sel_one_hot_i[44];
  assign data_masked[5736] = data_i[5736] & sel_one_hot_i[44];
  assign data_masked[5735] = data_i[5735] & sel_one_hot_i[44];
  assign data_masked[5734] = data_i[5734] & sel_one_hot_i[44];
  assign data_masked[5733] = data_i[5733] & sel_one_hot_i[44];
  assign data_masked[5732] = data_i[5732] & sel_one_hot_i[44];
  assign data_masked[5731] = data_i[5731] & sel_one_hot_i[44];
  assign data_masked[5730] = data_i[5730] & sel_one_hot_i[44];
  assign data_masked[5729] = data_i[5729] & sel_one_hot_i[44];
  assign data_masked[5728] = data_i[5728] & sel_one_hot_i[44];
  assign data_masked[5727] = data_i[5727] & sel_one_hot_i[44];
  assign data_masked[5726] = data_i[5726] & sel_one_hot_i[44];
  assign data_masked[5725] = data_i[5725] & sel_one_hot_i[44];
  assign data_masked[5724] = data_i[5724] & sel_one_hot_i[44];
  assign data_masked[5723] = data_i[5723] & sel_one_hot_i[44];
  assign data_masked[5722] = data_i[5722] & sel_one_hot_i[44];
  assign data_masked[5721] = data_i[5721] & sel_one_hot_i[44];
  assign data_masked[5720] = data_i[5720] & sel_one_hot_i[44];
  assign data_masked[5719] = data_i[5719] & sel_one_hot_i[44];
  assign data_masked[5718] = data_i[5718] & sel_one_hot_i[44];
  assign data_masked[5717] = data_i[5717] & sel_one_hot_i[44];
  assign data_masked[5716] = data_i[5716] & sel_one_hot_i[44];
  assign data_masked[5715] = data_i[5715] & sel_one_hot_i[44];
  assign data_masked[5714] = data_i[5714] & sel_one_hot_i[44];
  assign data_masked[5713] = data_i[5713] & sel_one_hot_i[44];
  assign data_masked[5712] = data_i[5712] & sel_one_hot_i[44];
  assign data_masked[5711] = data_i[5711] & sel_one_hot_i[44];
  assign data_masked[5710] = data_i[5710] & sel_one_hot_i[44];
  assign data_masked[5709] = data_i[5709] & sel_one_hot_i[44];
  assign data_masked[5708] = data_i[5708] & sel_one_hot_i[44];
  assign data_masked[5707] = data_i[5707] & sel_one_hot_i[44];
  assign data_masked[5706] = data_i[5706] & sel_one_hot_i[44];
  assign data_masked[5705] = data_i[5705] & sel_one_hot_i[44];
  assign data_masked[5704] = data_i[5704] & sel_one_hot_i[44];
  assign data_masked[5703] = data_i[5703] & sel_one_hot_i[44];
  assign data_masked[5702] = data_i[5702] & sel_one_hot_i[44];
  assign data_masked[5701] = data_i[5701] & sel_one_hot_i[44];
  assign data_masked[5700] = data_i[5700] & sel_one_hot_i[44];
  assign data_masked[5699] = data_i[5699] & sel_one_hot_i[44];
  assign data_masked[5698] = data_i[5698] & sel_one_hot_i[44];
  assign data_masked[5697] = data_i[5697] & sel_one_hot_i[44];
  assign data_masked[5696] = data_i[5696] & sel_one_hot_i[44];
  assign data_masked[5695] = data_i[5695] & sel_one_hot_i[44];
  assign data_masked[5694] = data_i[5694] & sel_one_hot_i[44];
  assign data_masked[5693] = data_i[5693] & sel_one_hot_i[44];
  assign data_masked[5692] = data_i[5692] & sel_one_hot_i[44];
  assign data_masked[5691] = data_i[5691] & sel_one_hot_i[44];
  assign data_masked[5690] = data_i[5690] & sel_one_hot_i[44];
  assign data_masked[5689] = data_i[5689] & sel_one_hot_i[44];
  assign data_masked[5688] = data_i[5688] & sel_one_hot_i[44];
  assign data_masked[5687] = data_i[5687] & sel_one_hot_i[44];
  assign data_masked[5686] = data_i[5686] & sel_one_hot_i[44];
  assign data_masked[5685] = data_i[5685] & sel_one_hot_i[44];
  assign data_masked[5684] = data_i[5684] & sel_one_hot_i[44];
  assign data_masked[5683] = data_i[5683] & sel_one_hot_i[44];
  assign data_masked[5682] = data_i[5682] & sel_one_hot_i[44];
  assign data_masked[5681] = data_i[5681] & sel_one_hot_i[44];
  assign data_masked[5680] = data_i[5680] & sel_one_hot_i[44];
  assign data_masked[5679] = data_i[5679] & sel_one_hot_i[44];
  assign data_masked[5678] = data_i[5678] & sel_one_hot_i[44];
  assign data_masked[5677] = data_i[5677] & sel_one_hot_i[44];
  assign data_masked[5676] = data_i[5676] & sel_one_hot_i[44];
  assign data_masked[5675] = data_i[5675] & sel_one_hot_i[44];
  assign data_masked[5674] = data_i[5674] & sel_one_hot_i[44];
  assign data_masked[5673] = data_i[5673] & sel_one_hot_i[44];
  assign data_masked[5672] = data_i[5672] & sel_one_hot_i[44];
  assign data_masked[5671] = data_i[5671] & sel_one_hot_i[44];
  assign data_masked[5670] = data_i[5670] & sel_one_hot_i[44];
  assign data_masked[5669] = data_i[5669] & sel_one_hot_i[44];
  assign data_masked[5668] = data_i[5668] & sel_one_hot_i[44];
  assign data_masked[5667] = data_i[5667] & sel_one_hot_i[44];
  assign data_masked[5666] = data_i[5666] & sel_one_hot_i[44];
  assign data_masked[5665] = data_i[5665] & sel_one_hot_i[44];
  assign data_masked[5664] = data_i[5664] & sel_one_hot_i[44];
  assign data_masked[5663] = data_i[5663] & sel_one_hot_i[44];
  assign data_masked[5662] = data_i[5662] & sel_one_hot_i[44];
  assign data_masked[5661] = data_i[5661] & sel_one_hot_i[44];
  assign data_masked[5660] = data_i[5660] & sel_one_hot_i[44];
  assign data_masked[5659] = data_i[5659] & sel_one_hot_i[44];
  assign data_masked[5658] = data_i[5658] & sel_one_hot_i[44];
  assign data_masked[5657] = data_i[5657] & sel_one_hot_i[44];
  assign data_masked[5656] = data_i[5656] & sel_one_hot_i[44];
  assign data_masked[5655] = data_i[5655] & sel_one_hot_i[44];
  assign data_masked[5654] = data_i[5654] & sel_one_hot_i[44];
  assign data_masked[5653] = data_i[5653] & sel_one_hot_i[44];
  assign data_masked[5652] = data_i[5652] & sel_one_hot_i[44];
  assign data_masked[5651] = data_i[5651] & sel_one_hot_i[44];
  assign data_masked[5650] = data_i[5650] & sel_one_hot_i[44];
  assign data_masked[5649] = data_i[5649] & sel_one_hot_i[44];
  assign data_masked[5648] = data_i[5648] & sel_one_hot_i[44];
  assign data_masked[5647] = data_i[5647] & sel_one_hot_i[44];
  assign data_masked[5646] = data_i[5646] & sel_one_hot_i[44];
  assign data_masked[5645] = data_i[5645] & sel_one_hot_i[44];
  assign data_masked[5644] = data_i[5644] & sel_one_hot_i[44];
  assign data_masked[5643] = data_i[5643] & sel_one_hot_i[44];
  assign data_masked[5642] = data_i[5642] & sel_one_hot_i[44];
  assign data_masked[5641] = data_i[5641] & sel_one_hot_i[44];
  assign data_masked[5640] = data_i[5640] & sel_one_hot_i[44];
  assign data_masked[5639] = data_i[5639] & sel_one_hot_i[44];
  assign data_masked[5638] = data_i[5638] & sel_one_hot_i[44];
  assign data_masked[5637] = data_i[5637] & sel_one_hot_i[44];
  assign data_masked[5636] = data_i[5636] & sel_one_hot_i[44];
  assign data_masked[5635] = data_i[5635] & sel_one_hot_i[44];
  assign data_masked[5634] = data_i[5634] & sel_one_hot_i[44];
  assign data_masked[5633] = data_i[5633] & sel_one_hot_i[44];
  assign data_masked[5632] = data_i[5632] & sel_one_hot_i[44];
  assign data_masked[5887] = data_i[5887] & sel_one_hot_i[45];
  assign data_masked[5886] = data_i[5886] & sel_one_hot_i[45];
  assign data_masked[5885] = data_i[5885] & sel_one_hot_i[45];
  assign data_masked[5884] = data_i[5884] & sel_one_hot_i[45];
  assign data_masked[5883] = data_i[5883] & sel_one_hot_i[45];
  assign data_masked[5882] = data_i[5882] & sel_one_hot_i[45];
  assign data_masked[5881] = data_i[5881] & sel_one_hot_i[45];
  assign data_masked[5880] = data_i[5880] & sel_one_hot_i[45];
  assign data_masked[5879] = data_i[5879] & sel_one_hot_i[45];
  assign data_masked[5878] = data_i[5878] & sel_one_hot_i[45];
  assign data_masked[5877] = data_i[5877] & sel_one_hot_i[45];
  assign data_masked[5876] = data_i[5876] & sel_one_hot_i[45];
  assign data_masked[5875] = data_i[5875] & sel_one_hot_i[45];
  assign data_masked[5874] = data_i[5874] & sel_one_hot_i[45];
  assign data_masked[5873] = data_i[5873] & sel_one_hot_i[45];
  assign data_masked[5872] = data_i[5872] & sel_one_hot_i[45];
  assign data_masked[5871] = data_i[5871] & sel_one_hot_i[45];
  assign data_masked[5870] = data_i[5870] & sel_one_hot_i[45];
  assign data_masked[5869] = data_i[5869] & sel_one_hot_i[45];
  assign data_masked[5868] = data_i[5868] & sel_one_hot_i[45];
  assign data_masked[5867] = data_i[5867] & sel_one_hot_i[45];
  assign data_masked[5866] = data_i[5866] & sel_one_hot_i[45];
  assign data_masked[5865] = data_i[5865] & sel_one_hot_i[45];
  assign data_masked[5864] = data_i[5864] & sel_one_hot_i[45];
  assign data_masked[5863] = data_i[5863] & sel_one_hot_i[45];
  assign data_masked[5862] = data_i[5862] & sel_one_hot_i[45];
  assign data_masked[5861] = data_i[5861] & sel_one_hot_i[45];
  assign data_masked[5860] = data_i[5860] & sel_one_hot_i[45];
  assign data_masked[5859] = data_i[5859] & sel_one_hot_i[45];
  assign data_masked[5858] = data_i[5858] & sel_one_hot_i[45];
  assign data_masked[5857] = data_i[5857] & sel_one_hot_i[45];
  assign data_masked[5856] = data_i[5856] & sel_one_hot_i[45];
  assign data_masked[5855] = data_i[5855] & sel_one_hot_i[45];
  assign data_masked[5854] = data_i[5854] & sel_one_hot_i[45];
  assign data_masked[5853] = data_i[5853] & sel_one_hot_i[45];
  assign data_masked[5852] = data_i[5852] & sel_one_hot_i[45];
  assign data_masked[5851] = data_i[5851] & sel_one_hot_i[45];
  assign data_masked[5850] = data_i[5850] & sel_one_hot_i[45];
  assign data_masked[5849] = data_i[5849] & sel_one_hot_i[45];
  assign data_masked[5848] = data_i[5848] & sel_one_hot_i[45];
  assign data_masked[5847] = data_i[5847] & sel_one_hot_i[45];
  assign data_masked[5846] = data_i[5846] & sel_one_hot_i[45];
  assign data_masked[5845] = data_i[5845] & sel_one_hot_i[45];
  assign data_masked[5844] = data_i[5844] & sel_one_hot_i[45];
  assign data_masked[5843] = data_i[5843] & sel_one_hot_i[45];
  assign data_masked[5842] = data_i[5842] & sel_one_hot_i[45];
  assign data_masked[5841] = data_i[5841] & sel_one_hot_i[45];
  assign data_masked[5840] = data_i[5840] & sel_one_hot_i[45];
  assign data_masked[5839] = data_i[5839] & sel_one_hot_i[45];
  assign data_masked[5838] = data_i[5838] & sel_one_hot_i[45];
  assign data_masked[5837] = data_i[5837] & sel_one_hot_i[45];
  assign data_masked[5836] = data_i[5836] & sel_one_hot_i[45];
  assign data_masked[5835] = data_i[5835] & sel_one_hot_i[45];
  assign data_masked[5834] = data_i[5834] & sel_one_hot_i[45];
  assign data_masked[5833] = data_i[5833] & sel_one_hot_i[45];
  assign data_masked[5832] = data_i[5832] & sel_one_hot_i[45];
  assign data_masked[5831] = data_i[5831] & sel_one_hot_i[45];
  assign data_masked[5830] = data_i[5830] & sel_one_hot_i[45];
  assign data_masked[5829] = data_i[5829] & sel_one_hot_i[45];
  assign data_masked[5828] = data_i[5828] & sel_one_hot_i[45];
  assign data_masked[5827] = data_i[5827] & sel_one_hot_i[45];
  assign data_masked[5826] = data_i[5826] & sel_one_hot_i[45];
  assign data_masked[5825] = data_i[5825] & sel_one_hot_i[45];
  assign data_masked[5824] = data_i[5824] & sel_one_hot_i[45];
  assign data_masked[5823] = data_i[5823] & sel_one_hot_i[45];
  assign data_masked[5822] = data_i[5822] & sel_one_hot_i[45];
  assign data_masked[5821] = data_i[5821] & sel_one_hot_i[45];
  assign data_masked[5820] = data_i[5820] & sel_one_hot_i[45];
  assign data_masked[5819] = data_i[5819] & sel_one_hot_i[45];
  assign data_masked[5818] = data_i[5818] & sel_one_hot_i[45];
  assign data_masked[5817] = data_i[5817] & sel_one_hot_i[45];
  assign data_masked[5816] = data_i[5816] & sel_one_hot_i[45];
  assign data_masked[5815] = data_i[5815] & sel_one_hot_i[45];
  assign data_masked[5814] = data_i[5814] & sel_one_hot_i[45];
  assign data_masked[5813] = data_i[5813] & sel_one_hot_i[45];
  assign data_masked[5812] = data_i[5812] & sel_one_hot_i[45];
  assign data_masked[5811] = data_i[5811] & sel_one_hot_i[45];
  assign data_masked[5810] = data_i[5810] & sel_one_hot_i[45];
  assign data_masked[5809] = data_i[5809] & sel_one_hot_i[45];
  assign data_masked[5808] = data_i[5808] & sel_one_hot_i[45];
  assign data_masked[5807] = data_i[5807] & sel_one_hot_i[45];
  assign data_masked[5806] = data_i[5806] & sel_one_hot_i[45];
  assign data_masked[5805] = data_i[5805] & sel_one_hot_i[45];
  assign data_masked[5804] = data_i[5804] & sel_one_hot_i[45];
  assign data_masked[5803] = data_i[5803] & sel_one_hot_i[45];
  assign data_masked[5802] = data_i[5802] & sel_one_hot_i[45];
  assign data_masked[5801] = data_i[5801] & sel_one_hot_i[45];
  assign data_masked[5800] = data_i[5800] & sel_one_hot_i[45];
  assign data_masked[5799] = data_i[5799] & sel_one_hot_i[45];
  assign data_masked[5798] = data_i[5798] & sel_one_hot_i[45];
  assign data_masked[5797] = data_i[5797] & sel_one_hot_i[45];
  assign data_masked[5796] = data_i[5796] & sel_one_hot_i[45];
  assign data_masked[5795] = data_i[5795] & sel_one_hot_i[45];
  assign data_masked[5794] = data_i[5794] & sel_one_hot_i[45];
  assign data_masked[5793] = data_i[5793] & sel_one_hot_i[45];
  assign data_masked[5792] = data_i[5792] & sel_one_hot_i[45];
  assign data_masked[5791] = data_i[5791] & sel_one_hot_i[45];
  assign data_masked[5790] = data_i[5790] & sel_one_hot_i[45];
  assign data_masked[5789] = data_i[5789] & sel_one_hot_i[45];
  assign data_masked[5788] = data_i[5788] & sel_one_hot_i[45];
  assign data_masked[5787] = data_i[5787] & sel_one_hot_i[45];
  assign data_masked[5786] = data_i[5786] & sel_one_hot_i[45];
  assign data_masked[5785] = data_i[5785] & sel_one_hot_i[45];
  assign data_masked[5784] = data_i[5784] & sel_one_hot_i[45];
  assign data_masked[5783] = data_i[5783] & sel_one_hot_i[45];
  assign data_masked[5782] = data_i[5782] & sel_one_hot_i[45];
  assign data_masked[5781] = data_i[5781] & sel_one_hot_i[45];
  assign data_masked[5780] = data_i[5780] & sel_one_hot_i[45];
  assign data_masked[5779] = data_i[5779] & sel_one_hot_i[45];
  assign data_masked[5778] = data_i[5778] & sel_one_hot_i[45];
  assign data_masked[5777] = data_i[5777] & sel_one_hot_i[45];
  assign data_masked[5776] = data_i[5776] & sel_one_hot_i[45];
  assign data_masked[5775] = data_i[5775] & sel_one_hot_i[45];
  assign data_masked[5774] = data_i[5774] & sel_one_hot_i[45];
  assign data_masked[5773] = data_i[5773] & sel_one_hot_i[45];
  assign data_masked[5772] = data_i[5772] & sel_one_hot_i[45];
  assign data_masked[5771] = data_i[5771] & sel_one_hot_i[45];
  assign data_masked[5770] = data_i[5770] & sel_one_hot_i[45];
  assign data_masked[5769] = data_i[5769] & sel_one_hot_i[45];
  assign data_masked[5768] = data_i[5768] & sel_one_hot_i[45];
  assign data_masked[5767] = data_i[5767] & sel_one_hot_i[45];
  assign data_masked[5766] = data_i[5766] & sel_one_hot_i[45];
  assign data_masked[5765] = data_i[5765] & sel_one_hot_i[45];
  assign data_masked[5764] = data_i[5764] & sel_one_hot_i[45];
  assign data_masked[5763] = data_i[5763] & sel_one_hot_i[45];
  assign data_masked[5762] = data_i[5762] & sel_one_hot_i[45];
  assign data_masked[5761] = data_i[5761] & sel_one_hot_i[45];
  assign data_masked[5760] = data_i[5760] & sel_one_hot_i[45];
  assign data_masked[6015] = data_i[6015] & sel_one_hot_i[46];
  assign data_masked[6014] = data_i[6014] & sel_one_hot_i[46];
  assign data_masked[6013] = data_i[6013] & sel_one_hot_i[46];
  assign data_masked[6012] = data_i[6012] & sel_one_hot_i[46];
  assign data_masked[6011] = data_i[6011] & sel_one_hot_i[46];
  assign data_masked[6010] = data_i[6010] & sel_one_hot_i[46];
  assign data_masked[6009] = data_i[6009] & sel_one_hot_i[46];
  assign data_masked[6008] = data_i[6008] & sel_one_hot_i[46];
  assign data_masked[6007] = data_i[6007] & sel_one_hot_i[46];
  assign data_masked[6006] = data_i[6006] & sel_one_hot_i[46];
  assign data_masked[6005] = data_i[6005] & sel_one_hot_i[46];
  assign data_masked[6004] = data_i[6004] & sel_one_hot_i[46];
  assign data_masked[6003] = data_i[6003] & sel_one_hot_i[46];
  assign data_masked[6002] = data_i[6002] & sel_one_hot_i[46];
  assign data_masked[6001] = data_i[6001] & sel_one_hot_i[46];
  assign data_masked[6000] = data_i[6000] & sel_one_hot_i[46];
  assign data_masked[5999] = data_i[5999] & sel_one_hot_i[46];
  assign data_masked[5998] = data_i[5998] & sel_one_hot_i[46];
  assign data_masked[5997] = data_i[5997] & sel_one_hot_i[46];
  assign data_masked[5996] = data_i[5996] & sel_one_hot_i[46];
  assign data_masked[5995] = data_i[5995] & sel_one_hot_i[46];
  assign data_masked[5994] = data_i[5994] & sel_one_hot_i[46];
  assign data_masked[5993] = data_i[5993] & sel_one_hot_i[46];
  assign data_masked[5992] = data_i[5992] & sel_one_hot_i[46];
  assign data_masked[5991] = data_i[5991] & sel_one_hot_i[46];
  assign data_masked[5990] = data_i[5990] & sel_one_hot_i[46];
  assign data_masked[5989] = data_i[5989] & sel_one_hot_i[46];
  assign data_masked[5988] = data_i[5988] & sel_one_hot_i[46];
  assign data_masked[5987] = data_i[5987] & sel_one_hot_i[46];
  assign data_masked[5986] = data_i[5986] & sel_one_hot_i[46];
  assign data_masked[5985] = data_i[5985] & sel_one_hot_i[46];
  assign data_masked[5984] = data_i[5984] & sel_one_hot_i[46];
  assign data_masked[5983] = data_i[5983] & sel_one_hot_i[46];
  assign data_masked[5982] = data_i[5982] & sel_one_hot_i[46];
  assign data_masked[5981] = data_i[5981] & sel_one_hot_i[46];
  assign data_masked[5980] = data_i[5980] & sel_one_hot_i[46];
  assign data_masked[5979] = data_i[5979] & sel_one_hot_i[46];
  assign data_masked[5978] = data_i[5978] & sel_one_hot_i[46];
  assign data_masked[5977] = data_i[5977] & sel_one_hot_i[46];
  assign data_masked[5976] = data_i[5976] & sel_one_hot_i[46];
  assign data_masked[5975] = data_i[5975] & sel_one_hot_i[46];
  assign data_masked[5974] = data_i[5974] & sel_one_hot_i[46];
  assign data_masked[5973] = data_i[5973] & sel_one_hot_i[46];
  assign data_masked[5972] = data_i[5972] & sel_one_hot_i[46];
  assign data_masked[5971] = data_i[5971] & sel_one_hot_i[46];
  assign data_masked[5970] = data_i[5970] & sel_one_hot_i[46];
  assign data_masked[5969] = data_i[5969] & sel_one_hot_i[46];
  assign data_masked[5968] = data_i[5968] & sel_one_hot_i[46];
  assign data_masked[5967] = data_i[5967] & sel_one_hot_i[46];
  assign data_masked[5966] = data_i[5966] & sel_one_hot_i[46];
  assign data_masked[5965] = data_i[5965] & sel_one_hot_i[46];
  assign data_masked[5964] = data_i[5964] & sel_one_hot_i[46];
  assign data_masked[5963] = data_i[5963] & sel_one_hot_i[46];
  assign data_masked[5962] = data_i[5962] & sel_one_hot_i[46];
  assign data_masked[5961] = data_i[5961] & sel_one_hot_i[46];
  assign data_masked[5960] = data_i[5960] & sel_one_hot_i[46];
  assign data_masked[5959] = data_i[5959] & sel_one_hot_i[46];
  assign data_masked[5958] = data_i[5958] & sel_one_hot_i[46];
  assign data_masked[5957] = data_i[5957] & sel_one_hot_i[46];
  assign data_masked[5956] = data_i[5956] & sel_one_hot_i[46];
  assign data_masked[5955] = data_i[5955] & sel_one_hot_i[46];
  assign data_masked[5954] = data_i[5954] & sel_one_hot_i[46];
  assign data_masked[5953] = data_i[5953] & sel_one_hot_i[46];
  assign data_masked[5952] = data_i[5952] & sel_one_hot_i[46];
  assign data_masked[5951] = data_i[5951] & sel_one_hot_i[46];
  assign data_masked[5950] = data_i[5950] & sel_one_hot_i[46];
  assign data_masked[5949] = data_i[5949] & sel_one_hot_i[46];
  assign data_masked[5948] = data_i[5948] & sel_one_hot_i[46];
  assign data_masked[5947] = data_i[5947] & sel_one_hot_i[46];
  assign data_masked[5946] = data_i[5946] & sel_one_hot_i[46];
  assign data_masked[5945] = data_i[5945] & sel_one_hot_i[46];
  assign data_masked[5944] = data_i[5944] & sel_one_hot_i[46];
  assign data_masked[5943] = data_i[5943] & sel_one_hot_i[46];
  assign data_masked[5942] = data_i[5942] & sel_one_hot_i[46];
  assign data_masked[5941] = data_i[5941] & sel_one_hot_i[46];
  assign data_masked[5940] = data_i[5940] & sel_one_hot_i[46];
  assign data_masked[5939] = data_i[5939] & sel_one_hot_i[46];
  assign data_masked[5938] = data_i[5938] & sel_one_hot_i[46];
  assign data_masked[5937] = data_i[5937] & sel_one_hot_i[46];
  assign data_masked[5936] = data_i[5936] & sel_one_hot_i[46];
  assign data_masked[5935] = data_i[5935] & sel_one_hot_i[46];
  assign data_masked[5934] = data_i[5934] & sel_one_hot_i[46];
  assign data_masked[5933] = data_i[5933] & sel_one_hot_i[46];
  assign data_masked[5932] = data_i[5932] & sel_one_hot_i[46];
  assign data_masked[5931] = data_i[5931] & sel_one_hot_i[46];
  assign data_masked[5930] = data_i[5930] & sel_one_hot_i[46];
  assign data_masked[5929] = data_i[5929] & sel_one_hot_i[46];
  assign data_masked[5928] = data_i[5928] & sel_one_hot_i[46];
  assign data_masked[5927] = data_i[5927] & sel_one_hot_i[46];
  assign data_masked[5926] = data_i[5926] & sel_one_hot_i[46];
  assign data_masked[5925] = data_i[5925] & sel_one_hot_i[46];
  assign data_masked[5924] = data_i[5924] & sel_one_hot_i[46];
  assign data_masked[5923] = data_i[5923] & sel_one_hot_i[46];
  assign data_masked[5922] = data_i[5922] & sel_one_hot_i[46];
  assign data_masked[5921] = data_i[5921] & sel_one_hot_i[46];
  assign data_masked[5920] = data_i[5920] & sel_one_hot_i[46];
  assign data_masked[5919] = data_i[5919] & sel_one_hot_i[46];
  assign data_masked[5918] = data_i[5918] & sel_one_hot_i[46];
  assign data_masked[5917] = data_i[5917] & sel_one_hot_i[46];
  assign data_masked[5916] = data_i[5916] & sel_one_hot_i[46];
  assign data_masked[5915] = data_i[5915] & sel_one_hot_i[46];
  assign data_masked[5914] = data_i[5914] & sel_one_hot_i[46];
  assign data_masked[5913] = data_i[5913] & sel_one_hot_i[46];
  assign data_masked[5912] = data_i[5912] & sel_one_hot_i[46];
  assign data_masked[5911] = data_i[5911] & sel_one_hot_i[46];
  assign data_masked[5910] = data_i[5910] & sel_one_hot_i[46];
  assign data_masked[5909] = data_i[5909] & sel_one_hot_i[46];
  assign data_masked[5908] = data_i[5908] & sel_one_hot_i[46];
  assign data_masked[5907] = data_i[5907] & sel_one_hot_i[46];
  assign data_masked[5906] = data_i[5906] & sel_one_hot_i[46];
  assign data_masked[5905] = data_i[5905] & sel_one_hot_i[46];
  assign data_masked[5904] = data_i[5904] & sel_one_hot_i[46];
  assign data_masked[5903] = data_i[5903] & sel_one_hot_i[46];
  assign data_masked[5902] = data_i[5902] & sel_one_hot_i[46];
  assign data_masked[5901] = data_i[5901] & sel_one_hot_i[46];
  assign data_masked[5900] = data_i[5900] & sel_one_hot_i[46];
  assign data_masked[5899] = data_i[5899] & sel_one_hot_i[46];
  assign data_masked[5898] = data_i[5898] & sel_one_hot_i[46];
  assign data_masked[5897] = data_i[5897] & sel_one_hot_i[46];
  assign data_masked[5896] = data_i[5896] & sel_one_hot_i[46];
  assign data_masked[5895] = data_i[5895] & sel_one_hot_i[46];
  assign data_masked[5894] = data_i[5894] & sel_one_hot_i[46];
  assign data_masked[5893] = data_i[5893] & sel_one_hot_i[46];
  assign data_masked[5892] = data_i[5892] & sel_one_hot_i[46];
  assign data_masked[5891] = data_i[5891] & sel_one_hot_i[46];
  assign data_masked[5890] = data_i[5890] & sel_one_hot_i[46];
  assign data_masked[5889] = data_i[5889] & sel_one_hot_i[46];
  assign data_masked[5888] = data_i[5888] & sel_one_hot_i[46];
  assign data_masked[6143] = data_i[6143] & sel_one_hot_i[47];
  assign data_masked[6142] = data_i[6142] & sel_one_hot_i[47];
  assign data_masked[6141] = data_i[6141] & sel_one_hot_i[47];
  assign data_masked[6140] = data_i[6140] & sel_one_hot_i[47];
  assign data_masked[6139] = data_i[6139] & sel_one_hot_i[47];
  assign data_masked[6138] = data_i[6138] & sel_one_hot_i[47];
  assign data_masked[6137] = data_i[6137] & sel_one_hot_i[47];
  assign data_masked[6136] = data_i[6136] & sel_one_hot_i[47];
  assign data_masked[6135] = data_i[6135] & sel_one_hot_i[47];
  assign data_masked[6134] = data_i[6134] & sel_one_hot_i[47];
  assign data_masked[6133] = data_i[6133] & sel_one_hot_i[47];
  assign data_masked[6132] = data_i[6132] & sel_one_hot_i[47];
  assign data_masked[6131] = data_i[6131] & sel_one_hot_i[47];
  assign data_masked[6130] = data_i[6130] & sel_one_hot_i[47];
  assign data_masked[6129] = data_i[6129] & sel_one_hot_i[47];
  assign data_masked[6128] = data_i[6128] & sel_one_hot_i[47];
  assign data_masked[6127] = data_i[6127] & sel_one_hot_i[47];
  assign data_masked[6126] = data_i[6126] & sel_one_hot_i[47];
  assign data_masked[6125] = data_i[6125] & sel_one_hot_i[47];
  assign data_masked[6124] = data_i[6124] & sel_one_hot_i[47];
  assign data_masked[6123] = data_i[6123] & sel_one_hot_i[47];
  assign data_masked[6122] = data_i[6122] & sel_one_hot_i[47];
  assign data_masked[6121] = data_i[6121] & sel_one_hot_i[47];
  assign data_masked[6120] = data_i[6120] & sel_one_hot_i[47];
  assign data_masked[6119] = data_i[6119] & sel_one_hot_i[47];
  assign data_masked[6118] = data_i[6118] & sel_one_hot_i[47];
  assign data_masked[6117] = data_i[6117] & sel_one_hot_i[47];
  assign data_masked[6116] = data_i[6116] & sel_one_hot_i[47];
  assign data_masked[6115] = data_i[6115] & sel_one_hot_i[47];
  assign data_masked[6114] = data_i[6114] & sel_one_hot_i[47];
  assign data_masked[6113] = data_i[6113] & sel_one_hot_i[47];
  assign data_masked[6112] = data_i[6112] & sel_one_hot_i[47];
  assign data_masked[6111] = data_i[6111] & sel_one_hot_i[47];
  assign data_masked[6110] = data_i[6110] & sel_one_hot_i[47];
  assign data_masked[6109] = data_i[6109] & sel_one_hot_i[47];
  assign data_masked[6108] = data_i[6108] & sel_one_hot_i[47];
  assign data_masked[6107] = data_i[6107] & sel_one_hot_i[47];
  assign data_masked[6106] = data_i[6106] & sel_one_hot_i[47];
  assign data_masked[6105] = data_i[6105] & sel_one_hot_i[47];
  assign data_masked[6104] = data_i[6104] & sel_one_hot_i[47];
  assign data_masked[6103] = data_i[6103] & sel_one_hot_i[47];
  assign data_masked[6102] = data_i[6102] & sel_one_hot_i[47];
  assign data_masked[6101] = data_i[6101] & sel_one_hot_i[47];
  assign data_masked[6100] = data_i[6100] & sel_one_hot_i[47];
  assign data_masked[6099] = data_i[6099] & sel_one_hot_i[47];
  assign data_masked[6098] = data_i[6098] & sel_one_hot_i[47];
  assign data_masked[6097] = data_i[6097] & sel_one_hot_i[47];
  assign data_masked[6096] = data_i[6096] & sel_one_hot_i[47];
  assign data_masked[6095] = data_i[6095] & sel_one_hot_i[47];
  assign data_masked[6094] = data_i[6094] & sel_one_hot_i[47];
  assign data_masked[6093] = data_i[6093] & sel_one_hot_i[47];
  assign data_masked[6092] = data_i[6092] & sel_one_hot_i[47];
  assign data_masked[6091] = data_i[6091] & sel_one_hot_i[47];
  assign data_masked[6090] = data_i[6090] & sel_one_hot_i[47];
  assign data_masked[6089] = data_i[6089] & sel_one_hot_i[47];
  assign data_masked[6088] = data_i[6088] & sel_one_hot_i[47];
  assign data_masked[6087] = data_i[6087] & sel_one_hot_i[47];
  assign data_masked[6086] = data_i[6086] & sel_one_hot_i[47];
  assign data_masked[6085] = data_i[6085] & sel_one_hot_i[47];
  assign data_masked[6084] = data_i[6084] & sel_one_hot_i[47];
  assign data_masked[6083] = data_i[6083] & sel_one_hot_i[47];
  assign data_masked[6082] = data_i[6082] & sel_one_hot_i[47];
  assign data_masked[6081] = data_i[6081] & sel_one_hot_i[47];
  assign data_masked[6080] = data_i[6080] & sel_one_hot_i[47];
  assign data_masked[6079] = data_i[6079] & sel_one_hot_i[47];
  assign data_masked[6078] = data_i[6078] & sel_one_hot_i[47];
  assign data_masked[6077] = data_i[6077] & sel_one_hot_i[47];
  assign data_masked[6076] = data_i[6076] & sel_one_hot_i[47];
  assign data_masked[6075] = data_i[6075] & sel_one_hot_i[47];
  assign data_masked[6074] = data_i[6074] & sel_one_hot_i[47];
  assign data_masked[6073] = data_i[6073] & sel_one_hot_i[47];
  assign data_masked[6072] = data_i[6072] & sel_one_hot_i[47];
  assign data_masked[6071] = data_i[6071] & sel_one_hot_i[47];
  assign data_masked[6070] = data_i[6070] & sel_one_hot_i[47];
  assign data_masked[6069] = data_i[6069] & sel_one_hot_i[47];
  assign data_masked[6068] = data_i[6068] & sel_one_hot_i[47];
  assign data_masked[6067] = data_i[6067] & sel_one_hot_i[47];
  assign data_masked[6066] = data_i[6066] & sel_one_hot_i[47];
  assign data_masked[6065] = data_i[6065] & sel_one_hot_i[47];
  assign data_masked[6064] = data_i[6064] & sel_one_hot_i[47];
  assign data_masked[6063] = data_i[6063] & sel_one_hot_i[47];
  assign data_masked[6062] = data_i[6062] & sel_one_hot_i[47];
  assign data_masked[6061] = data_i[6061] & sel_one_hot_i[47];
  assign data_masked[6060] = data_i[6060] & sel_one_hot_i[47];
  assign data_masked[6059] = data_i[6059] & sel_one_hot_i[47];
  assign data_masked[6058] = data_i[6058] & sel_one_hot_i[47];
  assign data_masked[6057] = data_i[6057] & sel_one_hot_i[47];
  assign data_masked[6056] = data_i[6056] & sel_one_hot_i[47];
  assign data_masked[6055] = data_i[6055] & sel_one_hot_i[47];
  assign data_masked[6054] = data_i[6054] & sel_one_hot_i[47];
  assign data_masked[6053] = data_i[6053] & sel_one_hot_i[47];
  assign data_masked[6052] = data_i[6052] & sel_one_hot_i[47];
  assign data_masked[6051] = data_i[6051] & sel_one_hot_i[47];
  assign data_masked[6050] = data_i[6050] & sel_one_hot_i[47];
  assign data_masked[6049] = data_i[6049] & sel_one_hot_i[47];
  assign data_masked[6048] = data_i[6048] & sel_one_hot_i[47];
  assign data_masked[6047] = data_i[6047] & sel_one_hot_i[47];
  assign data_masked[6046] = data_i[6046] & sel_one_hot_i[47];
  assign data_masked[6045] = data_i[6045] & sel_one_hot_i[47];
  assign data_masked[6044] = data_i[6044] & sel_one_hot_i[47];
  assign data_masked[6043] = data_i[6043] & sel_one_hot_i[47];
  assign data_masked[6042] = data_i[6042] & sel_one_hot_i[47];
  assign data_masked[6041] = data_i[6041] & sel_one_hot_i[47];
  assign data_masked[6040] = data_i[6040] & sel_one_hot_i[47];
  assign data_masked[6039] = data_i[6039] & sel_one_hot_i[47];
  assign data_masked[6038] = data_i[6038] & sel_one_hot_i[47];
  assign data_masked[6037] = data_i[6037] & sel_one_hot_i[47];
  assign data_masked[6036] = data_i[6036] & sel_one_hot_i[47];
  assign data_masked[6035] = data_i[6035] & sel_one_hot_i[47];
  assign data_masked[6034] = data_i[6034] & sel_one_hot_i[47];
  assign data_masked[6033] = data_i[6033] & sel_one_hot_i[47];
  assign data_masked[6032] = data_i[6032] & sel_one_hot_i[47];
  assign data_masked[6031] = data_i[6031] & sel_one_hot_i[47];
  assign data_masked[6030] = data_i[6030] & sel_one_hot_i[47];
  assign data_masked[6029] = data_i[6029] & sel_one_hot_i[47];
  assign data_masked[6028] = data_i[6028] & sel_one_hot_i[47];
  assign data_masked[6027] = data_i[6027] & sel_one_hot_i[47];
  assign data_masked[6026] = data_i[6026] & sel_one_hot_i[47];
  assign data_masked[6025] = data_i[6025] & sel_one_hot_i[47];
  assign data_masked[6024] = data_i[6024] & sel_one_hot_i[47];
  assign data_masked[6023] = data_i[6023] & sel_one_hot_i[47];
  assign data_masked[6022] = data_i[6022] & sel_one_hot_i[47];
  assign data_masked[6021] = data_i[6021] & sel_one_hot_i[47];
  assign data_masked[6020] = data_i[6020] & sel_one_hot_i[47];
  assign data_masked[6019] = data_i[6019] & sel_one_hot_i[47];
  assign data_masked[6018] = data_i[6018] & sel_one_hot_i[47];
  assign data_masked[6017] = data_i[6017] & sel_one_hot_i[47];
  assign data_masked[6016] = data_i[6016] & sel_one_hot_i[47];
  assign data_masked[6271] = data_i[6271] & sel_one_hot_i[48];
  assign data_masked[6270] = data_i[6270] & sel_one_hot_i[48];
  assign data_masked[6269] = data_i[6269] & sel_one_hot_i[48];
  assign data_masked[6268] = data_i[6268] & sel_one_hot_i[48];
  assign data_masked[6267] = data_i[6267] & sel_one_hot_i[48];
  assign data_masked[6266] = data_i[6266] & sel_one_hot_i[48];
  assign data_masked[6265] = data_i[6265] & sel_one_hot_i[48];
  assign data_masked[6264] = data_i[6264] & sel_one_hot_i[48];
  assign data_masked[6263] = data_i[6263] & sel_one_hot_i[48];
  assign data_masked[6262] = data_i[6262] & sel_one_hot_i[48];
  assign data_masked[6261] = data_i[6261] & sel_one_hot_i[48];
  assign data_masked[6260] = data_i[6260] & sel_one_hot_i[48];
  assign data_masked[6259] = data_i[6259] & sel_one_hot_i[48];
  assign data_masked[6258] = data_i[6258] & sel_one_hot_i[48];
  assign data_masked[6257] = data_i[6257] & sel_one_hot_i[48];
  assign data_masked[6256] = data_i[6256] & sel_one_hot_i[48];
  assign data_masked[6255] = data_i[6255] & sel_one_hot_i[48];
  assign data_masked[6254] = data_i[6254] & sel_one_hot_i[48];
  assign data_masked[6253] = data_i[6253] & sel_one_hot_i[48];
  assign data_masked[6252] = data_i[6252] & sel_one_hot_i[48];
  assign data_masked[6251] = data_i[6251] & sel_one_hot_i[48];
  assign data_masked[6250] = data_i[6250] & sel_one_hot_i[48];
  assign data_masked[6249] = data_i[6249] & sel_one_hot_i[48];
  assign data_masked[6248] = data_i[6248] & sel_one_hot_i[48];
  assign data_masked[6247] = data_i[6247] & sel_one_hot_i[48];
  assign data_masked[6246] = data_i[6246] & sel_one_hot_i[48];
  assign data_masked[6245] = data_i[6245] & sel_one_hot_i[48];
  assign data_masked[6244] = data_i[6244] & sel_one_hot_i[48];
  assign data_masked[6243] = data_i[6243] & sel_one_hot_i[48];
  assign data_masked[6242] = data_i[6242] & sel_one_hot_i[48];
  assign data_masked[6241] = data_i[6241] & sel_one_hot_i[48];
  assign data_masked[6240] = data_i[6240] & sel_one_hot_i[48];
  assign data_masked[6239] = data_i[6239] & sel_one_hot_i[48];
  assign data_masked[6238] = data_i[6238] & sel_one_hot_i[48];
  assign data_masked[6237] = data_i[6237] & sel_one_hot_i[48];
  assign data_masked[6236] = data_i[6236] & sel_one_hot_i[48];
  assign data_masked[6235] = data_i[6235] & sel_one_hot_i[48];
  assign data_masked[6234] = data_i[6234] & sel_one_hot_i[48];
  assign data_masked[6233] = data_i[6233] & sel_one_hot_i[48];
  assign data_masked[6232] = data_i[6232] & sel_one_hot_i[48];
  assign data_masked[6231] = data_i[6231] & sel_one_hot_i[48];
  assign data_masked[6230] = data_i[6230] & sel_one_hot_i[48];
  assign data_masked[6229] = data_i[6229] & sel_one_hot_i[48];
  assign data_masked[6228] = data_i[6228] & sel_one_hot_i[48];
  assign data_masked[6227] = data_i[6227] & sel_one_hot_i[48];
  assign data_masked[6226] = data_i[6226] & sel_one_hot_i[48];
  assign data_masked[6225] = data_i[6225] & sel_one_hot_i[48];
  assign data_masked[6224] = data_i[6224] & sel_one_hot_i[48];
  assign data_masked[6223] = data_i[6223] & sel_one_hot_i[48];
  assign data_masked[6222] = data_i[6222] & sel_one_hot_i[48];
  assign data_masked[6221] = data_i[6221] & sel_one_hot_i[48];
  assign data_masked[6220] = data_i[6220] & sel_one_hot_i[48];
  assign data_masked[6219] = data_i[6219] & sel_one_hot_i[48];
  assign data_masked[6218] = data_i[6218] & sel_one_hot_i[48];
  assign data_masked[6217] = data_i[6217] & sel_one_hot_i[48];
  assign data_masked[6216] = data_i[6216] & sel_one_hot_i[48];
  assign data_masked[6215] = data_i[6215] & sel_one_hot_i[48];
  assign data_masked[6214] = data_i[6214] & sel_one_hot_i[48];
  assign data_masked[6213] = data_i[6213] & sel_one_hot_i[48];
  assign data_masked[6212] = data_i[6212] & sel_one_hot_i[48];
  assign data_masked[6211] = data_i[6211] & sel_one_hot_i[48];
  assign data_masked[6210] = data_i[6210] & sel_one_hot_i[48];
  assign data_masked[6209] = data_i[6209] & sel_one_hot_i[48];
  assign data_masked[6208] = data_i[6208] & sel_one_hot_i[48];
  assign data_masked[6207] = data_i[6207] & sel_one_hot_i[48];
  assign data_masked[6206] = data_i[6206] & sel_one_hot_i[48];
  assign data_masked[6205] = data_i[6205] & sel_one_hot_i[48];
  assign data_masked[6204] = data_i[6204] & sel_one_hot_i[48];
  assign data_masked[6203] = data_i[6203] & sel_one_hot_i[48];
  assign data_masked[6202] = data_i[6202] & sel_one_hot_i[48];
  assign data_masked[6201] = data_i[6201] & sel_one_hot_i[48];
  assign data_masked[6200] = data_i[6200] & sel_one_hot_i[48];
  assign data_masked[6199] = data_i[6199] & sel_one_hot_i[48];
  assign data_masked[6198] = data_i[6198] & sel_one_hot_i[48];
  assign data_masked[6197] = data_i[6197] & sel_one_hot_i[48];
  assign data_masked[6196] = data_i[6196] & sel_one_hot_i[48];
  assign data_masked[6195] = data_i[6195] & sel_one_hot_i[48];
  assign data_masked[6194] = data_i[6194] & sel_one_hot_i[48];
  assign data_masked[6193] = data_i[6193] & sel_one_hot_i[48];
  assign data_masked[6192] = data_i[6192] & sel_one_hot_i[48];
  assign data_masked[6191] = data_i[6191] & sel_one_hot_i[48];
  assign data_masked[6190] = data_i[6190] & sel_one_hot_i[48];
  assign data_masked[6189] = data_i[6189] & sel_one_hot_i[48];
  assign data_masked[6188] = data_i[6188] & sel_one_hot_i[48];
  assign data_masked[6187] = data_i[6187] & sel_one_hot_i[48];
  assign data_masked[6186] = data_i[6186] & sel_one_hot_i[48];
  assign data_masked[6185] = data_i[6185] & sel_one_hot_i[48];
  assign data_masked[6184] = data_i[6184] & sel_one_hot_i[48];
  assign data_masked[6183] = data_i[6183] & sel_one_hot_i[48];
  assign data_masked[6182] = data_i[6182] & sel_one_hot_i[48];
  assign data_masked[6181] = data_i[6181] & sel_one_hot_i[48];
  assign data_masked[6180] = data_i[6180] & sel_one_hot_i[48];
  assign data_masked[6179] = data_i[6179] & sel_one_hot_i[48];
  assign data_masked[6178] = data_i[6178] & sel_one_hot_i[48];
  assign data_masked[6177] = data_i[6177] & sel_one_hot_i[48];
  assign data_masked[6176] = data_i[6176] & sel_one_hot_i[48];
  assign data_masked[6175] = data_i[6175] & sel_one_hot_i[48];
  assign data_masked[6174] = data_i[6174] & sel_one_hot_i[48];
  assign data_masked[6173] = data_i[6173] & sel_one_hot_i[48];
  assign data_masked[6172] = data_i[6172] & sel_one_hot_i[48];
  assign data_masked[6171] = data_i[6171] & sel_one_hot_i[48];
  assign data_masked[6170] = data_i[6170] & sel_one_hot_i[48];
  assign data_masked[6169] = data_i[6169] & sel_one_hot_i[48];
  assign data_masked[6168] = data_i[6168] & sel_one_hot_i[48];
  assign data_masked[6167] = data_i[6167] & sel_one_hot_i[48];
  assign data_masked[6166] = data_i[6166] & sel_one_hot_i[48];
  assign data_masked[6165] = data_i[6165] & sel_one_hot_i[48];
  assign data_masked[6164] = data_i[6164] & sel_one_hot_i[48];
  assign data_masked[6163] = data_i[6163] & sel_one_hot_i[48];
  assign data_masked[6162] = data_i[6162] & sel_one_hot_i[48];
  assign data_masked[6161] = data_i[6161] & sel_one_hot_i[48];
  assign data_masked[6160] = data_i[6160] & sel_one_hot_i[48];
  assign data_masked[6159] = data_i[6159] & sel_one_hot_i[48];
  assign data_masked[6158] = data_i[6158] & sel_one_hot_i[48];
  assign data_masked[6157] = data_i[6157] & sel_one_hot_i[48];
  assign data_masked[6156] = data_i[6156] & sel_one_hot_i[48];
  assign data_masked[6155] = data_i[6155] & sel_one_hot_i[48];
  assign data_masked[6154] = data_i[6154] & sel_one_hot_i[48];
  assign data_masked[6153] = data_i[6153] & sel_one_hot_i[48];
  assign data_masked[6152] = data_i[6152] & sel_one_hot_i[48];
  assign data_masked[6151] = data_i[6151] & sel_one_hot_i[48];
  assign data_masked[6150] = data_i[6150] & sel_one_hot_i[48];
  assign data_masked[6149] = data_i[6149] & sel_one_hot_i[48];
  assign data_masked[6148] = data_i[6148] & sel_one_hot_i[48];
  assign data_masked[6147] = data_i[6147] & sel_one_hot_i[48];
  assign data_masked[6146] = data_i[6146] & sel_one_hot_i[48];
  assign data_masked[6145] = data_i[6145] & sel_one_hot_i[48];
  assign data_masked[6144] = data_i[6144] & sel_one_hot_i[48];
  assign data_masked[6399] = data_i[6399] & sel_one_hot_i[49];
  assign data_masked[6398] = data_i[6398] & sel_one_hot_i[49];
  assign data_masked[6397] = data_i[6397] & sel_one_hot_i[49];
  assign data_masked[6396] = data_i[6396] & sel_one_hot_i[49];
  assign data_masked[6395] = data_i[6395] & sel_one_hot_i[49];
  assign data_masked[6394] = data_i[6394] & sel_one_hot_i[49];
  assign data_masked[6393] = data_i[6393] & sel_one_hot_i[49];
  assign data_masked[6392] = data_i[6392] & sel_one_hot_i[49];
  assign data_masked[6391] = data_i[6391] & sel_one_hot_i[49];
  assign data_masked[6390] = data_i[6390] & sel_one_hot_i[49];
  assign data_masked[6389] = data_i[6389] & sel_one_hot_i[49];
  assign data_masked[6388] = data_i[6388] & sel_one_hot_i[49];
  assign data_masked[6387] = data_i[6387] & sel_one_hot_i[49];
  assign data_masked[6386] = data_i[6386] & sel_one_hot_i[49];
  assign data_masked[6385] = data_i[6385] & sel_one_hot_i[49];
  assign data_masked[6384] = data_i[6384] & sel_one_hot_i[49];
  assign data_masked[6383] = data_i[6383] & sel_one_hot_i[49];
  assign data_masked[6382] = data_i[6382] & sel_one_hot_i[49];
  assign data_masked[6381] = data_i[6381] & sel_one_hot_i[49];
  assign data_masked[6380] = data_i[6380] & sel_one_hot_i[49];
  assign data_masked[6379] = data_i[6379] & sel_one_hot_i[49];
  assign data_masked[6378] = data_i[6378] & sel_one_hot_i[49];
  assign data_masked[6377] = data_i[6377] & sel_one_hot_i[49];
  assign data_masked[6376] = data_i[6376] & sel_one_hot_i[49];
  assign data_masked[6375] = data_i[6375] & sel_one_hot_i[49];
  assign data_masked[6374] = data_i[6374] & sel_one_hot_i[49];
  assign data_masked[6373] = data_i[6373] & sel_one_hot_i[49];
  assign data_masked[6372] = data_i[6372] & sel_one_hot_i[49];
  assign data_masked[6371] = data_i[6371] & sel_one_hot_i[49];
  assign data_masked[6370] = data_i[6370] & sel_one_hot_i[49];
  assign data_masked[6369] = data_i[6369] & sel_one_hot_i[49];
  assign data_masked[6368] = data_i[6368] & sel_one_hot_i[49];
  assign data_masked[6367] = data_i[6367] & sel_one_hot_i[49];
  assign data_masked[6366] = data_i[6366] & sel_one_hot_i[49];
  assign data_masked[6365] = data_i[6365] & sel_one_hot_i[49];
  assign data_masked[6364] = data_i[6364] & sel_one_hot_i[49];
  assign data_masked[6363] = data_i[6363] & sel_one_hot_i[49];
  assign data_masked[6362] = data_i[6362] & sel_one_hot_i[49];
  assign data_masked[6361] = data_i[6361] & sel_one_hot_i[49];
  assign data_masked[6360] = data_i[6360] & sel_one_hot_i[49];
  assign data_masked[6359] = data_i[6359] & sel_one_hot_i[49];
  assign data_masked[6358] = data_i[6358] & sel_one_hot_i[49];
  assign data_masked[6357] = data_i[6357] & sel_one_hot_i[49];
  assign data_masked[6356] = data_i[6356] & sel_one_hot_i[49];
  assign data_masked[6355] = data_i[6355] & sel_one_hot_i[49];
  assign data_masked[6354] = data_i[6354] & sel_one_hot_i[49];
  assign data_masked[6353] = data_i[6353] & sel_one_hot_i[49];
  assign data_masked[6352] = data_i[6352] & sel_one_hot_i[49];
  assign data_masked[6351] = data_i[6351] & sel_one_hot_i[49];
  assign data_masked[6350] = data_i[6350] & sel_one_hot_i[49];
  assign data_masked[6349] = data_i[6349] & sel_one_hot_i[49];
  assign data_masked[6348] = data_i[6348] & sel_one_hot_i[49];
  assign data_masked[6347] = data_i[6347] & sel_one_hot_i[49];
  assign data_masked[6346] = data_i[6346] & sel_one_hot_i[49];
  assign data_masked[6345] = data_i[6345] & sel_one_hot_i[49];
  assign data_masked[6344] = data_i[6344] & sel_one_hot_i[49];
  assign data_masked[6343] = data_i[6343] & sel_one_hot_i[49];
  assign data_masked[6342] = data_i[6342] & sel_one_hot_i[49];
  assign data_masked[6341] = data_i[6341] & sel_one_hot_i[49];
  assign data_masked[6340] = data_i[6340] & sel_one_hot_i[49];
  assign data_masked[6339] = data_i[6339] & sel_one_hot_i[49];
  assign data_masked[6338] = data_i[6338] & sel_one_hot_i[49];
  assign data_masked[6337] = data_i[6337] & sel_one_hot_i[49];
  assign data_masked[6336] = data_i[6336] & sel_one_hot_i[49];
  assign data_masked[6335] = data_i[6335] & sel_one_hot_i[49];
  assign data_masked[6334] = data_i[6334] & sel_one_hot_i[49];
  assign data_masked[6333] = data_i[6333] & sel_one_hot_i[49];
  assign data_masked[6332] = data_i[6332] & sel_one_hot_i[49];
  assign data_masked[6331] = data_i[6331] & sel_one_hot_i[49];
  assign data_masked[6330] = data_i[6330] & sel_one_hot_i[49];
  assign data_masked[6329] = data_i[6329] & sel_one_hot_i[49];
  assign data_masked[6328] = data_i[6328] & sel_one_hot_i[49];
  assign data_masked[6327] = data_i[6327] & sel_one_hot_i[49];
  assign data_masked[6326] = data_i[6326] & sel_one_hot_i[49];
  assign data_masked[6325] = data_i[6325] & sel_one_hot_i[49];
  assign data_masked[6324] = data_i[6324] & sel_one_hot_i[49];
  assign data_masked[6323] = data_i[6323] & sel_one_hot_i[49];
  assign data_masked[6322] = data_i[6322] & sel_one_hot_i[49];
  assign data_masked[6321] = data_i[6321] & sel_one_hot_i[49];
  assign data_masked[6320] = data_i[6320] & sel_one_hot_i[49];
  assign data_masked[6319] = data_i[6319] & sel_one_hot_i[49];
  assign data_masked[6318] = data_i[6318] & sel_one_hot_i[49];
  assign data_masked[6317] = data_i[6317] & sel_one_hot_i[49];
  assign data_masked[6316] = data_i[6316] & sel_one_hot_i[49];
  assign data_masked[6315] = data_i[6315] & sel_one_hot_i[49];
  assign data_masked[6314] = data_i[6314] & sel_one_hot_i[49];
  assign data_masked[6313] = data_i[6313] & sel_one_hot_i[49];
  assign data_masked[6312] = data_i[6312] & sel_one_hot_i[49];
  assign data_masked[6311] = data_i[6311] & sel_one_hot_i[49];
  assign data_masked[6310] = data_i[6310] & sel_one_hot_i[49];
  assign data_masked[6309] = data_i[6309] & sel_one_hot_i[49];
  assign data_masked[6308] = data_i[6308] & sel_one_hot_i[49];
  assign data_masked[6307] = data_i[6307] & sel_one_hot_i[49];
  assign data_masked[6306] = data_i[6306] & sel_one_hot_i[49];
  assign data_masked[6305] = data_i[6305] & sel_one_hot_i[49];
  assign data_masked[6304] = data_i[6304] & sel_one_hot_i[49];
  assign data_masked[6303] = data_i[6303] & sel_one_hot_i[49];
  assign data_masked[6302] = data_i[6302] & sel_one_hot_i[49];
  assign data_masked[6301] = data_i[6301] & sel_one_hot_i[49];
  assign data_masked[6300] = data_i[6300] & sel_one_hot_i[49];
  assign data_masked[6299] = data_i[6299] & sel_one_hot_i[49];
  assign data_masked[6298] = data_i[6298] & sel_one_hot_i[49];
  assign data_masked[6297] = data_i[6297] & sel_one_hot_i[49];
  assign data_masked[6296] = data_i[6296] & sel_one_hot_i[49];
  assign data_masked[6295] = data_i[6295] & sel_one_hot_i[49];
  assign data_masked[6294] = data_i[6294] & sel_one_hot_i[49];
  assign data_masked[6293] = data_i[6293] & sel_one_hot_i[49];
  assign data_masked[6292] = data_i[6292] & sel_one_hot_i[49];
  assign data_masked[6291] = data_i[6291] & sel_one_hot_i[49];
  assign data_masked[6290] = data_i[6290] & sel_one_hot_i[49];
  assign data_masked[6289] = data_i[6289] & sel_one_hot_i[49];
  assign data_masked[6288] = data_i[6288] & sel_one_hot_i[49];
  assign data_masked[6287] = data_i[6287] & sel_one_hot_i[49];
  assign data_masked[6286] = data_i[6286] & sel_one_hot_i[49];
  assign data_masked[6285] = data_i[6285] & sel_one_hot_i[49];
  assign data_masked[6284] = data_i[6284] & sel_one_hot_i[49];
  assign data_masked[6283] = data_i[6283] & sel_one_hot_i[49];
  assign data_masked[6282] = data_i[6282] & sel_one_hot_i[49];
  assign data_masked[6281] = data_i[6281] & sel_one_hot_i[49];
  assign data_masked[6280] = data_i[6280] & sel_one_hot_i[49];
  assign data_masked[6279] = data_i[6279] & sel_one_hot_i[49];
  assign data_masked[6278] = data_i[6278] & sel_one_hot_i[49];
  assign data_masked[6277] = data_i[6277] & sel_one_hot_i[49];
  assign data_masked[6276] = data_i[6276] & sel_one_hot_i[49];
  assign data_masked[6275] = data_i[6275] & sel_one_hot_i[49];
  assign data_masked[6274] = data_i[6274] & sel_one_hot_i[49];
  assign data_masked[6273] = data_i[6273] & sel_one_hot_i[49];
  assign data_masked[6272] = data_i[6272] & sel_one_hot_i[49];
  assign data_masked[6527] = data_i[6527] & sel_one_hot_i[50];
  assign data_masked[6526] = data_i[6526] & sel_one_hot_i[50];
  assign data_masked[6525] = data_i[6525] & sel_one_hot_i[50];
  assign data_masked[6524] = data_i[6524] & sel_one_hot_i[50];
  assign data_masked[6523] = data_i[6523] & sel_one_hot_i[50];
  assign data_masked[6522] = data_i[6522] & sel_one_hot_i[50];
  assign data_masked[6521] = data_i[6521] & sel_one_hot_i[50];
  assign data_masked[6520] = data_i[6520] & sel_one_hot_i[50];
  assign data_masked[6519] = data_i[6519] & sel_one_hot_i[50];
  assign data_masked[6518] = data_i[6518] & sel_one_hot_i[50];
  assign data_masked[6517] = data_i[6517] & sel_one_hot_i[50];
  assign data_masked[6516] = data_i[6516] & sel_one_hot_i[50];
  assign data_masked[6515] = data_i[6515] & sel_one_hot_i[50];
  assign data_masked[6514] = data_i[6514] & sel_one_hot_i[50];
  assign data_masked[6513] = data_i[6513] & sel_one_hot_i[50];
  assign data_masked[6512] = data_i[6512] & sel_one_hot_i[50];
  assign data_masked[6511] = data_i[6511] & sel_one_hot_i[50];
  assign data_masked[6510] = data_i[6510] & sel_one_hot_i[50];
  assign data_masked[6509] = data_i[6509] & sel_one_hot_i[50];
  assign data_masked[6508] = data_i[6508] & sel_one_hot_i[50];
  assign data_masked[6507] = data_i[6507] & sel_one_hot_i[50];
  assign data_masked[6506] = data_i[6506] & sel_one_hot_i[50];
  assign data_masked[6505] = data_i[6505] & sel_one_hot_i[50];
  assign data_masked[6504] = data_i[6504] & sel_one_hot_i[50];
  assign data_masked[6503] = data_i[6503] & sel_one_hot_i[50];
  assign data_masked[6502] = data_i[6502] & sel_one_hot_i[50];
  assign data_masked[6501] = data_i[6501] & sel_one_hot_i[50];
  assign data_masked[6500] = data_i[6500] & sel_one_hot_i[50];
  assign data_masked[6499] = data_i[6499] & sel_one_hot_i[50];
  assign data_masked[6498] = data_i[6498] & sel_one_hot_i[50];
  assign data_masked[6497] = data_i[6497] & sel_one_hot_i[50];
  assign data_masked[6496] = data_i[6496] & sel_one_hot_i[50];
  assign data_masked[6495] = data_i[6495] & sel_one_hot_i[50];
  assign data_masked[6494] = data_i[6494] & sel_one_hot_i[50];
  assign data_masked[6493] = data_i[6493] & sel_one_hot_i[50];
  assign data_masked[6492] = data_i[6492] & sel_one_hot_i[50];
  assign data_masked[6491] = data_i[6491] & sel_one_hot_i[50];
  assign data_masked[6490] = data_i[6490] & sel_one_hot_i[50];
  assign data_masked[6489] = data_i[6489] & sel_one_hot_i[50];
  assign data_masked[6488] = data_i[6488] & sel_one_hot_i[50];
  assign data_masked[6487] = data_i[6487] & sel_one_hot_i[50];
  assign data_masked[6486] = data_i[6486] & sel_one_hot_i[50];
  assign data_masked[6485] = data_i[6485] & sel_one_hot_i[50];
  assign data_masked[6484] = data_i[6484] & sel_one_hot_i[50];
  assign data_masked[6483] = data_i[6483] & sel_one_hot_i[50];
  assign data_masked[6482] = data_i[6482] & sel_one_hot_i[50];
  assign data_masked[6481] = data_i[6481] & sel_one_hot_i[50];
  assign data_masked[6480] = data_i[6480] & sel_one_hot_i[50];
  assign data_masked[6479] = data_i[6479] & sel_one_hot_i[50];
  assign data_masked[6478] = data_i[6478] & sel_one_hot_i[50];
  assign data_masked[6477] = data_i[6477] & sel_one_hot_i[50];
  assign data_masked[6476] = data_i[6476] & sel_one_hot_i[50];
  assign data_masked[6475] = data_i[6475] & sel_one_hot_i[50];
  assign data_masked[6474] = data_i[6474] & sel_one_hot_i[50];
  assign data_masked[6473] = data_i[6473] & sel_one_hot_i[50];
  assign data_masked[6472] = data_i[6472] & sel_one_hot_i[50];
  assign data_masked[6471] = data_i[6471] & sel_one_hot_i[50];
  assign data_masked[6470] = data_i[6470] & sel_one_hot_i[50];
  assign data_masked[6469] = data_i[6469] & sel_one_hot_i[50];
  assign data_masked[6468] = data_i[6468] & sel_one_hot_i[50];
  assign data_masked[6467] = data_i[6467] & sel_one_hot_i[50];
  assign data_masked[6466] = data_i[6466] & sel_one_hot_i[50];
  assign data_masked[6465] = data_i[6465] & sel_one_hot_i[50];
  assign data_masked[6464] = data_i[6464] & sel_one_hot_i[50];
  assign data_masked[6463] = data_i[6463] & sel_one_hot_i[50];
  assign data_masked[6462] = data_i[6462] & sel_one_hot_i[50];
  assign data_masked[6461] = data_i[6461] & sel_one_hot_i[50];
  assign data_masked[6460] = data_i[6460] & sel_one_hot_i[50];
  assign data_masked[6459] = data_i[6459] & sel_one_hot_i[50];
  assign data_masked[6458] = data_i[6458] & sel_one_hot_i[50];
  assign data_masked[6457] = data_i[6457] & sel_one_hot_i[50];
  assign data_masked[6456] = data_i[6456] & sel_one_hot_i[50];
  assign data_masked[6455] = data_i[6455] & sel_one_hot_i[50];
  assign data_masked[6454] = data_i[6454] & sel_one_hot_i[50];
  assign data_masked[6453] = data_i[6453] & sel_one_hot_i[50];
  assign data_masked[6452] = data_i[6452] & sel_one_hot_i[50];
  assign data_masked[6451] = data_i[6451] & sel_one_hot_i[50];
  assign data_masked[6450] = data_i[6450] & sel_one_hot_i[50];
  assign data_masked[6449] = data_i[6449] & sel_one_hot_i[50];
  assign data_masked[6448] = data_i[6448] & sel_one_hot_i[50];
  assign data_masked[6447] = data_i[6447] & sel_one_hot_i[50];
  assign data_masked[6446] = data_i[6446] & sel_one_hot_i[50];
  assign data_masked[6445] = data_i[6445] & sel_one_hot_i[50];
  assign data_masked[6444] = data_i[6444] & sel_one_hot_i[50];
  assign data_masked[6443] = data_i[6443] & sel_one_hot_i[50];
  assign data_masked[6442] = data_i[6442] & sel_one_hot_i[50];
  assign data_masked[6441] = data_i[6441] & sel_one_hot_i[50];
  assign data_masked[6440] = data_i[6440] & sel_one_hot_i[50];
  assign data_masked[6439] = data_i[6439] & sel_one_hot_i[50];
  assign data_masked[6438] = data_i[6438] & sel_one_hot_i[50];
  assign data_masked[6437] = data_i[6437] & sel_one_hot_i[50];
  assign data_masked[6436] = data_i[6436] & sel_one_hot_i[50];
  assign data_masked[6435] = data_i[6435] & sel_one_hot_i[50];
  assign data_masked[6434] = data_i[6434] & sel_one_hot_i[50];
  assign data_masked[6433] = data_i[6433] & sel_one_hot_i[50];
  assign data_masked[6432] = data_i[6432] & sel_one_hot_i[50];
  assign data_masked[6431] = data_i[6431] & sel_one_hot_i[50];
  assign data_masked[6430] = data_i[6430] & sel_one_hot_i[50];
  assign data_masked[6429] = data_i[6429] & sel_one_hot_i[50];
  assign data_masked[6428] = data_i[6428] & sel_one_hot_i[50];
  assign data_masked[6427] = data_i[6427] & sel_one_hot_i[50];
  assign data_masked[6426] = data_i[6426] & sel_one_hot_i[50];
  assign data_masked[6425] = data_i[6425] & sel_one_hot_i[50];
  assign data_masked[6424] = data_i[6424] & sel_one_hot_i[50];
  assign data_masked[6423] = data_i[6423] & sel_one_hot_i[50];
  assign data_masked[6422] = data_i[6422] & sel_one_hot_i[50];
  assign data_masked[6421] = data_i[6421] & sel_one_hot_i[50];
  assign data_masked[6420] = data_i[6420] & sel_one_hot_i[50];
  assign data_masked[6419] = data_i[6419] & sel_one_hot_i[50];
  assign data_masked[6418] = data_i[6418] & sel_one_hot_i[50];
  assign data_masked[6417] = data_i[6417] & sel_one_hot_i[50];
  assign data_masked[6416] = data_i[6416] & sel_one_hot_i[50];
  assign data_masked[6415] = data_i[6415] & sel_one_hot_i[50];
  assign data_masked[6414] = data_i[6414] & sel_one_hot_i[50];
  assign data_masked[6413] = data_i[6413] & sel_one_hot_i[50];
  assign data_masked[6412] = data_i[6412] & sel_one_hot_i[50];
  assign data_masked[6411] = data_i[6411] & sel_one_hot_i[50];
  assign data_masked[6410] = data_i[6410] & sel_one_hot_i[50];
  assign data_masked[6409] = data_i[6409] & sel_one_hot_i[50];
  assign data_masked[6408] = data_i[6408] & sel_one_hot_i[50];
  assign data_masked[6407] = data_i[6407] & sel_one_hot_i[50];
  assign data_masked[6406] = data_i[6406] & sel_one_hot_i[50];
  assign data_masked[6405] = data_i[6405] & sel_one_hot_i[50];
  assign data_masked[6404] = data_i[6404] & sel_one_hot_i[50];
  assign data_masked[6403] = data_i[6403] & sel_one_hot_i[50];
  assign data_masked[6402] = data_i[6402] & sel_one_hot_i[50];
  assign data_masked[6401] = data_i[6401] & sel_one_hot_i[50];
  assign data_masked[6400] = data_i[6400] & sel_one_hot_i[50];
  assign data_masked[6655] = data_i[6655] & sel_one_hot_i[51];
  assign data_masked[6654] = data_i[6654] & sel_one_hot_i[51];
  assign data_masked[6653] = data_i[6653] & sel_one_hot_i[51];
  assign data_masked[6652] = data_i[6652] & sel_one_hot_i[51];
  assign data_masked[6651] = data_i[6651] & sel_one_hot_i[51];
  assign data_masked[6650] = data_i[6650] & sel_one_hot_i[51];
  assign data_masked[6649] = data_i[6649] & sel_one_hot_i[51];
  assign data_masked[6648] = data_i[6648] & sel_one_hot_i[51];
  assign data_masked[6647] = data_i[6647] & sel_one_hot_i[51];
  assign data_masked[6646] = data_i[6646] & sel_one_hot_i[51];
  assign data_masked[6645] = data_i[6645] & sel_one_hot_i[51];
  assign data_masked[6644] = data_i[6644] & sel_one_hot_i[51];
  assign data_masked[6643] = data_i[6643] & sel_one_hot_i[51];
  assign data_masked[6642] = data_i[6642] & sel_one_hot_i[51];
  assign data_masked[6641] = data_i[6641] & sel_one_hot_i[51];
  assign data_masked[6640] = data_i[6640] & sel_one_hot_i[51];
  assign data_masked[6639] = data_i[6639] & sel_one_hot_i[51];
  assign data_masked[6638] = data_i[6638] & sel_one_hot_i[51];
  assign data_masked[6637] = data_i[6637] & sel_one_hot_i[51];
  assign data_masked[6636] = data_i[6636] & sel_one_hot_i[51];
  assign data_masked[6635] = data_i[6635] & sel_one_hot_i[51];
  assign data_masked[6634] = data_i[6634] & sel_one_hot_i[51];
  assign data_masked[6633] = data_i[6633] & sel_one_hot_i[51];
  assign data_masked[6632] = data_i[6632] & sel_one_hot_i[51];
  assign data_masked[6631] = data_i[6631] & sel_one_hot_i[51];
  assign data_masked[6630] = data_i[6630] & sel_one_hot_i[51];
  assign data_masked[6629] = data_i[6629] & sel_one_hot_i[51];
  assign data_masked[6628] = data_i[6628] & sel_one_hot_i[51];
  assign data_masked[6627] = data_i[6627] & sel_one_hot_i[51];
  assign data_masked[6626] = data_i[6626] & sel_one_hot_i[51];
  assign data_masked[6625] = data_i[6625] & sel_one_hot_i[51];
  assign data_masked[6624] = data_i[6624] & sel_one_hot_i[51];
  assign data_masked[6623] = data_i[6623] & sel_one_hot_i[51];
  assign data_masked[6622] = data_i[6622] & sel_one_hot_i[51];
  assign data_masked[6621] = data_i[6621] & sel_one_hot_i[51];
  assign data_masked[6620] = data_i[6620] & sel_one_hot_i[51];
  assign data_masked[6619] = data_i[6619] & sel_one_hot_i[51];
  assign data_masked[6618] = data_i[6618] & sel_one_hot_i[51];
  assign data_masked[6617] = data_i[6617] & sel_one_hot_i[51];
  assign data_masked[6616] = data_i[6616] & sel_one_hot_i[51];
  assign data_masked[6615] = data_i[6615] & sel_one_hot_i[51];
  assign data_masked[6614] = data_i[6614] & sel_one_hot_i[51];
  assign data_masked[6613] = data_i[6613] & sel_one_hot_i[51];
  assign data_masked[6612] = data_i[6612] & sel_one_hot_i[51];
  assign data_masked[6611] = data_i[6611] & sel_one_hot_i[51];
  assign data_masked[6610] = data_i[6610] & sel_one_hot_i[51];
  assign data_masked[6609] = data_i[6609] & sel_one_hot_i[51];
  assign data_masked[6608] = data_i[6608] & sel_one_hot_i[51];
  assign data_masked[6607] = data_i[6607] & sel_one_hot_i[51];
  assign data_masked[6606] = data_i[6606] & sel_one_hot_i[51];
  assign data_masked[6605] = data_i[6605] & sel_one_hot_i[51];
  assign data_masked[6604] = data_i[6604] & sel_one_hot_i[51];
  assign data_masked[6603] = data_i[6603] & sel_one_hot_i[51];
  assign data_masked[6602] = data_i[6602] & sel_one_hot_i[51];
  assign data_masked[6601] = data_i[6601] & sel_one_hot_i[51];
  assign data_masked[6600] = data_i[6600] & sel_one_hot_i[51];
  assign data_masked[6599] = data_i[6599] & sel_one_hot_i[51];
  assign data_masked[6598] = data_i[6598] & sel_one_hot_i[51];
  assign data_masked[6597] = data_i[6597] & sel_one_hot_i[51];
  assign data_masked[6596] = data_i[6596] & sel_one_hot_i[51];
  assign data_masked[6595] = data_i[6595] & sel_one_hot_i[51];
  assign data_masked[6594] = data_i[6594] & sel_one_hot_i[51];
  assign data_masked[6593] = data_i[6593] & sel_one_hot_i[51];
  assign data_masked[6592] = data_i[6592] & sel_one_hot_i[51];
  assign data_masked[6591] = data_i[6591] & sel_one_hot_i[51];
  assign data_masked[6590] = data_i[6590] & sel_one_hot_i[51];
  assign data_masked[6589] = data_i[6589] & sel_one_hot_i[51];
  assign data_masked[6588] = data_i[6588] & sel_one_hot_i[51];
  assign data_masked[6587] = data_i[6587] & sel_one_hot_i[51];
  assign data_masked[6586] = data_i[6586] & sel_one_hot_i[51];
  assign data_masked[6585] = data_i[6585] & sel_one_hot_i[51];
  assign data_masked[6584] = data_i[6584] & sel_one_hot_i[51];
  assign data_masked[6583] = data_i[6583] & sel_one_hot_i[51];
  assign data_masked[6582] = data_i[6582] & sel_one_hot_i[51];
  assign data_masked[6581] = data_i[6581] & sel_one_hot_i[51];
  assign data_masked[6580] = data_i[6580] & sel_one_hot_i[51];
  assign data_masked[6579] = data_i[6579] & sel_one_hot_i[51];
  assign data_masked[6578] = data_i[6578] & sel_one_hot_i[51];
  assign data_masked[6577] = data_i[6577] & sel_one_hot_i[51];
  assign data_masked[6576] = data_i[6576] & sel_one_hot_i[51];
  assign data_masked[6575] = data_i[6575] & sel_one_hot_i[51];
  assign data_masked[6574] = data_i[6574] & sel_one_hot_i[51];
  assign data_masked[6573] = data_i[6573] & sel_one_hot_i[51];
  assign data_masked[6572] = data_i[6572] & sel_one_hot_i[51];
  assign data_masked[6571] = data_i[6571] & sel_one_hot_i[51];
  assign data_masked[6570] = data_i[6570] & sel_one_hot_i[51];
  assign data_masked[6569] = data_i[6569] & sel_one_hot_i[51];
  assign data_masked[6568] = data_i[6568] & sel_one_hot_i[51];
  assign data_masked[6567] = data_i[6567] & sel_one_hot_i[51];
  assign data_masked[6566] = data_i[6566] & sel_one_hot_i[51];
  assign data_masked[6565] = data_i[6565] & sel_one_hot_i[51];
  assign data_masked[6564] = data_i[6564] & sel_one_hot_i[51];
  assign data_masked[6563] = data_i[6563] & sel_one_hot_i[51];
  assign data_masked[6562] = data_i[6562] & sel_one_hot_i[51];
  assign data_masked[6561] = data_i[6561] & sel_one_hot_i[51];
  assign data_masked[6560] = data_i[6560] & sel_one_hot_i[51];
  assign data_masked[6559] = data_i[6559] & sel_one_hot_i[51];
  assign data_masked[6558] = data_i[6558] & sel_one_hot_i[51];
  assign data_masked[6557] = data_i[6557] & sel_one_hot_i[51];
  assign data_masked[6556] = data_i[6556] & sel_one_hot_i[51];
  assign data_masked[6555] = data_i[6555] & sel_one_hot_i[51];
  assign data_masked[6554] = data_i[6554] & sel_one_hot_i[51];
  assign data_masked[6553] = data_i[6553] & sel_one_hot_i[51];
  assign data_masked[6552] = data_i[6552] & sel_one_hot_i[51];
  assign data_masked[6551] = data_i[6551] & sel_one_hot_i[51];
  assign data_masked[6550] = data_i[6550] & sel_one_hot_i[51];
  assign data_masked[6549] = data_i[6549] & sel_one_hot_i[51];
  assign data_masked[6548] = data_i[6548] & sel_one_hot_i[51];
  assign data_masked[6547] = data_i[6547] & sel_one_hot_i[51];
  assign data_masked[6546] = data_i[6546] & sel_one_hot_i[51];
  assign data_masked[6545] = data_i[6545] & sel_one_hot_i[51];
  assign data_masked[6544] = data_i[6544] & sel_one_hot_i[51];
  assign data_masked[6543] = data_i[6543] & sel_one_hot_i[51];
  assign data_masked[6542] = data_i[6542] & sel_one_hot_i[51];
  assign data_masked[6541] = data_i[6541] & sel_one_hot_i[51];
  assign data_masked[6540] = data_i[6540] & sel_one_hot_i[51];
  assign data_masked[6539] = data_i[6539] & sel_one_hot_i[51];
  assign data_masked[6538] = data_i[6538] & sel_one_hot_i[51];
  assign data_masked[6537] = data_i[6537] & sel_one_hot_i[51];
  assign data_masked[6536] = data_i[6536] & sel_one_hot_i[51];
  assign data_masked[6535] = data_i[6535] & sel_one_hot_i[51];
  assign data_masked[6534] = data_i[6534] & sel_one_hot_i[51];
  assign data_masked[6533] = data_i[6533] & sel_one_hot_i[51];
  assign data_masked[6532] = data_i[6532] & sel_one_hot_i[51];
  assign data_masked[6531] = data_i[6531] & sel_one_hot_i[51];
  assign data_masked[6530] = data_i[6530] & sel_one_hot_i[51];
  assign data_masked[6529] = data_i[6529] & sel_one_hot_i[51];
  assign data_masked[6528] = data_i[6528] & sel_one_hot_i[51];
  assign data_masked[6783] = data_i[6783] & sel_one_hot_i[52];
  assign data_masked[6782] = data_i[6782] & sel_one_hot_i[52];
  assign data_masked[6781] = data_i[6781] & sel_one_hot_i[52];
  assign data_masked[6780] = data_i[6780] & sel_one_hot_i[52];
  assign data_masked[6779] = data_i[6779] & sel_one_hot_i[52];
  assign data_masked[6778] = data_i[6778] & sel_one_hot_i[52];
  assign data_masked[6777] = data_i[6777] & sel_one_hot_i[52];
  assign data_masked[6776] = data_i[6776] & sel_one_hot_i[52];
  assign data_masked[6775] = data_i[6775] & sel_one_hot_i[52];
  assign data_masked[6774] = data_i[6774] & sel_one_hot_i[52];
  assign data_masked[6773] = data_i[6773] & sel_one_hot_i[52];
  assign data_masked[6772] = data_i[6772] & sel_one_hot_i[52];
  assign data_masked[6771] = data_i[6771] & sel_one_hot_i[52];
  assign data_masked[6770] = data_i[6770] & sel_one_hot_i[52];
  assign data_masked[6769] = data_i[6769] & sel_one_hot_i[52];
  assign data_masked[6768] = data_i[6768] & sel_one_hot_i[52];
  assign data_masked[6767] = data_i[6767] & sel_one_hot_i[52];
  assign data_masked[6766] = data_i[6766] & sel_one_hot_i[52];
  assign data_masked[6765] = data_i[6765] & sel_one_hot_i[52];
  assign data_masked[6764] = data_i[6764] & sel_one_hot_i[52];
  assign data_masked[6763] = data_i[6763] & sel_one_hot_i[52];
  assign data_masked[6762] = data_i[6762] & sel_one_hot_i[52];
  assign data_masked[6761] = data_i[6761] & sel_one_hot_i[52];
  assign data_masked[6760] = data_i[6760] & sel_one_hot_i[52];
  assign data_masked[6759] = data_i[6759] & sel_one_hot_i[52];
  assign data_masked[6758] = data_i[6758] & sel_one_hot_i[52];
  assign data_masked[6757] = data_i[6757] & sel_one_hot_i[52];
  assign data_masked[6756] = data_i[6756] & sel_one_hot_i[52];
  assign data_masked[6755] = data_i[6755] & sel_one_hot_i[52];
  assign data_masked[6754] = data_i[6754] & sel_one_hot_i[52];
  assign data_masked[6753] = data_i[6753] & sel_one_hot_i[52];
  assign data_masked[6752] = data_i[6752] & sel_one_hot_i[52];
  assign data_masked[6751] = data_i[6751] & sel_one_hot_i[52];
  assign data_masked[6750] = data_i[6750] & sel_one_hot_i[52];
  assign data_masked[6749] = data_i[6749] & sel_one_hot_i[52];
  assign data_masked[6748] = data_i[6748] & sel_one_hot_i[52];
  assign data_masked[6747] = data_i[6747] & sel_one_hot_i[52];
  assign data_masked[6746] = data_i[6746] & sel_one_hot_i[52];
  assign data_masked[6745] = data_i[6745] & sel_one_hot_i[52];
  assign data_masked[6744] = data_i[6744] & sel_one_hot_i[52];
  assign data_masked[6743] = data_i[6743] & sel_one_hot_i[52];
  assign data_masked[6742] = data_i[6742] & sel_one_hot_i[52];
  assign data_masked[6741] = data_i[6741] & sel_one_hot_i[52];
  assign data_masked[6740] = data_i[6740] & sel_one_hot_i[52];
  assign data_masked[6739] = data_i[6739] & sel_one_hot_i[52];
  assign data_masked[6738] = data_i[6738] & sel_one_hot_i[52];
  assign data_masked[6737] = data_i[6737] & sel_one_hot_i[52];
  assign data_masked[6736] = data_i[6736] & sel_one_hot_i[52];
  assign data_masked[6735] = data_i[6735] & sel_one_hot_i[52];
  assign data_masked[6734] = data_i[6734] & sel_one_hot_i[52];
  assign data_masked[6733] = data_i[6733] & sel_one_hot_i[52];
  assign data_masked[6732] = data_i[6732] & sel_one_hot_i[52];
  assign data_masked[6731] = data_i[6731] & sel_one_hot_i[52];
  assign data_masked[6730] = data_i[6730] & sel_one_hot_i[52];
  assign data_masked[6729] = data_i[6729] & sel_one_hot_i[52];
  assign data_masked[6728] = data_i[6728] & sel_one_hot_i[52];
  assign data_masked[6727] = data_i[6727] & sel_one_hot_i[52];
  assign data_masked[6726] = data_i[6726] & sel_one_hot_i[52];
  assign data_masked[6725] = data_i[6725] & sel_one_hot_i[52];
  assign data_masked[6724] = data_i[6724] & sel_one_hot_i[52];
  assign data_masked[6723] = data_i[6723] & sel_one_hot_i[52];
  assign data_masked[6722] = data_i[6722] & sel_one_hot_i[52];
  assign data_masked[6721] = data_i[6721] & sel_one_hot_i[52];
  assign data_masked[6720] = data_i[6720] & sel_one_hot_i[52];
  assign data_masked[6719] = data_i[6719] & sel_one_hot_i[52];
  assign data_masked[6718] = data_i[6718] & sel_one_hot_i[52];
  assign data_masked[6717] = data_i[6717] & sel_one_hot_i[52];
  assign data_masked[6716] = data_i[6716] & sel_one_hot_i[52];
  assign data_masked[6715] = data_i[6715] & sel_one_hot_i[52];
  assign data_masked[6714] = data_i[6714] & sel_one_hot_i[52];
  assign data_masked[6713] = data_i[6713] & sel_one_hot_i[52];
  assign data_masked[6712] = data_i[6712] & sel_one_hot_i[52];
  assign data_masked[6711] = data_i[6711] & sel_one_hot_i[52];
  assign data_masked[6710] = data_i[6710] & sel_one_hot_i[52];
  assign data_masked[6709] = data_i[6709] & sel_one_hot_i[52];
  assign data_masked[6708] = data_i[6708] & sel_one_hot_i[52];
  assign data_masked[6707] = data_i[6707] & sel_one_hot_i[52];
  assign data_masked[6706] = data_i[6706] & sel_one_hot_i[52];
  assign data_masked[6705] = data_i[6705] & sel_one_hot_i[52];
  assign data_masked[6704] = data_i[6704] & sel_one_hot_i[52];
  assign data_masked[6703] = data_i[6703] & sel_one_hot_i[52];
  assign data_masked[6702] = data_i[6702] & sel_one_hot_i[52];
  assign data_masked[6701] = data_i[6701] & sel_one_hot_i[52];
  assign data_masked[6700] = data_i[6700] & sel_one_hot_i[52];
  assign data_masked[6699] = data_i[6699] & sel_one_hot_i[52];
  assign data_masked[6698] = data_i[6698] & sel_one_hot_i[52];
  assign data_masked[6697] = data_i[6697] & sel_one_hot_i[52];
  assign data_masked[6696] = data_i[6696] & sel_one_hot_i[52];
  assign data_masked[6695] = data_i[6695] & sel_one_hot_i[52];
  assign data_masked[6694] = data_i[6694] & sel_one_hot_i[52];
  assign data_masked[6693] = data_i[6693] & sel_one_hot_i[52];
  assign data_masked[6692] = data_i[6692] & sel_one_hot_i[52];
  assign data_masked[6691] = data_i[6691] & sel_one_hot_i[52];
  assign data_masked[6690] = data_i[6690] & sel_one_hot_i[52];
  assign data_masked[6689] = data_i[6689] & sel_one_hot_i[52];
  assign data_masked[6688] = data_i[6688] & sel_one_hot_i[52];
  assign data_masked[6687] = data_i[6687] & sel_one_hot_i[52];
  assign data_masked[6686] = data_i[6686] & sel_one_hot_i[52];
  assign data_masked[6685] = data_i[6685] & sel_one_hot_i[52];
  assign data_masked[6684] = data_i[6684] & sel_one_hot_i[52];
  assign data_masked[6683] = data_i[6683] & sel_one_hot_i[52];
  assign data_masked[6682] = data_i[6682] & sel_one_hot_i[52];
  assign data_masked[6681] = data_i[6681] & sel_one_hot_i[52];
  assign data_masked[6680] = data_i[6680] & sel_one_hot_i[52];
  assign data_masked[6679] = data_i[6679] & sel_one_hot_i[52];
  assign data_masked[6678] = data_i[6678] & sel_one_hot_i[52];
  assign data_masked[6677] = data_i[6677] & sel_one_hot_i[52];
  assign data_masked[6676] = data_i[6676] & sel_one_hot_i[52];
  assign data_masked[6675] = data_i[6675] & sel_one_hot_i[52];
  assign data_masked[6674] = data_i[6674] & sel_one_hot_i[52];
  assign data_masked[6673] = data_i[6673] & sel_one_hot_i[52];
  assign data_masked[6672] = data_i[6672] & sel_one_hot_i[52];
  assign data_masked[6671] = data_i[6671] & sel_one_hot_i[52];
  assign data_masked[6670] = data_i[6670] & sel_one_hot_i[52];
  assign data_masked[6669] = data_i[6669] & sel_one_hot_i[52];
  assign data_masked[6668] = data_i[6668] & sel_one_hot_i[52];
  assign data_masked[6667] = data_i[6667] & sel_one_hot_i[52];
  assign data_masked[6666] = data_i[6666] & sel_one_hot_i[52];
  assign data_masked[6665] = data_i[6665] & sel_one_hot_i[52];
  assign data_masked[6664] = data_i[6664] & sel_one_hot_i[52];
  assign data_masked[6663] = data_i[6663] & sel_one_hot_i[52];
  assign data_masked[6662] = data_i[6662] & sel_one_hot_i[52];
  assign data_masked[6661] = data_i[6661] & sel_one_hot_i[52];
  assign data_masked[6660] = data_i[6660] & sel_one_hot_i[52];
  assign data_masked[6659] = data_i[6659] & sel_one_hot_i[52];
  assign data_masked[6658] = data_i[6658] & sel_one_hot_i[52];
  assign data_masked[6657] = data_i[6657] & sel_one_hot_i[52];
  assign data_masked[6656] = data_i[6656] & sel_one_hot_i[52];
  assign data_masked[6911] = data_i[6911] & sel_one_hot_i[53];
  assign data_masked[6910] = data_i[6910] & sel_one_hot_i[53];
  assign data_masked[6909] = data_i[6909] & sel_one_hot_i[53];
  assign data_masked[6908] = data_i[6908] & sel_one_hot_i[53];
  assign data_masked[6907] = data_i[6907] & sel_one_hot_i[53];
  assign data_masked[6906] = data_i[6906] & sel_one_hot_i[53];
  assign data_masked[6905] = data_i[6905] & sel_one_hot_i[53];
  assign data_masked[6904] = data_i[6904] & sel_one_hot_i[53];
  assign data_masked[6903] = data_i[6903] & sel_one_hot_i[53];
  assign data_masked[6902] = data_i[6902] & sel_one_hot_i[53];
  assign data_masked[6901] = data_i[6901] & sel_one_hot_i[53];
  assign data_masked[6900] = data_i[6900] & sel_one_hot_i[53];
  assign data_masked[6899] = data_i[6899] & sel_one_hot_i[53];
  assign data_masked[6898] = data_i[6898] & sel_one_hot_i[53];
  assign data_masked[6897] = data_i[6897] & sel_one_hot_i[53];
  assign data_masked[6896] = data_i[6896] & sel_one_hot_i[53];
  assign data_masked[6895] = data_i[6895] & sel_one_hot_i[53];
  assign data_masked[6894] = data_i[6894] & sel_one_hot_i[53];
  assign data_masked[6893] = data_i[6893] & sel_one_hot_i[53];
  assign data_masked[6892] = data_i[6892] & sel_one_hot_i[53];
  assign data_masked[6891] = data_i[6891] & sel_one_hot_i[53];
  assign data_masked[6890] = data_i[6890] & sel_one_hot_i[53];
  assign data_masked[6889] = data_i[6889] & sel_one_hot_i[53];
  assign data_masked[6888] = data_i[6888] & sel_one_hot_i[53];
  assign data_masked[6887] = data_i[6887] & sel_one_hot_i[53];
  assign data_masked[6886] = data_i[6886] & sel_one_hot_i[53];
  assign data_masked[6885] = data_i[6885] & sel_one_hot_i[53];
  assign data_masked[6884] = data_i[6884] & sel_one_hot_i[53];
  assign data_masked[6883] = data_i[6883] & sel_one_hot_i[53];
  assign data_masked[6882] = data_i[6882] & sel_one_hot_i[53];
  assign data_masked[6881] = data_i[6881] & sel_one_hot_i[53];
  assign data_masked[6880] = data_i[6880] & sel_one_hot_i[53];
  assign data_masked[6879] = data_i[6879] & sel_one_hot_i[53];
  assign data_masked[6878] = data_i[6878] & sel_one_hot_i[53];
  assign data_masked[6877] = data_i[6877] & sel_one_hot_i[53];
  assign data_masked[6876] = data_i[6876] & sel_one_hot_i[53];
  assign data_masked[6875] = data_i[6875] & sel_one_hot_i[53];
  assign data_masked[6874] = data_i[6874] & sel_one_hot_i[53];
  assign data_masked[6873] = data_i[6873] & sel_one_hot_i[53];
  assign data_masked[6872] = data_i[6872] & sel_one_hot_i[53];
  assign data_masked[6871] = data_i[6871] & sel_one_hot_i[53];
  assign data_masked[6870] = data_i[6870] & sel_one_hot_i[53];
  assign data_masked[6869] = data_i[6869] & sel_one_hot_i[53];
  assign data_masked[6868] = data_i[6868] & sel_one_hot_i[53];
  assign data_masked[6867] = data_i[6867] & sel_one_hot_i[53];
  assign data_masked[6866] = data_i[6866] & sel_one_hot_i[53];
  assign data_masked[6865] = data_i[6865] & sel_one_hot_i[53];
  assign data_masked[6864] = data_i[6864] & sel_one_hot_i[53];
  assign data_masked[6863] = data_i[6863] & sel_one_hot_i[53];
  assign data_masked[6862] = data_i[6862] & sel_one_hot_i[53];
  assign data_masked[6861] = data_i[6861] & sel_one_hot_i[53];
  assign data_masked[6860] = data_i[6860] & sel_one_hot_i[53];
  assign data_masked[6859] = data_i[6859] & sel_one_hot_i[53];
  assign data_masked[6858] = data_i[6858] & sel_one_hot_i[53];
  assign data_masked[6857] = data_i[6857] & sel_one_hot_i[53];
  assign data_masked[6856] = data_i[6856] & sel_one_hot_i[53];
  assign data_masked[6855] = data_i[6855] & sel_one_hot_i[53];
  assign data_masked[6854] = data_i[6854] & sel_one_hot_i[53];
  assign data_masked[6853] = data_i[6853] & sel_one_hot_i[53];
  assign data_masked[6852] = data_i[6852] & sel_one_hot_i[53];
  assign data_masked[6851] = data_i[6851] & sel_one_hot_i[53];
  assign data_masked[6850] = data_i[6850] & sel_one_hot_i[53];
  assign data_masked[6849] = data_i[6849] & sel_one_hot_i[53];
  assign data_masked[6848] = data_i[6848] & sel_one_hot_i[53];
  assign data_masked[6847] = data_i[6847] & sel_one_hot_i[53];
  assign data_masked[6846] = data_i[6846] & sel_one_hot_i[53];
  assign data_masked[6845] = data_i[6845] & sel_one_hot_i[53];
  assign data_masked[6844] = data_i[6844] & sel_one_hot_i[53];
  assign data_masked[6843] = data_i[6843] & sel_one_hot_i[53];
  assign data_masked[6842] = data_i[6842] & sel_one_hot_i[53];
  assign data_masked[6841] = data_i[6841] & sel_one_hot_i[53];
  assign data_masked[6840] = data_i[6840] & sel_one_hot_i[53];
  assign data_masked[6839] = data_i[6839] & sel_one_hot_i[53];
  assign data_masked[6838] = data_i[6838] & sel_one_hot_i[53];
  assign data_masked[6837] = data_i[6837] & sel_one_hot_i[53];
  assign data_masked[6836] = data_i[6836] & sel_one_hot_i[53];
  assign data_masked[6835] = data_i[6835] & sel_one_hot_i[53];
  assign data_masked[6834] = data_i[6834] & sel_one_hot_i[53];
  assign data_masked[6833] = data_i[6833] & sel_one_hot_i[53];
  assign data_masked[6832] = data_i[6832] & sel_one_hot_i[53];
  assign data_masked[6831] = data_i[6831] & sel_one_hot_i[53];
  assign data_masked[6830] = data_i[6830] & sel_one_hot_i[53];
  assign data_masked[6829] = data_i[6829] & sel_one_hot_i[53];
  assign data_masked[6828] = data_i[6828] & sel_one_hot_i[53];
  assign data_masked[6827] = data_i[6827] & sel_one_hot_i[53];
  assign data_masked[6826] = data_i[6826] & sel_one_hot_i[53];
  assign data_masked[6825] = data_i[6825] & sel_one_hot_i[53];
  assign data_masked[6824] = data_i[6824] & sel_one_hot_i[53];
  assign data_masked[6823] = data_i[6823] & sel_one_hot_i[53];
  assign data_masked[6822] = data_i[6822] & sel_one_hot_i[53];
  assign data_masked[6821] = data_i[6821] & sel_one_hot_i[53];
  assign data_masked[6820] = data_i[6820] & sel_one_hot_i[53];
  assign data_masked[6819] = data_i[6819] & sel_one_hot_i[53];
  assign data_masked[6818] = data_i[6818] & sel_one_hot_i[53];
  assign data_masked[6817] = data_i[6817] & sel_one_hot_i[53];
  assign data_masked[6816] = data_i[6816] & sel_one_hot_i[53];
  assign data_masked[6815] = data_i[6815] & sel_one_hot_i[53];
  assign data_masked[6814] = data_i[6814] & sel_one_hot_i[53];
  assign data_masked[6813] = data_i[6813] & sel_one_hot_i[53];
  assign data_masked[6812] = data_i[6812] & sel_one_hot_i[53];
  assign data_masked[6811] = data_i[6811] & sel_one_hot_i[53];
  assign data_masked[6810] = data_i[6810] & sel_one_hot_i[53];
  assign data_masked[6809] = data_i[6809] & sel_one_hot_i[53];
  assign data_masked[6808] = data_i[6808] & sel_one_hot_i[53];
  assign data_masked[6807] = data_i[6807] & sel_one_hot_i[53];
  assign data_masked[6806] = data_i[6806] & sel_one_hot_i[53];
  assign data_masked[6805] = data_i[6805] & sel_one_hot_i[53];
  assign data_masked[6804] = data_i[6804] & sel_one_hot_i[53];
  assign data_masked[6803] = data_i[6803] & sel_one_hot_i[53];
  assign data_masked[6802] = data_i[6802] & sel_one_hot_i[53];
  assign data_masked[6801] = data_i[6801] & sel_one_hot_i[53];
  assign data_masked[6800] = data_i[6800] & sel_one_hot_i[53];
  assign data_masked[6799] = data_i[6799] & sel_one_hot_i[53];
  assign data_masked[6798] = data_i[6798] & sel_one_hot_i[53];
  assign data_masked[6797] = data_i[6797] & sel_one_hot_i[53];
  assign data_masked[6796] = data_i[6796] & sel_one_hot_i[53];
  assign data_masked[6795] = data_i[6795] & sel_one_hot_i[53];
  assign data_masked[6794] = data_i[6794] & sel_one_hot_i[53];
  assign data_masked[6793] = data_i[6793] & sel_one_hot_i[53];
  assign data_masked[6792] = data_i[6792] & sel_one_hot_i[53];
  assign data_masked[6791] = data_i[6791] & sel_one_hot_i[53];
  assign data_masked[6790] = data_i[6790] & sel_one_hot_i[53];
  assign data_masked[6789] = data_i[6789] & sel_one_hot_i[53];
  assign data_masked[6788] = data_i[6788] & sel_one_hot_i[53];
  assign data_masked[6787] = data_i[6787] & sel_one_hot_i[53];
  assign data_masked[6786] = data_i[6786] & sel_one_hot_i[53];
  assign data_masked[6785] = data_i[6785] & sel_one_hot_i[53];
  assign data_masked[6784] = data_i[6784] & sel_one_hot_i[53];
  assign data_masked[7039] = data_i[7039] & sel_one_hot_i[54];
  assign data_masked[7038] = data_i[7038] & sel_one_hot_i[54];
  assign data_masked[7037] = data_i[7037] & sel_one_hot_i[54];
  assign data_masked[7036] = data_i[7036] & sel_one_hot_i[54];
  assign data_masked[7035] = data_i[7035] & sel_one_hot_i[54];
  assign data_masked[7034] = data_i[7034] & sel_one_hot_i[54];
  assign data_masked[7033] = data_i[7033] & sel_one_hot_i[54];
  assign data_masked[7032] = data_i[7032] & sel_one_hot_i[54];
  assign data_masked[7031] = data_i[7031] & sel_one_hot_i[54];
  assign data_masked[7030] = data_i[7030] & sel_one_hot_i[54];
  assign data_masked[7029] = data_i[7029] & sel_one_hot_i[54];
  assign data_masked[7028] = data_i[7028] & sel_one_hot_i[54];
  assign data_masked[7027] = data_i[7027] & sel_one_hot_i[54];
  assign data_masked[7026] = data_i[7026] & sel_one_hot_i[54];
  assign data_masked[7025] = data_i[7025] & sel_one_hot_i[54];
  assign data_masked[7024] = data_i[7024] & sel_one_hot_i[54];
  assign data_masked[7023] = data_i[7023] & sel_one_hot_i[54];
  assign data_masked[7022] = data_i[7022] & sel_one_hot_i[54];
  assign data_masked[7021] = data_i[7021] & sel_one_hot_i[54];
  assign data_masked[7020] = data_i[7020] & sel_one_hot_i[54];
  assign data_masked[7019] = data_i[7019] & sel_one_hot_i[54];
  assign data_masked[7018] = data_i[7018] & sel_one_hot_i[54];
  assign data_masked[7017] = data_i[7017] & sel_one_hot_i[54];
  assign data_masked[7016] = data_i[7016] & sel_one_hot_i[54];
  assign data_masked[7015] = data_i[7015] & sel_one_hot_i[54];
  assign data_masked[7014] = data_i[7014] & sel_one_hot_i[54];
  assign data_masked[7013] = data_i[7013] & sel_one_hot_i[54];
  assign data_masked[7012] = data_i[7012] & sel_one_hot_i[54];
  assign data_masked[7011] = data_i[7011] & sel_one_hot_i[54];
  assign data_masked[7010] = data_i[7010] & sel_one_hot_i[54];
  assign data_masked[7009] = data_i[7009] & sel_one_hot_i[54];
  assign data_masked[7008] = data_i[7008] & sel_one_hot_i[54];
  assign data_masked[7007] = data_i[7007] & sel_one_hot_i[54];
  assign data_masked[7006] = data_i[7006] & sel_one_hot_i[54];
  assign data_masked[7005] = data_i[7005] & sel_one_hot_i[54];
  assign data_masked[7004] = data_i[7004] & sel_one_hot_i[54];
  assign data_masked[7003] = data_i[7003] & sel_one_hot_i[54];
  assign data_masked[7002] = data_i[7002] & sel_one_hot_i[54];
  assign data_masked[7001] = data_i[7001] & sel_one_hot_i[54];
  assign data_masked[7000] = data_i[7000] & sel_one_hot_i[54];
  assign data_masked[6999] = data_i[6999] & sel_one_hot_i[54];
  assign data_masked[6998] = data_i[6998] & sel_one_hot_i[54];
  assign data_masked[6997] = data_i[6997] & sel_one_hot_i[54];
  assign data_masked[6996] = data_i[6996] & sel_one_hot_i[54];
  assign data_masked[6995] = data_i[6995] & sel_one_hot_i[54];
  assign data_masked[6994] = data_i[6994] & sel_one_hot_i[54];
  assign data_masked[6993] = data_i[6993] & sel_one_hot_i[54];
  assign data_masked[6992] = data_i[6992] & sel_one_hot_i[54];
  assign data_masked[6991] = data_i[6991] & sel_one_hot_i[54];
  assign data_masked[6990] = data_i[6990] & sel_one_hot_i[54];
  assign data_masked[6989] = data_i[6989] & sel_one_hot_i[54];
  assign data_masked[6988] = data_i[6988] & sel_one_hot_i[54];
  assign data_masked[6987] = data_i[6987] & sel_one_hot_i[54];
  assign data_masked[6986] = data_i[6986] & sel_one_hot_i[54];
  assign data_masked[6985] = data_i[6985] & sel_one_hot_i[54];
  assign data_masked[6984] = data_i[6984] & sel_one_hot_i[54];
  assign data_masked[6983] = data_i[6983] & sel_one_hot_i[54];
  assign data_masked[6982] = data_i[6982] & sel_one_hot_i[54];
  assign data_masked[6981] = data_i[6981] & sel_one_hot_i[54];
  assign data_masked[6980] = data_i[6980] & sel_one_hot_i[54];
  assign data_masked[6979] = data_i[6979] & sel_one_hot_i[54];
  assign data_masked[6978] = data_i[6978] & sel_one_hot_i[54];
  assign data_masked[6977] = data_i[6977] & sel_one_hot_i[54];
  assign data_masked[6976] = data_i[6976] & sel_one_hot_i[54];
  assign data_masked[6975] = data_i[6975] & sel_one_hot_i[54];
  assign data_masked[6974] = data_i[6974] & sel_one_hot_i[54];
  assign data_masked[6973] = data_i[6973] & sel_one_hot_i[54];
  assign data_masked[6972] = data_i[6972] & sel_one_hot_i[54];
  assign data_masked[6971] = data_i[6971] & sel_one_hot_i[54];
  assign data_masked[6970] = data_i[6970] & sel_one_hot_i[54];
  assign data_masked[6969] = data_i[6969] & sel_one_hot_i[54];
  assign data_masked[6968] = data_i[6968] & sel_one_hot_i[54];
  assign data_masked[6967] = data_i[6967] & sel_one_hot_i[54];
  assign data_masked[6966] = data_i[6966] & sel_one_hot_i[54];
  assign data_masked[6965] = data_i[6965] & sel_one_hot_i[54];
  assign data_masked[6964] = data_i[6964] & sel_one_hot_i[54];
  assign data_masked[6963] = data_i[6963] & sel_one_hot_i[54];
  assign data_masked[6962] = data_i[6962] & sel_one_hot_i[54];
  assign data_masked[6961] = data_i[6961] & sel_one_hot_i[54];
  assign data_masked[6960] = data_i[6960] & sel_one_hot_i[54];
  assign data_masked[6959] = data_i[6959] & sel_one_hot_i[54];
  assign data_masked[6958] = data_i[6958] & sel_one_hot_i[54];
  assign data_masked[6957] = data_i[6957] & sel_one_hot_i[54];
  assign data_masked[6956] = data_i[6956] & sel_one_hot_i[54];
  assign data_masked[6955] = data_i[6955] & sel_one_hot_i[54];
  assign data_masked[6954] = data_i[6954] & sel_one_hot_i[54];
  assign data_masked[6953] = data_i[6953] & sel_one_hot_i[54];
  assign data_masked[6952] = data_i[6952] & sel_one_hot_i[54];
  assign data_masked[6951] = data_i[6951] & sel_one_hot_i[54];
  assign data_masked[6950] = data_i[6950] & sel_one_hot_i[54];
  assign data_masked[6949] = data_i[6949] & sel_one_hot_i[54];
  assign data_masked[6948] = data_i[6948] & sel_one_hot_i[54];
  assign data_masked[6947] = data_i[6947] & sel_one_hot_i[54];
  assign data_masked[6946] = data_i[6946] & sel_one_hot_i[54];
  assign data_masked[6945] = data_i[6945] & sel_one_hot_i[54];
  assign data_masked[6944] = data_i[6944] & sel_one_hot_i[54];
  assign data_masked[6943] = data_i[6943] & sel_one_hot_i[54];
  assign data_masked[6942] = data_i[6942] & sel_one_hot_i[54];
  assign data_masked[6941] = data_i[6941] & sel_one_hot_i[54];
  assign data_masked[6940] = data_i[6940] & sel_one_hot_i[54];
  assign data_masked[6939] = data_i[6939] & sel_one_hot_i[54];
  assign data_masked[6938] = data_i[6938] & sel_one_hot_i[54];
  assign data_masked[6937] = data_i[6937] & sel_one_hot_i[54];
  assign data_masked[6936] = data_i[6936] & sel_one_hot_i[54];
  assign data_masked[6935] = data_i[6935] & sel_one_hot_i[54];
  assign data_masked[6934] = data_i[6934] & sel_one_hot_i[54];
  assign data_masked[6933] = data_i[6933] & sel_one_hot_i[54];
  assign data_masked[6932] = data_i[6932] & sel_one_hot_i[54];
  assign data_masked[6931] = data_i[6931] & sel_one_hot_i[54];
  assign data_masked[6930] = data_i[6930] & sel_one_hot_i[54];
  assign data_masked[6929] = data_i[6929] & sel_one_hot_i[54];
  assign data_masked[6928] = data_i[6928] & sel_one_hot_i[54];
  assign data_masked[6927] = data_i[6927] & sel_one_hot_i[54];
  assign data_masked[6926] = data_i[6926] & sel_one_hot_i[54];
  assign data_masked[6925] = data_i[6925] & sel_one_hot_i[54];
  assign data_masked[6924] = data_i[6924] & sel_one_hot_i[54];
  assign data_masked[6923] = data_i[6923] & sel_one_hot_i[54];
  assign data_masked[6922] = data_i[6922] & sel_one_hot_i[54];
  assign data_masked[6921] = data_i[6921] & sel_one_hot_i[54];
  assign data_masked[6920] = data_i[6920] & sel_one_hot_i[54];
  assign data_masked[6919] = data_i[6919] & sel_one_hot_i[54];
  assign data_masked[6918] = data_i[6918] & sel_one_hot_i[54];
  assign data_masked[6917] = data_i[6917] & sel_one_hot_i[54];
  assign data_masked[6916] = data_i[6916] & sel_one_hot_i[54];
  assign data_masked[6915] = data_i[6915] & sel_one_hot_i[54];
  assign data_masked[6914] = data_i[6914] & sel_one_hot_i[54];
  assign data_masked[6913] = data_i[6913] & sel_one_hot_i[54];
  assign data_masked[6912] = data_i[6912] & sel_one_hot_i[54];
  assign data_masked[7167] = data_i[7167] & sel_one_hot_i[55];
  assign data_masked[7166] = data_i[7166] & sel_one_hot_i[55];
  assign data_masked[7165] = data_i[7165] & sel_one_hot_i[55];
  assign data_masked[7164] = data_i[7164] & sel_one_hot_i[55];
  assign data_masked[7163] = data_i[7163] & sel_one_hot_i[55];
  assign data_masked[7162] = data_i[7162] & sel_one_hot_i[55];
  assign data_masked[7161] = data_i[7161] & sel_one_hot_i[55];
  assign data_masked[7160] = data_i[7160] & sel_one_hot_i[55];
  assign data_masked[7159] = data_i[7159] & sel_one_hot_i[55];
  assign data_masked[7158] = data_i[7158] & sel_one_hot_i[55];
  assign data_masked[7157] = data_i[7157] & sel_one_hot_i[55];
  assign data_masked[7156] = data_i[7156] & sel_one_hot_i[55];
  assign data_masked[7155] = data_i[7155] & sel_one_hot_i[55];
  assign data_masked[7154] = data_i[7154] & sel_one_hot_i[55];
  assign data_masked[7153] = data_i[7153] & sel_one_hot_i[55];
  assign data_masked[7152] = data_i[7152] & sel_one_hot_i[55];
  assign data_masked[7151] = data_i[7151] & sel_one_hot_i[55];
  assign data_masked[7150] = data_i[7150] & sel_one_hot_i[55];
  assign data_masked[7149] = data_i[7149] & sel_one_hot_i[55];
  assign data_masked[7148] = data_i[7148] & sel_one_hot_i[55];
  assign data_masked[7147] = data_i[7147] & sel_one_hot_i[55];
  assign data_masked[7146] = data_i[7146] & sel_one_hot_i[55];
  assign data_masked[7145] = data_i[7145] & sel_one_hot_i[55];
  assign data_masked[7144] = data_i[7144] & sel_one_hot_i[55];
  assign data_masked[7143] = data_i[7143] & sel_one_hot_i[55];
  assign data_masked[7142] = data_i[7142] & sel_one_hot_i[55];
  assign data_masked[7141] = data_i[7141] & sel_one_hot_i[55];
  assign data_masked[7140] = data_i[7140] & sel_one_hot_i[55];
  assign data_masked[7139] = data_i[7139] & sel_one_hot_i[55];
  assign data_masked[7138] = data_i[7138] & sel_one_hot_i[55];
  assign data_masked[7137] = data_i[7137] & sel_one_hot_i[55];
  assign data_masked[7136] = data_i[7136] & sel_one_hot_i[55];
  assign data_masked[7135] = data_i[7135] & sel_one_hot_i[55];
  assign data_masked[7134] = data_i[7134] & sel_one_hot_i[55];
  assign data_masked[7133] = data_i[7133] & sel_one_hot_i[55];
  assign data_masked[7132] = data_i[7132] & sel_one_hot_i[55];
  assign data_masked[7131] = data_i[7131] & sel_one_hot_i[55];
  assign data_masked[7130] = data_i[7130] & sel_one_hot_i[55];
  assign data_masked[7129] = data_i[7129] & sel_one_hot_i[55];
  assign data_masked[7128] = data_i[7128] & sel_one_hot_i[55];
  assign data_masked[7127] = data_i[7127] & sel_one_hot_i[55];
  assign data_masked[7126] = data_i[7126] & sel_one_hot_i[55];
  assign data_masked[7125] = data_i[7125] & sel_one_hot_i[55];
  assign data_masked[7124] = data_i[7124] & sel_one_hot_i[55];
  assign data_masked[7123] = data_i[7123] & sel_one_hot_i[55];
  assign data_masked[7122] = data_i[7122] & sel_one_hot_i[55];
  assign data_masked[7121] = data_i[7121] & sel_one_hot_i[55];
  assign data_masked[7120] = data_i[7120] & sel_one_hot_i[55];
  assign data_masked[7119] = data_i[7119] & sel_one_hot_i[55];
  assign data_masked[7118] = data_i[7118] & sel_one_hot_i[55];
  assign data_masked[7117] = data_i[7117] & sel_one_hot_i[55];
  assign data_masked[7116] = data_i[7116] & sel_one_hot_i[55];
  assign data_masked[7115] = data_i[7115] & sel_one_hot_i[55];
  assign data_masked[7114] = data_i[7114] & sel_one_hot_i[55];
  assign data_masked[7113] = data_i[7113] & sel_one_hot_i[55];
  assign data_masked[7112] = data_i[7112] & sel_one_hot_i[55];
  assign data_masked[7111] = data_i[7111] & sel_one_hot_i[55];
  assign data_masked[7110] = data_i[7110] & sel_one_hot_i[55];
  assign data_masked[7109] = data_i[7109] & sel_one_hot_i[55];
  assign data_masked[7108] = data_i[7108] & sel_one_hot_i[55];
  assign data_masked[7107] = data_i[7107] & sel_one_hot_i[55];
  assign data_masked[7106] = data_i[7106] & sel_one_hot_i[55];
  assign data_masked[7105] = data_i[7105] & sel_one_hot_i[55];
  assign data_masked[7104] = data_i[7104] & sel_one_hot_i[55];
  assign data_masked[7103] = data_i[7103] & sel_one_hot_i[55];
  assign data_masked[7102] = data_i[7102] & sel_one_hot_i[55];
  assign data_masked[7101] = data_i[7101] & sel_one_hot_i[55];
  assign data_masked[7100] = data_i[7100] & sel_one_hot_i[55];
  assign data_masked[7099] = data_i[7099] & sel_one_hot_i[55];
  assign data_masked[7098] = data_i[7098] & sel_one_hot_i[55];
  assign data_masked[7097] = data_i[7097] & sel_one_hot_i[55];
  assign data_masked[7096] = data_i[7096] & sel_one_hot_i[55];
  assign data_masked[7095] = data_i[7095] & sel_one_hot_i[55];
  assign data_masked[7094] = data_i[7094] & sel_one_hot_i[55];
  assign data_masked[7093] = data_i[7093] & sel_one_hot_i[55];
  assign data_masked[7092] = data_i[7092] & sel_one_hot_i[55];
  assign data_masked[7091] = data_i[7091] & sel_one_hot_i[55];
  assign data_masked[7090] = data_i[7090] & sel_one_hot_i[55];
  assign data_masked[7089] = data_i[7089] & sel_one_hot_i[55];
  assign data_masked[7088] = data_i[7088] & sel_one_hot_i[55];
  assign data_masked[7087] = data_i[7087] & sel_one_hot_i[55];
  assign data_masked[7086] = data_i[7086] & sel_one_hot_i[55];
  assign data_masked[7085] = data_i[7085] & sel_one_hot_i[55];
  assign data_masked[7084] = data_i[7084] & sel_one_hot_i[55];
  assign data_masked[7083] = data_i[7083] & sel_one_hot_i[55];
  assign data_masked[7082] = data_i[7082] & sel_one_hot_i[55];
  assign data_masked[7081] = data_i[7081] & sel_one_hot_i[55];
  assign data_masked[7080] = data_i[7080] & sel_one_hot_i[55];
  assign data_masked[7079] = data_i[7079] & sel_one_hot_i[55];
  assign data_masked[7078] = data_i[7078] & sel_one_hot_i[55];
  assign data_masked[7077] = data_i[7077] & sel_one_hot_i[55];
  assign data_masked[7076] = data_i[7076] & sel_one_hot_i[55];
  assign data_masked[7075] = data_i[7075] & sel_one_hot_i[55];
  assign data_masked[7074] = data_i[7074] & sel_one_hot_i[55];
  assign data_masked[7073] = data_i[7073] & sel_one_hot_i[55];
  assign data_masked[7072] = data_i[7072] & sel_one_hot_i[55];
  assign data_masked[7071] = data_i[7071] & sel_one_hot_i[55];
  assign data_masked[7070] = data_i[7070] & sel_one_hot_i[55];
  assign data_masked[7069] = data_i[7069] & sel_one_hot_i[55];
  assign data_masked[7068] = data_i[7068] & sel_one_hot_i[55];
  assign data_masked[7067] = data_i[7067] & sel_one_hot_i[55];
  assign data_masked[7066] = data_i[7066] & sel_one_hot_i[55];
  assign data_masked[7065] = data_i[7065] & sel_one_hot_i[55];
  assign data_masked[7064] = data_i[7064] & sel_one_hot_i[55];
  assign data_masked[7063] = data_i[7063] & sel_one_hot_i[55];
  assign data_masked[7062] = data_i[7062] & sel_one_hot_i[55];
  assign data_masked[7061] = data_i[7061] & sel_one_hot_i[55];
  assign data_masked[7060] = data_i[7060] & sel_one_hot_i[55];
  assign data_masked[7059] = data_i[7059] & sel_one_hot_i[55];
  assign data_masked[7058] = data_i[7058] & sel_one_hot_i[55];
  assign data_masked[7057] = data_i[7057] & sel_one_hot_i[55];
  assign data_masked[7056] = data_i[7056] & sel_one_hot_i[55];
  assign data_masked[7055] = data_i[7055] & sel_one_hot_i[55];
  assign data_masked[7054] = data_i[7054] & sel_one_hot_i[55];
  assign data_masked[7053] = data_i[7053] & sel_one_hot_i[55];
  assign data_masked[7052] = data_i[7052] & sel_one_hot_i[55];
  assign data_masked[7051] = data_i[7051] & sel_one_hot_i[55];
  assign data_masked[7050] = data_i[7050] & sel_one_hot_i[55];
  assign data_masked[7049] = data_i[7049] & sel_one_hot_i[55];
  assign data_masked[7048] = data_i[7048] & sel_one_hot_i[55];
  assign data_masked[7047] = data_i[7047] & sel_one_hot_i[55];
  assign data_masked[7046] = data_i[7046] & sel_one_hot_i[55];
  assign data_masked[7045] = data_i[7045] & sel_one_hot_i[55];
  assign data_masked[7044] = data_i[7044] & sel_one_hot_i[55];
  assign data_masked[7043] = data_i[7043] & sel_one_hot_i[55];
  assign data_masked[7042] = data_i[7042] & sel_one_hot_i[55];
  assign data_masked[7041] = data_i[7041] & sel_one_hot_i[55];
  assign data_masked[7040] = data_i[7040] & sel_one_hot_i[55];
  assign data_masked[7295] = data_i[7295] & sel_one_hot_i[56];
  assign data_masked[7294] = data_i[7294] & sel_one_hot_i[56];
  assign data_masked[7293] = data_i[7293] & sel_one_hot_i[56];
  assign data_masked[7292] = data_i[7292] & sel_one_hot_i[56];
  assign data_masked[7291] = data_i[7291] & sel_one_hot_i[56];
  assign data_masked[7290] = data_i[7290] & sel_one_hot_i[56];
  assign data_masked[7289] = data_i[7289] & sel_one_hot_i[56];
  assign data_masked[7288] = data_i[7288] & sel_one_hot_i[56];
  assign data_masked[7287] = data_i[7287] & sel_one_hot_i[56];
  assign data_masked[7286] = data_i[7286] & sel_one_hot_i[56];
  assign data_masked[7285] = data_i[7285] & sel_one_hot_i[56];
  assign data_masked[7284] = data_i[7284] & sel_one_hot_i[56];
  assign data_masked[7283] = data_i[7283] & sel_one_hot_i[56];
  assign data_masked[7282] = data_i[7282] & sel_one_hot_i[56];
  assign data_masked[7281] = data_i[7281] & sel_one_hot_i[56];
  assign data_masked[7280] = data_i[7280] & sel_one_hot_i[56];
  assign data_masked[7279] = data_i[7279] & sel_one_hot_i[56];
  assign data_masked[7278] = data_i[7278] & sel_one_hot_i[56];
  assign data_masked[7277] = data_i[7277] & sel_one_hot_i[56];
  assign data_masked[7276] = data_i[7276] & sel_one_hot_i[56];
  assign data_masked[7275] = data_i[7275] & sel_one_hot_i[56];
  assign data_masked[7274] = data_i[7274] & sel_one_hot_i[56];
  assign data_masked[7273] = data_i[7273] & sel_one_hot_i[56];
  assign data_masked[7272] = data_i[7272] & sel_one_hot_i[56];
  assign data_masked[7271] = data_i[7271] & sel_one_hot_i[56];
  assign data_masked[7270] = data_i[7270] & sel_one_hot_i[56];
  assign data_masked[7269] = data_i[7269] & sel_one_hot_i[56];
  assign data_masked[7268] = data_i[7268] & sel_one_hot_i[56];
  assign data_masked[7267] = data_i[7267] & sel_one_hot_i[56];
  assign data_masked[7266] = data_i[7266] & sel_one_hot_i[56];
  assign data_masked[7265] = data_i[7265] & sel_one_hot_i[56];
  assign data_masked[7264] = data_i[7264] & sel_one_hot_i[56];
  assign data_masked[7263] = data_i[7263] & sel_one_hot_i[56];
  assign data_masked[7262] = data_i[7262] & sel_one_hot_i[56];
  assign data_masked[7261] = data_i[7261] & sel_one_hot_i[56];
  assign data_masked[7260] = data_i[7260] & sel_one_hot_i[56];
  assign data_masked[7259] = data_i[7259] & sel_one_hot_i[56];
  assign data_masked[7258] = data_i[7258] & sel_one_hot_i[56];
  assign data_masked[7257] = data_i[7257] & sel_one_hot_i[56];
  assign data_masked[7256] = data_i[7256] & sel_one_hot_i[56];
  assign data_masked[7255] = data_i[7255] & sel_one_hot_i[56];
  assign data_masked[7254] = data_i[7254] & sel_one_hot_i[56];
  assign data_masked[7253] = data_i[7253] & sel_one_hot_i[56];
  assign data_masked[7252] = data_i[7252] & sel_one_hot_i[56];
  assign data_masked[7251] = data_i[7251] & sel_one_hot_i[56];
  assign data_masked[7250] = data_i[7250] & sel_one_hot_i[56];
  assign data_masked[7249] = data_i[7249] & sel_one_hot_i[56];
  assign data_masked[7248] = data_i[7248] & sel_one_hot_i[56];
  assign data_masked[7247] = data_i[7247] & sel_one_hot_i[56];
  assign data_masked[7246] = data_i[7246] & sel_one_hot_i[56];
  assign data_masked[7245] = data_i[7245] & sel_one_hot_i[56];
  assign data_masked[7244] = data_i[7244] & sel_one_hot_i[56];
  assign data_masked[7243] = data_i[7243] & sel_one_hot_i[56];
  assign data_masked[7242] = data_i[7242] & sel_one_hot_i[56];
  assign data_masked[7241] = data_i[7241] & sel_one_hot_i[56];
  assign data_masked[7240] = data_i[7240] & sel_one_hot_i[56];
  assign data_masked[7239] = data_i[7239] & sel_one_hot_i[56];
  assign data_masked[7238] = data_i[7238] & sel_one_hot_i[56];
  assign data_masked[7237] = data_i[7237] & sel_one_hot_i[56];
  assign data_masked[7236] = data_i[7236] & sel_one_hot_i[56];
  assign data_masked[7235] = data_i[7235] & sel_one_hot_i[56];
  assign data_masked[7234] = data_i[7234] & sel_one_hot_i[56];
  assign data_masked[7233] = data_i[7233] & sel_one_hot_i[56];
  assign data_masked[7232] = data_i[7232] & sel_one_hot_i[56];
  assign data_masked[7231] = data_i[7231] & sel_one_hot_i[56];
  assign data_masked[7230] = data_i[7230] & sel_one_hot_i[56];
  assign data_masked[7229] = data_i[7229] & sel_one_hot_i[56];
  assign data_masked[7228] = data_i[7228] & sel_one_hot_i[56];
  assign data_masked[7227] = data_i[7227] & sel_one_hot_i[56];
  assign data_masked[7226] = data_i[7226] & sel_one_hot_i[56];
  assign data_masked[7225] = data_i[7225] & sel_one_hot_i[56];
  assign data_masked[7224] = data_i[7224] & sel_one_hot_i[56];
  assign data_masked[7223] = data_i[7223] & sel_one_hot_i[56];
  assign data_masked[7222] = data_i[7222] & sel_one_hot_i[56];
  assign data_masked[7221] = data_i[7221] & sel_one_hot_i[56];
  assign data_masked[7220] = data_i[7220] & sel_one_hot_i[56];
  assign data_masked[7219] = data_i[7219] & sel_one_hot_i[56];
  assign data_masked[7218] = data_i[7218] & sel_one_hot_i[56];
  assign data_masked[7217] = data_i[7217] & sel_one_hot_i[56];
  assign data_masked[7216] = data_i[7216] & sel_one_hot_i[56];
  assign data_masked[7215] = data_i[7215] & sel_one_hot_i[56];
  assign data_masked[7214] = data_i[7214] & sel_one_hot_i[56];
  assign data_masked[7213] = data_i[7213] & sel_one_hot_i[56];
  assign data_masked[7212] = data_i[7212] & sel_one_hot_i[56];
  assign data_masked[7211] = data_i[7211] & sel_one_hot_i[56];
  assign data_masked[7210] = data_i[7210] & sel_one_hot_i[56];
  assign data_masked[7209] = data_i[7209] & sel_one_hot_i[56];
  assign data_masked[7208] = data_i[7208] & sel_one_hot_i[56];
  assign data_masked[7207] = data_i[7207] & sel_one_hot_i[56];
  assign data_masked[7206] = data_i[7206] & sel_one_hot_i[56];
  assign data_masked[7205] = data_i[7205] & sel_one_hot_i[56];
  assign data_masked[7204] = data_i[7204] & sel_one_hot_i[56];
  assign data_masked[7203] = data_i[7203] & sel_one_hot_i[56];
  assign data_masked[7202] = data_i[7202] & sel_one_hot_i[56];
  assign data_masked[7201] = data_i[7201] & sel_one_hot_i[56];
  assign data_masked[7200] = data_i[7200] & sel_one_hot_i[56];
  assign data_masked[7199] = data_i[7199] & sel_one_hot_i[56];
  assign data_masked[7198] = data_i[7198] & sel_one_hot_i[56];
  assign data_masked[7197] = data_i[7197] & sel_one_hot_i[56];
  assign data_masked[7196] = data_i[7196] & sel_one_hot_i[56];
  assign data_masked[7195] = data_i[7195] & sel_one_hot_i[56];
  assign data_masked[7194] = data_i[7194] & sel_one_hot_i[56];
  assign data_masked[7193] = data_i[7193] & sel_one_hot_i[56];
  assign data_masked[7192] = data_i[7192] & sel_one_hot_i[56];
  assign data_masked[7191] = data_i[7191] & sel_one_hot_i[56];
  assign data_masked[7190] = data_i[7190] & sel_one_hot_i[56];
  assign data_masked[7189] = data_i[7189] & sel_one_hot_i[56];
  assign data_masked[7188] = data_i[7188] & sel_one_hot_i[56];
  assign data_masked[7187] = data_i[7187] & sel_one_hot_i[56];
  assign data_masked[7186] = data_i[7186] & sel_one_hot_i[56];
  assign data_masked[7185] = data_i[7185] & sel_one_hot_i[56];
  assign data_masked[7184] = data_i[7184] & sel_one_hot_i[56];
  assign data_masked[7183] = data_i[7183] & sel_one_hot_i[56];
  assign data_masked[7182] = data_i[7182] & sel_one_hot_i[56];
  assign data_masked[7181] = data_i[7181] & sel_one_hot_i[56];
  assign data_masked[7180] = data_i[7180] & sel_one_hot_i[56];
  assign data_masked[7179] = data_i[7179] & sel_one_hot_i[56];
  assign data_masked[7178] = data_i[7178] & sel_one_hot_i[56];
  assign data_masked[7177] = data_i[7177] & sel_one_hot_i[56];
  assign data_masked[7176] = data_i[7176] & sel_one_hot_i[56];
  assign data_masked[7175] = data_i[7175] & sel_one_hot_i[56];
  assign data_masked[7174] = data_i[7174] & sel_one_hot_i[56];
  assign data_masked[7173] = data_i[7173] & sel_one_hot_i[56];
  assign data_masked[7172] = data_i[7172] & sel_one_hot_i[56];
  assign data_masked[7171] = data_i[7171] & sel_one_hot_i[56];
  assign data_masked[7170] = data_i[7170] & sel_one_hot_i[56];
  assign data_masked[7169] = data_i[7169] & sel_one_hot_i[56];
  assign data_masked[7168] = data_i[7168] & sel_one_hot_i[56];
  assign data_masked[7423] = data_i[7423] & sel_one_hot_i[57];
  assign data_masked[7422] = data_i[7422] & sel_one_hot_i[57];
  assign data_masked[7421] = data_i[7421] & sel_one_hot_i[57];
  assign data_masked[7420] = data_i[7420] & sel_one_hot_i[57];
  assign data_masked[7419] = data_i[7419] & sel_one_hot_i[57];
  assign data_masked[7418] = data_i[7418] & sel_one_hot_i[57];
  assign data_masked[7417] = data_i[7417] & sel_one_hot_i[57];
  assign data_masked[7416] = data_i[7416] & sel_one_hot_i[57];
  assign data_masked[7415] = data_i[7415] & sel_one_hot_i[57];
  assign data_masked[7414] = data_i[7414] & sel_one_hot_i[57];
  assign data_masked[7413] = data_i[7413] & sel_one_hot_i[57];
  assign data_masked[7412] = data_i[7412] & sel_one_hot_i[57];
  assign data_masked[7411] = data_i[7411] & sel_one_hot_i[57];
  assign data_masked[7410] = data_i[7410] & sel_one_hot_i[57];
  assign data_masked[7409] = data_i[7409] & sel_one_hot_i[57];
  assign data_masked[7408] = data_i[7408] & sel_one_hot_i[57];
  assign data_masked[7407] = data_i[7407] & sel_one_hot_i[57];
  assign data_masked[7406] = data_i[7406] & sel_one_hot_i[57];
  assign data_masked[7405] = data_i[7405] & sel_one_hot_i[57];
  assign data_masked[7404] = data_i[7404] & sel_one_hot_i[57];
  assign data_masked[7403] = data_i[7403] & sel_one_hot_i[57];
  assign data_masked[7402] = data_i[7402] & sel_one_hot_i[57];
  assign data_masked[7401] = data_i[7401] & sel_one_hot_i[57];
  assign data_masked[7400] = data_i[7400] & sel_one_hot_i[57];
  assign data_masked[7399] = data_i[7399] & sel_one_hot_i[57];
  assign data_masked[7398] = data_i[7398] & sel_one_hot_i[57];
  assign data_masked[7397] = data_i[7397] & sel_one_hot_i[57];
  assign data_masked[7396] = data_i[7396] & sel_one_hot_i[57];
  assign data_masked[7395] = data_i[7395] & sel_one_hot_i[57];
  assign data_masked[7394] = data_i[7394] & sel_one_hot_i[57];
  assign data_masked[7393] = data_i[7393] & sel_one_hot_i[57];
  assign data_masked[7392] = data_i[7392] & sel_one_hot_i[57];
  assign data_masked[7391] = data_i[7391] & sel_one_hot_i[57];
  assign data_masked[7390] = data_i[7390] & sel_one_hot_i[57];
  assign data_masked[7389] = data_i[7389] & sel_one_hot_i[57];
  assign data_masked[7388] = data_i[7388] & sel_one_hot_i[57];
  assign data_masked[7387] = data_i[7387] & sel_one_hot_i[57];
  assign data_masked[7386] = data_i[7386] & sel_one_hot_i[57];
  assign data_masked[7385] = data_i[7385] & sel_one_hot_i[57];
  assign data_masked[7384] = data_i[7384] & sel_one_hot_i[57];
  assign data_masked[7383] = data_i[7383] & sel_one_hot_i[57];
  assign data_masked[7382] = data_i[7382] & sel_one_hot_i[57];
  assign data_masked[7381] = data_i[7381] & sel_one_hot_i[57];
  assign data_masked[7380] = data_i[7380] & sel_one_hot_i[57];
  assign data_masked[7379] = data_i[7379] & sel_one_hot_i[57];
  assign data_masked[7378] = data_i[7378] & sel_one_hot_i[57];
  assign data_masked[7377] = data_i[7377] & sel_one_hot_i[57];
  assign data_masked[7376] = data_i[7376] & sel_one_hot_i[57];
  assign data_masked[7375] = data_i[7375] & sel_one_hot_i[57];
  assign data_masked[7374] = data_i[7374] & sel_one_hot_i[57];
  assign data_masked[7373] = data_i[7373] & sel_one_hot_i[57];
  assign data_masked[7372] = data_i[7372] & sel_one_hot_i[57];
  assign data_masked[7371] = data_i[7371] & sel_one_hot_i[57];
  assign data_masked[7370] = data_i[7370] & sel_one_hot_i[57];
  assign data_masked[7369] = data_i[7369] & sel_one_hot_i[57];
  assign data_masked[7368] = data_i[7368] & sel_one_hot_i[57];
  assign data_masked[7367] = data_i[7367] & sel_one_hot_i[57];
  assign data_masked[7366] = data_i[7366] & sel_one_hot_i[57];
  assign data_masked[7365] = data_i[7365] & sel_one_hot_i[57];
  assign data_masked[7364] = data_i[7364] & sel_one_hot_i[57];
  assign data_masked[7363] = data_i[7363] & sel_one_hot_i[57];
  assign data_masked[7362] = data_i[7362] & sel_one_hot_i[57];
  assign data_masked[7361] = data_i[7361] & sel_one_hot_i[57];
  assign data_masked[7360] = data_i[7360] & sel_one_hot_i[57];
  assign data_masked[7359] = data_i[7359] & sel_one_hot_i[57];
  assign data_masked[7358] = data_i[7358] & sel_one_hot_i[57];
  assign data_masked[7357] = data_i[7357] & sel_one_hot_i[57];
  assign data_masked[7356] = data_i[7356] & sel_one_hot_i[57];
  assign data_masked[7355] = data_i[7355] & sel_one_hot_i[57];
  assign data_masked[7354] = data_i[7354] & sel_one_hot_i[57];
  assign data_masked[7353] = data_i[7353] & sel_one_hot_i[57];
  assign data_masked[7352] = data_i[7352] & sel_one_hot_i[57];
  assign data_masked[7351] = data_i[7351] & sel_one_hot_i[57];
  assign data_masked[7350] = data_i[7350] & sel_one_hot_i[57];
  assign data_masked[7349] = data_i[7349] & sel_one_hot_i[57];
  assign data_masked[7348] = data_i[7348] & sel_one_hot_i[57];
  assign data_masked[7347] = data_i[7347] & sel_one_hot_i[57];
  assign data_masked[7346] = data_i[7346] & sel_one_hot_i[57];
  assign data_masked[7345] = data_i[7345] & sel_one_hot_i[57];
  assign data_masked[7344] = data_i[7344] & sel_one_hot_i[57];
  assign data_masked[7343] = data_i[7343] & sel_one_hot_i[57];
  assign data_masked[7342] = data_i[7342] & sel_one_hot_i[57];
  assign data_masked[7341] = data_i[7341] & sel_one_hot_i[57];
  assign data_masked[7340] = data_i[7340] & sel_one_hot_i[57];
  assign data_masked[7339] = data_i[7339] & sel_one_hot_i[57];
  assign data_masked[7338] = data_i[7338] & sel_one_hot_i[57];
  assign data_masked[7337] = data_i[7337] & sel_one_hot_i[57];
  assign data_masked[7336] = data_i[7336] & sel_one_hot_i[57];
  assign data_masked[7335] = data_i[7335] & sel_one_hot_i[57];
  assign data_masked[7334] = data_i[7334] & sel_one_hot_i[57];
  assign data_masked[7333] = data_i[7333] & sel_one_hot_i[57];
  assign data_masked[7332] = data_i[7332] & sel_one_hot_i[57];
  assign data_masked[7331] = data_i[7331] & sel_one_hot_i[57];
  assign data_masked[7330] = data_i[7330] & sel_one_hot_i[57];
  assign data_masked[7329] = data_i[7329] & sel_one_hot_i[57];
  assign data_masked[7328] = data_i[7328] & sel_one_hot_i[57];
  assign data_masked[7327] = data_i[7327] & sel_one_hot_i[57];
  assign data_masked[7326] = data_i[7326] & sel_one_hot_i[57];
  assign data_masked[7325] = data_i[7325] & sel_one_hot_i[57];
  assign data_masked[7324] = data_i[7324] & sel_one_hot_i[57];
  assign data_masked[7323] = data_i[7323] & sel_one_hot_i[57];
  assign data_masked[7322] = data_i[7322] & sel_one_hot_i[57];
  assign data_masked[7321] = data_i[7321] & sel_one_hot_i[57];
  assign data_masked[7320] = data_i[7320] & sel_one_hot_i[57];
  assign data_masked[7319] = data_i[7319] & sel_one_hot_i[57];
  assign data_masked[7318] = data_i[7318] & sel_one_hot_i[57];
  assign data_masked[7317] = data_i[7317] & sel_one_hot_i[57];
  assign data_masked[7316] = data_i[7316] & sel_one_hot_i[57];
  assign data_masked[7315] = data_i[7315] & sel_one_hot_i[57];
  assign data_masked[7314] = data_i[7314] & sel_one_hot_i[57];
  assign data_masked[7313] = data_i[7313] & sel_one_hot_i[57];
  assign data_masked[7312] = data_i[7312] & sel_one_hot_i[57];
  assign data_masked[7311] = data_i[7311] & sel_one_hot_i[57];
  assign data_masked[7310] = data_i[7310] & sel_one_hot_i[57];
  assign data_masked[7309] = data_i[7309] & sel_one_hot_i[57];
  assign data_masked[7308] = data_i[7308] & sel_one_hot_i[57];
  assign data_masked[7307] = data_i[7307] & sel_one_hot_i[57];
  assign data_masked[7306] = data_i[7306] & sel_one_hot_i[57];
  assign data_masked[7305] = data_i[7305] & sel_one_hot_i[57];
  assign data_masked[7304] = data_i[7304] & sel_one_hot_i[57];
  assign data_masked[7303] = data_i[7303] & sel_one_hot_i[57];
  assign data_masked[7302] = data_i[7302] & sel_one_hot_i[57];
  assign data_masked[7301] = data_i[7301] & sel_one_hot_i[57];
  assign data_masked[7300] = data_i[7300] & sel_one_hot_i[57];
  assign data_masked[7299] = data_i[7299] & sel_one_hot_i[57];
  assign data_masked[7298] = data_i[7298] & sel_one_hot_i[57];
  assign data_masked[7297] = data_i[7297] & sel_one_hot_i[57];
  assign data_masked[7296] = data_i[7296] & sel_one_hot_i[57];
  assign data_masked[7551] = data_i[7551] & sel_one_hot_i[58];
  assign data_masked[7550] = data_i[7550] & sel_one_hot_i[58];
  assign data_masked[7549] = data_i[7549] & sel_one_hot_i[58];
  assign data_masked[7548] = data_i[7548] & sel_one_hot_i[58];
  assign data_masked[7547] = data_i[7547] & sel_one_hot_i[58];
  assign data_masked[7546] = data_i[7546] & sel_one_hot_i[58];
  assign data_masked[7545] = data_i[7545] & sel_one_hot_i[58];
  assign data_masked[7544] = data_i[7544] & sel_one_hot_i[58];
  assign data_masked[7543] = data_i[7543] & sel_one_hot_i[58];
  assign data_masked[7542] = data_i[7542] & sel_one_hot_i[58];
  assign data_masked[7541] = data_i[7541] & sel_one_hot_i[58];
  assign data_masked[7540] = data_i[7540] & sel_one_hot_i[58];
  assign data_masked[7539] = data_i[7539] & sel_one_hot_i[58];
  assign data_masked[7538] = data_i[7538] & sel_one_hot_i[58];
  assign data_masked[7537] = data_i[7537] & sel_one_hot_i[58];
  assign data_masked[7536] = data_i[7536] & sel_one_hot_i[58];
  assign data_masked[7535] = data_i[7535] & sel_one_hot_i[58];
  assign data_masked[7534] = data_i[7534] & sel_one_hot_i[58];
  assign data_masked[7533] = data_i[7533] & sel_one_hot_i[58];
  assign data_masked[7532] = data_i[7532] & sel_one_hot_i[58];
  assign data_masked[7531] = data_i[7531] & sel_one_hot_i[58];
  assign data_masked[7530] = data_i[7530] & sel_one_hot_i[58];
  assign data_masked[7529] = data_i[7529] & sel_one_hot_i[58];
  assign data_masked[7528] = data_i[7528] & sel_one_hot_i[58];
  assign data_masked[7527] = data_i[7527] & sel_one_hot_i[58];
  assign data_masked[7526] = data_i[7526] & sel_one_hot_i[58];
  assign data_masked[7525] = data_i[7525] & sel_one_hot_i[58];
  assign data_masked[7524] = data_i[7524] & sel_one_hot_i[58];
  assign data_masked[7523] = data_i[7523] & sel_one_hot_i[58];
  assign data_masked[7522] = data_i[7522] & sel_one_hot_i[58];
  assign data_masked[7521] = data_i[7521] & sel_one_hot_i[58];
  assign data_masked[7520] = data_i[7520] & sel_one_hot_i[58];
  assign data_masked[7519] = data_i[7519] & sel_one_hot_i[58];
  assign data_masked[7518] = data_i[7518] & sel_one_hot_i[58];
  assign data_masked[7517] = data_i[7517] & sel_one_hot_i[58];
  assign data_masked[7516] = data_i[7516] & sel_one_hot_i[58];
  assign data_masked[7515] = data_i[7515] & sel_one_hot_i[58];
  assign data_masked[7514] = data_i[7514] & sel_one_hot_i[58];
  assign data_masked[7513] = data_i[7513] & sel_one_hot_i[58];
  assign data_masked[7512] = data_i[7512] & sel_one_hot_i[58];
  assign data_masked[7511] = data_i[7511] & sel_one_hot_i[58];
  assign data_masked[7510] = data_i[7510] & sel_one_hot_i[58];
  assign data_masked[7509] = data_i[7509] & sel_one_hot_i[58];
  assign data_masked[7508] = data_i[7508] & sel_one_hot_i[58];
  assign data_masked[7507] = data_i[7507] & sel_one_hot_i[58];
  assign data_masked[7506] = data_i[7506] & sel_one_hot_i[58];
  assign data_masked[7505] = data_i[7505] & sel_one_hot_i[58];
  assign data_masked[7504] = data_i[7504] & sel_one_hot_i[58];
  assign data_masked[7503] = data_i[7503] & sel_one_hot_i[58];
  assign data_masked[7502] = data_i[7502] & sel_one_hot_i[58];
  assign data_masked[7501] = data_i[7501] & sel_one_hot_i[58];
  assign data_masked[7500] = data_i[7500] & sel_one_hot_i[58];
  assign data_masked[7499] = data_i[7499] & sel_one_hot_i[58];
  assign data_masked[7498] = data_i[7498] & sel_one_hot_i[58];
  assign data_masked[7497] = data_i[7497] & sel_one_hot_i[58];
  assign data_masked[7496] = data_i[7496] & sel_one_hot_i[58];
  assign data_masked[7495] = data_i[7495] & sel_one_hot_i[58];
  assign data_masked[7494] = data_i[7494] & sel_one_hot_i[58];
  assign data_masked[7493] = data_i[7493] & sel_one_hot_i[58];
  assign data_masked[7492] = data_i[7492] & sel_one_hot_i[58];
  assign data_masked[7491] = data_i[7491] & sel_one_hot_i[58];
  assign data_masked[7490] = data_i[7490] & sel_one_hot_i[58];
  assign data_masked[7489] = data_i[7489] & sel_one_hot_i[58];
  assign data_masked[7488] = data_i[7488] & sel_one_hot_i[58];
  assign data_masked[7487] = data_i[7487] & sel_one_hot_i[58];
  assign data_masked[7486] = data_i[7486] & sel_one_hot_i[58];
  assign data_masked[7485] = data_i[7485] & sel_one_hot_i[58];
  assign data_masked[7484] = data_i[7484] & sel_one_hot_i[58];
  assign data_masked[7483] = data_i[7483] & sel_one_hot_i[58];
  assign data_masked[7482] = data_i[7482] & sel_one_hot_i[58];
  assign data_masked[7481] = data_i[7481] & sel_one_hot_i[58];
  assign data_masked[7480] = data_i[7480] & sel_one_hot_i[58];
  assign data_masked[7479] = data_i[7479] & sel_one_hot_i[58];
  assign data_masked[7478] = data_i[7478] & sel_one_hot_i[58];
  assign data_masked[7477] = data_i[7477] & sel_one_hot_i[58];
  assign data_masked[7476] = data_i[7476] & sel_one_hot_i[58];
  assign data_masked[7475] = data_i[7475] & sel_one_hot_i[58];
  assign data_masked[7474] = data_i[7474] & sel_one_hot_i[58];
  assign data_masked[7473] = data_i[7473] & sel_one_hot_i[58];
  assign data_masked[7472] = data_i[7472] & sel_one_hot_i[58];
  assign data_masked[7471] = data_i[7471] & sel_one_hot_i[58];
  assign data_masked[7470] = data_i[7470] & sel_one_hot_i[58];
  assign data_masked[7469] = data_i[7469] & sel_one_hot_i[58];
  assign data_masked[7468] = data_i[7468] & sel_one_hot_i[58];
  assign data_masked[7467] = data_i[7467] & sel_one_hot_i[58];
  assign data_masked[7466] = data_i[7466] & sel_one_hot_i[58];
  assign data_masked[7465] = data_i[7465] & sel_one_hot_i[58];
  assign data_masked[7464] = data_i[7464] & sel_one_hot_i[58];
  assign data_masked[7463] = data_i[7463] & sel_one_hot_i[58];
  assign data_masked[7462] = data_i[7462] & sel_one_hot_i[58];
  assign data_masked[7461] = data_i[7461] & sel_one_hot_i[58];
  assign data_masked[7460] = data_i[7460] & sel_one_hot_i[58];
  assign data_masked[7459] = data_i[7459] & sel_one_hot_i[58];
  assign data_masked[7458] = data_i[7458] & sel_one_hot_i[58];
  assign data_masked[7457] = data_i[7457] & sel_one_hot_i[58];
  assign data_masked[7456] = data_i[7456] & sel_one_hot_i[58];
  assign data_masked[7455] = data_i[7455] & sel_one_hot_i[58];
  assign data_masked[7454] = data_i[7454] & sel_one_hot_i[58];
  assign data_masked[7453] = data_i[7453] & sel_one_hot_i[58];
  assign data_masked[7452] = data_i[7452] & sel_one_hot_i[58];
  assign data_masked[7451] = data_i[7451] & sel_one_hot_i[58];
  assign data_masked[7450] = data_i[7450] & sel_one_hot_i[58];
  assign data_masked[7449] = data_i[7449] & sel_one_hot_i[58];
  assign data_masked[7448] = data_i[7448] & sel_one_hot_i[58];
  assign data_masked[7447] = data_i[7447] & sel_one_hot_i[58];
  assign data_masked[7446] = data_i[7446] & sel_one_hot_i[58];
  assign data_masked[7445] = data_i[7445] & sel_one_hot_i[58];
  assign data_masked[7444] = data_i[7444] & sel_one_hot_i[58];
  assign data_masked[7443] = data_i[7443] & sel_one_hot_i[58];
  assign data_masked[7442] = data_i[7442] & sel_one_hot_i[58];
  assign data_masked[7441] = data_i[7441] & sel_one_hot_i[58];
  assign data_masked[7440] = data_i[7440] & sel_one_hot_i[58];
  assign data_masked[7439] = data_i[7439] & sel_one_hot_i[58];
  assign data_masked[7438] = data_i[7438] & sel_one_hot_i[58];
  assign data_masked[7437] = data_i[7437] & sel_one_hot_i[58];
  assign data_masked[7436] = data_i[7436] & sel_one_hot_i[58];
  assign data_masked[7435] = data_i[7435] & sel_one_hot_i[58];
  assign data_masked[7434] = data_i[7434] & sel_one_hot_i[58];
  assign data_masked[7433] = data_i[7433] & sel_one_hot_i[58];
  assign data_masked[7432] = data_i[7432] & sel_one_hot_i[58];
  assign data_masked[7431] = data_i[7431] & sel_one_hot_i[58];
  assign data_masked[7430] = data_i[7430] & sel_one_hot_i[58];
  assign data_masked[7429] = data_i[7429] & sel_one_hot_i[58];
  assign data_masked[7428] = data_i[7428] & sel_one_hot_i[58];
  assign data_masked[7427] = data_i[7427] & sel_one_hot_i[58];
  assign data_masked[7426] = data_i[7426] & sel_one_hot_i[58];
  assign data_masked[7425] = data_i[7425] & sel_one_hot_i[58];
  assign data_masked[7424] = data_i[7424] & sel_one_hot_i[58];
  assign data_masked[7679] = data_i[7679] & sel_one_hot_i[59];
  assign data_masked[7678] = data_i[7678] & sel_one_hot_i[59];
  assign data_masked[7677] = data_i[7677] & sel_one_hot_i[59];
  assign data_masked[7676] = data_i[7676] & sel_one_hot_i[59];
  assign data_masked[7675] = data_i[7675] & sel_one_hot_i[59];
  assign data_masked[7674] = data_i[7674] & sel_one_hot_i[59];
  assign data_masked[7673] = data_i[7673] & sel_one_hot_i[59];
  assign data_masked[7672] = data_i[7672] & sel_one_hot_i[59];
  assign data_masked[7671] = data_i[7671] & sel_one_hot_i[59];
  assign data_masked[7670] = data_i[7670] & sel_one_hot_i[59];
  assign data_masked[7669] = data_i[7669] & sel_one_hot_i[59];
  assign data_masked[7668] = data_i[7668] & sel_one_hot_i[59];
  assign data_masked[7667] = data_i[7667] & sel_one_hot_i[59];
  assign data_masked[7666] = data_i[7666] & sel_one_hot_i[59];
  assign data_masked[7665] = data_i[7665] & sel_one_hot_i[59];
  assign data_masked[7664] = data_i[7664] & sel_one_hot_i[59];
  assign data_masked[7663] = data_i[7663] & sel_one_hot_i[59];
  assign data_masked[7662] = data_i[7662] & sel_one_hot_i[59];
  assign data_masked[7661] = data_i[7661] & sel_one_hot_i[59];
  assign data_masked[7660] = data_i[7660] & sel_one_hot_i[59];
  assign data_masked[7659] = data_i[7659] & sel_one_hot_i[59];
  assign data_masked[7658] = data_i[7658] & sel_one_hot_i[59];
  assign data_masked[7657] = data_i[7657] & sel_one_hot_i[59];
  assign data_masked[7656] = data_i[7656] & sel_one_hot_i[59];
  assign data_masked[7655] = data_i[7655] & sel_one_hot_i[59];
  assign data_masked[7654] = data_i[7654] & sel_one_hot_i[59];
  assign data_masked[7653] = data_i[7653] & sel_one_hot_i[59];
  assign data_masked[7652] = data_i[7652] & sel_one_hot_i[59];
  assign data_masked[7651] = data_i[7651] & sel_one_hot_i[59];
  assign data_masked[7650] = data_i[7650] & sel_one_hot_i[59];
  assign data_masked[7649] = data_i[7649] & sel_one_hot_i[59];
  assign data_masked[7648] = data_i[7648] & sel_one_hot_i[59];
  assign data_masked[7647] = data_i[7647] & sel_one_hot_i[59];
  assign data_masked[7646] = data_i[7646] & sel_one_hot_i[59];
  assign data_masked[7645] = data_i[7645] & sel_one_hot_i[59];
  assign data_masked[7644] = data_i[7644] & sel_one_hot_i[59];
  assign data_masked[7643] = data_i[7643] & sel_one_hot_i[59];
  assign data_masked[7642] = data_i[7642] & sel_one_hot_i[59];
  assign data_masked[7641] = data_i[7641] & sel_one_hot_i[59];
  assign data_masked[7640] = data_i[7640] & sel_one_hot_i[59];
  assign data_masked[7639] = data_i[7639] & sel_one_hot_i[59];
  assign data_masked[7638] = data_i[7638] & sel_one_hot_i[59];
  assign data_masked[7637] = data_i[7637] & sel_one_hot_i[59];
  assign data_masked[7636] = data_i[7636] & sel_one_hot_i[59];
  assign data_masked[7635] = data_i[7635] & sel_one_hot_i[59];
  assign data_masked[7634] = data_i[7634] & sel_one_hot_i[59];
  assign data_masked[7633] = data_i[7633] & sel_one_hot_i[59];
  assign data_masked[7632] = data_i[7632] & sel_one_hot_i[59];
  assign data_masked[7631] = data_i[7631] & sel_one_hot_i[59];
  assign data_masked[7630] = data_i[7630] & sel_one_hot_i[59];
  assign data_masked[7629] = data_i[7629] & sel_one_hot_i[59];
  assign data_masked[7628] = data_i[7628] & sel_one_hot_i[59];
  assign data_masked[7627] = data_i[7627] & sel_one_hot_i[59];
  assign data_masked[7626] = data_i[7626] & sel_one_hot_i[59];
  assign data_masked[7625] = data_i[7625] & sel_one_hot_i[59];
  assign data_masked[7624] = data_i[7624] & sel_one_hot_i[59];
  assign data_masked[7623] = data_i[7623] & sel_one_hot_i[59];
  assign data_masked[7622] = data_i[7622] & sel_one_hot_i[59];
  assign data_masked[7621] = data_i[7621] & sel_one_hot_i[59];
  assign data_masked[7620] = data_i[7620] & sel_one_hot_i[59];
  assign data_masked[7619] = data_i[7619] & sel_one_hot_i[59];
  assign data_masked[7618] = data_i[7618] & sel_one_hot_i[59];
  assign data_masked[7617] = data_i[7617] & sel_one_hot_i[59];
  assign data_masked[7616] = data_i[7616] & sel_one_hot_i[59];
  assign data_masked[7615] = data_i[7615] & sel_one_hot_i[59];
  assign data_masked[7614] = data_i[7614] & sel_one_hot_i[59];
  assign data_masked[7613] = data_i[7613] & sel_one_hot_i[59];
  assign data_masked[7612] = data_i[7612] & sel_one_hot_i[59];
  assign data_masked[7611] = data_i[7611] & sel_one_hot_i[59];
  assign data_masked[7610] = data_i[7610] & sel_one_hot_i[59];
  assign data_masked[7609] = data_i[7609] & sel_one_hot_i[59];
  assign data_masked[7608] = data_i[7608] & sel_one_hot_i[59];
  assign data_masked[7607] = data_i[7607] & sel_one_hot_i[59];
  assign data_masked[7606] = data_i[7606] & sel_one_hot_i[59];
  assign data_masked[7605] = data_i[7605] & sel_one_hot_i[59];
  assign data_masked[7604] = data_i[7604] & sel_one_hot_i[59];
  assign data_masked[7603] = data_i[7603] & sel_one_hot_i[59];
  assign data_masked[7602] = data_i[7602] & sel_one_hot_i[59];
  assign data_masked[7601] = data_i[7601] & sel_one_hot_i[59];
  assign data_masked[7600] = data_i[7600] & sel_one_hot_i[59];
  assign data_masked[7599] = data_i[7599] & sel_one_hot_i[59];
  assign data_masked[7598] = data_i[7598] & sel_one_hot_i[59];
  assign data_masked[7597] = data_i[7597] & sel_one_hot_i[59];
  assign data_masked[7596] = data_i[7596] & sel_one_hot_i[59];
  assign data_masked[7595] = data_i[7595] & sel_one_hot_i[59];
  assign data_masked[7594] = data_i[7594] & sel_one_hot_i[59];
  assign data_masked[7593] = data_i[7593] & sel_one_hot_i[59];
  assign data_masked[7592] = data_i[7592] & sel_one_hot_i[59];
  assign data_masked[7591] = data_i[7591] & sel_one_hot_i[59];
  assign data_masked[7590] = data_i[7590] & sel_one_hot_i[59];
  assign data_masked[7589] = data_i[7589] & sel_one_hot_i[59];
  assign data_masked[7588] = data_i[7588] & sel_one_hot_i[59];
  assign data_masked[7587] = data_i[7587] & sel_one_hot_i[59];
  assign data_masked[7586] = data_i[7586] & sel_one_hot_i[59];
  assign data_masked[7585] = data_i[7585] & sel_one_hot_i[59];
  assign data_masked[7584] = data_i[7584] & sel_one_hot_i[59];
  assign data_masked[7583] = data_i[7583] & sel_one_hot_i[59];
  assign data_masked[7582] = data_i[7582] & sel_one_hot_i[59];
  assign data_masked[7581] = data_i[7581] & sel_one_hot_i[59];
  assign data_masked[7580] = data_i[7580] & sel_one_hot_i[59];
  assign data_masked[7579] = data_i[7579] & sel_one_hot_i[59];
  assign data_masked[7578] = data_i[7578] & sel_one_hot_i[59];
  assign data_masked[7577] = data_i[7577] & sel_one_hot_i[59];
  assign data_masked[7576] = data_i[7576] & sel_one_hot_i[59];
  assign data_masked[7575] = data_i[7575] & sel_one_hot_i[59];
  assign data_masked[7574] = data_i[7574] & sel_one_hot_i[59];
  assign data_masked[7573] = data_i[7573] & sel_one_hot_i[59];
  assign data_masked[7572] = data_i[7572] & sel_one_hot_i[59];
  assign data_masked[7571] = data_i[7571] & sel_one_hot_i[59];
  assign data_masked[7570] = data_i[7570] & sel_one_hot_i[59];
  assign data_masked[7569] = data_i[7569] & sel_one_hot_i[59];
  assign data_masked[7568] = data_i[7568] & sel_one_hot_i[59];
  assign data_masked[7567] = data_i[7567] & sel_one_hot_i[59];
  assign data_masked[7566] = data_i[7566] & sel_one_hot_i[59];
  assign data_masked[7565] = data_i[7565] & sel_one_hot_i[59];
  assign data_masked[7564] = data_i[7564] & sel_one_hot_i[59];
  assign data_masked[7563] = data_i[7563] & sel_one_hot_i[59];
  assign data_masked[7562] = data_i[7562] & sel_one_hot_i[59];
  assign data_masked[7561] = data_i[7561] & sel_one_hot_i[59];
  assign data_masked[7560] = data_i[7560] & sel_one_hot_i[59];
  assign data_masked[7559] = data_i[7559] & sel_one_hot_i[59];
  assign data_masked[7558] = data_i[7558] & sel_one_hot_i[59];
  assign data_masked[7557] = data_i[7557] & sel_one_hot_i[59];
  assign data_masked[7556] = data_i[7556] & sel_one_hot_i[59];
  assign data_masked[7555] = data_i[7555] & sel_one_hot_i[59];
  assign data_masked[7554] = data_i[7554] & sel_one_hot_i[59];
  assign data_masked[7553] = data_i[7553] & sel_one_hot_i[59];
  assign data_masked[7552] = data_i[7552] & sel_one_hot_i[59];
  assign data_masked[7807] = data_i[7807] & sel_one_hot_i[60];
  assign data_masked[7806] = data_i[7806] & sel_one_hot_i[60];
  assign data_masked[7805] = data_i[7805] & sel_one_hot_i[60];
  assign data_masked[7804] = data_i[7804] & sel_one_hot_i[60];
  assign data_masked[7803] = data_i[7803] & sel_one_hot_i[60];
  assign data_masked[7802] = data_i[7802] & sel_one_hot_i[60];
  assign data_masked[7801] = data_i[7801] & sel_one_hot_i[60];
  assign data_masked[7800] = data_i[7800] & sel_one_hot_i[60];
  assign data_masked[7799] = data_i[7799] & sel_one_hot_i[60];
  assign data_masked[7798] = data_i[7798] & sel_one_hot_i[60];
  assign data_masked[7797] = data_i[7797] & sel_one_hot_i[60];
  assign data_masked[7796] = data_i[7796] & sel_one_hot_i[60];
  assign data_masked[7795] = data_i[7795] & sel_one_hot_i[60];
  assign data_masked[7794] = data_i[7794] & sel_one_hot_i[60];
  assign data_masked[7793] = data_i[7793] & sel_one_hot_i[60];
  assign data_masked[7792] = data_i[7792] & sel_one_hot_i[60];
  assign data_masked[7791] = data_i[7791] & sel_one_hot_i[60];
  assign data_masked[7790] = data_i[7790] & sel_one_hot_i[60];
  assign data_masked[7789] = data_i[7789] & sel_one_hot_i[60];
  assign data_masked[7788] = data_i[7788] & sel_one_hot_i[60];
  assign data_masked[7787] = data_i[7787] & sel_one_hot_i[60];
  assign data_masked[7786] = data_i[7786] & sel_one_hot_i[60];
  assign data_masked[7785] = data_i[7785] & sel_one_hot_i[60];
  assign data_masked[7784] = data_i[7784] & sel_one_hot_i[60];
  assign data_masked[7783] = data_i[7783] & sel_one_hot_i[60];
  assign data_masked[7782] = data_i[7782] & sel_one_hot_i[60];
  assign data_masked[7781] = data_i[7781] & sel_one_hot_i[60];
  assign data_masked[7780] = data_i[7780] & sel_one_hot_i[60];
  assign data_masked[7779] = data_i[7779] & sel_one_hot_i[60];
  assign data_masked[7778] = data_i[7778] & sel_one_hot_i[60];
  assign data_masked[7777] = data_i[7777] & sel_one_hot_i[60];
  assign data_masked[7776] = data_i[7776] & sel_one_hot_i[60];
  assign data_masked[7775] = data_i[7775] & sel_one_hot_i[60];
  assign data_masked[7774] = data_i[7774] & sel_one_hot_i[60];
  assign data_masked[7773] = data_i[7773] & sel_one_hot_i[60];
  assign data_masked[7772] = data_i[7772] & sel_one_hot_i[60];
  assign data_masked[7771] = data_i[7771] & sel_one_hot_i[60];
  assign data_masked[7770] = data_i[7770] & sel_one_hot_i[60];
  assign data_masked[7769] = data_i[7769] & sel_one_hot_i[60];
  assign data_masked[7768] = data_i[7768] & sel_one_hot_i[60];
  assign data_masked[7767] = data_i[7767] & sel_one_hot_i[60];
  assign data_masked[7766] = data_i[7766] & sel_one_hot_i[60];
  assign data_masked[7765] = data_i[7765] & sel_one_hot_i[60];
  assign data_masked[7764] = data_i[7764] & sel_one_hot_i[60];
  assign data_masked[7763] = data_i[7763] & sel_one_hot_i[60];
  assign data_masked[7762] = data_i[7762] & sel_one_hot_i[60];
  assign data_masked[7761] = data_i[7761] & sel_one_hot_i[60];
  assign data_masked[7760] = data_i[7760] & sel_one_hot_i[60];
  assign data_masked[7759] = data_i[7759] & sel_one_hot_i[60];
  assign data_masked[7758] = data_i[7758] & sel_one_hot_i[60];
  assign data_masked[7757] = data_i[7757] & sel_one_hot_i[60];
  assign data_masked[7756] = data_i[7756] & sel_one_hot_i[60];
  assign data_masked[7755] = data_i[7755] & sel_one_hot_i[60];
  assign data_masked[7754] = data_i[7754] & sel_one_hot_i[60];
  assign data_masked[7753] = data_i[7753] & sel_one_hot_i[60];
  assign data_masked[7752] = data_i[7752] & sel_one_hot_i[60];
  assign data_masked[7751] = data_i[7751] & sel_one_hot_i[60];
  assign data_masked[7750] = data_i[7750] & sel_one_hot_i[60];
  assign data_masked[7749] = data_i[7749] & sel_one_hot_i[60];
  assign data_masked[7748] = data_i[7748] & sel_one_hot_i[60];
  assign data_masked[7747] = data_i[7747] & sel_one_hot_i[60];
  assign data_masked[7746] = data_i[7746] & sel_one_hot_i[60];
  assign data_masked[7745] = data_i[7745] & sel_one_hot_i[60];
  assign data_masked[7744] = data_i[7744] & sel_one_hot_i[60];
  assign data_masked[7743] = data_i[7743] & sel_one_hot_i[60];
  assign data_masked[7742] = data_i[7742] & sel_one_hot_i[60];
  assign data_masked[7741] = data_i[7741] & sel_one_hot_i[60];
  assign data_masked[7740] = data_i[7740] & sel_one_hot_i[60];
  assign data_masked[7739] = data_i[7739] & sel_one_hot_i[60];
  assign data_masked[7738] = data_i[7738] & sel_one_hot_i[60];
  assign data_masked[7737] = data_i[7737] & sel_one_hot_i[60];
  assign data_masked[7736] = data_i[7736] & sel_one_hot_i[60];
  assign data_masked[7735] = data_i[7735] & sel_one_hot_i[60];
  assign data_masked[7734] = data_i[7734] & sel_one_hot_i[60];
  assign data_masked[7733] = data_i[7733] & sel_one_hot_i[60];
  assign data_masked[7732] = data_i[7732] & sel_one_hot_i[60];
  assign data_masked[7731] = data_i[7731] & sel_one_hot_i[60];
  assign data_masked[7730] = data_i[7730] & sel_one_hot_i[60];
  assign data_masked[7729] = data_i[7729] & sel_one_hot_i[60];
  assign data_masked[7728] = data_i[7728] & sel_one_hot_i[60];
  assign data_masked[7727] = data_i[7727] & sel_one_hot_i[60];
  assign data_masked[7726] = data_i[7726] & sel_one_hot_i[60];
  assign data_masked[7725] = data_i[7725] & sel_one_hot_i[60];
  assign data_masked[7724] = data_i[7724] & sel_one_hot_i[60];
  assign data_masked[7723] = data_i[7723] & sel_one_hot_i[60];
  assign data_masked[7722] = data_i[7722] & sel_one_hot_i[60];
  assign data_masked[7721] = data_i[7721] & sel_one_hot_i[60];
  assign data_masked[7720] = data_i[7720] & sel_one_hot_i[60];
  assign data_masked[7719] = data_i[7719] & sel_one_hot_i[60];
  assign data_masked[7718] = data_i[7718] & sel_one_hot_i[60];
  assign data_masked[7717] = data_i[7717] & sel_one_hot_i[60];
  assign data_masked[7716] = data_i[7716] & sel_one_hot_i[60];
  assign data_masked[7715] = data_i[7715] & sel_one_hot_i[60];
  assign data_masked[7714] = data_i[7714] & sel_one_hot_i[60];
  assign data_masked[7713] = data_i[7713] & sel_one_hot_i[60];
  assign data_masked[7712] = data_i[7712] & sel_one_hot_i[60];
  assign data_masked[7711] = data_i[7711] & sel_one_hot_i[60];
  assign data_masked[7710] = data_i[7710] & sel_one_hot_i[60];
  assign data_masked[7709] = data_i[7709] & sel_one_hot_i[60];
  assign data_masked[7708] = data_i[7708] & sel_one_hot_i[60];
  assign data_masked[7707] = data_i[7707] & sel_one_hot_i[60];
  assign data_masked[7706] = data_i[7706] & sel_one_hot_i[60];
  assign data_masked[7705] = data_i[7705] & sel_one_hot_i[60];
  assign data_masked[7704] = data_i[7704] & sel_one_hot_i[60];
  assign data_masked[7703] = data_i[7703] & sel_one_hot_i[60];
  assign data_masked[7702] = data_i[7702] & sel_one_hot_i[60];
  assign data_masked[7701] = data_i[7701] & sel_one_hot_i[60];
  assign data_masked[7700] = data_i[7700] & sel_one_hot_i[60];
  assign data_masked[7699] = data_i[7699] & sel_one_hot_i[60];
  assign data_masked[7698] = data_i[7698] & sel_one_hot_i[60];
  assign data_masked[7697] = data_i[7697] & sel_one_hot_i[60];
  assign data_masked[7696] = data_i[7696] & sel_one_hot_i[60];
  assign data_masked[7695] = data_i[7695] & sel_one_hot_i[60];
  assign data_masked[7694] = data_i[7694] & sel_one_hot_i[60];
  assign data_masked[7693] = data_i[7693] & sel_one_hot_i[60];
  assign data_masked[7692] = data_i[7692] & sel_one_hot_i[60];
  assign data_masked[7691] = data_i[7691] & sel_one_hot_i[60];
  assign data_masked[7690] = data_i[7690] & sel_one_hot_i[60];
  assign data_masked[7689] = data_i[7689] & sel_one_hot_i[60];
  assign data_masked[7688] = data_i[7688] & sel_one_hot_i[60];
  assign data_masked[7687] = data_i[7687] & sel_one_hot_i[60];
  assign data_masked[7686] = data_i[7686] & sel_one_hot_i[60];
  assign data_masked[7685] = data_i[7685] & sel_one_hot_i[60];
  assign data_masked[7684] = data_i[7684] & sel_one_hot_i[60];
  assign data_masked[7683] = data_i[7683] & sel_one_hot_i[60];
  assign data_masked[7682] = data_i[7682] & sel_one_hot_i[60];
  assign data_masked[7681] = data_i[7681] & sel_one_hot_i[60];
  assign data_masked[7680] = data_i[7680] & sel_one_hot_i[60];
  assign data_masked[7935] = data_i[7935] & sel_one_hot_i[61];
  assign data_masked[7934] = data_i[7934] & sel_one_hot_i[61];
  assign data_masked[7933] = data_i[7933] & sel_one_hot_i[61];
  assign data_masked[7932] = data_i[7932] & sel_one_hot_i[61];
  assign data_masked[7931] = data_i[7931] & sel_one_hot_i[61];
  assign data_masked[7930] = data_i[7930] & sel_one_hot_i[61];
  assign data_masked[7929] = data_i[7929] & sel_one_hot_i[61];
  assign data_masked[7928] = data_i[7928] & sel_one_hot_i[61];
  assign data_masked[7927] = data_i[7927] & sel_one_hot_i[61];
  assign data_masked[7926] = data_i[7926] & sel_one_hot_i[61];
  assign data_masked[7925] = data_i[7925] & sel_one_hot_i[61];
  assign data_masked[7924] = data_i[7924] & sel_one_hot_i[61];
  assign data_masked[7923] = data_i[7923] & sel_one_hot_i[61];
  assign data_masked[7922] = data_i[7922] & sel_one_hot_i[61];
  assign data_masked[7921] = data_i[7921] & sel_one_hot_i[61];
  assign data_masked[7920] = data_i[7920] & sel_one_hot_i[61];
  assign data_masked[7919] = data_i[7919] & sel_one_hot_i[61];
  assign data_masked[7918] = data_i[7918] & sel_one_hot_i[61];
  assign data_masked[7917] = data_i[7917] & sel_one_hot_i[61];
  assign data_masked[7916] = data_i[7916] & sel_one_hot_i[61];
  assign data_masked[7915] = data_i[7915] & sel_one_hot_i[61];
  assign data_masked[7914] = data_i[7914] & sel_one_hot_i[61];
  assign data_masked[7913] = data_i[7913] & sel_one_hot_i[61];
  assign data_masked[7912] = data_i[7912] & sel_one_hot_i[61];
  assign data_masked[7911] = data_i[7911] & sel_one_hot_i[61];
  assign data_masked[7910] = data_i[7910] & sel_one_hot_i[61];
  assign data_masked[7909] = data_i[7909] & sel_one_hot_i[61];
  assign data_masked[7908] = data_i[7908] & sel_one_hot_i[61];
  assign data_masked[7907] = data_i[7907] & sel_one_hot_i[61];
  assign data_masked[7906] = data_i[7906] & sel_one_hot_i[61];
  assign data_masked[7905] = data_i[7905] & sel_one_hot_i[61];
  assign data_masked[7904] = data_i[7904] & sel_one_hot_i[61];
  assign data_masked[7903] = data_i[7903] & sel_one_hot_i[61];
  assign data_masked[7902] = data_i[7902] & sel_one_hot_i[61];
  assign data_masked[7901] = data_i[7901] & sel_one_hot_i[61];
  assign data_masked[7900] = data_i[7900] & sel_one_hot_i[61];
  assign data_masked[7899] = data_i[7899] & sel_one_hot_i[61];
  assign data_masked[7898] = data_i[7898] & sel_one_hot_i[61];
  assign data_masked[7897] = data_i[7897] & sel_one_hot_i[61];
  assign data_masked[7896] = data_i[7896] & sel_one_hot_i[61];
  assign data_masked[7895] = data_i[7895] & sel_one_hot_i[61];
  assign data_masked[7894] = data_i[7894] & sel_one_hot_i[61];
  assign data_masked[7893] = data_i[7893] & sel_one_hot_i[61];
  assign data_masked[7892] = data_i[7892] & sel_one_hot_i[61];
  assign data_masked[7891] = data_i[7891] & sel_one_hot_i[61];
  assign data_masked[7890] = data_i[7890] & sel_one_hot_i[61];
  assign data_masked[7889] = data_i[7889] & sel_one_hot_i[61];
  assign data_masked[7888] = data_i[7888] & sel_one_hot_i[61];
  assign data_masked[7887] = data_i[7887] & sel_one_hot_i[61];
  assign data_masked[7886] = data_i[7886] & sel_one_hot_i[61];
  assign data_masked[7885] = data_i[7885] & sel_one_hot_i[61];
  assign data_masked[7884] = data_i[7884] & sel_one_hot_i[61];
  assign data_masked[7883] = data_i[7883] & sel_one_hot_i[61];
  assign data_masked[7882] = data_i[7882] & sel_one_hot_i[61];
  assign data_masked[7881] = data_i[7881] & sel_one_hot_i[61];
  assign data_masked[7880] = data_i[7880] & sel_one_hot_i[61];
  assign data_masked[7879] = data_i[7879] & sel_one_hot_i[61];
  assign data_masked[7878] = data_i[7878] & sel_one_hot_i[61];
  assign data_masked[7877] = data_i[7877] & sel_one_hot_i[61];
  assign data_masked[7876] = data_i[7876] & sel_one_hot_i[61];
  assign data_masked[7875] = data_i[7875] & sel_one_hot_i[61];
  assign data_masked[7874] = data_i[7874] & sel_one_hot_i[61];
  assign data_masked[7873] = data_i[7873] & sel_one_hot_i[61];
  assign data_masked[7872] = data_i[7872] & sel_one_hot_i[61];
  assign data_masked[7871] = data_i[7871] & sel_one_hot_i[61];
  assign data_masked[7870] = data_i[7870] & sel_one_hot_i[61];
  assign data_masked[7869] = data_i[7869] & sel_one_hot_i[61];
  assign data_masked[7868] = data_i[7868] & sel_one_hot_i[61];
  assign data_masked[7867] = data_i[7867] & sel_one_hot_i[61];
  assign data_masked[7866] = data_i[7866] & sel_one_hot_i[61];
  assign data_masked[7865] = data_i[7865] & sel_one_hot_i[61];
  assign data_masked[7864] = data_i[7864] & sel_one_hot_i[61];
  assign data_masked[7863] = data_i[7863] & sel_one_hot_i[61];
  assign data_masked[7862] = data_i[7862] & sel_one_hot_i[61];
  assign data_masked[7861] = data_i[7861] & sel_one_hot_i[61];
  assign data_masked[7860] = data_i[7860] & sel_one_hot_i[61];
  assign data_masked[7859] = data_i[7859] & sel_one_hot_i[61];
  assign data_masked[7858] = data_i[7858] & sel_one_hot_i[61];
  assign data_masked[7857] = data_i[7857] & sel_one_hot_i[61];
  assign data_masked[7856] = data_i[7856] & sel_one_hot_i[61];
  assign data_masked[7855] = data_i[7855] & sel_one_hot_i[61];
  assign data_masked[7854] = data_i[7854] & sel_one_hot_i[61];
  assign data_masked[7853] = data_i[7853] & sel_one_hot_i[61];
  assign data_masked[7852] = data_i[7852] & sel_one_hot_i[61];
  assign data_masked[7851] = data_i[7851] & sel_one_hot_i[61];
  assign data_masked[7850] = data_i[7850] & sel_one_hot_i[61];
  assign data_masked[7849] = data_i[7849] & sel_one_hot_i[61];
  assign data_masked[7848] = data_i[7848] & sel_one_hot_i[61];
  assign data_masked[7847] = data_i[7847] & sel_one_hot_i[61];
  assign data_masked[7846] = data_i[7846] & sel_one_hot_i[61];
  assign data_masked[7845] = data_i[7845] & sel_one_hot_i[61];
  assign data_masked[7844] = data_i[7844] & sel_one_hot_i[61];
  assign data_masked[7843] = data_i[7843] & sel_one_hot_i[61];
  assign data_masked[7842] = data_i[7842] & sel_one_hot_i[61];
  assign data_masked[7841] = data_i[7841] & sel_one_hot_i[61];
  assign data_masked[7840] = data_i[7840] & sel_one_hot_i[61];
  assign data_masked[7839] = data_i[7839] & sel_one_hot_i[61];
  assign data_masked[7838] = data_i[7838] & sel_one_hot_i[61];
  assign data_masked[7837] = data_i[7837] & sel_one_hot_i[61];
  assign data_masked[7836] = data_i[7836] & sel_one_hot_i[61];
  assign data_masked[7835] = data_i[7835] & sel_one_hot_i[61];
  assign data_masked[7834] = data_i[7834] & sel_one_hot_i[61];
  assign data_masked[7833] = data_i[7833] & sel_one_hot_i[61];
  assign data_masked[7832] = data_i[7832] & sel_one_hot_i[61];
  assign data_masked[7831] = data_i[7831] & sel_one_hot_i[61];
  assign data_masked[7830] = data_i[7830] & sel_one_hot_i[61];
  assign data_masked[7829] = data_i[7829] & sel_one_hot_i[61];
  assign data_masked[7828] = data_i[7828] & sel_one_hot_i[61];
  assign data_masked[7827] = data_i[7827] & sel_one_hot_i[61];
  assign data_masked[7826] = data_i[7826] & sel_one_hot_i[61];
  assign data_masked[7825] = data_i[7825] & sel_one_hot_i[61];
  assign data_masked[7824] = data_i[7824] & sel_one_hot_i[61];
  assign data_masked[7823] = data_i[7823] & sel_one_hot_i[61];
  assign data_masked[7822] = data_i[7822] & sel_one_hot_i[61];
  assign data_masked[7821] = data_i[7821] & sel_one_hot_i[61];
  assign data_masked[7820] = data_i[7820] & sel_one_hot_i[61];
  assign data_masked[7819] = data_i[7819] & sel_one_hot_i[61];
  assign data_masked[7818] = data_i[7818] & sel_one_hot_i[61];
  assign data_masked[7817] = data_i[7817] & sel_one_hot_i[61];
  assign data_masked[7816] = data_i[7816] & sel_one_hot_i[61];
  assign data_masked[7815] = data_i[7815] & sel_one_hot_i[61];
  assign data_masked[7814] = data_i[7814] & sel_one_hot_i[61];
  assign data_masked[7813] = data_i[7813] & sel_one_hot_i[61];
  assign data_masked[7812] = data_i[7812] & sel_one_hot_i[61];
  assign data_masked[7811] = data_i[7811] & sel_one_hot_i[61];
  assign data_masked[7810] = data_i[7810] & sel_one_hot_i[61];
  assign data_masked[7809] = data_i[7809] & sel_one_hot_i[61];
  assign data_masked[7808] = data_i[7808] & sel_one_hot_i[61];
  assign data_masked[8063] = data_i[8063] & sel_one_hot_i[62];
  assign data_masked[8062] = data_i[8062] & sel_one_hot_i[62];
  assign data_masked[8061] = data_i[8061] & sel_one_hot_i[62];
  assign data_masked[8060] = data_i[8060] & sel_one_hot_i[62];
  assign data_masked[8059] = data_i[8059] & sel_one_hot_i[62];
  assign data_masked[8058] = data_i[8058] & sel_one_hot_i[62];
  assign data_masked[8057] = data_i[8057] & sel_one_hot_i[62];
  assign data_masked[8056] = data_i[8056] & sel_one_hot_i[62];
  assign data_masked[8055] = data_i[8055] & sel_one_hot_i[62];
  assign data_masked[8054] = data_i[8054] & sel_one_hot_i[62];
  assign data_masked[8053] = data_i[8053] & sel_one_hot_i[62];
  assign data_masked[8052] = data_i[8052] & sel_one_hot_i[62];
  assign data_masked[8051] = data_i[8051] & sel_one_hot_i[62];
  assign data_masked[8050] = data_i[8050] & sel_one_hot_i[62];
  assign data_masked[8049] = data_i[8049] & sel_one_hot_i[62];
  assign data_masked[8048] = data_i[8048] & sel_one_hot_i[62];
  assign data_masked[8047] = data_i[8047] & sel_one_hot_i[62];
  assign data_masked[8046] = data_i[8046] & sel_one_hot_i[62];
  assign data_masked[8045] = data_i[8045] & sel_one_hot_i[62];
  assign data_masked[8044] = data_i[8044] & sel_one_hot_i[62];
  assign data_masked[8043] = data_i[8043] & sel_one_hot_i[62];
  assign data_masked[8042] = data_i[8042] & sel_one_hot_i[62];
  assign data_masked[8041] = data_i[8041] & sel_one_hot_i[62];
  assign data_masked[8040] = data_i[8040] & sel_one_hot_i[62];
  assign data_masked[8039] = data_i[8039] & sel_one_hot_i[62];
  assign data_masked[8038] = data_i[8038] & sel_one_hot_i[62];
  assign data_masked[8037] = data_i[8037] & sel_one_hot_i[62];
  assign data_masked[8036] = data_i[8036] & sel_one_hot_i[62];
  assign data_masked[8035] = data_i[8035] & sel_one_hot_i[62];
  assign data_masked[8034] = data_i[8034] & sel_one_hot_i[62];
  assign data_masked[8033] = data_i[8033] & sel_one_hot_i[62];
  assign data_masked[8032] = data_i[8032] & sel_one_hot_i[62];
  assign data_masked[8031] = data_i[8031] & sel_one_hot_i[62];
  assign data_masked[8030] = data_i[8030] & sel_one_hot_i[62];
  assign data_masked[8029] = data_i[8029] & sel_one_hot_i[62];
  assign data_masked[8028] = data_i[8028] & sel_one_hot_i[62];
  assign data_masked[8027] = data_i[8027] & sel_one_hot_i[62];
  assign data_masked[8026] = data_i[8026] & sel_one_hot_i[62];
  assign data_masked[8025] = data_i[8025] & sel_one_hot_i[62];
  assign data_masked[8024] = data_i[8024] & sel_one_hot_i[62];
  assign data_masked[8023] = data_i[8023] & sel_one_hot_i[62];
  assign data_masked[8022] = data_i[8022] & sel_one_hot_i[62];
  assign data_masked[8021] = data_i[8021] & sel_one_hot_i[62];
  assign data_masked[8020] = data_i[8020] & sel_one_hot_i[62];
  assign data_masked[8019] = data_i[8019] & sel_one_hot_i[62];
  assign data_masked[8018] = data_i[8018] & sel_one_hot_i[62];
  assign data_masked[8017] = data_i[8017] & sel_one_hot_i[62];
  assign data_masked[8016] = data_i[8016] & sel_one_hot_i[62];
  assign data_masked[8015] = data_i[8015] & sel_one_hot_i[62];
  assign data_masked[8014] = data_i[8014] & sel_one_hot_i[62];
  assign data_masked[8013] = data_i[8013] & sel_one_hot_i[62];
  assign data_masked[8012] = data_i[8012] & sel_one_hot_i[62];
  assign data_masked[8011] = data_i[8011] & sel_one_hot_i[62];
  assign data_masked[8010] = data_i[8010] & sel_one_hot_i[62];
  assign data_masked[8009] = data_i[8009] & sel_one_hot_i[62];
  assign data_masked[8008] = data_i[8008] & sel_one_hot_i[62];
  assign data_masked[8007] = data_i[8007] & sel_one_hot_i[62];
  assign data_masked[8006] = data_i[8006] & sel_one_hot_i[62];
  assign data_masked[8005] = data_i[8005] & sel_one_hot_i[62];
  assign data_masked[8004] = data_i[8004] & sel_one_hot_i[62];
  assign data_masked[8003] = data_i[8003] & sel_one_hot_i[62];
  assign data_masked[8002] = data_i[8002] & sel_one_hot_i[62];
  assign data_masked[8001] = data_i[8001] & sel_one_hot_i[62];
  assign data_masked[8000] = data_i[8000] & sel_one_hot_i[62];
  assign data_masked[7999] = data_i[7999] & sel_one_hot_i[62];
  assign data_masked[7998] = data_i[7998] & sel_one_hot_i[62];
  assign data_masked[7997] = data_i[7997] & sel_one_hot_i[62];
  assign data_masked[7996] = data_i[7996] & sel_one_hot_i[62];
  assign data_masked[7995] = data_i[7995] & sel_one_hot_i[62];
  assign data_masked[7994] = data_i[7994] & sel_one_hot_i[62];
  assign data_masked[7993] = data_i[7993] & sel_one_hot_i[62];
  assign data_masked[7992] = data_i[7992] & sel_one_hot_i[62];
  assign data_masked[7991] = data_i[7991] & sel_one_hot_i[62];
  assign data_masked[7990] = data_i[7990] & sel_one_hot_i[62];
  assign data_masked[7989] = data_i[7989] & sel_one_hot_i[62];
  assign data_masked[7988] = data_i[7988] & sel_one_hot_i[62];
  assign data_masked[7987] = data_i[7987] & sel_one_hot_i[62];
  assign data_masked[7986] = data_i[7986] & sel_one_hot_i[62];
  assign data_masked[7985] = data_i[7985] & sel_one_hot_i[62];
  assign data_masked[7984] = data_i[7984] & sel_one_hot_i[62];
  assign data_masked[7983] = data_i[7983] & sel_one_hot_i[62];
  assign data_masked[7982] = data_i[7982] & sel_one_hot_i[62];
  assign data_masked[7981] = data_i[7981] & sel_one_hot_i[62];
  assign data_masked[7980] = data_i[7980] & sel_one_hot_i[62];
  assign data_masked[7979] = data_i[7979] & sel_one_hot_i[62];
  assign data_masked[7978] = data_i[7978] & sel_one_hot_i[62];
  assign data_masked[7977] = data_i[7977] & sel_one_hot_i[62];
  assign data_masked[7976] = data_i[7976] & sel_one_hot_i[62];
  assign data_masked[7975] = data_i[7975] & sel_one_hot_i[62];
  assign data_masked[7974] = data_i[7974] & sel_one_hot_i[62];
  assign data_masked[7973] = data_i[7973] & sel_one_hot_i[62];
  assign data_masked[7972] = data_i[7972] & sel_one_hot_i[62];
  assign data_masked[7971] = data_i[7971] & sel_one_hot_i[62];
  assign data_masked[7970] = data_i[7970] & sel_one_hot_i[62];
  assign data_masked[7969] = data_i[7969] & sel_one_hot_i[62];
  assign data_masked[7968] = data_i[7968] & sel_one_hot_i[62];
  assign data_masked[7967] = data_i[7967] & sel_one_hot_i[62];
  assign data_masked[7966] = data_i[7966] & sel_one_hot_i[62];
  assign data_masked[7965] = data_i[7965] & sel_one_hot_i[62];
  assign data_masked[7964] = data_i[7964] & sel_one_hot_i[62];
  assign data_masked[7963] = data_i[7963] & sel_one_hot_i[62];
  assign data_masked[7962] = data_i[7962] & sel_one_hot_i[62];
  assign data_masked[7961] = data_i[7961] & sel_one_hot_i[62];
  assign data_masked[7960] = data_i[7960] & sel_one_hot_i[62];
  assign data_masked[7959] = data_i[7959] & sel_one_hot_i[62];
  assign data_masked[7958] = data_i[7958] & sel_one_hot_i[62];
  assign data_masked[7957] = data_i[7957] & sel_one_hot_i[62];
  assign data_masked[7956] = data_i[7956] & sel_one_hot_i[62];
  assign data_masked[7955] = data_i[7955] & sel_one_hot_i[62];
  assign data_masked[7954] = data_i[7954] & sel_one_hot_i[62];
  assign data_masked[7953] = data_i[7953] & sel_one_hot_i[62];
  assign data_masked[7952] = data_i[7952] & sel_one_hot_i[62];
  assign data_masked[7951] = data_i[7951] & sel_one_hot_i[62];
  assign data_masked[7950] = data_i[7950] & sel_one_hot_i[62];
  assign data_masked[7949] = data_i[7949] & sel_one_hot_i[62];
  assign data_masked[7948] = data_i[7948] & sel_one_hot_i[62];
  assign data_masked[7947] = data_i[7947] & sel_one_hot_i[62];
  assign data_masked[7946] = data_i[7946] & sel_one_hot_i[62];
  assign data_masked[7945] = data_i[7945] & sel_one_hot_i[62];
  assign data_masked[7944] = data_i[7944] & sel_one_hot_i[62];
  assign data_masked[7943] = data_i[7943] & sel_one_hot_i[62];
  assign data_masked[7942] = data_i[7942] & sel_one_hot_i[62];
  assign data_masked[7941] = data_i[7941] & sel_one_hot_i[62];
  assign data_masked[7940] = data_i[7940] & sel_one_hot_i[62];
  assign data_masked[7939] = data_i[7939] & sel_one_hot_i[62];
  assign data_masked[7938] = data_i[7938] & sel_one_hot_i[62];
  assign data_masked[7937] = data_i[7937] & sel_one_hot_i[62];
  assign data_masked[7936] = data_i[7936] & sel_one_hot_i[62];
  assign data_masked[8191] = data_i[8191] & sel_one_hot_i[63];
  assign data_masked[8190] = data_i[8190] & sel_one_hot_i[63];
  assign data_masked[8189] = data_i[8189] & sel_one_hot_i[63];
  assign data_masked[8188] = data_i[8188] & sel_one_hot_i[63];
  assign data_masked[8187] = data_i[8187] & sel_one_hot_i[63];
  assign data_masked[8186] = data_i[8186] & sel_one_hot_i[63];
  assign data_masked[8185] = data_i[8185] & sel_one_hot_i[63];
  assign data_masked[8184] = data_i[8184] & sel_one_hot_i[63];
  assign data_masked[8183] = data_i[8183] & sel_one_hot_i[63];
  assign data_masked[8182] = data_i[8182] & sel_one_hot_i[63];
  assign data_masked[8181] = data_i[8181] & sel_one_hot_i[63];
  assign data_masked[8180] = data_i[8180] & sel_one_hot_i[63];
  assign data_masked[8179] = data_i[8179] & sel_one_hot_i[63];
  assign data_masked[8178] = data_i[8178] & sel_one_hot_i[63];
  assign data_masked[8177] = data_i[8177] & sel_one_hot_i[63];
  assign data_masked[8176] = data_i[8176] & sel_one_hot_i[63];
  assign data_masked[8175] = data_i[8175] & sel_one_hot_i[63];
  assign data_masked[8174] = data_i[8174] & sel_one_hot_i[63];
  assign data_masked[8173] = data_i[8173] & sel_one_hot_i[63];
  assign data_masked[8172] = data_i[8172] & sel_one_hot_i[63];
  assign data_masked[8171] = data_i[8171] & sel_one_hot_i[63];
  assign data_masked[8170] = data_i[8170] & sel_one_hot_i[63];
  assign data_masked[8169] = data_i[8169] & sel_one_hot_i[63];
  assign data_masked[8168] = data_i[8168] & sel_one_hot_i[63];
  assign data_masked[8167] = data_i[8167] & sel_one_hot_i[63];
  assign data_masked[8166] = data_i[8166] & sel_one_hot_i[63];
  assign data_masked[8165] = data_i[8165] & sel_one_hot_i[63];
  assign data_masked[8164] = data_i[8164] & sel_one_hot_i[63];
  assign data_masked[8163] = data_i[8163] & sel_one_hot_i[63];
  assign data_masked[8162] = data_i[8162] & sel_one_hot_i[63];
  assign data_masked[8161] = data_i[8161] & sel_one_hot_i[63];
  assign data_masked[8160] = data_i[8160] & sel_one_hot_i[63];
  assign data_masked[8159] = data_i[8159] & sel_one_hot_i[63];
  assign data_masked[8158] = data_i[8158] & sel_one_hot_i[63];
  assign data_masked[8157] = data_i[8157] & sel_one_hot_i[63];
  assign data_masked[8156] = data_i[8156] & sel_one_hot_i[63];
  assign data_masked[8155] = data_i[8155] & sel_one_hot_i[63];
  assign data_masked[8154] = data_i[8154] & sel_one_hot_i[63];
  assign data_masked[8153] = data_i[8153] & sel_one_hot_i[63];
  assign data_masked[8152] = data_i[8152] & sel_one_hot_i[63];
  assign data_masked[8151] = data_i[8151] & sel_one_hot_i[63];
  assign data_masked[8150] = data_i[8150] & sel_one_hot_i[63];
  assign data_masked[8149] = data_i[8149] & sel_one_hot_i[63];
  assign data_masked[8148] = data_i[8148] & sel_one_hot_i[63];
  assign data_masked[8147] = data_i[8147] & sel_one_hot_i[63];
  assign data_masked[8146] = data_i[8146] & sel_one_hot_i[63];
  assign data_masked[8145] = data_i[8145] & sel_one_hot_i[63];
  assign data_masked[8144] = data_i[8144] & sel_one_hot_i[63];
  assign data_masked[8143] = data_i[8143] & sel_one_hot_i[63];
  assign data_masked[8142] = data_i[8142] & sel_one_hot_i[63];
  assign data_masked[8141] = data_i[8141] & sel_one_hot_i[63];
  assign data_masked[8140] = data_i[8140] & sel_one_hot_i[63];
  assign data_masked[8139] = data_i[8139] & sel_one_hot_i[63];
  assign data_masked[8138] = data_i[8138] & sel_one_hot_i[63];
  assign data_masked[8137] = data_i[8137] & sel_one_hot_i[63];
  assign data_masked[8136] = data_i[8136] & sel_one_hot_i[63];
  assign data_masked[8135] = data_i[8135] & sel_one_hot_i[63];
  assign data_masked[8134] = data_i[8134] & sel_one_hot_i[63];
  assign data_masked[8133] = data_i[8133] & sel_one_hot_i[63];
  assign data_masked[8132] = data_i[8132] & sel_one_hot_i[63];
  assign data_masked[8131] = data_i[8131] & sel_one_hot_i[63];
  assign data_masked[8130] = data_i[8130] & sel_one_hot_i[63];
  assign data_masked[8129] = data_i[8129] & sel_one_hot_i[63];
  assign data_masked[8128] = data_i[8128] & sel_one_hot_i[63];
  assign data_masked[8127] = data_i[8127] & sel_one_hot_i[63];
  assign data_masked[8126] = data_i[8126] & sel_one_hot_i[63];
  assign data_masked[8125] = data_i[8125] & sel_one_hot_i[63];
  assign data_masked[8124] = data_i[8124] & sel_one_hot_i[63];
  assign data_masked[8123] = data_i[8123] & sel_one_hot_i[63];
  assign data_masked[8122] = data_i[8122] & sel_one_hot_i[63];
  assign data_masked[8121] = data_i[8121] & sel_one_hot_i[63];
  assign data_masked[8120] = data_i[8120] & sel_one_hot_i[63];
  assign data_masked[8119] = data_i[8119] & sel_one_hot_i[63];
  assign data_masked[8118] = data_i[8118] & sel_one_hot_i[63];
  assign data_masked[8117] = data_i[8117] & sel_one_hot_i[63];
  assign data_masked[8116] = data_i[8116] & sel_one_hot_i[63];
  assign data_masked[8115] = data_i[8115] & sel_one_hot_i[63];
  assign data_masked[8114] = data_i[8114] & sel_one_hot_i[63];
  assign data_masked[8113] = data_i[8113] & sel_one_hot_i[63];
  assign data_masked[8112] = data_i[8112] & sel_one_hot_i[63];
  assign data_masked[8111] = data_i[8111] & sel_one_hot_i[63];
  assign data_masked[8110] = data_i[8110] & sel_one_hot_i[63];
  assign data_masked[8109] = data_i[8109] & sel_one_hot_i[63];
  assign data_masked[8108] = data_i[8108] & sel_one_hot_i[63];
  assign data_masked[8107] = data_i[8107] & sel_one_hot_i[63];
  assign data_masked[8106] = data_i[8106] & sel_one_hot_i[63];
  assign data_masked[8105] = data_i[8105] & sel_one_hot_i[63];
  assign data_masked[8104] = data_i[8104] & sel_one_hot_i[63];
  assign data_masked[8103] = data_i[8103] & sel_one_hot_i[63];
  assign data_masked[8102] = data_i[8102] & sel_one_hot_i[63];
  assign data_masked[8101] = data_i[8101] & sel_one_hot_i[63];
  assign data_masked[8100] = data_i[8100] & sel_one_hot_i[63];
  assign data_masked[8099] = data_i[8099] & sel_one_hot_i[63];
  assign data_masked[8098] = data_i[8098] & sel_one_hot_i[63];
  assign data_masked[8097] = data_i[8097] & sel_one_hot_i[63];
  assign data_masked[8096] = data_i[8096] & sel_one_hot_i[63];
  assign data_masked[8095] = data_i[8095] & sel_one_hot_i[63];
  assign data_masked[8094] = data_i[8094] & sel_one_hot_i[63];
  assign data_masked[8093] = data_i[8093] & sel_one_hot_i[63];
  assign data_masked[8092] = data_i[8092] & sel_one_hot_i[63];
  assign data_masked[8091] = data_i[8091] & sel_one_hot_i[63];
  assign data_masked[8090] = data_i[8090] & sel_one_hot_i[63];
  assign data_masked[8089] = data_i[8089] & sel_one_hot_i[63];
  assign data_masked[8088] = data_i[8088] & sel_one_hot_i[63];
  assign data_masked[8087] = data_i[8087] & sel_one_hot_i[63];
  assign data_masked[8086] = data_i[8086] & sel_one_hot_i[63];
  assign data_masked[8085] = data_i[8085] & sel_one_hot_i[63];
  assign data_masked[8084] = data_i[8084] & sel_one_hot_i[63];
  assign data_masked[8083] = data_i[8083] & sel_one_hot_i[63];
  assign data_masked[8082] = data_i[8082] & sel_one_hot_i[63];
  assign data_masked[8081] = data_i[8081] & sel_one_hot_i[63];
  assign data_masked[8080] = data_i[8080] & sel_one_hot_i[63];
  assign data_masked[8079] = data_i[8079] & sel_one_hot_i[63];
  assign data_masked[8078] = data_i[8078] & sel_one_hot_i[63];
  assign data_masked[8077] = data_i[8077] & sel_one_hot_i[63];
  assign data_masked[8076] = data_i[8076] & sel_one_hot_i[63];
  assign data_masked[8075] = data_i[8075] & sel_one_hot_i[63];
  assign data_masked[8074] = data_i[8074] & sel_one_hot_i[63];
  assign data_masked[8073] = data_i[8073] & sel_one_hot_i[63];
  assign data_masked[8072] = data_i[8072] & sel_one_hot_i[63];
  assign data_masked[8071] = data_i[8071] & sel_one_hot_i[63];
  assign data_masked[8070] = data_i[8070] & sel_one_hot_i[63];
  assign data_masked[8069] = data_i[8069] & sel_one_hot_i[63];
  assign data_masked[8068] = data_i[8068] & sel_one_hot_i[63];
  assign data_masked[8067] = data_i[8067] & sel_one_hot_i[63];
  assign data_masked[8066] = data_i[8066] & sel_one_hot_i[63];
  assign data_masked[8065] = data_i[8065] & sel_one_hot_i[63];
  assign data_masked[8064] = data_i[8064] & sel_one_hot_i[63];
  assign data_masked[8319] = data_i[8319] & sel_one_hot_i[64];
  assign data_masked[8318] = data_i[8318] & sel_one_hot_i[64];
  assign data_masked[8317] = data_i[8317] & sel_one_hot_i[64];
  assign data_masked[8316] = data_i[8316] & sel_one_hot_i[64];
  assign data_masked[8315] = data_i[8315] & sel_one_hot_i[64];
  assign data_masked[8314] = data_i[8314] & sel_one_hot_i[64];
  assign data_masked[8313] = data_i[8313] & sel_one_hot_i[64];
  assign data_masked[8312] = data_i[8312] & sel_one_hot_i[64];
  assign data_masked[8311] = data_i[8311] & sel_one_hot_i[64];
  assign data_masked[8310] = data_i[8310] & sel_one_hot_i[64];
  assign data_masked[8309] = data_i[8309] & sel_one_hot_i[64];
  assign data_masked[8308] = data_i[8308] & sel_one_hot_i[64];
  assign data_masked[8307] = data_i[8307] & sel_one_hot_i[64];
  assign data_masked[8306] = data_i[8306] & sel_one_hot_i[64];
  assign data_masked[8305] = data_i[8305] & sel_one_hot_i[64];
  assign data_masked[8304] = data_i[8304] & sel_one_hot_i[64];
  assign data_masked[8303] = data_i[8303] & sel_one_hot_i[64];
  assign data_masked[8302] = data_i[8302] & sel_one_hot_i[64];
  assign data_masked[8301] = data_i[8301] & sel_one_hot_i[64];
  assign data_masked[8300] = data_i[8300] & sel_one_hot_i[64];
  assign data_masked[8299] = data_i[8299] & sel_one_hot_i[64];
  assign data_masked[8298] = data_i[8298] & sel_one_hot_i[64];
  assign data_masked[8297] = data_i[8297] & sel_one_hot_i[64];
  assign data_masked[8296] = data_i[8296] & sel_one_hot_i[64];
  assign data_masked[8295] = data_i[8295] & sel_one_hot_i[64];
  assign data_masked[8294] = data_i[8294] & sel_one_hot_i[64];
  assign data_masked[8293] = data_i[8293] & sel_one_hot_i[64];
  assign data_masked[8292] = data_i[8292] & sel_one_hot_i[64];
  assign data_masked[8291] = data_i[8291] & sel_one_hot_i[64];
  assign data_masked[8290] = data_i[8290] & sel_one_hot_i[64];
  assign data_masked[8289] = data_i[8289] & sel_one_hot_i[64];
  assign data_masked[8288] = data_i[8288] & sel_one_hot_i[64];
  assign data_masked[8287] = data_i[8287] & sel_one_hot_i[64];
  assign data_masked[8286] = data_i[8286] & sel_one_hot_i[64];
  assign data_masked[8285] = data_i[8285] & sel_one_hot_i[64];
  assign data_masked[8284] = data_i[8284] & sel_one_hot_i[64];
  assign data_masked[8283] = data_i[8283] & sel_one_hot_i[64];
  assign data_masked[8282] = data_i[8282] & sel_one_hot_i[64];
  assign data_masked[8281] = data_i[8281] & sel_one_hot_i[64];
  assign data_masked[8280] = data_i[8280] & sel_one_hot_i[64];
  assign data_masked[8279] = data_i[8279] & sel_one_hot_i[64];
  assign data_masked[8278] = data_i[8278] & sel_one_hot_i[64];
  assign data_masked[8277] = data_i[8277] & sel_one_hot_i[64];
  assign data_masked[8276] = data_i[8276] & sel_one_hot_i[64];
  assign data_masked[8275] = data_i[8275] & sel_one_hot_i[64];
  assign data_masked[8274] = data_i[8274] & sel_one_hot_i[64];
  assign data_masked[8273] = data_i[8273] & sel_one_hot_i[64];
  assign data_masked[8272] = data_i[8272] & sel_one_hot_i[64];
  assign data_masked[8271] = data_i[8271] & sel_one_hot_i[64];
  assign data_masked[8270] = data_i[8270] & sel_one_hot_i[64];
  assign data_masked[8269] = data_i[8269] & sel_one_hot_i[64];
  assign data_masked[8268] = data_i[8268] & sel_one_hot_i[64];
  assign data_masked[8267] = data_i[8267] & sel_one_hot_i[64];
  assign data_masked[8266] = data_i[8266] & sel_one_hot_i[64];
  assign data_masked[8265] = data_i[8265] & sel_one_hot_i[64];
  assign data_masked[8264] = data_i[8264] & sel_one_hot_i[64];
  assign data_masked[8263] = data_i[8263] & sel_one_hot_i[64];
  assign data_masked[8262] = data_i[8262] & sel_one_hot_i[64];
  assign data_masked[8261] = data_i[8261] & sel_one_hot_i[64];
  assign data_masked[8260] = data_i[8260] & sel_one_hot_i[64];
  assign data_masked[8259] = data_i[8259] & sel_one_hot_i[64];
  assign data_masked[8258] = data_i[8258] & sel_one_hot_i[64];
  assign data_masked[8257] = data_i[8257] & sel_one_hot_i[64];
  assign data_masked[8256] = data_i[8256] & sel_one_hot_i[64];
  assign data_masked[8255] = data_i[8255] & sel_one_hot_i[64];
  assign data_masked[8254] = data_i[8254] & sel_one_hot_i[64];
  assign data_masked[8253] = data_i[8253] & sel_one_hot_i[64];
  assign data_masked[8252] = data_i[8252] & sel_one_hot_i[64];
  assign data_masked[8251] = data_i[8251] & sel_one_hot_i[64];
  assign data_masked[8250] = data_i[8250] & sel_one_hot_i[64];
  assign data_masked[8249] = data_i[8249] & sel_one_hot_i[64];
  assign data_masked[8248] = data_i[8248] & sel_one_hot_i[64];
  assign data_masked[8247] = data_i[8247] & sel_one_hot_i[64];
  assign data_masked[8246] = data_i[8246] & sel_one_hot_i[64];
  assign data_masked[8245] = data_i[8245] & sel_one_hot_i[64];
  assign data_masked[8244] = data_i[8244] & sel_one_hot_i[64];
  assign data_masked[8243] = data_i[8243] & sel_one_hot_i[64];
  assign data_masked[8242] = data_i[8242] & sel_one_hot_i[64];
  assign data_masked[8241] = data_i[8241] & sel_one_hot_i[64];
  assign data_masked[8240] = data_i[8240] & sel_one_hot_i[64];
  assign data_masked[8239] = data_i[8239] & sel_one_hot_i[64];
  assign data_masked[8238] = data_i[8238] & sel_one_hot_i[64];
  assign data_masked[8237] = data_i[8237] & sel_one_hot_i[64];
  assign data_masked[8236] = data_i[8236] & sel_one_hot_i[64];
  assign data_masked[8235] = data_i[8235] & sel_one_hot_i[64];
  assign data_masked[8234] = data_i[8234] & sel_one_hot_i[64];
  assign data_masked[8233] = data_i[8233] & sel_one_hot_i[64];
  assign data_masked[8232] = data_i[8232] & sel_one_hot_i[64];
  assign data_masked[8231] = data_i[8231] & sel_one_hot_i[64];
  assign data_masked[8230] = data_i[8230] & sel_one_hot_i[64];
  assign data_masked[8229] = data_i[8229] & sel_one_hot_i[64];
  assign data_masked[8228] = data_i[8228] & sel_one_hot_i[64];
  assign data_masked[8227] = data_i[8227] & sel_one_hot_i[64];
  assign data_masked[8226] = data_i[8226] & sel_one_hot_i[64];
  assign data_masked[8225] = data_i[8225] & sel_one_hot_i[64];
  assign data_masked[8224] = data_i[8224] & sel_one_hot_i[64];
  assign data_masked[8223] = data_i[8223] & sel_one_hot_i[64];
  assign data_masked[8222] = data_i[8222] & sel_one_hot_i[64];
  assign data_masked[8221] = data_i[8221] & sel_one_hot_i[64];
  assign data_masked[8220] = data_i[8220] & sel_one_hot_i[64];
  assign data_masked[8219] = data_i[8219] & sel_one_hot_i[64];
  assign data_masked[8218] = data_i[8218] & sel_one_hot_i[64];
  assign data_masked[8217] = data_i[8217] & sel_one_hot_i[64];
  assign data_masked[8216] = data_i[8216] & sel_one_hot_i[64];
  assign data_masked[8215] = data_i[8215] & sel_one_hot_i[64];
  assign data_masked[8214] = data_i[8214] & sel_one_hot_i[64];
  assign data_masked[8213] = data_i[8213] & sel_one_hot_i[64];
  assign data_masked[8212] = data_i[8212] & sel_one_hot_i[64];
  assign data_masked[8211] = data_i[8211] & sel_one_hot_i[64];
  assign data_masked[8210] = data_i[8210] & sel_one_hot_i[64];
  assign data_masked[8209] = data_i[8209] & sel_one_hot_i[64];
  assign data_masked[8208] = data_i[8208] & sel_one_hot_i[64];
  assign data_masked[8207] = data_i[8207] & sel_one_hot_i[64];
  assign data_masked[8206] = data_i[8206] & sel_one_hot_i[64];
  assign data_masked[8205] = data_i[8205] & sel_one_hot_i[64];
  assign data_masked[8204] = data_i[8204] & sel_one_hot_i[64];
  assign data_masked[8203] = data_i[8203] & sel_one_hot_i[64];
  assign data_masked[8202] = data_i[8202] & sel_one_hot_i[64];
  assign data_masked[8201] = data_i[8201] & sel_one_hot_i[64];
  assign data_masked[8200] = data_i[8200] & sel_one_hot_i[64];
  assign data_masked[8199] = data_i[8199] & sel_one_hot_i[64];
  assign data_masked[8198] = data_i[8198] & sel_one_hot_i[64];
  assign data_masked[8197] = data_i[8197] & sel_one_hot_i[64];
  assign data_masked[8196] = data_i[8196] & sel_one_hot_i[64];
  assign data_masked[8195] = data_i[8195] & sel_one_hot_i[64];
  assign data_masked[8194] = data_i[8194] & sel_one_hot_i[64];
  assign data_masked[8193] = data_i[8193] & sel_one_hot_i[64];
  assign data_masked[8192] = data_i[8192] & sel_one_hot_i[64];
  assign data_masked[8447] = data_i[8447] & sel_one_hot_i[65];
  assign data_masked[8446] = data_i[8446] & sel_one_hot_i[65];
  assign data_masked[8445] = data_i[8445] & sel_one_hot_i[65];
  assign data_masked[8444] = data_i[8444] & sel_one_hot_i[65];
  assign data_masked[8443] = data_i[8443] & sel_one_hot_i[65];
  assign data_masked[8442] = data_i[8442] & sel_one_hot_i[65];
  assign data_masked[8441] = data_i[8441] & sel_one_hot_i[65];
  assign data_masked[8440] = data_i[8440] & sel_one_hot_i[65];
  assign data_masked[8439] = data_i[8439] & sel_one_hot_i[65];
  assign data_masked[8438] = data_i[8438] & sel_one_hot_i[65];
  assign data_masked[8437] = data_i[8437] & sel_one_hot_i[65];
  assign data_masked[8436] = data_i[8436] & sel_one_hot_i[65];
  assign data_masked[8435] = data_i[8435] & sel_one_hot_i[65];
  assign data_masked[8434] = data_i[8434] & sel_one_hot_i[65];
  assign data_masked[8433] = data_i[8433] & sel_one_hot_i[65];
  assign data_masked[8432] = data_i[8432] & sel_one_hot_i[65];
  assign data_masked[8431] = data_i[8431] & sel_one_hot_i[65];
  assign data_masked[8430] = data_i[8430] & sel_one_hot_i[65];
  assign data_masked[8429] = data_i[8429] & sel_one_hot_i[65];
  assign data_masked[8428] = data_i[8428] & sel_one_hot_i[65];
  assign data_masked[8427] = data_i[8427] & sel_one_hot_i[65];
  assign data_masked[8426] = data_i[8426] & sel_one_hot_i[65];
  assign data_masked[8425] = data_i[8425] & sel_one_hot_i[65];
  assign data_masked[8424] = data_i[8424] & sel_one_hot_i[65];
  assign data_masked[8423] = data_i[8423] & sel_one_hot_i[65];
  assign data_masked[8422] = data_i[8422] & sel_one_hot_i[65];
  assign data_masked[8421] = data_i[8421] & sel_one_hot_i[65];
  assign data_masked[8420] = data_i[8420] & sel_one_hot_i[65];
  assign data_masked[8419] = data_i[8419] & sel_one_hot_i[65];
  assign data_masked[8418] = data_i[8418] & sel_one_hot_i[65];
  assign data_masked[8417] = data_i[8417] & sel_one_hot_i[65];
  assign data_masked[8416] = data_i[8416] & sel_one_hot_i[65];
  assign data_masked[8415] = data_i[8415] & sel_one_hot_i[65];
  assign data_masked[8414] = data_i[8414] & sel_one_hot_i[65];
  assign data_masked[8413] = data_i[8413] & sel_one_hot_i[65];
  assign data_masked[8412] = data_i[8412] & sel_one_hot_i[65];
  assign data_masked[8411] = data_i[8411] & sel_one_hot_i[65];
  assign data_masked[8410] = data_i[8410] & sel_one_hot_i[65];
  assign data_masked[8409] = data_i[8409] & sel_one_hot_i[65];
  assign data_masked[8408] = data_i[8408] & sel_one_hot_i[65];
  assign data_masked[8407] = data_i[8407] & sel_one_hot_i[65];
  assign data_masked[8406] = data_i[8406] & sel_one_hot_i[65];
  assign data_masked[8405] = data_i[8405] & sel_one_hot_i[65];
  assign data_masked[8404] = data_i[8404] & sel_one_hot_i[65];
  assign data_masked[8403] = data_i[8403] & sel_one_hot_i[65];
  assign data_masked[8402] = data_i[8402] & sel_one_hot_i[65];
  assign data_masked[8401] = data_i[8401] & sel_one_hot_i[65];
  assign data_masked[8400] = data_i[8400] & sel_one_hot_i[65];
  assign data_masked[8399] = data_i[8399] & sel_one_hot_i[65];
  assign data_masked[8398] = data_i[8398] & sel_one_hot_i[65];
  assign data_masked[8397] = data_i[8397] & sel_one_hot_i[65];
  assign data_masked[8396] = data_i[8396] & sel_one_hot_i[65];
  assign data_masked[8395] = data_i[8395] & sel_one_hot_i[65];
  assign data_masked[8394] = data_i[8394] & sel_one_hot_i[65];
  assign data_masked[8393] = data_i[8393] & sel_one_hot_i[65];
  assign data_masked[8392] = data_i[8392] & sel_one_hot_i[65];
  assign data_masked[8391] = data_i[8391] & sel_one_hot_i[65];
  assign data_masked[8390] = data_i[8390] & sel_one_hot_i[65];
  assign data_masked[8389] = data_i[8389] & sel_one_hot_i[65];
  assign data_masked[8388] = data_i[8388] & sel_one_hot_i[65];
  assign data_masked[8387] = data_i[8387] & sel_one_hot_i[65];
  assign data_masked[8386] = data_i[8386] & sel_one_hot_i[65];
  assign data_masked[8385] = data_i[8385] & sel_one_hot_i[65];
  assign data_masked[8384] = data_i[8384] & sel_one_hot_i[65];
  assign data_masked[8383] = data_i[8383] & sel_one_hot_i[65];
  assign data_masked[8382] = data_i[8382] & sel_one_hot_i[65];
  assign data_masked[8381] = data_i[8381] & sel_one_hot_i[65];
  assign data_masked[8380] = data_i[8380] & sel_one_hot_i[65];
  assign data_masked[8379] = data_i[8379] & sel_one_hot_i[65];
  assign data_masked[8378] = data_i[8378] & sel_one_hot_i[65];
  assign data_masked[8377] = data_i[8377] & sel_one_hot_i[65];
  assign data_masked[8376] = data_i[8376] & sel_one_hot_i[65];
  assign data_masked[8375] = data_i[8375] & sel_one_hot_i[65];
  assign data_masked[8374] = data_i[8374] & sel_one_hot_i[65];
  assign data_masked[8373] = data_i[8373] & sel_one_hot_i[65];
  assign data_masked[8372] = data_i[8372] & sel_one_hot_i[65];
  assign data_masked[8371] = data_i[8371] & sel_one_hot_i[65];
  assign data_masked[8370] = data_i[8370] & sel_one_hot_i[65];
  assign data_masked[8369] = data_i[8369] & sel_one_hot_i[65];
  assign data_masked[8368] = data_i[8368] & sel_one_hot_i[65];
  assign data_masked[8367] = data_i[8367] & sel_one_hot_i[65];
  assign data_masked[8366] = data_i[8366] & sel_one_hot_i[65];
  assign data_masked[8365] = data_i[8365] & sel_one_hot_i[65];
  assign data_masked[8364] = data_i[8364] & sel_one_hot_i[65];
  assign data_masked[8363] = data_i[8363] & sel_one_hot_i[65];
  assign data_masked[8362] = data_i[8362] & sel_one_hot_i[65];
  assign data_masked[8361] = data_i[8361] & sel_one_hot_i[65];
  assign data_masked[8360] = data_i[8360] & sel_one_hot_i[65];
  assign data_masked[8359] = data_i[8359] & sel_one_hot_i[65];
  assign data_masked[8358] = data_i[8358] & sel_one_hot_i[65];
  assign data_masked[8357] = data_i[8357] & sel_one_hot_i[65];
  assign data_masked[8356] = data_i[8356] & sel_one_hot_i[65];
  assign data_masked[8355] = data_i[8355] & sel_one_hot_i[65];
  assign data_masked[8354] = data_i[8354] & sel_one_hot_i[65];
  assign data_masked[8353] = data_i[8353] & sel_one_hot_i[65];
  assign data_masked[8352] = data_i[8352] & sel_one_hot_i[65];
  assign data_masked[8351] = data_i[8351] & sel_one_hot_i[65];
  assign data_masked[8350] = data_i[8350] & sel_one_hot_i[65];
  assign data_masked[8349] = data_i[8349] & sel_one_hot_i[65];
  assign data_masked[8348] = data_i[8348] & sel_one_hot_i[65];
  assign data_masked[8347] = data_i[8347] & sel_one_hot_i[65];
  assign data_masked[8346] = data_i[8346] & sel_one_hot_i[65];
  assign data_masked[8345] = data_i[8345] & sel_one_hot_i[65];
  assign data_masked[8344] = data_i[8344] & sel_one_hot_i[65];
  assign data_masked[8343] = data_i[8343] & sel_one_hot_i[65];
  assign data_masked[8342] = data_i[8342] & sel_one_hot_i[65];
  assign data_masked[8341] = data_i[8341] & sel_one_hot_i[65];
  assign data_masked[8340] = data_i[8340] & sel_one_hot_i[65];
  assign data_masked[8339] = data_i[8339] & sel_one_hot_i[65];
  assign data_masked[8338] = data_i[8338] & sel_one_hot_i[65];
  assign data_masked[8337] = data_i[8337] & sel_one_hot_i[65];
  assign data_masked[8336] = data_i[8336] & sel_one_hot_i[65];
  assign data_masked[8335] = data_i[8335] & sel_one_hot_i[65];
  assign data_masked[8334] = data_i[8334] & sel_one_hot_i[65];
  assign data_masked[8333] = data_i[8333] & sel_one_hot_i[65];
  assign data_masked[8332] = data_i[8332] & sel_one_hot_i[65];
  assign data_masked[8331] = data_i[8331] & sel_one_hot_i[65];
  assign data_masked[8330] = data_i[8330] & sel_one_hot_i[65];
  assign data_masked[8329] = data_i[8329] & sel_one_hot_i[65];
  assign data_masked[8328] = data_i[8328] & sel_one_hot_i[65];
  assign data_masked[8327] = data_i[8327] & sel_one_hot_i[65];
  assign data_masked[8326] = data_i[8326] & sel_one_hot_i[65];
  assign data_masked[8325] = data_i[8325] & sel_one_hot_i[65];
  assign data_masked[8324] = data_i[8324] & sel_one_hot_i[65];
  assign data_masked[8323] = data_i[8323] & sel_one_hot_i[65];
  assign data_masked[8322] = data_i[8322] & sel_one_hot_i[65];
  assign data_masked[8321] = data_i[8321] & sel_one_hot_i[65];
  assign data_masked[8320] = data_i[8320] & sel_one_hot_i[65];
  assign data_masked[8575] = data_i[8575] & sel_one_hot_i[66];
  assign data_masked[8574] = data_i[8574] & sel_one_hot_i[66];
  assign data_masked[8573] = data_i[8573] & sel_one_hot_i[66];
  assign data_masked[8572] = data_i[8572] & sel_one_hot_i[66];
  assign data_masked[8571] = data_i[8571] & sel_one_hot_i[66];
  assign data_masked[8570] = data_i[8570] & sel_one_hot_i[66];
  assign data_masked[8569] = data_i[8569] & sel_one_hot_i[66];
  assign data_masked[8568] = data_i[8568] & sel_one_hot_i[66];
  assign data_masked[8567] = data_i[8567] & sel_one_hot_i[66];
  assign data_masked[8566] = data_i[8566] & sel_one_hot_i[66];
  assign data_masked[8565] = data_i[8565] & sel_one_hot_i[66];
  assign data_masked[8564] = data_i[8564] & sel_one_hot_i[66];
  assign data_masked[8563] = data_i[8563] & sel_one_hot_i[66];
  assign data_masked[8562] = data_i[8562] & sel_one_hot_i[66];
  assign data_masked[8561] = data_i[8561] & sel_one_hot_i[66];
  assign data_masked[8560] = data_i[8560] & sel_one_hot_i[66];
  assign data_masked[8559] = data_i[8559] & sel_one_hot_i[66];
  assign data_masked[8558] = data_i[8558] & sel_one_hot_i[66];
  assign data_masked[8557] = data_i[8557] & sel_one_hot_i[66];
  assign data_masked[8556] = data_i[8556] & sel_one_hot_i[66];
  assign data_masked[8555] = data_i[8555] & sel_one_hot_i[66];
  assign data_masked[8554] = data_i[8554] & sel_one_hot_i[66];
  assign data_masked[8553] = data_i[8553] & sel_one_hot_i[66];
  assign data_masked[8552] = data_i[8552] & sel_one_hot_i[66];
  assign data_masked[8551] = data_i[8551] & sel_one_hot_i[66];
  assign data_masked[8550] = data_i[8550] & sel_one_hot_i[66];
  assign data_masked[8549] = data_i[8549] & sel_one_hot_i[66];
  assign data_masked[8548] = data_i[8548] & sel_one_hot_i[66];
  assign data_masked[8547] = data_i[8547] & sel_one_hot_i[66];
  assign data_masked[8546] = data_i[8546] & sel_one_hot_i[66];
  assign data_masked[8545] = data_i[8545] & sel_one_hot_i[66];
  assign data_masked[8544] = data_i[8544] & sel_one_hot_i[66];
  assign data_masked[8543] = data_i[8543] & sel_one_hot_i[66];
  assign data_masked[8542] = data_i[8542] & sel_one_hot_i[66];
  assign data_masked[8541] = data_i[8541] & sel_one_hot_i[66];
  assign data_masked[8540] = data_i[8540] & sel_one_hot_i[66];
  assign data_masked[8539] = data_i[8539] & sel_one_hot_i[66];
  assign data_masked[8538] = data_i[8538] & sel_one_hot_i[66];
  assign data_masked[8537] = data_i[8537] & sel_one_hot_i[66];
  assign data_masked[8536] = data_i[8536] & sel_one_hot_i[66];
  assign data_masked[8535] = data_i[8535] & sel_one_hot_i[66];
  assign data_masked[8534] = data_i[8534] & sel_one_hot_i[66];
  assign data_masked[8533] = data_i[8533] & sel_one_hot_i[66];
  assign data_masked[8532] = data_i[8532] & sel_one_hot_i[66];
  assign data_masked[8531] = data_i[8531] & sel_one_hot_i[66];
  assign data_masked[8530] = data_i[8530] & sel_one_hot_i[66];
  assign data_masked[8529] = data_i[8529] & sel_one_hot_i[66];
  assign data_masked[8528] = data_i[8528] & sel_one_hot_i[66];
  assign data_masked[8527] = data_i[8527] & sel_one_hot_i[66];
  assign data_masked[8526] = data_i[8526] & sel_one_hot_i[66];
  assign data_masked[8525] = data_i[8525] & sel_one_hot_i[66];
  assign data_masked[8524] = data_i[8524] & sel_one_hot_i[66];
  assign data_masked[8523] = data_i[8523] & sel_one_hot_i[66];
  assign data_masked[8522] = data_i[8522] & sel_one_hot_i[66];
  assign data_masked[8521] = data_i[8521] & sel_one_hot_i[66];
  assign data_masked[8520] = data_i[8520] & sel_one_hot_i[66];
  assign data_masked[8519] = data_i[8519] & sel_one_hot_i[66];
  assign data_masked[8518] = data_i[8518] & sel_one_hot_i[66];
  assign data_masked[8517] = data_i[8517] & sel_one_hot_i[66];
  assign data_masked[8516] = data_i[8516] & sel_one_hot_i[66];
  assign data_masked[8515] = data_i[8515] & sel_one_hot_i[66];
  assign data_masked[8514] = data_i[8514] & sel_one_hot_i[66];
  assign data_masked[8513] = data_i[8513] & sel_one_hot_i[66];
  assign data_masked[8512] = data_i[8512] & sel_one_hot_i[66];
  assign data_masked[8511] = data_i[8511] & sel_one_hot_i[66];
  assign data_masked[8510] = data_i[8510] & sel_one_hot_i[66];
  assign data_masked[8509] = data_i[8509] & sel_one_hot_i[66];
  assign data_masked[8508] = data_i[8508] & sel_one_hot_i[66];
  assign data_masked[8507] = data_i[8507] & sel_one_hot_i[66];
  assign data_masked[8506] = data_i[8506] & sel_one_hot_i[66];
  assign data_masked[8505] = data_i[8505] & sel_one_hot_i[66];
  assign data_masked[8504] = data_i[8504] & sel_one_hot_i[66];
  assign data_masked[8503] = data_i[8503] & sel_one_hot_i[66];
  assign data_masked[8502] = data_i[8502] & sel_one_hot_i[66];
  assign data_masked[8501] = data_i[8501] & sel_one_hot_i[66];
  assign data_masked[8500] = data_i[8500] & sel_one_hot_i[66];
  assign data_masked[8499] = data_i[8499] & sel_one_hot_i[66];
  assign data_masked[8498] = data_i[8498] & sel_one_hot_i[66];
  assign data_masked[8497] = data_i[8497] & sel_one_hot_i[66];
  assign data_masked[8496] = data_i[8496] & sel_one_hot_i[66];
  assign data_masked[8495] = data_i[8495] & sel_one_hot_i[66];
  assign data_masked[8494] = data_i[8494] & sel_one_hot_i[66];
  assign data_masked[8493] = data_i[8493] & sel_one_hot_i[66];
  assign data_masked[8492] = data_i[8492] & sel_one_hot_i[66];
  assign data_masked[8491] = data_i[8491] & sel_one_hot_i[66];
  assign data_masked[8490] = data_i[8490] & sel_one_hot_i[66];
  assign data_masked[8489] = data_i[8489] & sel_one_hot_i[66];
  assign data_masked[8488] = data_i[8488] & sel_one_hot_i[66];
  assign data_masked[8487] = data_i[8487] & sel_one_hot_i[66];
  assign data_masked[8486] = data_i[8486] & sel_one_hot_i[66];
  assign data_masked[8485] = data_i[8485] & sel_one_hot_i[66];
  assign data_masked[8484] = data_i[8484] & sel_one_hot_i[66];
  assign data_masked[8483] = data_i[8483] & sel_one_hot_i[66];
  assign data_masked[8482] = data_i[8482] & sel_one_hot_i[66];
  assign data_masked[8481] = data_i[8481] & sel_one_hot_i[66];
  assign data_masked[8480] = data_i[8480] & sel_one_hot_i[66];
  assign data_masked[8479] = data_i[8479] & sel_one_hot_i[66];
  assign data_masked[8478] = data_i[8478] & sel_one_hot_i[66];
  assign data_masked[8477] = data_i[8477] & sel_one_hot_i[66];
  assign data_masked[8476] = data_i[8476] & sel_one_hot_i[66];
  assign data_masked[8475] = data_i[8475] & sel_one_hot_i[66];
  assign data_masked[8474] = data_i[8474] & sel_one_hot_i[66];
  assign data_masked[8473] = data_i[8473] & sel_one_hot_i[66];
  assign data_masked[8472] = data_i[8472] & sel_one_hot_i[66];
  assign data_masked[8471] = data_i[8471] & sel_one_hot_i[66];
  assign data_masked[8470] = data_i[8470] & sel_one_hot_i[66];
  assign data_masked[8469] = data_i[8469] & sel_one_hot_i[66];
  assign data_masked[8468] = data_i[8468] & sel_one_hot_i[66];
  assign data_masked[8467] = data_i[8467] & sel_one_hot_i[66];
  assign data_masked[8466] = data_i[8466] & sel_one_hot_i[66];
  assign data_masked[8465] = data_i[8465] & sel_one_hot_i[66];
  assign data_masked[8464] = data_i[8464] & sel_one_hot_i[66];
  assign data_masked[8463] = data_i[8463] & sel_one_hot_i[66];
  assign data_masked[8462] = data_i[8462] & sel_one_hot_i[66];
  assign data_masked[8461] = data_i[8461] & sel_one_hot_i[66];
  assign data_masked[8460] = data_i[8460] & sel_one_hot_i[66];
  assign data_masked[8459] = data_i[8459] & sel_one_hot_i[66];
  assign data_masked[8458] = data_i[8458] & sel_one_hot_i[66];
  assign data_masked[8457] = data_i[8457] & sel_one_hot_i[66];
  assign data_masked[8456] = data_i[8456] & sel_one_hot_i[66];
  assign data_masked[8455] = data_i[8455] & sel_one_hot_i[66];
  assign data_masked[8454] = data_i[8454] & sel_one_hot_i[66];
  assign data_masked[8453] = data_i[8453] & sel_one_hot_i[66];
  assign data_masked[8452] = data_i[8452] & sel_one_hot_i[66];
  assign data_masked[8451] = data_i[8451] & sel_one_hot_i[66];
  assign data_masked[8450] = data_i[8450] & sel_one_hot_i[66];
  assign data_masked[8449] = data_i[8449] & sel_one_hot_i[66];
  assign data_masked[8448] = data_i[8448] & sel_one_hot_i[66];
  assign data_masked[8703] = data_i[8703] & sel_one_hot_i[67];
  assign data_masked[8702] = data_i[8702] & sel_one_hot_i[67];
  assign data_masked[8701] = data_i[8701] & sel_one_hot_i[67];
  assign data_masked[8700] = data_i[8700] & sel_one_hot_i[67];
  assign data_masked[8699] = data_i[8699] & sel_one_hot_i[67];
  assign data_masked[8698] = data_i[8698] & sel_one_hot_i[67];
  assign data_masked[8697] = data_i[8697] & sel_one_hot_i[67];
  assign data_masked[8696] = data_i[8696] & sel_one_hot_i[67];
  assign data_masked[8695] = data_i[8695] & sel_one_hot_i[67];
  assign data_masked[8694] = data_i[8694] & sel_one_hot_i[67];
  assign data_masked[8693] = data_i[8693] & sel_one_hot_i[67];
  assign data_masked[8692] = data_i[8692] & sel_one_hot_i[67];
  assign data_masked[8691] = data_i[8691] & sel_one_hot_i[67];
  assign data_masked[8690] = data_i[8690] & sel_one_hot_i[67];
  assign data_masked[8689] = data_i[8689] & sel_one_hot_i[67];
  assign data_masked[8688] = data_i[8688] & sel_one_hot_i[67];
  assign data_masked[8687] = data_i[8687] & sel_one_hot_i[67];
  assign data_masked[8686] = data_i[8686] & sel_one_hot_i[67];
  assign data_masked[8685] = data_i[8685] & sel_one_hot_i[67];
  assign data_masked[8684] = data_i[8684] & sel_one_hot_i[67];
  assign data_masked[8683] = data_i[8683] & sel_one_hot_i[67];
  assign data_masked[8682] = data_i[8682] & sel_one_hot_i[67];
  assign data_masked[8681] = data_i[8681] & sel_one_hot_i[67];
  assign data_masked[8680] = data_i[8680] & sel_one_hot_i[67];
  assign data_masked[8679] = data_i[8679] & sel_one_hot_i[67];
  assign data_masked[8678] = data_i[8678] & sel_one_hot_i[67];
  assign data_masked[8677] = data_i[8677] & sel_one_hot_i[67];
  assign data_masked[8676] = data_i[8676] & sel_one_hot_i[67];
  assign data_masked[8675] = data_i[8675] & sel_one_hot_i[67];
  assign data_masked[8674] = data_i[8674] & sel_one_hot_i[67];
  assign data_masked[8673] = data_i[8673] & sel_one_hot_i[67];
  assign data_masked[8672] = data_i[8672] & sel_one_hot_i[67];
  assign data_masked[8671] = data_i[8671] & sel_one_hot_i[67];
  assign data_masked[8670] = data_i[8670] & sel_one_hot_i[67];
  assign data_masked[8669] = data_i[8669] & sel_one_hot_i[67];
  assign data_masked[8668] = data_i[8668] & sel_one_hot_i[67];
  assign data_masked[8667] = data_i[8667] & sel_one_hot_i[67];
  assign data_masked[8666] = data_i[8666] & sel_one_hot_i[67];
  assign data_masked[8665] = data_i[8665] & sel_one_hot_i[67];
  assign data_masked[8664] = data_i[8664] & sel_one_hot_i[67];
  assign data_masked[8663] = data_i[8663] & sel_one_hot_i[67];
  assign data_masked[8662] = data_i[8662] & sel_one_hot_i[67];
  assign data_masked[8661] = data_i[8661] & sel_one_hot_i[67];
  assign data_masked[8660] = data_i[8660] & sel_one_hot_i[67];
  assign data_masked[8659] = data_i[8659] & sel_one_hot_i[67];
  assign data_masked[8658] = data_i[8658] & sel_one_hot_i[67];
  assign data_masked[8657] = data_i[8657] & sel_one_hot_i[67];
  assign data_masked[8656] = data_i[8656] & sel_one_hot_i[67];
  assign data_masked[8655] = data_i[8655] & sel_one_hot_i[67];
  assign data_masked[8654] = data_i[8654] & sel_one_hot_i[67];
  assign data_masked[8653] = data_i[8653] & sel_one_hot_i[67];
  assign data_masked[8652] = data_i[8652] & sel_one_hot_i[67];
  assign data_masked[8651] = data_i[8651] & sel_one_hot_i[67];
  assign data_masked[8650] = data_i[8650] & sel_one_hot_i[67];
  assign data_masked[8649] = data_i[8649] & sel_one_hot_i[67];
  assign data_masked[8648] = data_i[8648] & sel_one_hot_i[67];
  assign data_masked[8647] = data_i[8647] & sel_one_hot_i[67];
  assign data_masked[8646] = data_i[8646] & sel_one_hot_i[67];
  assign data_masked[8645] = data_i[8645] & sel_one_hot_i[67];
  assign data_masked[8644] = data_i[8644] & sel_one_hot_i[67];
  assign data_masked[8643] = data_i[8643] & sel_one_hot_i[67];
  assign data_masked[8642] = data_i[8642] & sel_one_hot_i[67];
  assign data_masked[8641] = data_i[8641] & sel_one_hot_i[67];
  assign data_masked[8640] = data_i[8640] & sel_one_hot_i[67];
  assign data_masked[8639] = data_i[8639] & sel_one_hot_i[67];
  assign data_masked[8638] = data_i[8638] & sel_one_hot_i[67];
  assign data_masked[8637] = data_i[8637] & sel_one_hot_i[67];
  assign data_masked[8636] = data_i[8636] & sel_one_hot_i[67];
  assign data_masked[8635] = data_i[8635] & sel_one_hot_i[67];
  assign data_masked[8634] = data_i[8634] & sel_one_hot_i[67];
  assign data_masked[8633] = data_i[8633] & sel_one_hot_i[67];
  assign data_masked[8632] = data_i[8632] & sel_one_hot_i[67];
  assign data_masked[8631] = data_i[8631] & sel_one_hot_i[67];
  assign data_masked[8630] = data_i[8630] & sel_one_hot_i[67];
  assign data_masked[8629] = data_i[8629] & sel_one_hot_i[67];
  assign data_masked[8628] = data_i[8628] & sel_one_hot_i[67];
  assign data_masked[8627] = data_i[8627] & sel_one_hot_i[67];
  assign data_masked[8626] = data_i[8626] & sel_one_hot_i[67];
  assign data_masked[8625] = data_i[8625] & sel_one_hot_i[67];
  assign data_masked[8624] = data_i[8624] & sel_one_hot_i[67];
  assign data_masked[8623] = data_i[8623] & sel_one_hot_i[67];
  assign data_masked[8622] = data_i[8622] & sel_one_hot_i[67];
  assign data_masked[8621] = data_i[8621] & sel_one_hot_i[67];
  assign data_masked[8620] = data_i[8620] & sel_one_hot_i[67];
  assign data_masked[8619] = data_i[8619] & sel_one_hot_i[67];
  assign data_masked[8618] = data_i[8618] & sel_one_hot_i[67];
  assign data_masked[8617] = data_i[8617] & sel_one_hot_i[67];
  assign data_masked[8616] = data_i[8616] & sel_one_hot_i[67];
  assign data_masked[8615] = data_i[8615] & sel_one_hot_i[67];
  assign data_masked[8614] = data_i[8614] & sel_one_hot_i[67];
  assign data_masked[8613] = data_i[8613] & sel_one_hot_i[67];
  assign data_masked[8612] = data_i[8612] & sel_one_hot_i[67];
  assign data_masked[8611] = data_i[8611] & sel_one_hot_i[67];
  assign data_masked[8610] = data_i[8610] & sel_one_hot_i[67];
  assign data_masked[8609] = data_i[8609] & sel_one_hot_i[67];
  assign data_masked[8608] = data_i[8608] & sel_one_hot_i[67];
  assign data_masked[8607] = data_i[8607] & sel_one_hot_i[67];
  assign data_masked[8606] = data_i[8606] & sel_one_hot_i[67];
  assign data_masked[8605] = data_i[8605] & sel_one_hot_i[67];
  assign data_masked[8604] = data_i[8604] & sel_one_hot_i[67];
  assign data_masked[8603] = data_i[8603] & sel_one_hot_i[67];
  assign data_masked[8602] = data_i[8602] & sel_one_hot_i[67];
  assign data_masked[8601] = data_i[8601] & sel_one_hot_i[67];
  assign data_masked[8600] = data_i[8600] & sel_one_hot_i[67];
  assign data_masked[8599] = data_i[8599] & sel_one_hot_i[67];
  assign data_masked[8598] = data_i[8598] & sel_one_hot_i[67];
  assign data_masked[8597] = data_i[8597] & sel_one_hot_i[67];
  assign data_masked[8596] = data_i[8596] & sel_one_hot_i[67];
  assign data_masked[8595] = data_i[8595] & sel_one_hot_i[67];
  assign data_masked[8594] = data_i[8594] & sel_one_hot_i[67];
  assign data_masked[8593] = data_i[8593] & sel_one_hot_i[67];
  assign data_masked[8592] = data_i[8592] & sel_one_hot_i[67];
  assign data_masked[8591] = data_i[8591] & sel_one_hot_i[67];
  assign data_masked[8590] = data_i[8590] & sel_one_hot_i[67];
  assign data_masked[8589] = data_i[8589] & sel_one_hot_i[67];
  assign data_masked[8588] = data_i[8588] & sel_one_hot_i[67];
  assign data_masked[8587] = data_i[8587] & sel_one_hot_i[67];
  assign data_masked[8586] = data_i[8586] & sel_one_hot_i[67];
  assign data_masked[8585] = data_i[8585] & sel_one_hot_i[67];
  assign data_masked[8584] = data_i[8584] & sel_one_hot_i[67];
  assign data_masked[8583] = data_i[8583] & sel_one_hot_i[67];
  assign data_masked[8582] = data_i[8582] & sel_one_hot_i[67];
  assign data_masked[8581] = data_i[8581] & sel_one_hot_i[67];
  assign data_masked[8580] = data_i[8580] & sel_one_hot_i[67];
  assign data_masked[8579] = data_i[8579] & sel_one_hot_i[67];
  assign data_masked[8578] = data_i[8578] & sel_one_hot_i[67];
  assign data_masked[8577] = data_i[8577] & sel_one_hot_i[67];
  assign data_masked[8576] = data_i[8576] & sel_one_hot_i[67];
  assign data_masked[8831] = data_i[8831] & sel_one_hot_i[68];
  assign data_masked[8830] = data_i[8830] & sel_one_hot_i[68];
  assign data_masked[8829] = data_i[8829] & sel_one_hot_i[68];
  assign data_masked[8828] = data_i[8828] & sel_one_hot_i[68];
  assign data_masked[8827] = data_i[8827] & sel_one_hot_i[68];
  assign data_masked[8826] = data_i[8826] & sel_one_hot_i[68];
  assign data_masked[8825] = data_i[8825] & sel_one_hot_i[68];
  assign data_masked[8824] = data_i[8824] & sel_one_hot_i[68];
  assign data_masked[8823] = data_i[8823] & sel_one_hot_i[68];
  assign data_masked[8822] = data_i[8822] & sel_one_hot_i[68];
  assign data_masked[8821] = data_i[8821] & sel_one_hot_i[68];
  assign data_masked[8820] = data_i[8820] & sel_one_hot_i[68];
  assign data_masked[8819] = data_i[8819] & sel_one_hot_i[68];
  assign data_masked[8818] = data_i[8818] & sel_one_hot_i[68];
  assign data_masked[8817] = data_i[8817] & sel_one_hot_i[68];
  assign data_masked[8816] = data_i[8816] & sel_one_hot_i[68];
  assign data_masked[8815] = data_i[8815] & sel_one_hot_i[68];
  assign data_masked[8814] = data_i[8814] & sel_one_hot_i[68];
  assign data_masked[8813] = data_i[8813] & sel_one_hot_i[68];
  assign data_masked[8812] = data_i[8812] & sel_one_hot_i[68];
  assign data_masked[8811] = data_i[8811] & sel_one_hot_i[68];
  assign data_masked[8810] = data_i[8810] & sel_one_hot_i[68];
  assign data_masked[8809] = data_i[8809] & sel_one_hot_i[68];
  assign data_masked[8808] = data_i[8808] & sel_one_hot_i[68];
  assign data_masked[8807] = data_i[8807] & sel_one_hot_i[68];
  assign data_masked[8806] = data_i[8806] & sel_one_hot_i[68];
  assign data_masked[8805] = data_i[8805] & sel_one_hot_i[68];
  assign data_masked[8804] = data_i[8804] & sel_one_hot_i[68];
  assign data_masked[8803] = data_i[8803] & sel_one_hot_i[68];
  assign data_masked[8802] = data_i[8802] & sel_one_hot_i[68];
  assign data_masked[8801] = data_i[8801] & sel_one_hot_i[68];
  assign data_masked[8800] = data_i[8800] & sel_one_hot_i[68];
  assign data_masked[8799] = data_i[8799] & sel_one_hot_i[68];
  assign data_masked[8798] = data_i[8798] & sel_one_hot_i[68];
  assign data_masked[8797] = data_i[8797] & sel_one_hot_i[68];
  assign data_masked[8796] = data_i[8796] & sel_one_hot_i[68];
  assign data_masked[8795] = data_i[8795] & sel_one_hot_i[68];
  assign data_masked[8794] = data_i[8794] & sel_one_hot_i[68];
  assign data_masked[8793] = data_i[8793] & sel_one_hot_i[68];
  assign data_masked[8792] = data_i[8792] & sel_one_hot_i[68];
  assign data_masked[8791] = data_i[8791] & sel_one_hot_i[68];
  assign data_masked[8790] = data_i[8790] & sel_one_hot_i[68];
  assign data_masked[8789] = data_i[8789] & sel_one_hot_i[68];
  assign data_masked[8788] = data_i[8788] & sel_one_hot_i[68];
  assign data_masked[8787] = data_i[8787] & sel_one_hot_i[68];
  assign data_masked[8786] = data_i[8786] & sel_one_hot_i[68];
  assign data_masked[8785] = data_i[8785] & sel_one_hot_i[68];
  assign data_masked[8784] = data_i[8784] & sel_one_hot_i[68];
  assign data_masked[8783] = data_i[8783] & sel_one_hot_i[68];
  assign data_masked[8782] = data_i[8782] & sel_one_hot_i[68];
  assign data_masked[8781] = data_i[8781] & sel_one_hot_i[68];
  assign data_masked[8780] = data_i[8780] & sel_one_hot_i[68];
  assign data_masked[8779] = data_i[8779] & sel_one_hot_i[68];
  assign data_masked[8778] = data_i[8778] & sel_one_hot_i[68];
  assign data_masked[8777] = data_i[8777] & sel_one_hot_i[68];
  assign data_masked[8776] = data_i[8776] & sel_one_hot_i[68];
  assign data_masked[8775] = data_i[8775] & sel_one_hot_i[68];
  assign data_masked[8774] = data_i[8774] & sel_one_hot_i[68];
  assign data_masked[8773] = data_i[8773] & sel_one_hot_i[68];
  assign data_masked[8772] = data_i[8772] & sel_one_hot_i[68];
  assign data_masked[8771] = data_i[8771] & sel_one_hot_i[68];
  assign data_masked[8770] = data_i[8770] & sel_one_hot_i[68];
  assign data_masked[8769] = data_i[8769] & sel_one_hot_i[68];
  assign data_masked[8768] = data_i[8768] & sel_one_hot_i[68];
  assign data_masked[8767] = data_i[8767] & sel_one_hot_i[68];
  assign data_masked[8766] = data_i[8766] & sel_one_hot_i[68];
  assign data_masked[8765] = data_i[8765] & sel_one_hot_i[68];
  assign data_masked[8764] = data_i[8764] & sel_one_hot_i[68];
  assign data_masked[8763] = data_i[8763] & sel_one_hot_i[68];
  assign data_masked[8762] = data_i[8762] & sel_one_hot_i[68];
  assign data_masked[8761] = data_i[8761] & sel_one_hot_i[68];
  assign data_masked[8760] = data_i[8760] & sel_one_hot_i[68];
  assign data_masked[8759] = data_i[8759] & sel_one_hot_i[68];
  assign data_masked[8758] = data_i[8758] & sel_one_hot_i[68];
  assign data_masked[8757] = data_i[8757] & sel_one_hot_i[68];
  assign data_masked[8756] = data_i[8756] & sel_one_hot_i[68];
  assign data_masked[8755] = data_i[8755] & sel_one_hot_i[68];
  assign data_masked[8754] = data_i[8754] & sel_one_hot_i[68];
  assign data_masked[8753] = data_i[8753] & sel_one_hot_i[68];
  assign data_masked[8752] = data_i[8752] & sel_one_hot_i[68];
  assign data_masked[8751] = data_i[8751] & sel_one_hot_i[68];
  assign data_masked[8750] = data_i[8750] & sel_one_hot_i[68];
  assign data_masked[8749] = data_i[8749] & sel_one_hot_i[68];
  assign data_masked[8748] = data_i[8748] & sel_one_hot_i[68];
  assign data_masked[8747] = data_i[8747] & sel_one_hot_i[68];
  assign data_masked[8746] = data_i[8746] & sel_one_hot_i[68];
  assign data_masked[8745] = data_i[8745] & sel_one_hot_i[68];
  assign data_masked[8744] = data_i[8744] & sel_one_hot_i[68];
  assign data_masked[8743] = data_i[8743] & sel_one_hot_i[68];
  assign data_masked[8742] = data_i[8742] & sel_one_hot_i[68];
  assign data_masked[8741] = data_i[8741] & sel_one_hot_i[68];
  assign data_masked[8740] = data_i[8740] & sel_one_hot_i[68];
  assign data_masked[8739] = data_i[8739] & sel_one_hot_i[68];
  assign data_masked[8738] = data_i[8738] & sel_one_hot_i[68];
  assign data_masked[8737] = data_i[8737] & sel_one_hot_i[68];
  assign data_masked[8736] = data_i[8736] & sel_one_hot_i[68];
  assign data_masked[8735] = data_i[8735] & sel_one_hot_i[68];
  assign data_masked[8734] = data_i[8734] & sel_one_hot_i[68];
  assign data_masked[8733] = data_i[8733] & sel_one_hot_i[68];
  assign data_masked[8732] = data_i[8732] & sel_one_hot_i[68];
  assign data_masked[8731] = data_i[8731] & sel_one_hot_i[68];
  assign data_masked[8730] = data_i[8730] & sel_one_hot_i[68];
  assign data_masked[8729] = data_i[8729] & sel_one_hot_i[68];
  assign data_masked[8728] = data_i[8728] & sel_one_hot_i[68];
  assign data_masked[8727] = data_i[8727] & sel_one_hot_i[68];
  assign data_masked[8726] = data_i[8726] & sel_one_hot_i[68];
  assign data_masked[8725] = data_i[8725] & sel_one_hot_i[68];
  assign data_masked[8724] = data_i[8724] & sel_one_hot_i[68];
  assign data_masked[8723] = data_i[8723] & sel_one_hot_i[68];
  assign data_masked[8722] = data_i[8722] & sel_one_hot_i[68];
  assign data_masked[8721] = data_i[8721] & sel_one_hot_i[68];
  assign data_masked[8720] = data_i[8720] & sel_one_hot_i[68];
  assign data_masked[8719] = data_i[8719] & sel_one_hot_i[68];
  assign data_masked[8718] = data_i[8718] & sel_one_hot_i[68];
  assign data_masked[8717] = data_i[8717] & sel_one_hot_i[68];
  assign data_masked[8716] = data_i[8716] & sel_one_hot_i[68];
  assign data_masked[8715] = data_i[8715] & sel_one_hot_i[68];
  assign data_masked[8714] = data_i[8714] & sel_one_hot_i[68];
  assign data_masked[8713] = data_i[8713] & sel_one_hot_i[68];
  assign data_masked[8712] = data_i[8712] & sel_one_hot_i[68];
  assign data_masked[8711] = data_i[8711] & sel_one_hot_i[68];
  assign data_masked[8710] = data_i[8710] & sel_one_hot_i[68];
  assign data_masked[8709] = data_i[8709] & sel_one_hot_i[68];
  assign data_masked[8708] = data_i[8708] & sel_one_hot_i[68];
  assign data_masked[8707] = data_i[8707] & sel_one_hot_i[68];
  assign data_masked[8706] = data_i[8706] & sel_one_hot_i[68];
  assign data_masked[8705] = data_i[8705] & sel_one_hot_i[68];
  assign data_masked[8704] = data_i[8704] & sel_one_hot_i[68];
  assign data_masked[8959] = data_i[8959] & sel_one_hot_i[69];
  assign data_masked[8958] = data_i[8958] & sel_one_hot_i[69];
  assign data_masked[8957] = data_i[8957] & sel_one_hot_i[69];
  assign data_masked[8956] = data_i[8956] & sel_one_hot_i[69];
  assign data_masked[8955] = data_i[8955] & sel_one_hot_i[69];
  assign data_masked[8954] = data_i[8954] & sel_one_hot_i[69];
  assign data_masked[8953] = data_i[8953] & sel_one_hot_i[69];
  assign data_masked[8952] = data_i[8952] & sel_one_hot_i[69];
  assign data_masked[8951] = data_i[8951] & sel_one_hot_i[69];
  assign data_masked[8950] = data_i[8950] & sel_one_hot_i[69];
  assign data_masked[8949] = data_i[8949] & sel_one_hot_i[69];
  assign data_masked[8948] = data_i[8948] & sel_one_hot_i[69];
  assign data_masked[8947] = data_i[8947] & sel_one_hot_i[69];
  assign data_masked[8946] = data_i[8946] & sel_one_hot_i[69];
  assign data_masked[8945] = data_i[8945] & sel_one_hot_i[69];
  assign data_masked[8944] = data_i[8944] & sel_one_hot_i[69];
  assign data_masked[8943] = data_i[8943] & sel_one_hot_i[69];
  assign data_masked[8942] = data_i[8942] & sel_one_hot_i[69];
  assign data_masked[8941] = data_i[8941] & sel_one_hot_i[69];
  assign data_masked[8940] = data_i[8940] & sel_one_hot_i[69];
  assign data_masked[8939] = data_i[8939] & sel_one_hot_i[69];
  assign data_masked[8938] = data_i[8938] & sel_one_hot_i[69];
  assign data_masked[8937] = data_i[8937] & sel_one_hot_i[69];
  assign data_masked[8936] = data_i[8936] & sel_one_hot_i[69];
  assign data_masked[8935] = data_i[8935] & sel_one_hot_i[69];
  assign data_masked[8934] = data_i[8934] & sel_one_hot_i[69];
  assign data_masked[8933] = data_i[8933] & sel_one_hot_i[69];
  assign data_masked[8932] = data_i[8932] & sel_one_hot_i[69];
  assign data_masked[8931] = data_i[8931] & sel_one_hot_i[69];
  assign data_masked[8930] = data_i[8930] & sel_one_hot_i[69];
  assign data_masked[8929] = data_i[8929] & sel_one_hot_i[69];
  assign data_masked[8928] = data_i[8928] & sel_one_hot_i[69];
  assign data_masked[8927] = data_i[8927] & sel_one_hot_i[69];
  assign data_masked[8926] = data_i[8926] & sel_one_hot_i[69];
  assign data_masked[8925] = data_i[8925] & sel_one_hot_i[69];
  assign data_masked[8924] = data_i[8924] & sel_one_hot_i[69];
  assign data_masked[8923] = data_i[8923] & sel_one_hot_i[69];
  assign data_masked[8922] = data_i[8922] & sel_one_hot_i[69];
  assign data_masked[8921] = data_i[8921] & sel_one_hot_i[69];
  assign data_masked[8920] = data_i[8920] & sel_one_hot_i[69];
  assign data_masked[8919] = data_i[8919] & sel_one_hot_i[69];
  assign data_masked[8918] = data_i[8918] & sel_one_hot_i[69];
  assign data_masked[8917] = data_i[8917] & sel_one_hot_i[69];
  assign data_masked[8916] = data_i[8916] & sel_one_hot_i[69];
  assign data_masked[8915] = data_i[8915] & sel_one_hot_i[69];
  assign data_masked[8914] = data_i[8914] & sel_one_hot_i[69];
  assign data_masked[8913] = data_i[8913] & sel_one_hot_i[69];
  assign data_masked[8912] = data_i[8912] & sel_one_hot_i[69];
  assign data_masked[8911] = data_i[8911] & sel_one_hot_i[69];
  assign data_masked[8910] = data_i[8910] & sel_one_hot_i[69];
  assign data_masked[8909] = data_i[8909] & sel_one_hot_i[69];
  assign data_masked[8908] = data_i[8908] & sel_one_hot_i[69];
  assign data_masked[8907] = data_i[8907] & sel_one_hot_i[69];
  assign data_masked[8906] = data_i[8906] & sel_one_hot_i[69];
  assign data_masked[8905] = data_i[8905] & sel_one_hot_i[69];
  assign data_masked[8904] = data_i[8904] & sel_one_hot_i[69];
  assign data_masked[8903] = data_i[8903] & sel_one_hot_i[69];
  assign data_masked[8902] = data_i[8902] & sel_one_hot_i[69];
  assign data_masked[8901] = data_i[8901] & sel_one_hot_i[69];
  assign data_masked[8900] = data_i[8900] & sel_one_hot_i[69];
  assign data_masked[8899] = data_i[8899] & sel_one_hot_i[69];
  assign data_masked[8898] = data_i[8898] & sel_one_hot_i[69];
  assign data_masked[8897] = data_i[8897] & sel_one_hot_i[69];
  assign data_masked[8896] = data_i[8896] & sel_one_hot_i[69];
  assign data_masked[8895] = data_i[8895] & sel_one_hot_i[69];
  assign data_masked[8894] = data_i[8894] & sel_one_hot_i[69];
  assign data_masked[8893] = data_i[8893] & sel_one_hot_i[69];
  assign data_masked[8892] = data_i[8892] & sel_one_hot_i[69];
  assign data_masked[8891] = data_i[8891] & sel_one_hot_i[69];
  assign data_masked[8890] = data_i[8890] & sel_one_hot_i[69];
  assign data_masked[8889] = data_i[8889] & sel_one_hot_i[69];
  assign data_masked[8888] = data_i[8888] & sel_one_hot_i[69];
  assign data_masked[8887] = data_i[8887] & sel_one_hot_i[69];
  assign data_masked[8886] = data_i[8886] & sel_one_hot_i[69];
  assign data_masked[8885] = data_i[8885] & sel_one_hot_i[69];
  assign data_masked[8884] = data_i[8884] & sel_one_hot_i[69];
  assign data_masked[8883] = data_i[8883] & sel_one_hot_i[69];
  assign data_masked[8882] = data_i[8882] & sel_one_hot_i[69];
  assign data_masked[8881] = data_i[8881] & sel_one_hot_i[69];
  assign data_masked[8880] = data_i[8880] & sel_one_hot_i[69];
  assign data_masked[8879] = data_i[8879] & sel_one_hot_i[69];
  assign data_masked[8878] = data_i[8878] & sel_one_hot_i[69];
  assign data_masked[8877] = data_i[8877] & sel_one_hot_i[69];
  assign data_masked[8876] = data_i[8876] & sel_one_hot_i[69];
  assign data_masked[8875] = data_i[8875] & sel_one_hot_i[69];
  assign data_masked[8874] = data_i[8874] & sel_one_hot_i[69];
  assign data_masked[8873] = data_i[8873] & sel_one_hot_i[69];
  assign data_masked[8872] = data_i[8872] & sel_one_hot_i[69];
  assign data_masked[8871] = data_i[8871] & sel_one_hot_i[69];
  assign data_masked[8870] = data_i[8870] & sel_one_hot_i[69];
  assign data_masked[8869] = data_i[8869] & sel_one_hot_i[69];
  assign data_masked[8868] = data_i[8868] & sel_one_hot_i[69];
  assign data_masked[8867] = data_i[8867] & sel_one_hot_i[69];
  assign data_masked[8866] = data_i[8866] & sel_one_hot_i[69];
  assign data_masked[8865] = data_i[8865] & sel_one_hot_i[69];
  assign data_masked[8864] = data_i[8864] & sel_one_hot_i[69];
  assign data_masked[8863] = data_i[8863] & sel_one_hot_i[69];
  assign data_masked[8862] = data_i[8862] & sel_one_hot_i[69];
  assign data_masked[8861] = data_i[8861] & sel_one_hot_i[69];
  assign data_masked[8860] = data_i[8860] & sel_one_hot_i[69];
  assign data_masked[8859] = data_i[8859] & sel_one_hot_i[69];
  assign data_masked[8858] = data_i[8858] & sel_one_hot_i[69];
  assign data_masked[8857] = data_i[8857] & sel_one_hot_i[69];
  assign data_masked[8856] = data_i[8856] & sel_one_hot_i[69];
  assign data_masked[8855] = data_i[8855] & sel_one_hot_i[69];
  assign data_masked[8854] = data_i[8854] & sel_one_hot_i[69];
  assign data_masked[8853] = data_i[8853] & sel_one_hot_i[69];
  assign data_masked[8852] = data_i[8852] & sel_one_hot_i[69];
  assign data_masked[8851] = data_i[8851] & sel_one_hot_i[69];
  assign data_masked[8850] = data_i[8850] & sel_one_hot_i[69];
  assign data_masked[8849] = data_i[8849] & sel_one_hot_i[69];
  assign data_masked[8848] = data_i[8848] & sel_one_hot_i[69];
  assign data_masked[8847] = data_i[8847] & sel_one_hot_i[69];
  assign data_masked[8846] = data_i[8846] & sel_one_hot_i[69];
  assign data_masked[8845] = data_i[8845] & sel_one_hot_i[69];
  assign data_masked[8844] = data_i[8844] & sel_one_hot_i[69];
  assign data_masked[8843] = data_i[8843] & sel_one_hot_i[69];
  assign data_masked[8842] = data_i[8842] & sel_one_hot_i[69];
  assign data_masked[8841] = data_i[8841] & sel_one_hot_i[69];
  assign data_masked[8840] = data_i[8840] & sel_one_hot_i[69];
  assign data_masked[8839] = data_i[8839] & sel_one_hot_i[69];
  assign data_masked[8838] = data_i[8838] & sel_one_hot_i[69];
  assign data_masked[8837] = data_i[8837] & sel_one_hot_i[69];
  assign data_masked[8836] = data_i[8836] & sel_one_hot_i[69];
  assign data_masked[8835] = data_i[8835] & sel_one_hot_i[69];
  assign data_masked[8834] = data_i[8834] & sel_one_hot_i[69];
  assign data_masked[8833] = data_i[8833] & sel_one_hot_i[69];
  assign data_masked[8832] = data_i[8832] & sel_one_hot_i[69];
  assign data_masked[9087] = data_i[9087] & sel_one_hot_i[70];
  assign data_masked[9086] = data_i[9086] & sel_one_hot_i[70];
  assign data_masked[9085] = data_i[9085] & sel_one_hot_i[70];
  assign data_masked[9084] = data_i[9084] & sel_one_hot_i[70];
  assign data_masked[9083] = data_i[9083] & sel_one_hot_i[70];
  assign data_masked[9082] = data_i[9082] & sel_one_hot_i[70];
  assign data_masked[9081] = data_i[9081] & sel_one_hot_i[70];
  assign data_masked[9080] = data_i[9080] & sel_one_hot_i[70];
  assign data_masked[9079] = data_i[9079] & sel_one_hot_i[70];
  assign data_masked[9078] = data_i[9078] & sel_one_hot_i[70];
  assign data_masked[9077] = data_i[9077] & sel_one_hot_i[70];
  assign data_masked[9076] = data_i[9076] & sel_one_hot_i[70];
  assign data_masked[9075] = data_i[9075] & sel_one_hot_i[70];
  assign data_masked[9074] = data_i[9074] & sel_one_hot_i[70];
  assign data_masked[9073] = data_i[9073] & sel_one_hot_i[70];
  assign data_masked[9072] = data_i[9072] & sel_one_hot_i[70];
  assign data_masked[9071] = data_i[9071] & sel_one_hot_i[70];
  assign data_masked[9070] = data_i[9070] & sel_one_hot_i[70];
  assign data_masked[9069] = data_i[9069] & sel_one_hot_i[70];
  assign data_masked[9068] = data_i[9068] & sel_one_hot_i[70];
  assign data_masked[9067] = data_i[9067] & sel_one_hot_i[70];
  assign data_masked[9066] = data_i[9066] & sel_one_hot_i[70];
  assign data_masked[9065] = data_i[9065] & sel_one_hot_i[70];
  assign data_masked[9064] = data_i[9064] & sel_one_hot_i[70];
  assign data_masked[9063] = data_i[9063] & sel_one_hot_i[70];
  assign data_masked[9062] = data_i[9062] & sel_one_hot_i[70];
  assign data_masked[9061] = data_i[9061] & sel_one_hot_i[70];
  assign data_masked[9060] = data_i[9060] & sel_one_hot_i[70];
  assign data_masked[9059] = data_i[9059] & sel_one_hot_i[70];
  assign data_masked[9058] = data_i[9058] & sel_one_hot_i[70];
  assign data_masked[9057] = data_i[9057] & sel_one_hot_i[70];
  assign data_masked[9056] = data_i[9056] & sel_one_hot_i[70];
  assign data_masked[9055] = data_i[9055] & sel_one_hot_i[70];
  assign data_masked[9054] = data_i[9054] & sel_one_hot_i[70];
  assign data_masked[9053] = data_i[9053] & sel_one_hot_i[70];
  assign data_masked[9052] = data_i[9052] & sel_one_hot_i[70];
  assign data_masked[9051] = data_i[9051] & sel_one_hot_i[70];
  assign data_masked[9050] = data_i[9050] & sel_one_hot_i[70];
  assign data_masked[9049] = data_i[9049] & sel_one_hot_i[70];
  assign data_masked[9048] = data_i[9048] & sel_one_hot_i[70];
  assign data_masked[9047] = data_i[9047] & sel_one_hot_i[70];
  assign data_masked[9046] = data_i[9046] & sel_one_hot_i[70];
  assign data_masked[9045] = data_i[9045] & sel_one_hot_i[70];
  assign data_masked[9044] = data_i[9044] & sel_one_hot_i[70];
  assign data_masked[9043] = data_i[9043] & sel_one_hot_i[70];
  assign data_masked[9042] = data_i[9042] & sel_one_hot_i[70];
  assign data_masked[9041] = data_i[9041] & sel_one_hot_i[70];
  assign data_masked[9040] = data_i[9040] & sel_one_hot_i[70];
  assign data_masked[9039] = data_i[9039] & sel_one_hot_i[70];
  assign data_masked[9038] = data_i[9038] & sel_one_hot_i[70];
  assign data_masked[9037] = data_i[9037] & sel_one_hot_i[70];
  assign data_masked[9036] = data_i[9036] & sel_one_hot_i[70];
  assign data_masked[9035] = data_i[9035] & sel_one_hot_i[70];
  assign data_masked[9034] = data_i[9034] & sel_one_hot_i[70];
  assign data_masked[9033] = data_i[9033] & sel_one_hot_i[70];
  assign data_masked[9032] = data_i[9032] & sel_one_hot_i[70];
  assign data_masked[9031] = data_i[9031] & sel_one_hot_i[70];
  assign data_masked[9030] = data_i[9030] & sel_one_hot_i[70];
  assign data_masked[9029] = data_i[9029] & sel_one_hot_i[70];
  assign data_masked[9028] = data_i[9028] & sel_one_hot_i[70];
  assign data_masked[9027] = data_i[9027] & sel_one_hot_i[70];
  assign data_masked[9026] = data_i[9026] & sel_one_hot_i[70];
  assign data_masked[9025] = data_i[9025] & sel_one_hot_i[70];
  assign data_masked[9024] = data_i[9024] & sel_one_hot_i[70];
  assign data_masked[9023] = data_i[9023] & sel_one_hot_i[70];
  assign data_masked[9022] = data_i[9022] & sel_one_hot_i[70];
  assign data_masked[9021] = data_i[9021] & sel_one_hot_i[70];
  assign data_masked[9020] = data_i[9020] & sel_one_hot_i[70];
  assign data_masked[9019] = data_i[9019] & sel_one_hot_i[70];
  assign data_masked[9018] = data_i[9018] & sel_one_hot_i[70];
  assign data_masked[9017] = data_i[9017] & sel_one_hot_i[70];
  assign data_masked[9016] = data_i[9016] & sel_one_hot_i[70];
  assign data_masked[9015] = data_i[9015] & sel_one_hot_i[70];
  assign data_masked[9014] = data_i[9014] & sel_one_hot_i[70];
  assign data_masked[9013] = data_i[9013] & sel_one_hot_i[70];
  assign data_masked[9012] = data_i[9012] & sel_one_hot_i[70];
  assign data_masked[9011] = data_i[9011] & sel_one_hot_i[70];
  assign data_masked[9010] = data_i[9010] & sel_one_hot_i[70];
  assign data_masked[9009] = data_i[9009] & sel_one_hot_i[70];
  assign data_masked[9008] = data_i[9008] & sel_one_hot_i[70];
  assign data_masked[9007] = data_i[9007] & sel_one_hot_i[70];
  assign data_masked[9006] = data_i[9006] & sel_one_hot_i[70];
  assign data_masked[9005] = data_i[9005] & sel_one_hot_i[70];
  assign data_masked[9004] = data_i[9004] & sel_one_hot_i[70];
  assign data_masked[9003] = data_i[9003] & sel_one_hot_i[70];
  assign data_masked[9002] = data_i[9002] & sel_one_hot_i[70];
  assign data_masked[9001] = data_i[9001] & sel_one_hot_i[70];
  assign data_masked[9000] = data_i[9000] & sel_one_hot_i[70];
  assign data_masked[8999] = data_i[8999] & sel_one_hot_i[70];
  assign data_masked[8998] = data_i[8998] & sel_one_hot_i[70];
  assign data_masked[8997] = data_i[8997] & sel_one_hot_i[70];
  assign data_masked[8996] = data_i[8996] & sel_one_hot_i[70];
  assign data_masked[8995] = data_i[8995] & sel_one_hot_i[70];
  assign data_masked[8994] = data_i[8994] & sel_one_hot_i[70];
  assign data_masked[8993] = data_i[8993] & sel_one_hot_i[70];
  assign data_masked[8992] = data_i[8992] & sel_one_hot_i[70];
  assign data_masked[8991] = data_i[8991] & sel_one_hot_i[70];
  assign data_masked[8990] = data_i[8990] & sel_one_hot_i[70];
  assign data_masked[8989] = data_i[8989] & sel_one_hot_i[70];
  assign data_masked[8988] = data_i[8988] & sel_one_hot_i[70];
  assign data_masked[8987] = data_i[8987] & sel_one_hot_i[70];
  assign data_masked[8986] = data_i[8986] & sel_one_hot_i[70];
  assign data_masked[8985] = data_i[8985] & sel_one_hot_i[70];
  assign data_masked[8984] = data_i[8984] & sel_one_hot_i[70];
  assign data_masked[8983] = data_i[8983] & sel_one_hot_i[70];
  assign data_masked[8982] = data_i[8982] & sel_one_hot_i[70];
  assign data_masked[8981] = data_i[8981] & sel_one_hot_i[70];
  assign data_masked[8980] = data_i[8980] & sel_one_hot_i[70];
  assign data_masked[8979] = data_i[8979] & sel_one_hot_i[70];
  assign data_masked[8978] = data_i[8978] & sel_one_hot_i[70];
  assign data_masked[8977] = data_i[8977] & sel_one_hot_i[70];
  assign data_masked[8976] = data_i[8976] & sel_one_hot_i[70];
  assign data_masked[8975] = data_i[8975] & sel_one_hot_i[70];
  assign data_masked[8974] = data_i[8974] & sel_one_hot_i[70];
  assign data_masked[8973] = data_i[8973] & sel_one_hot_i[70];
  assign data_masked[8972] = data_i[8972] & sel_one_hot_i[70];
  assign data_masked[8971] = data_i[8971] & sel_one_hot_i[70];
  assign data_masked[8970] = data_i[8970] & sel_one_hot_i[70];
  assign data_masked[8969] = data_i[8969] & sel_one_hot_i[70];
  assign data_masked[8968] = data_i[8968] & sel_one_hot_i[70];
  assign data_masked[8967] = data_i[8967] & sel_one_hot_i[70];
  assign data_masked[8966] = data_i[8966] & sel_one_hot_i[70];
  assign data_masked[8965] = data_i[8965] & sel_one_hot_i[70];
  assign data_masked[8964] = data_i[8964] & sel_one_hot_i[70];
  assign data_masked[8963] = data_i[8963] & sel_one_hot_i[70];
  assign data_masked[8962] = data_i[8962] & sel_one_hot_i[70];
  assign data_masked[8961] = data_i[8961] & sel_one_hot_i[70];
  assign data_masked[8960] = data_i[8960] & sel_one_hot_i[70];
  assign data_masked[9215] = data_i[9215] & sel_one_hot_i[71];
  assign data_masked[9214] = data_i[9214] & sel_one_hot_i[71];
  assign data_masked[9213] = data_i[9213] & sel_one_hot_i[71];
  assign data_masked[9212] = data_i[9212] & sel_one_hot_i[71];
  assign data_masked[9211] = data_i[9211] & sel_one_hot_i[71];
  assign data_masked[9210] = data_i[9210] & sel_one_hot_i[71];
  assign data_masked[9209] = data_i[9209] & sel_one_hot_i[71];
  assign data_masked[9208] = data_i[9208] & sel_one_hot_i[71];
  assign data_masked[9207] = data_i[9207] & sel_one_hot_i[71];
  assign data_masked[9206] = data_i[9206] & sel_one_hot_i[71];
  assign data_masked[9205] = data_i[9205] & sel_one_hot_i[71];
  assign data_masked[9204] = data_i[9204] & sel_one_hot_i[71];
  assign data_masked[9203] = data_i[9203] & sel_one_hot_i[71];
  assign data_masked[9202] = data_i[9202] & sel_one_hot_i[71];
  assign data_masked[9201] = data_i[9201] & sel_one_hot_i[71];
  assign data_masked[9200] = data_i[9200] & sel_one_hot_i[71];
  assign data_masked[9199] = data_i[9199] & sel_one_hot_i[71];
  assign data_masked[9198] = data_i[9198] & sel_one_hot_i[71];
  assign data_masked[9197] = data_i[9197] & sel_one_hot_i[71];
  assign data_masked[9196] = data_i[9196] & sel_one_hot_i[71];
  assign data_masked[9195] = data_i[9195] & sel_one_hot_i[71];
  assign data_masked[9194] = data_i[9194] & sel_one_hot_i[71];
  assign data_masked[9193] = data_i[9193] & sel_one_hot_i[71];
  assign data_masked[9192] = data_i[9192] & sel_one_hot_i[71];
  assign data_masked[9191] = data_i[9191] & sel_one_hot_i[71];
  assign data_masked[9190] = data_i[9190] & sel_one_hot_i[71];
  assign data_masked[9189] = data_i[9189] & sel_one_hot_i[71];
  assign data_masked[9188] = data_i[9188] & sel_one_hot_i[71];
  assign data_masked[9187] = data_i[9187] & sel_one_hot_i[71];
  assign data_masked[9186] = data_i[9186] & sel_one_hot_i[71];
  assign data_masked[9185] = data_i[9185] & sel_one_hot_i[71];
  assign data_masked[9184] = data_i[9184] & sel_one_hot_i[71];
  assign data_masked[9183] = data_i[9183] & sel_one_hot_i[71];
  assign data_masked[9182] = data_i[9182] & sel_one_hot_i[71];
  assign data_masked[9181] = data_i[9181] & sel_one_hot_i[71];
  assign data_masked[9180] = data_i[9180] & sel_one_hot_i[71];
  assign data_masked[9179] = data_i[9179] & sel_one_hot_i[71];
  assign data_masked[9178] = data_i[9178] & sel_one_hot_i[71];
  assign data_masked[9177] = data_i[9177] & sel_one_hot_i[71];
  assign data_masked[9176] = data_i[9176] & sel_one_hot_i[71];
  assign data_masked[9175] = data_i[9175] & sel_one_hot_i[71];
  assign data_masked[9174] = data_i[9174] & sel_one_hot_i[71];
  assign data_masked[9173] = data_i[9173] & sel_one_hot_i[71];
  assign data_masked[9172] = data_i[9172] & sel_one_hot_i[71];
  assign data_masked[9171] = data_i[9171] & sel_one_hot_i[71];
  assign data_masked[9170] = data_i[9170] & sel_one_hot_i[71];
  assign data_masked[9169] = data_i[9169] & sel_one_hot_i[71];
  assign data_masked[9168] = data_i[9168] & sel_one_hot_i[71];
  assign data_masked[9167] = data_i[9167] & sel_one_hot_i[71];
  assign data_masked[9166] = data_i[9166] & sel_one_hot_i[71];
  assign data_masked[9165] = data_i[9165] & sel_one_hot_i[71];
  assign data_masked[9164] = data_i[9164] & sel_one_hot_i[71];
  assign data_masked[9163] = data_i[9163] & sel_one_hot_i[71];
  assign data_masked[9162] = data_i[9162] & sel_one_hot_i[71];
  assign data_masked[9161] = data_i[9161] & sel_one_hot_i[71];
  assign data_masked[9160] = data_i[9160] & sel_one_hot_i[71];
  assign data_masked[9159] = data_i[9159] & sel_one_hot_i[71];
  assign data_masked[9158] = data_i[9158] & sel_one_hot_i[71];
  assign data_masked[9157] = data_i[9157] & sel_one_hot_i[71];
  assign data_masked[9156] = data_i[9156] & sel_one_hot_i[71];
  assign data_masked[9155] = data_i[9155] & sel_one_hot_i[71];
  assign data_masked[9154] = data_i[9154] & sel_one_hot_i[71];
  assign data_masked[9153] = data_i[9153] & sel_one_hot_i[71];
  assign data_masked[9152] = data_i[9152] & sel_one_hot_i[71];
  assign data_masked[9151] = data_i[9151] & sel_one_hot_i[71];
  assign data_masked[9150] = data_i[9150] & sel_one_hot_i[71];
  assign data_masked[9149] = data_i[9149] & sel_one_hot_i[71];
  assign data_masked[9148] = data_i[9148] & sel_one_hot_i[71];
  assign data_masked[9147] = data_i[9147] & sel_one_hot_i[71];
  assign data_masked[9146] = data_i[9146] & sel_one_hot_i[71];
  assign data_masked[9145] = data_i[9145] & sel_one_hot_i[71];
  assign data_masked[9144] = data_i[9144] & sel_one_hot_i[71];
  assign data_masked[9143] = data_i[9143] & sel_one_hot_i[71];
  assign data_masked[9142] = data_i[9142] & sel_one_hot_i[71];
  assign data_masked[9141] = data_i[9141] & sel_one_hot_i[71];
  assign data_masked[9140] = data_i[9140] & sel_one_hot_i[71];
  assign data_masked[9139] = data_i[9139] & sel_one_hot_i[71];
  assign data_masked[9138] = data_i[9138] & sel_one_hot_i[71];
  assign data_masked[9137] = data_i[9137] & sel_one_hot_i[71];
  assign data_masked[9136] = data_i[9136] & sel_one_hot_i[71];
  assign data_masked[9135] = data_i[9135] & sel_one_hot_i[71];
  assign data_masked[9134] = data_i[9134] & sel_one_hot_i[71];
  assign data_masked[9133] = data_i[9133] & sel_one_hot_i[71];
  assign data_masked[9132] = data_i[9132] & sel_one_hot_i[71];
  assign data_masked[9131] = data_i[9131] & sel_one_hot_i[71];
  assign data_masked[9130] = data_i[9130] & sel_one_hot_i[71];
  assign data_masked[9129] = data_i[9129] & sel_one_hot_i[71];
  assign data_masked[9128] = data_i[9128] & sel_one_hot_i[71];
  assign data_masked[9127] = data_i[9127] & sel_one_hot_i[71];
  assign data_masked[9126] = data_i[9126] & sel_one_hot_i[71];
  assign data_masked[9125] = data_i[9125] & sel_one_hot_i[71];
  assign data_masked[9124] = data_i[9124] & sel_one_hot_i[71];
  assign data_masked[9123] = data_i[9123] & sel_one_hot_i[71];
  assign data_masked[9122] = data_i[9122] & sel_one_hot_i[71];
  assign data_masked[9121] = data_i[9121] & sel_one_hot_i[71];
  assign data_masked[9120] = data_i[9120] & sel_one_hot_i[71];
  assign data_masked[9119] = data_i[9119] & sel_one_hot_i[71];
  assign data_masked[9118] = data_i[9118] & sel_one_hot_i[71];
  assign data_masked[9117] = data_i[9117] & sel_one_hot_i[71];
  assign data_masked[9116] = data_i[9116] & sel_one_hot_i[71];
  assign data_masked[9115] = data_i[9115] & sel_one_hot_i[71];
  assign data_masked[9114] = data_i[9114] & sel_one_hot_i[71];
  assign data_masked[9113] = data_i[9113] & sel_one_hot_i[71];
  assign data_masked[9112] = data_i[9112] & sel_one_hot_i[71];
  assign data_masked[9111] = data_i[9111] & sel_one_hot_i[71];
  assign data_masked[9110] = data_i[9110] & sel_one_hot_i[71];
  assign data_masked[9109] = data_i[9109] & sel_one_hot_i[71];
  assign data_masked[9108] = data_i[9108] & sel_one_hot_i[71];
  assign data_masked[9107] = data_i[9107] & sel_one_hot_i[71];
  assign data_masked[9106] = data_i[9106] & sel_one_hot_i[71];
  assign data_masked[9105] = data_i[9105] & sel_one_hot_i[71];
  assign data_masked[9104] = data_i[9104] & sel_one_hot_i[71];
  assign data_masked[9103] = data_i[9103] & sel_one_hot_i[71];
  assign data_masked[9102] = data_i[9102] & sel_one_hot_i[71];
  assign data_masked[9101] = data_i[9101] & sel_one_hot_i[71];
  assign data_masked[9100] = data_i[9100] & sel_one_hot_i[71];
  assign data_masked[9099] = data_i[9099] & sel_one_hot_i[71];
  assign data_masked[9098] = data_i[9098] & sel_one_hot_i[71];
  assign data_masked[9097] = data_i[9097] & sel_one_hot_i[71];
  assign data_masked[9096] = data_i[9096] & sel_one_hot_i[71];
  assign data_masked[9095] = data_i[9095] & sel_one_hot_i[71];
  assign data_masked[9094] = data_i[9094] & sel_one_hot_i[71];
  assign data_masked[9093] = data_i[9093] & sel_one_hot_i[71];
  assign data_masked[9092] = data_i[9092] & sel_one_hot_i[71];
  assign data_masked[9091] = data_i[9091] & sel_one_hot_i[71];
  assign data_masked[9090] = data_i[9090] & sel_one_hot_i[71];
  assign data_masked[9089] = data_i[9089] & sel_one_hot_i[71];
  assign data_masked[9088] = data_i[9088] & sel_one_hot_i[71];
  assign data_masked[9343] = data_i[9343] & sel_one_hot_i[72];
  assign data_masked[9342] = data_i[9342] & sel_one_hot_i[72];
  assign data_masked[9341] = data_i[9341] & sel_one_hot_i[72];
  assign data_masked[9340] = data_i[9340] & sel_one_hot_i[72];
  assign data_masked[9339] = data_i[9339] & sel_one_hot_i[72];
  assign data_masked[9338] = data_i[9338] & sel_one_hot_i[72];
  assign data_masked[9337] = data_i[9337] & sel_one_hot_i[72];
  assign data_masked[9336] = data_i[9336] & sel_one_hot_i[72];
  assign data_masked[9335] = data_i[9335] & sel_one_hot_i[72];
  assign data_masked[9334] = data_i[9334] & sel_one_hot_i[72];
  assign data_masked[9333] = data_i[9333] & sel_one_hot_i[72];
  assign data_masked[9332] = data_i[9332] & sel_one_hot_i[72];
  assign data_masked[9331] = data_i[9331] & sel_one_hot_i[72];
  assign data_masked[9330] = data_i[9330] & sel_one_hot_i[72];
  assign data_masked[9329] = data_i[9329] & sel_one_hot_i[72];
  assign data_masked[9328] = data_i[9328] & sel_one_hot_i[72];
  assign data_masked[9327] = data_i[9327] & sel_one_hot_i[72];
  assign data_masked[9326] = data_i[9326] & sel_one_hot_i[72];
  assign data_masked[9325] = data_i[9325] & sel_one_hot_i[72];
  assign data_masked[9324] = data_i[9324] & sel_one_hot_i[72];
  assign data_masked[9323] = data_i[9323] & sel_one_hot_i[72];
  assign data_masked[9322] = data_i[9322] & sel_one_hot_i[72];
  assign data_masked[9321] = data_i[9321] & sel_one_hot_i[72];
  assign data_masked[9320] = data_i[9320] & sel_one_hot_i[72];
  assign data_masked[9319] = data_i[9319] & sel_one_hot_i[72];
  assign data_masked[9318] = data_i[9318] & sel_one_hot_i[72];
  assign data_masked[9317] = data_i[9317] & sel_one_hot_i[72];
  assign data_masked[9316] = data_i[9316] & sel_one_hot_i[72];
  assign data_masked[9315] = data_i[9315] & sel_one_hot_i[72];
  assign data_masked[9314] = data_i[9314] & sel_one_hot_i[72];
  assign data_masked[9313] = data_i[9313] & sel_one_hot_i[72];
  assign data_masked[9312] = data_i[9312] & sel_one_hot_i[72];
  assign data_masked[9311] = data_i[9311] & sel_one_hot_i[72];
  assign data_masked[9310] = data_i[9310] & sel_one_hot_i[72];
  assign data_masked[9309] = data_i[9309] & sel_one_hot_i[72];
  assign data_masked[9308] = data_i[9308] & sel_one_hot_i[72];
  assign data_masked[9307] = data_i[9307] & sel_one_hot_i[72];
  assign data_masked[9306] = data_i[9306] & sel_one_hot_i[72];
  assign data_masked[9305] = data_i[9305] & sel_one_hot_i[72];
  assign data_masked[9304] = data_i[9304] & sel_one_hot_i[72];
  assign data_masked[9303] = data_i[9303] & sel_one_hot_i[72];
  assign data_masked[9302] = data_i[9302] & sel_one_hot_i[72];
  assign data_masked[9301] = data_i[9301] & sel_one_hot_i[72];
  assign data_masked[9300] = data_i[9300] & sel_one_hot_i[72];
  assign data_masked[9299] = data_i[9299] & sel_one_hot_i[72];
  assign data_masked[9298] = data_i[9298] & sel_one_hot_i[72];
  assign data_masked[9297] = data_i[9297] & sel_one_hot_i[72];
  assign data_masked[9296] = data_i[9296] & sel_one_hot_i[72];
  assign data_masked[9295] = data_i[9295] & sel_one_hot_i[72];
  assign data_masked[9294] = data_i[9294] & sel_one_hot_i[72];
  assign data_masked[9293] = data_i[9293] & sel_one_hot_i[72];
  assign data_masked[9292] = data_i[9292] & sel_one_hot_i[72];
  assign data_masked[9291] = data_i[9291] & sel_one_hot_i[72];
  assign data_masked[9290] = data_i[9290] & sel_one_hot_i[72];
  assign data_masked[9289] = data_i[9289] & sel_one_hot_i[72];
  assign data_masked[9288] = data_i[9288] & sel_one_hot_i[72];
  assign data_masked[9287] = data_i[9287] & sel_one_hot_i[72];
  assign data_masked[9286] = data_i[9286] & sel_one_hot_i[72];
  assign data_masked[9285] = data_i[9285] & sel_one_hot_i[72];
  assign data_masked[9284] = data_i[9284] & sel_one_hot_i[72];
  assign data_masked[9283] = data_i[9283] & sel_one_hot_i[72];
  assign data_masked[9282] = data_i[9282] & sel_one_hot_i[72];
  assign data_masked[9281] = data_i[9281] & sel_one_hot_i[72];
  assign data_masked[9280] = data_i[9280] & sel_one_hot_i[72];
  assign data_masked[9279] = data_i[9279] & sel_one_hot_i[72];
  assign data_masked[9278] = data_i[9278] & sel_one_hot_i[72];
  assign data_masked[9277] = data_i[9277] & sel_one_hot_i[72];
  assign data_masked[9276] = data_i[9276] & sel_one_hot_i[72];
  assign data_masked[9275] = data_i[9275] & sel_one_hot_i[72];
  assign data_masked[9274] = data_i[9274] & sel_one_hot_i[72];
  assign data_masked[9273] = data_i[9273] & sel_one_hot_i[72];
  assign data_masked[9272] = data_i[9272] & sel_one_hot_i[72];
  assign data_masked[9271] = data_i[9271] & sel_one_hot_i[72];
  assign data_masked[9270] = data_i[9270] & sel_one_hot_i[72];
  assign data_masked[9269] = data_i[9269] & sel_one_hot_i[72];
  assign data_masked[9268] = data_i[9268] & sel_one_hot_i[72];
  assign data_masked[9267] = data_i[9267] & sel_one_hot_i[72];
  assign data_masked[9266] = data_i[9266] & sel_one_hot_i[72];
  assign data_masked[9265] = data_i[9265] & sel_one_hot_i[72];
  assign data_masked[9264] = data_i[9264] & sel_one_hot_i[72];
  assign data_masked[9263] = data_i[9263] & sel_one_hot_i[72];
  assign data_masked[9262] = data_i[9262] & sel_one_hot_i[72];
  assign data_masked[9261] = data_i[9261] & sel_one_hot_i[72];
  assign data_masked[9260] = data_i[9260] & sel_one_hot_i[72];
  assign data_masked[9259] = data_i[9259] & sel_one_hot_i[72];
  assign data_masked[9258] = data_i[9258] & sel_one_hot_i[72];
  assign data_masked[9257] = data_i[9257] & sel_one_hot_i[72];
  assign data_masked[9256] = data_i[9256] & sel_one_hot_i[72];
  assign data_masked[9255] = data_i[9255] & sel_one_hot_i[72];
  assign data_masked[9254] = data_i[9254] & sel_one_hot_i[72];
  assign data_masked[9253] = data_i[9253] & sel_one_hot_i[72];
  assign data_masked[9252] = data_i[9252] & sel_one_hot_i[72];
  assign data_masked[9251] = data_i[9251] & sel_one_hot_i[72];
  assign data_masked[9250] = data_i[9250] & sel_one_hot_i[72];
  assign data_masked[9249] = data_i[9249] & sel_one_hot_i[72];
  assign data_masked[9248] = data_i[9248] & sel_one_hot_i[72];
  assign data_masked[9247] = data_i[9247] & sel_one_hot_i[72];
  assign data_masked[9246] = data_i[9246] & sel_one_hot_i[72];
  assign data_masked[9245] = data_i[9245] & sel_one_hot_i[72];
  assign data_masked[9244] = data_i[9244] & sel_one_hot_i[72];
  assign data_masked[9243] = data_i[9243] & sel_one_hot_i[72];
  assign data_masked[9242] = data_i[9242] & sel_one_hot_i[72];
  assign data_masked[9241] = data_i[9241] & sel_one_hot_i[72];
  assign data_masked[9240] = data_i[9240] & sel_one_hot_i[72];
  assign data_masked[9239] = data_i[9239] & sel_one_hot_i[72];
  assign data_masked[9238] = data_i[9238] & sel_one_hot_i[72];
  assign data_masked[9237] = data_i[9237] & sel_one_hot_i[72];
  assign data_masked[9236] = data_i[9236] & sel_one_hot_i[72];
  assign data_masked[9235] = data_i[9235] & sel_one_hot_i[72];
  assign data_masked[9234] = data_i[9234] & sel_one_hot_i[72];
  assign data_masked[9233] = data_i[9233] & sel_one_hot_i[72];
  assign data_masked[9232] = data_i[9232] & sel_one_hot_i[72];
  assign data_masked[9231] = data_i[9231] & sel_one_hot_i[72];
  assign data_masked[9230] = data_i[9230] & sel_one_hot_i[72];
  assign data_masked[9229] = data_i[9229] & sel_one_hot_i[72];
  assign data_masked[9228] = data_i[9228] & sel_one_hot_i[72];
  assign data_masked[9227] = data_i[9227] & sel_one_hot_i[72];
  assign data_masked[9226] = data_i[9226] & sel_one_hot_i[72];
  assign data_masked[9225] = data_i[9225] & sel_one_hot_i[72];
  assign data_masked[9224] = data_i[9224] & sel_one_hot_i[72];
  assign data_masked[9223] = data_i[9223] & sel_one_hot_i[72];
  assign data_masked[9222] = data_i[9222] & sel_one_hot_i[72];
  assign data_masked[9221] = data_i[9221] & sel_one_hot_i[72];
  assign data_masked[9220] = data_i[9220] & sel_one_hot_i[72];
  assign data_masked[9219] = data_i[9219] & sel_one_hot_i[72];
  assign data_masked[9218] = data_i[9218] & sel_one_hot_i[72];
  assign data_masked[9217] = data_i[9217] & sel_one_hot_i[72];
  assign data_masked[9216] = data_i[9216] & sel_one_hot_i[72];
  assign data_masked[9471] = data_i[9471] & sel_one_hot_i[73];
  assign data_masked[9470] = data_i[9470] & sel_one_hot_i[73];
  assign data_masked[9469] = data_i[9469] & sel_one_hot_i[73];
  assign data_masked[9468] = data_i[9468] & sel_one_hot_i[73];
  assign data_masked[9467] = data_i[9467] & sel_one_hot_i[73];
  assign data_masked[9466] = data_i[9466] & sel_one_hot_i[73];
  assign data_masked[9465] = data_i[9465] & sel_one_hot_i[73];
  assign data_masked[9464] = data_i[9464] & sel_one_hot_i[73];
  assign data_masked[9463] = data_i[9463] & sel_one_hot_i[73];
  assign data_masked[9462] = data_i[9462] & sel_one_hot_i[73];
  assign data_masked[9461] = data_i[9461] & sel_one_hot_i[73];
  assign data_masked[9460] = data_i[9460] & sel_one_hot_i[73];
  assign data_masked[9459] = data_i[9459] & sel_one_hot_i[73];
  assign data_masked[9458] = data_i[9458] & sel_one_hot_i[73];
  assign data_masked[9457] = data_i[9457] & sel_one_hot_i[73];
  assign data_masked[9456] = data_i[9456] & sel_one_hot_i[73];
  assign data_masked[9455] = data_i[9455] & sel_one_hot_i[73];
  assign data_masked[9454] = data_i[9454] & sel_one_hot_i[73];
  assign data_masked[9453] = data_i[9453] & sel_one_hot_i[73];
  assign data_masked[9452] = data_i[9452] & sel_one_hot_i[73];
  assign data_masked[9451] = data_i[9451] & sel_one_hot_i[73];
  assign data_masked[9450] = data_i[9450] & sel_one_hot_i[73];
  assign data_masked[9449] = data_i[9449] & sel_one_hot_i[73];
  assign data_masked[9448] = data_i[9448] & sel_one_hot_i[73];
  assign data_masked[9447] = data_i[9447] & sel_one_hot_i[73];
  assign data_masked[9446] = data_i[9446] & sel_one_hot_i[73];
  assign data_masked[9445] = data_i[9445] & sel_one_hot_i[73];
  assign data_masked[9444] = data_i[9444] & sel_one_hot_i[73];
  assign data_masked[9443] = data_i[9443] & sel_one_hot_i[73];
  assign data_masked[9442] = data_i[9442] & sel_one_hot_i[73];
  assign data_masked[9441] = data_i[9441] & sel_one_hot_i[73];
  assign data_masked[9440] = data_i[9440] & sel_one_hot_i[73];
  assign data_masked[9439] = data_i[9439] & sel_one_hot_i[73];
  assign data_masked[9438] = data_i[9438] & sel_one_hot_i[73];
  assign data_masked[9437] = data_i[9437] & sel_one_hot_i[73];
  assign data_masked[9436] = data_i[9436] & sel_one_hot_i[73];
  assign data_masked[9435] = data_i[9435] & sel_one_hot_i[73];
  assign data_masked[9434] = data_i[9434] & sel_one_hot_i[73];
  assign data_masked[9433] = data_i[9433] & sel_one_hot_i[73];
  assign data_masked[9432] = data_i[9432] & sel_one_hot_i[73];
  assign data_masked[9431] = data_i[9431] & sel_one_hot_i[73];
  assign data_masked[9430] = data_i[9430] & sel_one_hot_i[73];
  assign data_masked[9429] = data_i[9429] & sel_one_hot_i[73];
  assign data_masked[9428] = data_i[9428] & sel_one_hot_i[73];
  assign data_masked[9427] = data_i[9427] & sel_one_hot_i[73];
  assign data_masked[9426] = data_i[9426] & sel_one_hot_i[73];
  assign data_masked[9425] = data_i[9425] & sel_one_hot_i[73];
  assign data_masked[9424] = data_i[9424] & sel_one_hot_i[73];
  assign data_masked[9423] = data_i[9423] & sel_one_hot_i[73];
  assign data_masked[9422] = data_i[9422] & sel_one_hot_i[73];
  assign data_masked[9421] = data_i[9421] & sel_one_hot_i[73];
  assign data_masked[9420] = data_i[9420] & sel_one_hot_i[73];
  assign data_masked[9419] = data_i[9419] & sel_one_hot_i[73];
  assign data_masked[9418] = data_i[9418] & sel_one_hot_i[73];
  assign data_masked[9417] = data_i[9417] & sel_one_hot_i[73];
  assign data_masked[9416] = data_i[9416] & sel_one_hot_i[73];
  assign data_masked[9415] = data_i[9415] & sel_one_hot_i[73];
  assign data_masked[9414] = data_i[9414] & sel_one_hot_i[73];
  assign data_masked[9413] = data_i[9413] & sel_one_hot_i[73];
  assign data_masked[9412] = data_i[9412] & sel_one_hot_i[73];
  assign data_masked[9411] = data_i[9411] & sel_one_hot_i[73];
  assign data_masked[9410] = data_i[9410] & sel_one_hot_i[73];
  assign data_masked[9409] = data_i[9409] & sel_one_hot_i[73];
  assign data_masked[9408] = data_i[9408] & sel_one_hot_i[73];
  assign data_masked[9407] = data_i[9407] & sel_one_hot_i[73];
  assign data_masked[9406] = data_i[9406] & sel_one_hot_i[73];
  assign data_masked[9405] = data_i[9405] & sel_one_hot_i[73];
  assign data_masked[9404] = data_i[9404] & sel_one_hot_i[73];
  assign data_masked[9403] = data_i[9403] & sel_one_hot_i[73];
  assign data_masked[9402] = data_i[9402] & sel_one_hot_i[73];
  assign data_masked[9401] = data_i[9401] & sel_one_hot_i[73];
  assign data_masked[9400] = data_i[9400] & sel_one_hot_i[73];
  assign data_masked[9399] = data_i[9399] & sel_one_hot_i[73];
  assign data_masked[9398] = data_i[9398] & sel_one_hot_i[73];
  assign data_masked[9397] = data_i[9397] & sel_one_hot_i[73];
  assign data_masked[9396] = data_i[9396] & sel_one_hot_i[73];
  assign data_masked[9395] = data_i[9395] & sel_one_hot_i[73];
  assign data_masked[9394] = data_i[9394] & sel_one_hot_i[73];
  assign data_masked[9393] = data_i[9393] & sel_one_hot_i[73];
  assign data_masked[9392] = data_i[9392] & sel_one_hot_i[73];
  assign data_masked[9391] = data_i[9391] & sel_one_hot_i[73];
  assign data_masked[9390] = data_i[9390] & sel_one_hot_i[73];
  assign data_masked[9389] = data_i[9389] & sel_one_hot_i[73];
  assign data_masked[9388] = data_i[9388] & sel_one_hot_i[73];
  assign data_masked[9387] = data_i[9387] & sel_one_hot_i[73];
  assign data_masked[9386] = data_i[9386] & sel_one_hot_i[73];
  assign data_masked[9385] = data_i[9385] & sel_one_hot_i[73];
  assign data_masked[9384] = data_i[9384] & sel_one_hot_i[73];
  assign data_masked[9383] = data_i[9383] & sel_one_hot_i[73];
  assign data_masked[9382] = data_i[9382] & sel_one_hot_i[73];
  assign data_masked[9381] = data_i[9381] & sel_one_hot_i[73];
  assign data_masked[9380] = data_i[9380] & sel_one_hot_i[73];
  assign data_masked[9379] = data_i[9379] & sel_one_hot_i[73];
  assign data_masked[9378] = data_i[9378] & sel_one_hot_i[73];
  assign data_masked[9377] = data_i[9377] & sel_one_hot_i[73];
  assign data_masked[9376] = data_i[9376] & sel_one_hot_i[73];
  assign data_masked[9375] = data_i[9375] & sel_one_hot_i[73];
  assign data_masked[9374] = data_i[9374] & sel_one_hot_i[73];
  assign data_masked[9373] = data_i[9373] & sel_one_hot_i[73];
  assign data_masked[9372] = data_i[9372] & sel_one_hot_i[73];
  assign data_masked[9371] = data_i[9371] & sel_one_hot_i[73];
  assign data_masked[9370] = data_i[9370] & sel_one_hot_i[73];
  assign data_masked[9369] = data_i[9369] & sel_one_hot_i[73];
  assign data_masked[9368] = data_i[9368] & sel_one_hot_i[73];
  assign data_masked[9367] = data_i[9367] & sel_one_hot_i[73];
  assign data_masked[9366] = data_i[9366] & sel_one_hot_i[73];
  assign data_masked[9365] = data_i[9365] & sel_one_hot_i[73];
  assign data_masked[9364] = data_i[9364] & sel_one_hot_i[73];
  assign data_masked[9363] = data_i[9363] & sel_one_hot_i[73];
  assign data_masked[9362] = data_i[9362] & sel_one_hot_i[73];
  assign data_masked[9361] = data_i[9361] & sel_one_hot_i[73];
  assign data_masked[9360] = data_i[9360] & sel_one_hot_i[73];
  assign data_masked[9359] = data_i[9359] & sel_one_hot_i[73];
  assign data_masked[9358] = data_i[9358] & sel_one_hot_i[73];
  assign data_masked[9357] = data_i[9357] & sel_one_hot_i[73];
  assign data_masked[9356] = data_i[9356] & sel_one_hot_i[73];
  assign data_masked[9355] = data_i[9355] & sel_one_hot_i[73];
  assign data_masked[9354] = data_i[9354] & sel_one_hot_i[73];
  assign data_masked[9353] = data_i[9353] & sel_one_hot_i[73];
  assign data_masked[9352] = data_i[9352] & sel_one_hot_i[73];
  assign data_masked[9351] = data_i[9351] & sel_one_hot_i[73];
  assign data_masked[9350] = data_i[9350] & sel_one_hot_i[73];
  assign data_masked[9349] = data_i[9349] & sel_one_hot_i[73];
  assign data_masked[9348] = data_i[9348] & sel_one_hot_i[73];
  assign data_masked[9347] = data_i[9347] & sel_one_hot_i[73];
  assign data_masked[9346] = data_i[9346] & sel_one_hot_i[73];
  assign data_masked[9345] = data_i[9345] & sel_one_hot_i[73];
  assign data_masked[9344] = data_i[9344] & sel_one_hot_i[73];
  assign data_masked[9599] = data_i[9599] & sel_one_hot_i[74];
  assign data_masked[9598] = data_i[9598] & sel_one_hot_i[74];
  assign data_masked[9597] = data_i[9597] & sel_one_hot_i[74];
  assign data_masked[9596] = data_i[9596] & sel_one_hot_i[74];
  assign data_masked[9595] = data_i[9595] & sel_one_hot_i[74];
  assign data_masked[9594] = data_i[9594] & sel_one_hot_i[74];
  assign data_masked[9593] = data_i[9593] & sel_one_hot_i[74];
  assign data_masked[9592] = data_i[9592] & sel_one_hot_i[74];
  assign data_masked[9591] = data_i[9591] & sel_one_hot_i[74];
  assign data_masked[9590] = data_i[9590] & sel_one_hot_i[74];
  assign data_masked[9589] = data_i[9589] & sel_one_hot_i[74];
  assign data_masked[9588] = data_i[9588] & sel_one_hot_i[74];
  assign data_masked[9587] = data_i[9587] & sel_one_hot_i[74];
  assign data_masked[9586] = data_i[9586] & sel_one_hot_i[74];
  assign data_masked[9585] = data_i[9585] & sel_one_hot_i[74];
  assign data_masked[9584] = data_i[9584] & sel_one_hot_i[74];
  assign data_masked[9583] = data_i[9583] & sel_one_hot_i[74];
  assign data_masked[9582] = data_i[9582] & sel_one_hot_i[74];
  assign data_masked[9581] = data_i[9581] & sel_one_hot_i[74];
  assign data_masked[9580] = data_i[9580] & sel_one_hot_i[74];
  assign data_masked[9579] = data_i[9579] & sel_one_hot_i[74];
  assign data_masked[9578] = data_i[9578] & sel_one_hot_i[74];
  assign data_masked[9577] = data_i[9577] & sel_one_hot_i[74];
  assign data_masked[9576] = data_i[9576] & sel_one_hot_i[74];
  assign data_masked[9575] = data_i[9575] & sel_one_hot_i[74];
  assign data_masked[9574] = data_i[9574] & sel_one_hot_i[74];
  assign data_masked[9573] = data_i[9573] & sel_one_hot_i[74];
  assign data_masked[9572] = data_i[9572] & sel_one_hot_i[74];
  assign data_masked[9571] = data_i[9571] & sel_one_hot_i[74];
  assign data_masked[9570] = data_i[9570] & sel_one_hot_i[74];
  assign data_masked[9569] = data_i[9569] & sel_one_hot_i[74];
  assign data_masked[9568] = data_i[9568] & sel_one_hot_i[74];
  assign data_masked[9567] = data_i[9567] & sel_one_hot_i[74];
  assign data_masked[9566] = data_i[9566] & sel_one_hot_i[74];
  assign data_masked[9565] = data_i[9565] & sel_one_hot_i[74];
  assign data_masked[9564] = data_i[9564] & sel_one_hot_i[74];
  assign data_masked[9563] = data_i[9563] & sel_one_hot_i[74];
  assign data_masked[9562] = data_i[9562] & sel_one_hot_i[74];
  assign data_masked[9561] = data_i[9561] & sel_one_hot_i[74];
  assign data_masked[9560] = data_i[9560] & sel_one_hot_i[74];
  assign data_masked[9559] = data_i[9559] & sel_one_hot_i[74];
  assign data_masked[9558] = data_i[9558] & sel_one_hot_i[74];
  assign data_masked[9557] = data_i[9557] & sel_one_hot_i[74];
  assign data_masked[9556] = data_i[9556] & sel_one_hot_i[74];
  assign data_masked[9555] = data_i[9555] & sel_one_hot_i[74];
  assign data_masked[9554] = data_i[9554] & sel_one_hot_i[74];
  assign data_masked[9553] = data_i[9553] & sel_one_hot_i[74];
  assign data_masked[9552] = data_i[9552] & sel_one_hot_i[74];
  assign data_masked[9551] = data_i[9551] & sel_one_hot_i[74];
  assign data_masked[9550] = data_i[9550] & sel_one_hot_i[74];
  assign data_masked[9549] = data_i[9549] & sel_one_hot_i[74];
  assign data_masked[9548] = data_i[9548] & sel_one_hot_i[74];
  assign data_masked[9547] = data_i[9547] & sel_one_hot_i[74];
  assign data_masked[9546] = data_i[9546] & sel_one_hot_i[74];
  assign data_masked[9545] = data_i[9545] & sel_one_hot_i[74];
  assign data_masked[9544] = data_i[9544] & sel_one_hot_i[74];
  assign data_masked[9543] = data_i[9543] & sel_one_hot_i[74];
  assign data_masked[9542] = data_i[9542] & sel_one_hot_i[74];
  assign data_masked[9541] = data_i[9541] & sel_one_hot_i[74];
  assign data_masked[9540] = data_i[9540] & sel_one_hot_i[74];
  assign data_masked[9539] = data_i[9539] & sel_one_hot_i[74];
  assign data_masked[9538] = data_i[9538] & sel_one_hot_i[74];
  assign data_masked[9537] = data_i[9537] & sel_one_hot_i[74];
  assign data_masked[9536] = data_i[9536] & sel_one_hot_i[74];
  assign data_masked[9535] = data_i[9535] & sel_one_hot_i[74];
  assign data_masked[9534] = data_i[9534] & sel_one_hot_i[74];
  assign data_masked[9533] = data_i[9533] & sel_one_hot_i[74];
  assign data_masked[9532] = data_i[9532] & sel_one_hot_i[74];
  assign data_masked[9531] = data_i[9531] & sel_one_hot_i[74];
  assign data_masked[9530] = data_i[9530] & sel_one_hot_i[74];
  assign data_masked[9529] = data_i[9529] & sel_one_hot_i[74];
  assign data_masked[9528] = data_i[9528] & sel_one_hot_i[74];
  assign data_masked[9527] = data_i[9527] & sel_one_hot_i[74];
  assign data_masked[9526] = data_i[9526] & sel_one_hot_i[74];
  assign data_masked[9525] = data_i[9525] & sel_one_hot_i[74];
  assign data_masked[9524] = data_i[9524] & sel_one_hot_i[74];
  assign data_masked[9523] = data_i[9523] & sel_one_hot_i[74];
  assign data_masked[9522] = data_i[9522] & sel_one_hot_i[74];
  assign data_masked[9521] = data_i[9521] & sel_one_hot_i[74];
  assign data_masked[9520] = data_i[9520] & sel_one_hot_i[74];
  assign data_masked[9519] = data_i[9519] & sel_one_hot_i[74];
  assign data_masked[9518] = data_i[9518] & sel_one_hot_i[74];
  assign data_masked[9517] = data_i[9517] & sel_one_hot_i[74];
  assign data_masked[9516] = data_i[9516] & sel_one_hot_i[74];
  assign data_masked[9515] = data_i[9515] & sel_one_hot_i[74];
  assign data_masked[9514] = data_i[9514] & sel_one_hot_i[74];
  assign data_masked[9513] = data_i[9513] & sel_one_hot_i[74];
  assign data_masked[9512] = data_i[9512] & sel_one_hot_i[74];
  assign data_masked[9511] = data_i[9511] & sel_one_hot_i[74];
  assign data_masked[9510] = data_i[9510] & sel_one_hot_i[74];
  assign data_masked[9509] = data_i[9509] & sel_one_hot_i[74];
  assign data_masked[9508] = data_i[9508] & sel_one_hot_i[74];
  assign data_masked[9507] = data_i[9507] & sel_one_hot_i[74];
  assign data_masked[9506] = data_i[9506] & sel_one_hot_i[74];
  assign data_masked[9505] = data_i[9505] & sel_one_hot_i[74];
  assign data_masked[9504] = data_i[9504] & sel_one_hot_i[74];
  assign data_masked[9503] = data_i[9503] & sel_one_hot_i[74];
  assign data_masked[9502] = data_i[9502] & sel_one_hot_i[74];
  assign data_masked[9501] = data_i[9501] & sel_one_hot_i[74];
  assign data_masked[9500] = data_i[9500] & sel_one_hot_i[74];
  assign data_masked[9499] = data_i[9499] & sel_one_hot_i[74];
  assign data_masked[9498] = data_i[9498] & sel_one_hot_i[74];
  assign data_masked[9497] = data_i[9497] & sel_one_hot_i[74];
  assign data_masked[9496] = data_i[9496] & sel_one_hot_i[74];
  assign data_masked[9495] = data_i[9495] & sel_one_hot_i[74];
  assign data_masked[9494] = data_i[9494] & sel_one_hot_i[74];
  assign data_masked[9493] = data_i[9493] & sel_one_hot_i[74];
  assign data_masked[9492] = data_i[9492] & sel_one_hot_i[74];
  assign data_masked[9491] = data_i[9491] & sel_one_hot_i[74];
  assign data_masked[9490] = data_i[9490] & sel_one_hot_i[74];
  assign data_masked[9489] = data_i[9489] & sel_one_hot_i[74];
  assign data_masked[9488] = data_i[9488] & sel_one_hot_i[74];
  assign data_masked[9487] = data_i[9487] & sel_one_hot_i[74];
  assign data_masked[9486] = data_i[9486] & sel_one_hot_i[74];
  assign data_masked[9485] = data_i[9485] & sel_one_hot_i[74];
  assign data_masked[9484] = data_i[9484] & sel_one_hot_i[74];
  assign data_masked[9483] = data_i[9483] & sel_one_hot_i[74];
  assign data_masked[9482] = data_i[9482] & sel_one_hot_i[74];
  assign data_masked[9481] = data_i[9481] & sel_one_hot_i[74];
  assign data_masked[9480] = data_i[9480] & sel_one_hot_i[74];
  assign data_masked[9479] = data_i[9479] & sel_one_hot_i[74];
  assign data_masked[9478] = data_i[9478] & sel_one_hot_i[74];
  assign data_masked[9477] = data_i[9477] & sel_one_hot_i[74];
  assign data_masked[9476] = data_i[9476] & sel_one_hot_i[74];
  assign data_masked[9475] = data_i[9475] & sel_one_hot_i[74];
  assign data_masked[9474] = data_i[9474] & sel_one_hot_i[74];
  assign data_masked[9473] = data_i[9473] & sel_one_hot_i[74];
  assign data_masked[9472] = data_i[9472] & sel_one_hot_i[74];
  assign data_masked[9727] = data_i[9727] & sel_one_hot_i[75];
  assign data_masked[9726] = data_i[9726] & sel_one_hot_i[75];
  assign data_masked[9725] = data_i[9725] & sel_one_hot_i[75];
  assign data_masked[9724] = data_i[9724] & sel_one_hot_i[75];
  assign data_masked[9723] = data_i[9723] & sel_one_hot_i[75];
  assign data_masked[9722] = data_i[9722] & sel_one_hot_i[75];
  assign data_masked[9721] = data_i[9721] & sel_one_hot_i[75];
  assign data_masked[9720] = data_i[9720] & sel_one_hot_i[75];
  assign data_masked[9719] = data_i[9719] & sel_one_hot_i[75];
  assign data_masked[9718] = data_i[9718] & sel_one_hot_i[75];
  assign data_masked[9717] = data_i[9717] & sel_one_hot_i[75];
  assign data_masked[9716] = data_i[9716] & sel_one_hot_i[75];
  assign data_masked[9715] = data_i[9715] & sel_one_hot_i[75];
  assign data_masked[9714] = data_i[9714] & sel_one_hot_i[75];
  assign data_masked[9713] = data_i[9713] & sel_one_hot_i[75];
  assign data_masked[9712] = data_i[9712] & sel_one_hot_i[75];
  assign data_masked[9711] = data_i[9711] & sel_one_hot_i[75];
  assign data_masked[9710] = data_i[9710] & sel_one_hot_i[75];
  assign data_masked[9709] = data_i[9709] & sel_one_hot_i[75];
  assign data_masked[9708] = data_i[9708] & sel_one_hot_i[75];
  assign data_masked[9707] = data_i[9707] & sel_one_hot_i[75];
  assign data_masked[9706] = data_i[9706] & sel_one_hot_i[75];
  assign data_masked[9705] = data_i[9705] & sel_one_hot_i[75];
  assign data_masked[9704] = data_i[9704] & sel_one_hot_i[75];
  assign data_masked[9703] = data_i[9703] & sel_one_hot_i[75];
  assign data_masked[9702] = data_i[9702] & sel_one_hot_i[75];
  assign data_masked[9701] = data_i[9701] & sel_one_hot_i[75];
  assign data_masked[9700] = data_i[9700] & sel_one_hot_i[75];
  assign data_masked[9699] = data_i[9699] & sel_one_hot_i[75];
  assign data_masked[9698] = data_i[9698] & sel_one_hot_i[75];
  assign data_masked[9697] = data_i[9697] & sel_one_hot_i[75];
  assign data_masked[9696] = data_i[9696] & sel_one_hot_i[75];
  assign data_masked[9695] = data_i[9695] & sel_one_hot_i[75];
  assign data_masked[9694] = data_i[9694] & sel_one_hot_i[75];
  assign data_masked[9693] = data_i[9693] & sel_one_hot_i[75];
  assign data_masked[9692] = data_i[9692] & sel_one_hot_i[75];
  assign data_masked[9691] = data_i[9691] & sel_one_hot_i[75];
  assign data_masked[9690] = data_i[9690] & sel_one_hot_i[75];
  assign data_masked[9689] = data_i[9689] & sel_one_hot_i[75];
  assign data_masked[9688] = data_i[9688] & sel_one_hot_i[75];
  assign data_masked[9687] = data_i[9687] & sel_one_hot_i[75];
  assign data_masked[9686] = data_i[9686] & sel_one_hot_i[75];
  assign data_masked[9685] = data_i[9685] & sel_one_hot_i[75];
  assign data_masked[9684] = data_i[9684] & sel_one_hot_i[75];
  assign data_masked[9683] = data_i[9683] & sel_one_hot_i[75];
  assign data_masked[9682] = data_i[9682] & sel_one_hot_i[75];
  assign data_masked[9681] = data_i[9681] & sel_one_hot_i[75];
  assign data_masked[9680] = data_i[9680] & sel_one_hot_i[75];
  assign data_masked[9679] = data_i[9679] & sel_one_hot_i[75];
  assign data_masked[9678] = data_i[9678] & sel_one_hot_i[75];
  assign data_masked[9677] = data_i[9677] & sel_one_hot_i[75];
  assign data_masked[9676] = data_i[9676] & sel_one_hot_i[75];
  assign data_masked[9675] = data_i[9675] & sel_one_hot_i[75];
  assign data_masked[9674] = data_i[9674] & sel_one_hot_i[75];
  assign data_masked[9673] = data_i[9673] & sel_one_hot_i[75];
  assign data_masked[9672] = data_i[9672] & sel_one_hot_i[75];
  assign data_masked[9671] = data_i[9671] & sel_one_hot_i[75];
  assign data_masked[9670] = data_i[9670] & sel_one_hot_i[75];
  assign data_masked[9669] = data_i[9669] & sel_one_hot_i[75];
  assign data_masked[9668] = data_i[9668] & sel_one_hot_i[75];
  assign data_masked[9667] = data_i[9667] & sel_one_hot_i[75];
  assign data_masked[9666] = data_i[9666] & sel_one_hot_i[75];
  assign data_masked[9665] = data_i[9665] & sel_one_hot_i[75];
  assign data_masked[9664] = data_i[9664] & sel_one_hot_i[75];
  assign data_masked[9663] = data_i[9663] & sel_one_hot_i[75];
  assign data_masked[9662] = data_i[9662] & sel_one_hot_i[75];
  assign data_masked[9661] = data_i[9661] & sel_one_hot_i[75];
  assign data_masked[9660] = data_i[9660] & sel_one_hot_i[75];
  assign data_masked[9659] = data_i[9659] & sel_one_hot_i[75];
  assign data_masked[9658] = data_i[9658] & sel_one_hot_i[75];
  assign data_masked[9657] = data_i[9657] & sel_one_hot_i[75];
  assign data_masked[9656] = data_i[9656] & sel_one_hot_i[75];
  assign data_masked[9655] = data_i[9655] & sel_one_hot_i[75];
  assign data_masked[9654] = data_i[9654] & sel_one_hot_i[75];
  assign data_masked[9653] = data_i[9653] & sel_one_hot_i[75];
  assign data_masked[9652] = data_i[9652] & sel_one_hot_i[75];
  assign data_masked[9651] = data_i[9651] & sel_one_hot_i[75];
  assign data_masked[9650] = data_i[9650] & sel_one_hot_i[75];
  assign data_masked[9649] = data_i[9649] & sel_one_hot_i[75];
  assign data_masked[9648] = data_i[9648] & sel_one_hot_i[75];
  assign data_masked[9647] = data_i[9647] & sel_one_hot_i[75];
  assign data_masked[9646] = data_i[9646] & sel_one_hot_i[75];
  assign data_masked[9645] = data_i[9645] & sel_one_hot_i[75];
  assign data_masked[9644] = data_i[9644] & sel_one_hot_i[75];
  assign data_masked[9643] = data_i[9643] & sel_one_hot_i[75];
  assign data_masked[9642] = data_i[9642] & sel_one_hot_i[75];
  assign data_masked[9641] = data_i[9641] & sel_one_hot_i[75];
  assign data_masked[9640] = data_i[9640] & sel_one_hot_i[75];
  assign data_masked[9639] = data_i[9639] & sel_one_hot_i[75];
  assign data_masked[9638] = data_i[9638] & sel_one_hot_i[75];
  assign data_masked[9637] = data_i[9637] & sel_one_hot_i[75];
  assign data_masked[9636] = data_i[9636] & sel_one_hot_i[75];
  assign data_masked[9635] = data_i[9635] & sel_one_hot_i[75];
  assign data_masked[9634] = data_i[9634] & sel_one_hot_i[75];
  assign data_masked[9633] = data_i[9633] & sel_one_hot_i[75];
  assign data_masked[9632] = data_i[9632] & sel_one_hot_i[75];
  assign data_masked[9631] = data_i[9631] & sel_one_hot_i[75];
  assign data_masked[9630] = data_i[9630] & sel_one_hot_i[75];
  assign data_masked[9629] = data_i[9629] & sel_one_hot_i[75];
  assign data_masked[9628] = data_i[9628] & sel_one_hot_i[75];
  assign data_masked[9627] = data_i[9627] & sel_one_hot_i[75];
  assign data_masked[9626] = data_i[9626] & sel_one_hot_i[75];
  assign data_masked[9625] = data_i[9625] & sel_one_hot_i[75];
  assign data_masked[9624] = data_i[9624] & sel_one_hot_i[75];
  assign data_masked[9623] = data_i[9623] & sel_one_hot_i[75];
  assign data_masked[9622] = data_i[9622] & sel_one_hot_i[75];
  assign data_masked[9621] = data_i[9621] & sel_one_hot_i[75];
  assign data_masked[9620] = data_i[9620] & sel_one_hot_i[75];
  assign data_masked[9619] = data_i[9619] & sel_one_hot_i[75];
  assign data_masked[9618] = data_i[9618] & sel_one_hot_i[75];
  assign data_masked[9617] = data_i[9617] & sel_one_hot_i[75];
  assign data_masked[9616] = data_i[9616] & sel_one_hot_i[75];
  assign data_masked[9615] = data_i[9615] & sel_one_hot_i[75];
  assign data_masked[9614] = data_i[9614] & sel_one_hot_i[75];
  assign data_masked[9613] = data_i[9613] & sel_one_hot_i[75];
  assign data_masked[9612] = data_i[9612] & sel_one_hot_i[75];
  assign data_masked[9611] = data_i[9611] & sel_one_hot_i[75];
  assign data_masked[9610] = data_i[9610] & sel_one_hot_i[75];
  assign data_masked[9609] = data_i[9609] & sel_one_hot_i[75];
  assign data_masked[9608] = data_i[9608] & sel_one_hot_i[75];
  assign data_masked[9607] = data_i[9607] & sel_one_hot_i[75];
  assign data_masked[9606] = data_i[9606] & sel_one_hot_i[75];
  assign data_masked[9605] = data_i[9605] & sel_one_hot_i[75];
  assign data_masked[9604] = data_i[9604] & sel_one_hot_i[75];
  assign data_masked[9603] = data_i[9603] & sel_one_hot_i[75];
  assign data_masked[9602] = data_i[9602] & sel_one_hot_i[75];
  assign data_masked[9601] = data_i[9601] & sel_one_hot_i[75];
  assign data_masked[9600] = data_i[9600] & sel_one_hot_i[75];
  assign data_masked[9855] = data_i[9855] & sel_one_hot_i[76];
  assign data_masked[9854] = data_i[9854] & sel_one_hot_i[76];
  assign data_masked[9853] = data_i[9853] & sel_one_hot_i[76];
  assign data_masked[9852] = data_i[9852] & sel_one_hot_i[76];
  assign data_masked[9851] = data_i[9851] & sel_one_hot_i[76];
  assign data_masked[9850] = data_i[9850] & sel_one_hot_i[76];
  assign data_masked[9849] = data_i[9849] & sel_one_hot_i[76];
  assign data_masked[9848] = data_i[9848] & sel_one_hot_i[76];
  assign data_masked[9847] = data_i[9847] & sel_one_hot_i[76];
  assign data_masked[9846] = data_i[9846] & sel_one_hot_i[76];
  assign data_masked[9845] = data_i[9845] & sel_one_hot_i[76];
  assign data_masked[9844] = data_i[9844] & sel_one_hot_i[76];
  assign data_masked[9843] = data_i[9843] & sel_one_hot_i[76];
  assign data_masked[9842] = data_i[9842] & sel_one_hot_i[76];
  assign data_masked[9841] = data_i[9841] & sel_one_hot_i[76];
  assign data_masked[9840] = data_i[9840] & sel_one_hot_i[76];
  assign data_masked[9839] = data_i[9839] & sel_one_hot_i[76];
  assign data_masked[9838] = data_i[9838] & sel_one_hot_i[76];
  assign data_masked[9837] = data_i[9837] & sel_one_hot_i[76];
  assign data_masked[9836] = data_i[9836] & sel_one_hot_i[76];
  assign data_masked[9835] = data_i[9835] & sel_one_hot_i[76];
  assign data_masked[9834] = data_i[9834] & sel_one_hot_i[76];
  assign data_masked[9833] = data_i[9833] & sel_one_hot_i[76];
  assign data_masked[9832] = data_i[9832] & sel_one_hot_i[76];
  assign data_masked[9831] = data_i[9831] & sel_one_hot_i[76];
  assign data_masked[9830] = data_i[9830] & sel_one_hot_i[76];
  assign data_masked[9829] = data_i[9829] & sel_one_hot_i[76];
  assign data_masked[9828] = data_i[9828] & sel_one_hot_i[76];
  assign data_masked[9827] = data_i[9827] & sel_one_hot_i[76];
  assign data_masked[9826] = data_i[9826] & sel_one_hot_i[76];
  assign data_masked[9825] = data_i[9825] & sel_one_hot_i[76];
  assign data_masked[9824] = data_i[9824] & sel_one_hot_i[76];
  assign data_masked[9823] = data_i[9823] & sel_one_hot_i[76];
  assign data_masked[9822] = data_i[9822] & sel_one_hot_i[76];
  assign data_masked[9821] = data_i[9821] & sel_one_hot_i[76];
  assign data_masked[9820] = data_i[9820] & sel_one_hot_i[76];
  assign data_masked[9819] = data_i[9819] & sel_one_hot_i[76];
  assign data_masked[9818] = data_i[9818] & sel_one_hot_i[76];
  assign data_masked[9817] = data_i[9817] & sel_one_hot_i[76];
  assign data_masked[9816] = data_i[9816] & sel_one_hot_i[76];
  assign data_masked[9815] = data_i[9815] & sel_one_hot_i[76];
  assign data_masked[9814] = data_i[9814] & sel_one_hot_i[76];
  assign data_masked[9813] = data_i[9813] & sel_one_hot_i[76];
  assign data_masked[9812] = data_i[9812] & sel_one_hot_i[76];
  assign data_masked[9811] = data_i[9811] & sel_one_hot_i[76];
  assign data_masked[9810] = data_i[9810] & sel_one_hot_i[76];
  assign data_masked[9809] = data_i[9809] & sel_one_hot_i[76];
  assign data_masked[9808] = data_i[9808] & sel_one_hot_i[76];
  assign data_masked[9807] = data_i[9807] & sel_one_hot_i[76];
  assign data_masked[9806] = data_i[9806] & sel_one_hot_i[76];
  assign data_masked[9805] = data_i[9805] & sel_one_hot_i[76];
  assign data_masked[9804] = data_i[9804] & sel_one_hot_i[76];
  assign data_masked[9803] = data_i[9803] & sel_one_hot_i[76];
  assign data_masked[9802] = data_i[9802] & sel_one_hot_i[76];
  assign data_masked[9801] = data_i[9801] & sel_one_hot_i[76];
  assign data_masked[9800] = data_i[9800] & sel_one_hot_i[76];
  assign data_masked[9799] = data_i[9799] & sel_one_hot_i[76];
  assign data_masked[9798] = data_i[9798] & sel_one_hot_i[76];
  assign data_masked[9797] = data_i[9797] & sel_one_hot_i[76];
  assign data_masked[9796] = data_i[9796] & sel_one_hot_i[76];
  assign data_masked[9795] = data_i[9795] & sel_one_hot_i[76];
  assign data_masked[9794] = data_i[9794] & sel_one_hot_i[76];
  assign data_masked[9793] = data_i[9793] & sel_one_hot_i[76];
  assign data_masked[9792] = data_i[9792] & sel_one_hot_i[76];
  assign data_masked[9791] = data_i[9791] & sel_one_hot_i[76];
  assign data_masked[9790] = data_i[9790] & sel_one_hot_i[76];
  assign data_masked[9789] = data_i[9789] & sel_one_hot_i[76];
  assign data_masked[9788] = data_i[9788] & sel_one_hot_i[76];
  assign data_masked[9787] = data_i[9787] & sel_one_hot_i[76];
  assign data_masked[9786] = data_i[9786] & sel_one_hot_i[76];
  assign data_masked[9785] = data_i[9785] & sel_one_hot_i[76];
  assign data_masked[9784] = data_i[9784] & sel_one_hot_i[76];
  assign data_masked[9783] = data_i[9783] & sel_one_hot_i[76];
  assign data_masked[9782] = data_i[9782] & sel_one_hot_i[76];
  assign data_masked[9781] = data_i[9781] & sel_one_hot_i[76];
  assign data_masked[9780] = data_i[9780] & sel_one_hot_i[76];
  assign data_masked[9779] = data_i[9779] & sel_one_hot_i[76];
  assign data_masked[9778] = data_i[9778] & sel_one_hot_i[76];
  assign data_masked[9777] = data_i[9777] & sel_one_hot_i[76];
  assign data_masked[9776] = data_i[9776] & sel_one_hot_i[76];
  assign data_masked[9775] = data_i[9775] & sel_one_hot_i[76];
  assign data_masked[9774] = data_i[9774] & sel_one_hot_i[76];
  assign data_masked[9773] = data_i[9773] & sel_one_hot_i[76];
  assign data_masked[9772] = data_i[9772] & sel_one_hot_i[76];
  assign data_masked[9771] = data_i[9771] & sel_one_hot_i[76];
  assign data_masked[9770] = data_i[9770] & sel_one_hot_i[76];
  assign data_masked[9769] = data_i[9769] & sel_one_hot_i[76];
  assign data_masked[9768] = data_i[9768] & sel_one_hot_i[76];
  assign data_masked[9767] = data_i[9767] & sel_one_hot_i[76];
  assign data_masked[9766] = data_i[9766] & sel_one_hot_i[76];
  assign data_masked[9765] = data_i[9765] & sel_one_hot_i[76];
  assign data_masked[9764] = data_i[9764] & sel_one_hot_i[76];
  assign data_masked[9763] = data_i[9763] & sel_one_hot_i[76];
  assign data_masked[9762] = data_i[9762] & sel_one_hot_i[76];
  assign data_masked[9761] = data_i[9761] & sel_one_hot_i[76];
  assign data_masked[9760] = data_i[9760] & sel_one_hot_i[76];
  assign data_masked[9759] = data_i[9759] & sel_one_hot_i[76];
  assign data_masked[9758] = data_i[9758] & sel_one_hot_i[76];
  assign data_masked[9757] = data_i[9757] & sel_one_hot_i[76];
  assign data_masked[9756] = data_i[9756] & sel_one_hot_i[76];
  assign data_masked[9755] = data_i[9755] & sel_one_hot_i[76];
  assign data_masked[9754] = data_i[9754] & sel_one_hot_i[76];
  assign data_masked[9753] = data_i[9753] & sel_one_hot_i[76];
  assign data_masked[9752] = data_i[9752] & sel_one_hot_i[76];
  assign data_masked[9751] = data_i[9751] & sel_one_hot_i[76];
  assign data_masked[9750] = data_i[9750] & sel_one_hot_i[76];
  assign data_masked[9749] = data_i[9749] & sel_one_hot_i[76];
  assign data_masked[9748] = data_i[9748] & sel_one_hot_i[76];
  assign data_masked[9747] = data_i[9747] & sel_one_hot_i[76];
  assign data_masked[9746] = data_i[9746] & sel_one_hot_i[76];
  assign data_masked[9745] = data_i[9745] & sel_one_hot_i[76];
  assign data_masked[9744] = data_i[9744] & sel_one_hot_i[76];
  assign data_masked[9743] = data_i[9743] & sel_one_hot_i[76];
  assign data_masked[9742] = data_i[9742] & sel_one_hot_i[76];
  assign data_masked[9741] = data_i[9741] & sel_one_hot_i[76];
  assign data_masked[9740] = data_i[9740] & sel_one_hot_i[76];
  assign data_masked[9739] = data_i[9739] & sel_one_hot_i[76];
  assign data_masked[9738] = data_i[9738] & sel_one_hot_i[76];
  assign data_masked[9737] = data_i[9737] & sel_one_hot_i[76];
  assign data_masked[9736] = data_i[9736] & sel_one_hot_i[76];
  assign data_masked[9735] = data_i[9735] & sel_one_hot_i[76];
  assign data_masked[9734] = data_i[9734] & sel_one_hot_i[76];
  assign data_masked[9733] = data_i[9733] & sel_one_hot_i[76];
  assign data_masked[9732] = data_i[9732] & sel_one_hot_i[76];
  assign data_masked[9731] = data_i[9731] & sel_one_hot_i[76];
  assign data_masked[9730] = data_i[9730] & sel_one_hot_i[76];
  assign data_masked[9729] = data_i[9729] & sel_one_hot_i[76];
  assign data_masked[9728] = data_i[9728] & sel_one_hot_i[76];
  assign data_masked[9983] = data_i[9983] & sel_one_hot_i[77];
  assign data_masked[9982] = data_i[9982] & sel_one_hot_i[77];
  assign data_masked[9981] = data_i[9981] & sel_one_hot_i[77];
  assign data_masked[9980] = data_i[9980] & sel_one_hot_i[77];
  assign data_masked[9979] = data_i[9979] & sel_one_hot_i[77];
  assign data_masked[9978] = data_i[9978] & sel_one_hot_i[77];
  assign data_masked[9977] = data_i[9977] & sel_one_hot_i[77];
  assign data_masked[9976] = data_i[9976] & sel_one_hot_i[77];
  assign data_masked[9975] = data_i[9975] & sel_one_hot_i[77];
  assign data_masked[9974] = data_i[9974] & sel_one_hot_i[77];
  assign data_masked[9973] = data_i[9973] & sel_one_hot_i[77];
  assign data_masked[9972] = data_i[9972] & sel_one_hot_i[77];
  assign data_masked[9971] = data_i[9971] & sel_one_hot_i[77];
  assign data_masked[9970] = data_i[9970] & sel_one_hot_i[77];
  assign data_masked[9969] = data_i[9969] & sel_one_hot_i[77];
  assign data_masked[9968] = data_i[9968] & sel_one_hot_i[77];
  assign data_masked[9967] = data_i[9967] & sel_one_hot_i[77];
  assign data_masked[9966] = data_i[9966] & sel_one_hot_i[77];
  assign data_masked[9965] = data_i[9965] & sel_one_hot_i[77];
  assign data_masked[9964] = data_i[9964] & sel_one_hot_i[77];
  assign data_masked[9963] = data_i[9963] & sel_one_hot_i[77];
  assign data_masked[9962] = data_i[9962] & sel_one_hot_i[77];
  assign data_masked[9961] = data_i[9961] & sel_one_hot_i[77];
  assign data_masked[9960] = data_i[9960] & sel_one_hot_i[77];
  assign data_masked[9959] = data_i[9959] & sel_one_hot_i[77];
  assign data_masked[9958] = data_i[9958] & sel_one_hot_i[77];
  assign data_masked[9957] = data_i[9957] & sel_one_hot_i[77];
  assign data_masked[9956] = data_i[9956] & sel_one_hot_i[77];
  assign data_masked[9955] = data_i[9955] & sel_one_hot_i[77];
  assign data_masked[9954] = data_i[9954] & sel_one_hot_i[77];
  assign data_masked[9953] = data_i[9953] & sel_one_hot_i[77];
  assign data_masked[9952] = data_i[9952] & sel_one_hot_i[77];
  assign data_masked[9951] = data_i[9951] & sel_one_hot_i[77];
  assign data_masked[9950] = data_i[9950] & sel_one_hot_i[77];
  assign data_masked[9949] = data_i[9949] & sel_one_hot_i[77];
  assign data_masked[9948] = data_i[9948] & sel_one_hot_i[77];
  assign data_masked[9947] = data_i[9947] & sel_one_hot_i[77];
  assign data_masked[9946] = data_i[9946] & sel_one_hot_i[77];
  assign data_masked[9945] = data_i[9945] & sel_one_hot_i[77];
  assign data_masked[9944] = data_i[9944] & sel_one_hot_i[77];
  assign data_masked[9943] = data_i[9943] & sel_one_hot_i[77];
  assign data_masked[9942] = data_i[9942] & sel_one_hot_i[77];
  assign data_masked[9941] = data_i[9941] & sel_one_hot_i[77];
  assign data_masked[9940] = data_i[9940] & sel_one_hot_i[77];
  assign data_masked[9939] = data_i[9939] & sel_one_hot_i[77];
  assign data_masked[9938] = data_i[9938] & sel_one_hot_i[77];
  assign data_masked[9937] = data_i[9937] & sel_one_hot_i[77];
  assign data_masked[9936] = data_i[9936] & sel_one_hot_i[77];
  assign data_masked[9935] = data_i[9935] & sel_one_hot_i[77];
  assign data_masked[9934] = data_i[9934] & sel_one_hot_i[77];
  assign data_masked[9933] = data_i[9933] & sel_one_hot_i[77];
  assign data_masked[9932] = data_i[9932] & sel_one_hot_i[77];
  assign data_masked[9931] = data_i[9931] & sel_one_hot_i[77];
  assign data_masked[9930] = data_i[9930] & sel_one_hot_i[77];
  assign data_masked[9929] = data_i[9929] & sel_one_hot_i[77];
  assign data_masked[9928] = data_i[9928] & sel_one_hot_i[77];
  assign data_masked[9927] = data_i[9927] & sel_one_hot_i[77];
  assign data_masked[9926] = data_i[9926] & sel_one_hot_i[77];
  assign data_masked[9925] = data_i[9925] & sel_one_hot_i[77];
  assign data_masked[9924] = data_i[9924] & sel_one_hot_i[77];
  assign data_masked[9923] = data_i[9923] & sel_one_hot_i[77];
  assign data_masked[9922] = data_i[9922] & sel_one_hot_i[77];
  assign data_masked[9921] = data_i[9921] & sel_one_hot_i[77];
  assign data_masked[9920] = data_i[9920] & sel_one_hot_i[77];
  assign data_masked[9919] = data_i[9919] & sel_one_hot_i[77];
  assign data_masked[9918] = data_i[9918] & sel_one_hot_i[77];
  assign data_masked[9917] = data_i[9917] & sel_one_hot_i[77];
  assign data_masked[9916] = data_i[9916] & sel_one_hot_i[77];
  assign data_masked[9915] = data_i[9915] & sel_one_hot_i[77];
  assign data_masked[9914] = data_i[9914] & sel_one_hot_i[77];
  assign data_masked[9913] = data_i[9913] & sel_one_hot_i[77];
  assign data_masked[9912] = data_i[9912] & sel_one_hot_i[77];
  assign data_masked[9911] = data_i[9911] & sel_one_hot_i[77];
  assign data_masked[9910] = data_i[9910] & sel_one_hot_i[77];
  assign data_masked[9909] = data_i[9909] & sel_one_hot_i[77];
  assign data_masked[9908] = data_i[9908] & sel_one_hot_i[77];
  assign data_masked[9907] = data_i[9907] & sel_one_hot_i[77];
  assign data_masked[9906] = data_i[9906] & sel_one_hot_i[77];
  assign data_masked[9905] = data_i[9905] & sel_one_hot_i[77];
  assign data_masked[9904] = data_i[9904] & sel_one_hot_i[77];
  assign data_masked[9903] = data_i[9903] & sel_one_hot_i[77];
  assign data_masked[9902] = data_i[9902] & sel_one_hot_i[77];
  assign data_masked[9901] = data_i[9901] & sel_one_hot_i[77];
  assign data_masked[9900] = data_i[9900] & sel_one_hot_i[77];
  assign data_masked[9899] = data_i[9899] & sel_one_hot_i[77];
  assign data_masked[9898] = data_i[9898] & sel_one_hot_i[77];
  assign data_masked[9897] = data_i[9897] & sel_one_hot_i[77];
  assign data_masked[9896] = data_i[9896] & sel_one_hot_i[77];
  assign data_masked[9895] = data_i[9895] & sel_one_hot_i[77];
  assign data_masked[9894] = data_i[9894] & sel_one_hot_i[77];
  assign data_masked[9893] = data_i[9893] & sel_one_hot_i[77];
  assign data_masked[9892] = data_i[9892] & sel_one_hot_i[77];
  assign data_masked[9891] = data_i[9891] & sel_one_hot_i[77];
  assign data_masked[9890] = data_i[9890] & sel_one_hot_i[77];
  assign data_masked[9889] = data_i[9889] & sel_one_hot_i[77];
  assign data_masked[9888] = data_i[9888] & sel_one_hot_i[77];
  assign data_masked[9887] = data_i[9887] & sel_one_hot_i[77];
  assign data_masked[9886] = data_i[9886] & sel_one_hot_i[77];
  assign data_masked[9885] = data_i[9885] & sel_one_hot_i[77];
  assign data_masked[9884] = data_i[9884] & sel_one_hot_i[77];
  assign data_masked[9883] = data_i[9883] & sel_one_hot_i[77];
  assign data_masked[9882] = data_i[9882] & sel_one_hot_i[77];
  assign data_masked[9881] = data_i[9881] & sel_one_hot_i[77];
  assign data_masked[9880] = data_i[9880] & sel_one_hot_i[77];
  assign data_masked[9879] = data_i[9879] & sel_one_hot_i[77];
  assign data_masked[9878] = data_i[9878] & sel_one_hot_i[77];
  assign data_masked[9877] = data_i[9877] & sel_one_hot_i[77];
  assign data_masked[9876] = data_i[9876] & sel_one_hot_i[77];
  assign data_masked[9875] = data_i[9875] & sel_one_hot_i[77];
  assign data_masked[9874] = data_i[9874] & sel_one_hot_i[77];
  assign data_masked[9873] = data_i[9873] & sel_one_hot_i[77];
  assign data_masked[9872] = data_i[9872] & sel_one_hot_i[77];
  assign data_masked[9871] = data_i[9871] & sel_one_hot_i[77];
  assign data_masked[9870] = data_i[9870] & sel_one_hot_i[77];
  assign data_masked[9869] = data_i[9869] & sel_one_hot_i[77];
  assign data_masked[9868] = data_i[9868] & sel_one_hot_i[77];
  assign data_masked[9867] = data_i[9867] & sel_one_hot_i[77];
  assign data_masked[9866] = data_i[9866] & sel_one_hot_i[77];
  assign data_masked[9865] = data_i[9865] & sel_one_hot_i[77];
  assign data_masked[9864] = data_i[9864] & sel_one_hot_i[77];
  assign data_masked[9863] = data_i[9863] & sel_one_hot_i[77];
  assign data_masked[9862] = data_i[9862] & sel_one_hot_i[77];
  assign data_masked[9861] = data_i[9861] & sel_one_hot_i[77];
  assign data_masked[9860] = data_i[9860] & sel_one_hot_i[77];
  assign data_masked[9859] = data_i[9859] & sel_one_hot_i[77];
  assign data_masked[9858] = data_i[9858] & sel_one_hot_i[77];
  assign data_masked[9857] = data_i[9857] & sel_one_hot_i[77];
  assign data_masked[9856] = data_i[9856] & sel_one_hot_i[77];
  assign data_masked[10111] = data_i[10111] & sel_one_hot_i[78];
  assign data_masked[10110] = data_i[10110] & sel_one_hot_i[78];
  assign data_masked[10109] = data_i[10109] & sel_one_hot_i[78];
  assign data_masked[10108] = data_i[10108] & sel_one_hot_i[78];
  assign data_masked[10107] = data_i[10107] & sel_one_hot_i[78];
  assign data_masked[10106] = data_i[10106] & sel_one_hot_i[78];
  assign data_masked[10105] = data_i[10105] & sel_one_hot_i[78];
  assign data_masked[10104] = data_i[10104] & sel_one_hot_i[78];
  assign data_masked[10103] = data_i[10103] & sel_one_hot_i[78];
  assign data_masked[10102] = data_i[10102] & sel_one_hot_i[78];
  assign data_masked[10101] = data_i[10101] & sel_one_hot_i[78];
  assign data_masked[10100] = data_i[10100] & sel_one_hot_i[78];
  assign data_masked[10099] = data_i[10099] & sel_one_hot_i[78];
  assign data_masked[10098] = data_i[10098] & sel_one_hot_i[78];
  assign data_masked[10097] = data_i[10097] & sel_one_hot_i[78];
  assign data_masked[10096] = data_i[10096] & sel_one_hot_i[78];
  assign data_masked[10095] = data_i[10095] & sel_one_hot_i[78];
  assign data_masked[10094] = data_i[10094] & sel_one_hot_i[78];
  assign data_masked[10093] = data_i[10093] & sel_one_hot_i[78];
  assign data_masked[10092] = data_i[10092] & sel_one_hot_i[78];
  assign data_masked[10091] = data_i[10091] & sel_one_hot_i[78];
  assign data_masked[10090] = data_i[10090] & sel_one_hot_i[78];
  assign data_masked[10089] = data_i[10089] & sel_one_hot_i[78];
  assign data_masked[10088] = data_i[10088] & sel_one_hot_i[78];
  assign data_masked[10087] = data_i[10087] & sel_one_hot_i[78];
  assign data_masked[10086] = data_i[10086] & sel_one_hot_i[78];
  assign data_masked[10085] = data_i[10085] & sel_one_hot_i[78];
  assign data_masked[10084] = data_i[10084] & sel_one_hot_i[78];
  assign data_masked[10083] = data_i[10083] & sel_one_hot_i[78];
  assign data_masked[10082] = data_i[10082] & sel_one_hot_i[78];
  assign data_masked[10081] = data_i[10081] & sel_one_hot_i[78];
  assign data_masked[10080] = data_i[10080] & sel_one_hot_i[78];
  assign data_masked[10079] = data_i[10079] & sel_one_hot_i[78];
  assign data_masked[10078] = data_i[10078] & sel_one_hot_i[78];
  assign data_masked[10077] = data_i[10077] & sel_one_hot_i[78];
  assign data_masked[10076] = data_i[10076] & sel_one_hot_i[78];
  assign data_masked[10075] = data_i[10075] & sel_one_hot_i[78];
  assign data_masked[10074] = data_i[10074] & sel_one_hot_i[78];
  assign data_masked[10073] = data_i[10073] & sel_one_hot_i[78];
  assign data_masked[10072] = data_i[10072] & sel_one_hot_i[78];
  assign data_masked[10071] = data_i[10071] & sel_one_hot_i[78];
  assign data_masked[10070] = data_i[10070] & sel_one_hot_i[78];
  assign data_masked[10069] = data_i[10069] & sel_one_hot_i[78];
  assign data_masked[10068] = data_i[10068] & sel_one_hot_i[78];
  assign data_masked[10067] = data_i[10067] & sel_one_hot_i[78];
  assign data_masked[10066] = data_i[10066] & sel_one_hot_i[78];
  assign data_masked[10065] = data_i[10065] & sel_one_hot_i[78];
  assign data_masked[10064] = data_i[10064] & sel_one_hot_i[78];
  assign data_masked[10063] = data_i[10063] & sel_one_hot_i[78];
  assign data_masked[10062] = data_i[10062] & sel_one_hot_i[78];
  assign data_masked[10061] = data_i[10061] & sel_one_hot_i[78];
  assign data_masked[10060] = data_i[10060] & sel_one_hot_i[78];
  assign data_masked[10059] = data_i[10059] & sel_one_hot_i[78];
  assign data_masked[10058] = data_i[10058] & sel_one_hot_i[78];
  assign data_masked[10057] = data_i[10057] & sel_one_hot_i[78];
  assign data_masked[10056] = data_i[10056] & sel_one_hot_i[78];
  assign data_masked[10055] = data_i[10055] & sel_one_hot_i[78];
  assign data_masked[10054] = data_i[10054] & sel_one_hot_i[78];
  assign data_masked[10053] = data_i[10053] & sel_one_hot_i[78];
  assign data_masked[10052] = data_i[10052] & sel_one_hot_i[78];
  assign data_masked[10051] = data_i[10051] & sel_one_hot_i[78];
  assign data_masked[10050] = data_i[10050] & sel_one_hot_i[78];
  assign data_masked[10049] = data_i[10049] & sel_one_hot_i[78];
  assign data_masked[10048] = data_i[10048] & sel_one_hot_i[78];
  assign data_masked[10047] = data_i[10047] & sel_one_hot_i[78];
  assign data_masked[10046] = data_i[10046] & sel_one_hot_i[78];
  assign data_masked[10045] = data_i[10045] & sel_one_hot_i[78];
  assign data_masked[10044] = data_i[10044] & sel_one_hot_i[78];
  assign data_masked[10043] = data_i[10043] & sel_one_hot_i[78];
  assign data_masked[10042] = data_i[10042] & sel_one_hot_i[78];
  assign data_masked[10041] = data_i[10041] & sel_one_hot_i[78];
  assign data_masked[10040] = data_i[10040] & sel_one_hot_i[78];
  assign data_masked[10039] = data_i[10039] & sel_one_hot_i[78];
  assign data_masked[10038] = data_i[10038] & sel_one_hot_i[78];
  assign data_masked[10037] = data_i[10037] & sel_one_hot_i[78];
  assign data_masked[10036] = data_i[10036] & sel_one_hot_i[78];
  assign data_masked[10035] = data_i[10035] & sel_one_hot_i[78];
  assign data_masked[10034] = data_i[10034] & sel_one_hot_i[78];
  assign data_masked[10033] = data_i[10033] & sel_one_hot_i[78];
  assign data_masked[10032] = data_i[10032] & sel_one_hot_i[78];
  assign data_masked[10031] = data_i[10031] & sel_one_hot_i[78];
  assign data_masked[10030] = data_i[10030] & sel_one_hot_i[78];
  assign data_masked[10029] = data_i[10029] & sel_one_hot_i[78];
  assign data_masked[10028] = data_i[10028] & sel_one_hot_i[78];
  assign data_masked[10027] = data_i[10027] & sel_one_hot_i[78];
  assign data_masked[10026] = data_i[10026] & sel_one_hot_i[78];
  assign data_masked[10025] = data_i[10025] & sel_one_hot_i[78];
  assign data_masked[10024] = data_i[10024] & sel_one_hot_i[78];
  assign data_masked[10023] = data_i[10023] & sel_one_hot_i[78];
  assign data_masked[10022] = data_i[10022] & sel_one_hot_i[78];
  assign data_masked[10021] = data_i[10021] & sel_one_hot_i[78];
  assign data_masked[10020] = data_i[10020] & sel_one_hot_i[78];
  assign data_masked[10019] = data_i[10019] & sel_one_hot_i[78];
  assign data_masked[10018] = data_i[10018] & sel_one_hot_i[78];
  assign data_masked[10017] = data_i[10017] & sel_one_hot_i[78];
  assign data_masked[10016] = data_i[10016] & sel_one_hot_i[78];
  assign data_masked[10015] = data_i[10015] & sel_one_hot_i[78];
  assign data_masked[10014] = data_i[10014] & sel_one_hot_i[78];
  assign data_masked[10013] = data_i[10013] & sel_one_hot_i[78];
  assign data_masked[10012] = data_i[10012] & sel_one_hot_i[78];
  assign data_masked[10011] = data_i[10011] & sel_one_hot_i[78];
  assign data_masked[10010] = data_i[10010] & sel_one_hot_i[78];
  assign data_masked[10009] = data_i[10009] & sel_one_hot_i[78];
  assign data_masked[10008] = data_i[10008] & sel_one_hot_i[78];
  assign data_masked[10007] = data_i[10007] & sel_one_hot_i[78];
  assign data_masked[10006] = data_i[10006] & sel_one_hot_i[78];
  assign data_masked[10005] = data_i[10005] & sel_one_hot_i[78];
  assign data_masked[10004] = data_i[10004] & sel_one_hot_i[78];
  assign data_masked[10003] = data_i[10003] & sel_one_hot_i[78];
  assign data_masked[10002] = data_i[10002] & sel_one_hot_i[78];
  assign data_masked[10001] = data_i[10001] & sel_one_hot_i[78];
  assign data_masked[10000] = data_i[10000] & sel_one_hot_i[78];
  assign data_masked[9999] = data_i[9999] & sel_one_hot_i[78];
  assign data_masked[9998] = data_i[9998] & sel_one_hot_i[78];
  assign data_masked[9997] = data_i[9997] & sel_one_hot_i[78];
  assign data_masked[9996] = data_i[9996] & sel_one_hot_i[78];
  assign data_masked[9995] = data_i[9995] & sel_one_hot_i[78];
  assign data_masked[9994] = data_i[9994] & sel_one_hot_i[78];
  assign data_masked[9993] = data_i[9993] & sel_one_hot_i[78];
  assign data_masked[9992] = data_i[9992] & sel_one_hot_i[78];
  assign data_masked[9991] = data_i[9991] & sel_one_hot_i[78];
  assign data_masked[9990] = data_i[9990] & sel_one_hot_i[78];
  assign data_masked[9989] = data_i[9989] & sel_one_hot_i[78];
  assign data_masked[9988] = data_i[9988] & sel_one_hot_i[78];
  assign data_masked[9987] = data_i[9987] & sel_one_hot_i[78];
  assign data_masked[9986] = data_i[9986] & sel_one_hot_i[78];
  assign data_masked[9985] = data_i[9985] & sel_one_hot_i[78];
  assign data_masked[9984] = data_i[9984] & sel_one_hot_i[78];
  assign data_masked[10239] = data_i[10239] & sel_one_hot_i[79];
  assign data_masked[10238] = data_i[10238] & sel_one_hot_i[79];
  assign data_masked[10237] = data_i[10237] & sel_one_hot_i[79];
  assign data_masked[10236] = data_i[10236] & sel_one_hot_i[79];
  assign data_masked[10235] = data_i[10235] & sel_one_hot_i[79];
  assign data_masked[10234] = data_i[10234] & sel_one_hot_i[79];
  assign data_masked[10233] = data_i[10233] & sel_one_hot_i[79];
  assign data_masked[10232] = data_i[10232] & sel_one_hot_i[79];
  assign data_masked[10231] = data_i[10231] & sel_one_hot_i[79];
  assign data_masked[10230] = data_i[10230] & sel_one_hot_i[79];
  assign data_masked[10229] = data_i[10229] & sel_one_hot_i[79];
  assign data_masked[10228] = data_i[10228] & sel_one_hot_i[79];
  assign data_masked[10227] = data_i[10227] & sel_one_hot_i[79];
  assign data_masked[10226] = data_i[10226] & sel_one_hot_i[79];
  assign data_masked[10225] = data_i[10225] & sel_one_hot_i[79];
  assign data_masked[10224] = data_i[10224] & sel_one_hot_i[79];
  assign data_masked[10223] = data_i[10223] & sel_one_hot_i[79];
  assign data_masked[10222] = data_i[10222] & sel_one_hot_i[79];
  assign data_masked[10221] = data_i[10221] & sel_one_hot_i[79];
  assign data_masked[10220] = data_i[10220] & sel_one_hot_i[79];
  assign data_masked[10219] = data_i[10219] & sel_one_hot_i[79];
  assign data_masked[10218] = data_i[10218] & sel_one_hot_i[79];
  assign data_masked[10217] = data_i[10217] & sel_one_hot_i[79];
  assign data_masked[10216] = data_i[10216] & sel_one_hot_i[79];
  assign data_masked[10215] = data_i[10215] & sel_one_hot_i[79];
  assign data_masked[10214] = data_i[10214] & sel_one_hot_i[79];
  assign data_masked[10213] = data_i[10213] & sel_one_hot_i[79];
  assign data_masked[10212] = data_i[10212] & sel_one_hot_i[79];
  assign data_masked[10211] = data_i[10211] & sel_one_hot_i[79];
  assign data_masked[10210] = data_i[10210] & sel_one_hot_i[79];
  assign data_masked[10209] = data_i[10209] & sel_one_hot_i[79];
  assign data_masked[10208] = data_i[10208] & sel_one_hot_i[79];
  assign data_masked[10207] = data_i[10207] & sel_one_hot_i[79];
  assign data_masked[10206] = data_i[10206] & sel_one_hot_i[79];
  assign data_masked[10205] = data_i[10205] & sel_one_hot_i[79];
  assign data_masked[10204] = data_i[10204] & sel_one_hot_i[79];
  assign data_masked[10203] = data_i[10203] & sel_one_hot_i[79];
  assign data_masked[10202] = data_i[10202] & sel_one_hot_i[79];
  assign data_masked[10201] = data_i[10201] & sel_one_hot_i[79];
  assign data_masked[10200] = data_i[10200] & sel_one_hot_i[79];
  assign data_masked[10199] = data_i[10199] & sel_one_hot_i[79];
  assign data_masked[10198] = data_i[10198] & sel_one_hot_i[79];
  assign data_masked[10197] = data_i[10197] & sel_one_hot_i[79];
  assign data_masked[10196] = data_i[10196] & sel_one_hot_i[79];
  assign data_masked[10195] = data_i[10195] & sel_one_hot_i[79];
  assign data_masked[10194] = data_i[10194] & sel_one_hot_i[79];
  assign data_masked[10193] = data_i[10193] & sel_one_hot_i[79];
  assign data_masked[10192] = data_i[10192] & sel_one_hot_i[79];
  assign data_masked[10191] = data_i[10191] & sel_one_hot_i[79];
  assign data_masked[10190] = data_i[10190] & sel_one_hot_i[79];
  assign data_masked[10189] = data_i[10189] & sel_one_hot_i[79];
  assign data_masked[10188] = data_i[10188] & sel_one_hot_i[79];
  assign data_masked[10187] = data_i[10187] & sel_one_hot_i[79];
  assign data_masked[10186] = data_i[10186] & sel_one_hot_i[79];
  assign data_masked[10185] = data_i[10185] & sel_one_hot_i[79];
  assign data_masked[10184] = data_i[10184] & sel_one_hot_i[79];
  assign data_masked[10183] = data_i[10183] & sel_one_hot_i[79];
  assign data_masked[10182] = data_i[10182] & sel_one_hot_i[79];
  assign data_masked[10181] = data_i[10181] & sel_one_hot_i[79];
  assign data_masked[10180] = data_i[10180] & sel_one_hot_i[79];
  assign data_masked[10179] = data_i[10179] & sel_one_hot_i[79];
  assign data_masked[10178] = data_i[10178] & sel_one_hot_i[79];
  assign data_masked[10177] = data_i[10177] & sel_one_hot_i[79];
  assign data_masked[10176] = data_i[10176] & sel_one_hot_i[79];
  assign data_masked[10175] = data_i[10175] & sel_one_hot_i[79];
  assign data_masked[10174] = data_i[10174] & sel_one_hot_i[79];
  assign data_masked[10173] = data_i[10173] & sel_one_hot_i[79];
  assign data_masked[10172] = data_i[10172] & sel_one_hot_i[79];
  assign data_masked[10171] = data_i[10171] & sel_one_hot_i[79];
  assign data_masked[10170] = data_i[10170] & sel_one_hot_i[79];
  assign data_masked[10169] = data_i[10169] & sel_one_hot_i[79];
  assign data_masked[10168] = data_i[10168] & sel_one_hot_i[79];
  assign data_masked[10167] = data_i[10167] & sel_one_hot_i[79];
  assign data_masked[10166] = data_i[10166] & sel_one_hot_i[79];
  assign data_masked[10165] = data_i[10165] & sel_one_hot_i[79];
  assign data_masked[10164] = data_i[10164] & sel_one_hot_i[79];
  assign data_masked[10163] = data_i[10163] & sel_one_hot_i[79];
  assign data_masked[10162] = data_i[10162] & sel_one_hot_i[79];
  assign data_masked[10161] = data_i[10161] & sel_one_hot_i[79];
  assign data_masked[10160] = data_i[10160] & sel_one_hot_i[79];
  assign data_masked[10159] = data_i[10159] & sel_one_hot_i[79];
  assign data_masked[10158] = data_i[10158] & sel_one_hot_i[79];
  assign data_masked[10157] = data_i[10157] & sel_one_hot_i[79];
  assign data_masked[10156] = data_i[10156] & sel_one_hot_i[79];
  assign data_masked[10155] = data_i[10155] & sel_one_hot_i[79];
  assign data_masked[10154] = data_i[10154] & sel_one_hot_i[79];
  assign data_masked[10153] = data_i[10153] & sel_one_hot_i[79];
  assign data_masked[10152] = data_i[10152] & sel_one_hot_i[79];
  assign data_masked[10151] = data_i[10151] & sel_one_hot_i[79];
  assign data_masked[10150] = data_i[10150] & sel_one_hot_i[79];
  assign data_masked[10149] = data_i[10149] & sel_one_hot_i[79];
  assign data_masked[10148] = data_i[10148] & sel_one_hot_i[79];
  assign data_masked[10147] = data_i[10147] & sel_one_hot_i[79];
  assign data_masked[10146] = data_i[10146] & sel_one_hot_i[79];
  assign data_masked[10145] = data_i[10145] & sel_one_hot_i[79];
  assign data_masked[10144] = data_i[10144] & sel_one_hot_i[79];
  assign data_masked[10143] = data_i[10143] & sel_one_hot_i[79];
  assign data_masked[10142] = data_i[10142] & sel_one_hot_i[79];
  assign data_masked[10141] = data_i[10141] & sel_one_hot_i[79];
  assign data_masked[10140] = data_i[10140] & sel_one_hot_i[79];
  assign data_masked[10139] = data_i[10139] & sel_one_hot_i[79];
  assign data_masked[10138] = data_i[10138] & sel_one_hot_i[79];
  assign data_masked[10137] = data_i[10137] & sel_one_hot_i[79];
  assign data_masked[10136] = data_i[10136] & sel_one_hot_i[79];
  assign data_masked[10135] = data_i[10135] & sel_one_hot_i[79];
  assign data_masked[10134] = data_i[10134] & sel_one_hot_i[79];
  assign data_masked[10133] = data_i[10133] & sel_one_hot_i[79];
  assign data_masked[10132] = data_i[10132] & sel_one_hot_i[79];
  assign data_masked[10131] = data_i[10131] & sel_one_hot_i[79];
  assign data_masked[10130] = data_i[10130] & sel_one_hot_i[79];
  assign data_masked[10129] = data_i[10129] & sel_one_hot_i[79];
  assign data_masked[10128] = data_i[10128] & sel_one_hot_i[79];
  assign data_masked[10127] = data_i[10127] & sel_one_hot_i[79];
  assign data_masked[10126] = data_i[10126] & sel_one_hot_i[79];
  assign data_masked[10125] = data_i[10125] & sel_one_hot_i[79];
  assign data_masked[10124] = data_i[10124] & sel_one_hot_i[79];
  assign data_masked[10123] = data_i[10123] & sel_one_hot_i[79];
  assign data_masked[10122] = data_i[10122] & sel_one_hot_i[79];
  assign data_masked[10121] = data_i[10121] & sel_one_hot_i[79];
  assign data_masked[10120] = data_i[10120] & sel_one_hot_i[79];
  assign data_masked[10119] = data_i[10119] & sel_one_hot_i[79];
  assign data_masked[10118] = data_i[10118] & sel_one_hot_i[79];
  assign data_masked[10117] = data_i[10117] & sel_one_hot_i[79];
  assign data_masked[10116] = data_i[10116] & sel_one_hot_i[79];
  assign data_masked[10115] = data_i[10115] & sel_one_hot_i[79];
  assign data_masked[10114] = data_i[10114] & sel_one_hot_i[79];
  assign data_masked[10113] = data_i[10113] & sel_one_hot_i[79];
  assign data_masked[10112] = data_i[10112] & sel_one_hot_i[79];
  assign data_masked[10367] = data_i[10367] & sel_one_hot_i[80];
  assign data_masked[10366] = data_i[10366] & sel_one_hot_i[80];
  assign data_masked[10365] = data_i[10365] & sel_one_hot_i[80];
  assign data_masked[10364] = data_i[10364] & sel_one_hot_i[80];
  assign data_masked[10363] = data_i[10363] & sel_one_hot_i[80];
  assign data_masked[10362] = data_i[10362] & sel_one_hot_i[80];
  assign data_masked[10361] = data_i[10361] & sel_one_hot_i[80];
  assign data_masked[10360] = data_i[10360] & sel_one_hot_i[80];
  assign data_masked[10359] = data_i[10359] & sel_one_hot_i[80];
  assign data_masked[10358] = data_i[10358] & sel_one_hot_i[80];
  assign data_masked[10357] = data_i[10357] & sel_one_hot_i[80];
  assign data_masked[10356] = data_i[10356] & sel_one_hot_i[80];
  assign data_masked[10355] = data_i[10355] & sel_one_hot_i[80];
  assign data_masked[10354] = data_i[10354] & sel_one_hot_i[80];
  assign data_masked[10353] = data_i[10353] & sel_one_hot_i[80];
  assign data_masked[10352] = data_i[10352] & sel_one_hot_i[80];
  assign data_masked[10351] = data_i[10351] & sel_one_hot_i[80];
  assign data_masked[10350] = data_i[10350] & sel_one_hot_i[80];
  assign data_masked[10349] = data_i[10349] & sel_one_hot_i[80];
  assign data_masked[10348] = data_i[10348] & sel_one_hot_i[80];
  assign data_masked[10347] = data_i[10347] & sel_one_hot_i[80];
  assign data_masked[10346] = data_i[10346] & sel_one_hot_i[80];
  assign data_masked[10345] = data_i[10345] & sel_one_hot_i[80];
  assign data_masked[10344] = data_i[10344] & sel_one_hot_i[80];
  assign data_masked[10343] = data_i[10343] & sel_one_hot_i[80];
  assign data_masked[10342] = data_i[10342] & sel_one_hot_i[80];
  assign data_masked[10341] = data_i[10341] & sel_one_hot_i[80];
  assign data_masked[10340] = data_i[10340] & sel_one_hot_i[80];
  assign data_masked[10339] = data_i[10339] & sel_one_hot_i[80];
  assign data_masked[10338] = data_i[10338] & sel_one_hot_i[80];
  assign data_masked[10337] = data_i[10337] & sel_one_hot_i[80];
  assign data_masked[10336] = data_i[10336] & sel_one_hot_i[80];
  assign data_masked[10335] = data_i[10335] & sel_one_hot_i[80];
  assign data_masked[10334] = data_i[10334] & sel_one_hot_i[80];
  assign data_masked[10333] = data_i[10333] & sel_one_hot_i[80];
  assign data_masked[10332] = data_i[10332] & sel_one_hot_i[80];
  assign data_masked[10331] = data_i[10331] & sel_one_hot_i[80];
  assign data_masked[10330] = data_i[10330] & sel_one_hot_i[80];
  assign data_masked[10329] = data_i[10329] & sel_one_hot_i[80];
  assign data_masked[10328] = data_i[10328] & sel_one_hot_i[80];
  assign data_masked[10327] = data_i[10327] & sel_one_hot_i[80];
  assign data_masked[10326] = data_i[10326] & sel_one_hot_i[80];
  assign data_masked[10325] = data_i[10325] & sel_one_hot_i[80];
  assign data_masked[10324] = data_i[10324] & sel_one_hot_i[80];
  assign data_masked[10323] = data_i[10323] & sel_one_hot_i[80];
  assign data_masked[10322] = data_i[10322] & sel_one_hot_i[80];
  assign data_masked[10321] = data_i[10321] & sel_one_hot_i[80];
  assign data_masked[10320] = data_i[10320] & sel_one_hot_i[80];
  assign data_masked[10319] = data_i[10319] & sel_one_hot_i[80];
  assign data_masked[10318] = data_i[10318] & sel_one_hot_i[80];
  assign data_masked[10317] = data_i[10317] & sel_one_hot_i[80];
  assign data_masked[10316] = data_i[10316] & sel_one_hot_i[80];
  assign data_masked[10315] = data_i[10315] & sel_one_hot_i[80];
  assign data_masked[10314] = data_i[10314] & sel_one_hot_i[80];
  assign data_masked[10313] = data_i[10313] & sel_one_hot_i[80];
  assign data_masked[10312] = data_i[10312] & sel_one_hot_i[80];
  assign data_masked[10311] = data_i[10311] & sel_one_hot_i[80];
  assign data_masked[10310] = data_i[10310] & sel_one_hot_i[80];
  assign data_masked[10309] = data_i[10309] & sel_one_hot_i[80];
  assign data_masked[10308] = data_i[10308] & sel_one_hot_i[80];
  assign data_masked[10307] = data_i[10307] & sel_one_hot_i[80];
  assign data_masked[10306] = data_i[10306] & sel_one_hot_i[80];
  assign data_masked[10305] = data_i[10305] & sel_one_hot_i[80];
  assign data_masked[10304] = data_i[10304] & sel_one_hot_i[80];
  assign data_masked[10303] = data_i[10303] & sel_one_hot_i[80];
  assign data_masked[10302] = data_i[10302] & sel_one_hot_i[80];
  assign data_masked[10301] = data_i[10301] & sel_one_hot_i[80];
  assign data_masked[10300] = data_i[10300] & sel_one_hot_i[80];
  assign data_masked[10299] = data_i[10299] & sel_one_hot_i[80];
  assign data_masked[10298] = data_i[10298] & sel_one_hot_i[80];
  assign data_masked[10297] = data_i[10297] & sel_one_hot_i[80];
  assign data_masked[10296] = data_i[10296] & sel_one_hot_i[80];
  assign data_masked[10295] = data_i[10295] & sel_one_hot_i[80];
  assign data_masked[10294] = data_i[10294] & sel_one_hot_i[80];
  assign data_masked[10293] = data_i[10293] & sel_one_hot_i[80];
  assign data_masked[10292] = data_i[10292] & sel_one_hot_i[80];
  assign data_masked[10291] = data_i[10291] & sel_one_hot_i[80];
  assign data_masked[10290] = data_i[10290] & sel_one_hot_i[80];
  assign data_masked[10289] = data_i[10289] & sel_one_hot_i[80];
  assign data_masked[10288] = data_i[10288] & sel_one_hot_i[80];
  assign data_masked[10287] = data_i[10287] & sel_one_hot_i[80];
  assign data_masked[10286] = data_i[10286] & sel_one_hot_i[80];
  assign data_masked[10285] = data_i[10285] & sel_one_hot_i[80];
  assign data_masked[10284] = data_i[10284] & sel_one_hot_i[80];
  assign data_masked[10283] = data_i[10283] & sel_one_hot_i[80];
  assign data_masked[10282] = data_i[10282] & sel_one_hot_i[80];
  assign data_masked[10281] = data_i[10281] & sel_one_hot_i[80];
  assign data_masked[10280] = data_i[10280] & sel_one_hot_i[80];
  assign data_masked[10279] = data_i[10279] & sel_one_hot_i[80];
  assign data_masked[10278] = data_i[10278] & sel_one_hot_i[80];
  assign data_masked[10277] = data_i[10277] & sel_one_hot_i[80];
  assign data_masked[10276] = data_i[10276] & sel_one_hot_i[80];
  assign data_masked[10275] = data_i[10275] & sel_one_hot_i[80];
  assign data_masked[10274] = data_i[10274] & sel_one_hot_i[80];
  assign data_masked[10273] = data_i[10273] & sel_one_hot_i[80];
  assign data_masked[10272] = data_i[10272] & sel_one_hot_i[80];
  assign data_masked[10271] = data_i[10271] & sel_one_hot_i[80];
  assign data_masked[10270] = data_i[10270] & sel_one_hot_i[80];
  assign data_masked[10269] = data_i[10269] & sel_one_hot_i[80];
  assign data_masked[10268] = data_i[10268] & sel_one_hot_i[80];
  assign data_masked[10267] = data_i[10267] & sel_one_hot_i[80];
  assign data_masked[10266] = data_i[10266] & sel_one_hot_i[80];
  assign data_masked[10265] = data_i[10265] & sel_one_hot_i[80];
  assign data_masked[10264] = data_i[10264] & sel_one_hot_i[80];
  assign data_masked[10263] = data_i[10263] & sel_one_hot_i[80];
  assign data_masked[10262] = data_i[10262] & sel_one_hot_i[80];
  assign data_masked[10261] = data_i[10261] & sel_one_hot_i[80];
  assign data_masked[10260] = data_i[10260] & sel_one_hot_i[80];
  assign data_masked[10259] = data_i[10259] & sel_one_hot_i[80];
  assign data_masked[10258] = data_i[10258] & sel_one_hot_i[80];
  assign data_masked[10257] = data_i[10257] & sel_one_hot_i[80];
  assign data_masked[10256] = data_i[10256] & sel_one_hot_i[80];
  assign data_masked[10255] = data_i[10255] & sel_one_hot_i[80];
  assign data_masked[10254] = data_i[10254] & sel_one_hot_i[80];
  assign data_masked[10253] = data_i[10253] & sel_one_hot_i[80];
  assign data_masked[10252] = data_i[10252] & sel_one_hot_i[80];
  assign data_masked[10251] = data_i[10251] & sel_one_hot_i[80];
  assign data_masked[10250] = data_i[10250] & sel_one_hot_i[80];
  assign data_masked[10249] = data_i[10249] & sel_one_hot_i[80];
  assign data_masked[10248] = data_i[10248] & sel_one_hot_i[80];
  assign data_masked[10247] = data_i[10247] & sel_one_hot_i[80];
  assign data_masked[10246] = data_i[10246] & sel_one_hot_i[80];
  assign data_masked[10245] = data_i[10245] & sel_one_hot_i[80];
  assign data_masked[10244] = data_i[10244] & sel_one_hot_i[80];
  assign data_masked[10243] = data_i[10243] & sel_one_hot_i[80];
  assign data_masked[10242] = data_i[10242] & sel_one_hot_i[80];
  assign data_masked[10241] = data_i[10241] & sel_one_hot_i[80];
  assign data_masked[10240] = data_i[10240] & sel_one_hot_i[80];
  assign data_masked[10495] = data_i[10495] & sel_one_hot_i[81];
  assign data_masked[10494] = data_i[10494] & sel_one_hot_i[81];
  assign data_masked[10493] = data_i[10493] & sel_one_hot_i[81];
  assign data_masked[10492] = data_i[10492] & sel_one_hot_i[81];
  assign data_masked[10491] = data_i[10491] & sel_one_hot_i[81];
  assign data_masked[10490] = data_i[10490] & sel_one_hot_i[81];
  assign data_masked[10489] = data_i[10489] & sel_one_hot_i[81];
  assign data_masked[10488] = data_i[10488] & sel_one_hot_i[81];
  assign data_masked[10487] = data_i[10487] & sel_one_hot_i[81];
  assign data_masked[10486] = data_i[10486] & sel_one_hot_i[81];
  assign data_masked[10485] = data_i[10485] & sel_one_hot_i[81];
  assign data_masked[10484] = data_i[10484] & sel_one_hot_i[81];
  assign data_masked[10483] = data_i[10483] & sel_one_hot_i[81];
  assign data_masked[10482] = data_i[10482] & sel_one_hot_i[81];
  assign data_masked[10481] = data_i[10481] & sel_one_hot_i[81];
  assign data_masked[10480] = data_i[10480] & sel_one_hot_i[81];
  assign data_masked[10479] = data_i[10479] & sel_one_hot_i[81];
  assign data_masked[10478] = data_i[10478] & sel_one_hot_i[81];
  assign data_masked[10477] = data_i[10477] & sel_one_hot_i[81];
  assign data_masked[10476] = data_i[10476] & sel_one_hot_i[81];
  assign data_masked[10475] = data_i[10475] & sel_one_hot_i[81];
  assign data_masked[10474] = data_i[10474] & sel_one_hot_i[81];
  assign data_masked[10473] = data_i[10473] & sel_one_hot_i[81];
  assign data_masked[10472] = data_i[10472] & sel_one_hot_i[81];
  assign data_masked[10471] = data_i[10471] & sel_one_hot_i[81];
  assign data_masked[10470] = data_i[10470] & sel_one_hot_i[81];
  assign data_masked[10469] = data_i[10469] & sel_one_hot_i[81];
  assign data_masked[10468] = data_i[10468] & sel_one_hot_i[81];
  assign data_masked[10467] = data_i[10467] & sel_one_hot_i[81];
  assign data_masked[10466] = data_i[10466] & sel_one_hot_i[81];
  assign data_masked[10465] = data_i[10465] & sel_one_hot_i[81];
  assign data_masked[10464] = data_i[10464] & sel_one_hot_i[81];
  assign data_masked[10463] = data_i[10463] & sel_one_hot_i[81];
  assign data_masked[10462] = data_i[10462] & sel_one_hot_i[81];
  assign data_masked[10461] = data_i[10461] & sel_one_hot_i[81];
  assign data_masked[10460] = data_i[10460] & sel_one_hot_i[81];
  assign data_masked[10459] = data_i[10459] & sel_one_hot_i[81];
  assign data_masked[10458] = data_i[10458] & sel_one_hot_i[81];
  assign data_masked[10457] = data_i[10457] & sel_one_hot_i[81];
  assign data_masked[10456] = data_i[10456] & sel_one_hot_i[81];
  assign data_masked[10455] = data_i[10455] & sel_one_hot_i[81];
  assign data_masked[10454] = data_i[10454] & sel_one_hot_i[81];
  assign data_masked[10453] = data_i[10453] & sel_one_hot_i[81];
  assign data_masked[10452] = data_i[10452] & sel_one_hot_i[81];
  assign data_masked[10451] = data_i[10451] & sel_one_hot_i[81];
  assign data_masked[10450] = data_i[10450] & sel_one_hot_i[81];
  assign data_masked[10449] = data_i[10449] & sel_one_hot_i[81];
  assign data_masked[10448] = data_i[10448] & sel_one_hot_i[81];
  assign data_masked[10447] = data_i[10447] & sel_one_hot_i[81];
  assign data_masked[10446] = data_i[10446] & sel_one_hot_i[81];
  assign data_masked[10445] = data_i[10445] & sel_one_hot_i[81];
  assign data_masked[10444] = data_i[10444] & sel_one_hot_i[81];
  assign data_masked[10443] = data_i[10443] & sel_one_hot_i[81];
  assign data_masked[10442] = data_i[10442] & sel_one_hot_i[81];
  assign data_masked[10441] = data_i[10441] & sel_one_hot_i[81];
  assign data_masked[10440] = data_i[10440] & sel_one_hot_i[81];
  assign data_masked[10439] = data_i[10439] & sel_one_hot_i[81];
  assign data_masked[10438] = data_i[10438] & sel_one_hot_i[81];
  assign data_masked[10437] = data_i[10437] & sel_one_hot_i[81];
  assign data_masked[10436] = data_i[10436] & sel_one_hot_i[81];
  assign data_masked[10435] = data_i[10435] & sel_one_hot_i[81];
  assign data_masked[10434] = data_i[10434] & sel_one_hot_i[81];
  assign data_masked[10433] = data_i[10433] & sel_one_hot_i[81];
  assign data_masked[10432] = data_i[10432] & sel_one_hot_i[81];
  assign data_masked[10431] = data_i[10431] & sel_one_hot_i[81];
  assign data_masked[10430] = data_i[10430] & sel_one_hot_i[81];
  assign data_masked[10429] = data_i[10429] & sel_one_hot_i[81];
  assign data_masked[10428] = data_i[10428] & sel_one_hot_i[81];
  assign data_masked[10427] = data_i[10427] & sel_one_hot_i[81];
  assign data_masked[10426] = data_i[10426] & sel_one_hot_i[81];
  assign data_masked[10425] = data_i[10425] & sel_one_hot_i[81];
  assign data_masked[10424] = data_i[10424] & sel_one_hot_i[81];
  assign data_masked[10423] = data_i[10423] & sel_one_hot_i[81];
  assign data_masked[10422] = data_i[10422] & sel_one_hot_i[81];
  assign data_masked[10421] = data_i[10421] & sel_one_hot_i[81];
  assign data_masked[10420] = data_i[10420] & sel_one_hot_i[81];
  assign data_masked[10419] = data_i[10419] & sel_one_hot_i[81];
  assign data_masked[10418] = data_i[10418] & sel_one_hot_i[81];
  assign data_masked[10417] = data_i[10417] & sel_one_hot_i[81];
  assign data_masked[10416] = data_i[10416] & sel_one_hot_i[81];
  assign data_masked[10415] = data_i[10415] & sel_one_hot_i[81];
  assign data_masked[10414] = data_i[10414] & sel_one_hot_i[81];
  assign data_masked[10413] = data_i[10413] & sel_one_hot_i[81];
  assign data_masked[10412] = data_i[10412] & sel_one_hot_i[81];
  assign data_masked[10411] = data_i[10411] & sel_one_hot_i[81];
  assign data_masked[10410] = data_i[10410] & sel_one_hot_i[81];
  assign data_masked[10409] = data_i[10409] & sel_one_hot_i[81];
  assign data_masked[10408] = data_i[10408] & sel_one_hot_i[81];
  assign data_masked[10407] = data_i[10407] & sel_one_hot_i[81];
  assign data_masked[10406] = data_i[10406] & sel_one_hot_i[81];
  assign data_masked[10405] = data_i[10405] & sel_one_hot_i[81];
  assign data_masked[10404] = data_i[10404] & sel_one_hot_i[81];
  assign data_masked[10403] = data_i[10403] & sel_one_hot_i[81];
  assign data_masked[10402] = data_i[10402] & sel_one_hot_i[81];
  assign data_masked[10401] = data_i[10401] & sel_one_hot_i[81];
  assign data_masked[10400] = data_i[10400] & sel_one_hot_i[81];
  assign data_masked[10399] = data_i[10399] & sel_one_hot_i[81];
  assign data_masked[10398] = data_i[10398] & sel_one_hot_i[81];
  assign data_masked[10397] = data_i[10397] & sel_one_hot_i[81];
  assign data_masked[10396] = data_i[10396] & sel_one_hot_i[81];
  assign data_masked[10395] = data_i[10395] & sel_one_hot_i[81];
  assign data_masked[10394] = data_i[10394] & sel_one_hot_i[81];
  assign data_masked[10393] = data_i[10393] & sel_one_hot_i[81];
  assign data_masked[10392] = data_i[10392] & sel_one_hot_i[81];
  assign data_masked[10391] = data_i[10391] & sel_one_hot_i[81];
  assign data_masked[10390] = data_i[10390] & sel_one_hot_i[81];
  assign data_masked[10389] = data_i[10389] & sel_one_hot_i[81];
  assign data_masked[10388] = data_i[10388] & sel_one_hot_i[81];
  assign data_masked[10387] = data_i[10387] & sel_one_hot_i[81];
  assign data_masked[10386] = data_i[10386] & sel_one_hot_i[81];
  assign data_masked[10385] = data_i[10385] & sel_one_hot_i[81];
  assign data_masked[10384] = data_i[10384] & sel_one_hot_i[81];
  assign data_masked[10383] = data_i[10383] & sel_one_hot_i[81];
  assign data_masked[10382] = data_i[10382] & sel_one_hot_i[81];
  assign data_masked[10381] = data_i[10381] & sel_one_hot_i[81];
  assign data_masked[10380] = data_i[10380] & sel_one_hot_i[81];
  assign data_masked[10379] = data_i[10379] & sel_one_hot_i[81];
  assign data_masked[10378] = data_i[10378] & sel_one_hot_i[81];
  assign data_masked[10377] = data_i[10377] & sel_one_hot_i[81];
  assign data_masked[10376] = data_i[10376] & sel_one_hot_i[81];
  assign data_masked[10375] = data_i[10375] & sel_one_hot_i[81];
  assign data_masked[10374] = data_i[10374] & sel_one_hot_i[81];
  assign data_masked[10373] = data_i[10373] & sel_one_hot_i[81];
  assign data_masked[10372] = data_i[10372] & sel_one_hot_i[81];
  assign data_masked[10371] = data_i[10371] & sel_one_hot_i[81];
  assign data_masked[10370] = data_i[10370] & sel_one_hot_i[81];
  assign data_masked[10369] = data_i[10369] & sel_one_hot_i[81];
  assign data_masked[10368] = data_i[10368] & sel_one_hot_i[81];
  assign data_masked[10623] = data_i[10623] & sel_one_hot_i[82];
  assign data_masked[10622] = data_i[10622] & sel_one_hot_i[82];
  assign data_masked[10621] = data_i[10621] & sel_one_hot_i[82];
  assign data_masked[10620] = data_i[10620] & sel_one_hot_i[82];
  assign data_masked[10619] = data_i[10619] & sel_one_hot_i[82];
  assign data_masked[10618] = data_i[10618] & sel_one_hot_i[82];
  assign data_masked[10617] = data_i[10617] & sel_one_hot_i[82];
  assign data_masked[10616] = data_i[10616] & sel_one_hot_i[82];
  assign data_masked[10615] = data_i[10615] & sel_one_hot_i[82];
  assign data_masked[10614] = data_i[10614] & sel_one_hot_i[82];
  assign data_masked[10613] = data_i[10613] & sel_one_hot_i[82];
  assign data_masked[10612] = data_i[10612] & sel_one_hot_i[82];
  assign data_masked[10611] = data_i[10611] & sel_one_hot_i[82];
  assign data_masked[10610] = data_i[10610] & sel_one_hot_i[82];
  assign data_masked[10609] = data_i[10609] & sel_one_hot_i[82];
  assign data_masked[10608] = data_i[10608] & sel_one_hot_i[82];
  assign data_masked[10607] = data_i[10607] & sel_one_hot_i[82];
  assign data_masked[10606] = data_i[10606] & sel_one_hot_i[82];
  assign data_masked[10605] = data_i[10605] & sel_one_hot_i[82];
  assign data_masked[10604] = data_i[10604] & sel_one_hot_i[82];
  assign data_masked[10603] = data_i[10603] & sel_one_hot_i[82];
  assign data_masked[10602] = data_i[10602] & sel_one_hot_i[82];
  assign data_masked[10601] = data_i[10601] & sel_one_hot_i[82];
  assign data_masked[10600] = data_i[10600] & sel_one_hot_i[82];
  assign data_masked[10599] = data_i[10599] & sel_one_hot_i[82];
  assign data_masked[10598] = data_i[10598] & sel_one_hot_i[82];
  assign data_masked[10597] = data_i[10597] & sel_one_hot_i[82];
  assign data_masked[10596] = data_i[10596] & sel_one_hot_i[82];
  assign data_masked[10595] = data_i[10595] & sel_one_hot_i[82];
  assign data_masked[10594] = data_i[10594] & sel_one_hot_i[82];
  assign data_masked[10593] = data_i[10593] & sel_one_hot_i[82];
  assign data_masked[10592] = data_i[10592] & sel_one_hot_i[82];
  assign data_masked[10591] = data_i[10591] & sel_one_hot_i[82];
  assign data_masked[10590] = data_i[10590] & sel_one_hot_i[82];
  assign data_masked[10589] = data_i[10589] & sel_one_hot_i[82];
  assign data_masked[10588] = data_i[10588] & sel_one_hot_i[82];
  assign data_masked[10587] = data_i[10587] & sel_one_hot_i[82];
  assign data_masked[10586] = data_i[10586] & sel_one_hot_i[82];
  assign data_masked[10585] = data_i[10585] & sel_one_hot_i[82];
  assign data_masked[10584] = data_i[10584] & sel_one_hot_i[82];
  assign data_masked[10583] = data_i[10583] & sel_one_hot_i[82];
  assign data_masked[10582] = data_i[10582] & sel_one_hot_i[82];
  assign data_masked[10581] = data_i[10581] & sel_one_hot_i[82];
  assign data_masked[10580] = data_i[10580] & sel_one_hot_i[82];
  assign data_masked[10579] = data_i[10579] & sel_one_hot_i[82];
  assign data_masked[10578] = data_i[10578] & sel_one_hot_i[82];
  assign data_masked[10577] = data_i[10577] & sel_one_hot_i[82];
  assign data_masked[10576] = data_i[10576] & sel_one_hot_i[82];
  assign data_masked[10575] = data_i[10575] & sel_one_hot_i[82];
  assign data_masked[10574] = data_i[10574] & sel_one_hot_i[82];
  assign data_masked[10573] = data_i[10573] & sel_one_hot_i[82];
  assign data_masked[10572] = data_i[10572] & sel_one_hot_i[82];
  assign data_masked[10571] = data_i[10571] & sel_one_hot_i[82];
  assign data_masked[10570] = data_i[10570] & sel_one_hot_i[82];
  assign data_masked[10569] = data_i[10569] & sel_one_hot_i[82];
  assign data_masked[10568] = data_i[10568] & sel_one_hot_i[82];
  assign data_masked[10567] = data_i[10567] & sel_one_hot_i[82];
  assign data_masked[10566] = data_i[10566] & sel_one_hot_i[82];
  assign data_masked[10565] = data_i[10565] & sel_one_hot_i[82];
  assign data_masked[10564] = data_i[10564] & sel_one_hot_i[82];
  assign data_masked[10563] = data_i[10563] & sel_one_hot_i[82];
  assign data_masked[10562] = data_i[10562] & sel_one_hot_i[82];
  assign data_masked[10561] = data_i[10561] & sel_one_hot_i[82];
  assign data_masked[10560] = data_i[10560] & sel_one_hot_i[82];
  assign data_masked[10559] = data_i[10559] & sel_one_hot_i[82];
  assign data_masked[10558] = data_i[10558] & sel_one_hot_i[82];
  assign data_masked[10557] = data_i[10557] & sel_one_hot_i[82];
  assign data_masked[10556] = data_i[10556] & sel_one_hot_i[82];
  assign data_masked[10555] = data_i[10555] & sel_one_hot_i[82];
  assign data_masked[10554] = data_i[10554] & sel_one_hot_i[82];
  assign data_masked[10553] = data_i[10553] & sel_one_hot_i[82];
  assign data_masked[10552] = data_i[10552] & sel_one_hot_i[82];
  assign data_masked[10551] = data_i[10551] & sel_one_hot_i[82];
  assign data_masked[10550] = data_i[10550] & sel_one_hot_i[82];
  assign data_masked[10549] = data_i[10549] & sel_one_hot_i[82];
  assign data_masked[10548] = data_i[10548] & sel_one_hot_i[82];
  assign data_masked[10547] = data_i[10547] & sel_one_hot_i[82];
  assign data_masked[10546] = data_i[10546] & sel_one_hot_i[82];
  assign data_masked[10545] = data_i[10545] & sel_one_hot_i[82];
  assign data_masked[10544] = data_i[10544] & sel_one_hot_i[82];
  assign data_masked[10543] = data_i[10543] & sel_one_hot_i[82];
  assign data_masked[10542] = data_i[10542] & sel_one_hot_i[82];
  assign data_masked[10541] = data_i[10541] & sel_one_hot_i[82];
  assign data_masked[10540] = data_i[10540] & sel_one_hot_i[82];
  assign data_masked[10539] = data_i[10539] & sel_one_hot_i[82];
  assign data_masked[10538] = data_i[10538] & sel_one_hot_i[82];
  assign data_masked[10537] = data_i[10537] & sel_one_hot_i[82];
  assign data_masked[10536] = data_i[10536] & sel_one_hot_i[82];
  assign data_masked[10535] = data_i[10535] & sel_one_hot_i[82];
  assign data_masked[10534] = data_i[10534] & sel_one_hot_i[82];
  assign data_masked[10533] = data_i[10533] & sel_one_hot_i[82];
  assign data_masked[10532] = data_i[10532] & sel_one_hot_i[82];
  assign data_masked[10531] = data_i[10531] & sel_one_hot_i[82];
  assign data_masked[10530] = data_i[10530] & sel_one_hot_i[82];
  assign data_masked[10529] = data_i[10529] & sel_one_hot_i[82];
  assign data_masked[10528] = data_i[10528] & sel_one_hot_i[82];
  assign data_masked[10527] = data_i[10527] & sel_one_hot_i[82];
  assign data_masked[10526] = data_i[10526] & sel_one_hot_i[82];
  assign data_masked[10525] = data_i[10525] & sel_one_hot_i[82];
  assign data_masked[10524] = data_i[10524] & sel_one_hot_i[82];
  assign data_masked[10523] = data_i[10523] & sel_one_hot_i[82];
  assign data_masked[10522] = data_i[10522] & sel_one_hot_i[82];
  assign data_masked[10521] = data_i[10521] & sel_one_hot_i[82];
  assign data_masked[10520] = data_i[10520] & sel_one_hot_i[82];
  assign data_masked[10519] = data_i[10519] & sel_one_hot_i[82];
  assign data_masked[10518] = data_i[10518] & sel_one_hot_i[82];
  assign data_masked[10517] = data_i[10517] & sel_one_hot_i[82];
  assign data_masked[10516] = data_i[10516] & sel_one_hot_i[82];
  assign data_masked[10515] = data_i[10515] & sel_one_hot_i[82];
  assign data_masked[10514] = data_i[10514] & sel_one_hot_i[82];
  assign data_masked[10513] = data_i[10513] & sel_one_hot_i[82];
  assign data_masked[10512] = data_i[10512] & sel_one_hot_i[82];
  assign data_masked[10511] = data_i[10511] & sel_one_hot_i[82];
  assign data_masked[10510] = data_i[10510] & sel_one_hot_i[82];
  assign data_masked[10509] = data_i[10509] & sel_one_hot_i[82];
  assign data_masked[10508] = data_i[10508] & sel_one_hot_i[82];
  assign data_masked[10507] = data_i[10507] & sel_one_hot_i[82];
  assign data_masked[10506] = data_i[10506] & sel_one_hot_i[82];
  assign data_masked[10505] = data_i[10505] & sel_one_hot_i[82];
  assign data_masked[10504] = data_i[10504] & sel_one_hot_i[82];
  assign data_masked[10503] = data_i[10503] & sel_one_hot_i[82];
  assign data_masked[10502] = data_i[10502] & sel_one_hot_i[82];
  assign data_masked[10501] = data_i[10501] & sel_one_hot_i[82];
  assign data_masked[10500] = data_i[10500] & sel_one_hot_i[82];
  assign data_masked[10499] = data_i[10499] & sel_one_hot_i[82];
  assign data_masked[10498] = data_i[10498] & sel_one_hot_i[82];
  assign data_masked[10497] = data_i[10497] & sel_one_hot_i[82];
  assign data_masked[10496] = data_i[10496] & sel_one_hot_i[82];
  assign data_masked[10751] = data_i[10751] & sel_one_hot_i[83];
  assign data_masked[10750] = data_i[10750] & sel_one_hot_i[83];
  assign data_masked[10749] = data_i[10749] & sel_one_hot_i[83];
  assign data_masked[10748] = data_i[10748] & sel_one_hot_i[83];
  assign data_masked[10747] = data_i[10747] & sel_one_hot_i[83];
  assign data_masked[10746] = data_i[10746] & sel_one_hot_i[83];
  assign data_masked[10745] = data_i[10745] & sel_one_hot_i[83];
  assign data_masked[10744] = data_i[10744] & sel_one_hot_i[83];
  assign data_masked[10743] = data_i[10743] & sel_one_hot_i[83];
  assign data_masked[10742] = data_i[10742] & sel_one_hot_i[83];
  assign data_masked[10741] = data_i[10741] & sel_one_hot_i[83];
  assign data_masked[10740] = data_i[10740] & sel_one_hot_i[83];
  assign data_masked[10739] = data_i[10739] & sel_one_hot_i[83];
  assign data_masked[10738] = data_i[10738] & sel_one_hot_i[83];
  assign data_masked[10737] = data_i[10737] & sel_one_hot_i[83];
  assign data_masked[10736] = data_i[10736] & sel_one_hot_i[83];
  assign data_masked[10735] = data_i[10735] & sel_one_hot_i[83];
  assign data_masked[10734] = data_i[10734] & sel_one_hot_i[83];
  assign data_masked[10733] = data_i[10733] & sel_one_hot_i[83];
  assign data_masked[10732] = data_i[10732] & sel_one_hot_i[83];
  assign data_masked[10731] = data_i[10731] & sel_one_hot_i[83];
  assign data_masked[10730] = data_i[10730] & sel_one_hot_i[83];
  assign data_masked[10729] = data_i[10729] & sel_one_hot_i[83];
  assign data_masked[10728] = data_i[10728] & sel_one_hot_i[83];
  assign data_masked[10727] = data_i[10727] & sel_one_hot_i[83];
  assign data_masked[10726] = data_i[10726] & sel_one_hot_i[83];
  assign data_masked[10725] = data_i[10725] & sel_one_hot_i[83];
  assign data_masked[10724] = data_i[10724] & sel_one_hot_i[83];
  assign data_masked[10723] = data_i[10723] & sel_one_hot_i[83];
  assign data_masked[10722] = data_i[10722] & sel_one_hot_i[83];
  assign data_masked[10721] = data_i[10721] & sel_one_hot_i[83];
  assign data_masked[10720] = data_i[10720] & sel_one_hot_i[83];
  assign data_masked[10719] = data_i[10719] & sel_one_hot_i[83];
  assign data_masked[10718] = data_i[10718] & sel_one_hot_i[83];
  assign data_masked[10717] = data_i[10717] & sel_one_hot_i[83];
  assign data_masked[10716] = data_i[10716] & sel_one_hot_i[83];
  assign data_masked[10715] = data_i[10715] & sel_one_hot_i[83];
  assign data_masked[10714] = data_i[10714] & sel_one_hot_i[83];
  assign data_masked[10713] = data_i[10713] & sel_one_hot_i[83];
  assign data_masked[10712] = data_i[10712] & sel_one_hot_i[83];
  assign data_masked[10711] = data_i[10711] & sel_one_hot_i[83];
  assign data_masked[10710] = data_i[10710] & sel_one_hot_i[83];
  assign data_masked[10709] = data_i[10709] & sel_one_hot_i[83];
  assign data_masked[10708] = data_i[10708] & sel_one_hot_i[83];
  assign data_masked[10707] = data_i[10707] & sel_one_hot_i[83];
  assign data_masked[10706] = data_i[10706] & sel_one_hot_i[83];
  assign data_masked[10705] = data_i[10705] & sel_one_hot_i[83];
  assign data_masked[10704] = data_i[10704] & sel_one_hot_i[83];
  assign data_masked[10703] = data_i[10703] & sel_one_hot_i[83];
  assign data_masked[10702] = data_i[10702] & sel_one_hot_i[83];
  assign data_masked[10701] = data_i[10701] & sel_one_hot_i[83];
  assign data_masked[10700] = data_i[10700] & sel_one_hot_i[83];
  assign data_masked[10699] = data_i[10699] & sel_one_hot_i[83];
  assign data_masked[10698] = data_i[10698] & sel_one_hot_i[83];
  assign data_masked[10697] = data_i[10697] & sel_one_hot_i[83];
  assign data_masked[10696] = data_i[10696] & sel_one_hot_i[83];
  assign data_masked[10695] = data_i[10695] & sel_one_hot_i[83];
  assign data_masked[10694] = data_i[10694] & sel_one_hot_i[83];
  assign data_masked[10693] = data_i[10693] & sel_one_hot_i[83];
  assign data_masked[10692] = data_i[10692] & sel_one_hot_i[83];
  assign data_masked[10691] = data_i[10691] & sel_one_hot_i[83];
  assign data_masked[10690] = data_i[10690] & sel_one_hot_i[83];
  assign data_masked[10689] = data_i[10689] & sel_one_hot_i[83];
  assign data_masked[10688] = data_i[10688] & sel_one_hot_i[83];
  assign data_masked[10687] = data_i[10687] & sel_one_hot_i[83];
  assign data_masked[10686] = data_i[10686] & sel_one_hot_i[83];
  assign data_masked[10685] = data_i[10685] & sel_one_hot_i[83];
  assign data_masked[10684] = data_i[10684] & sel_one_hot_i[83];
  assign data_masked[10683] = data_i[10683] & sel_one_hot_i[83];
  assign data_masked[10682] = data_i[10682] & sel_one_hot_i[83];
  assign data_masked[10681] = data_i[10681] & sel_one_hot_i[83];
  assign data_masked[10680] = data_i[10680] & sel_one_hot_i[83];
  assign data_masked[10679] = data_i[10679] & sel_one_hot_i[83];
  assign data_masked[10678] = data_i[10678] & sel_one_hot_i[83];
  assign data_masked[10677] = data_i[10677] & sel_one_hot_i[83];
  assign data_masked[10676] = data_i[10676] & sel_one_hot_i[83];
  assign data_masked[10675] = data_i[10675] & sel_one_hot_i[83];
  assign data_masked[10674] = data_i[10674] & sel_one_hot_i[83];
  assign data_masked[10673] = data_i[10673] & sel_one_hot_i[83];
  assign data_masked[10672] = data_i[10672] & sel_one_hot_i[83];
  assign data_masked[10671] = data_i[10671] & sel_one_hot_i[83];
  assign data_masked[10670] = data_i[10670] & sel_one_hot_i[83];
  assign data_masked[10669] = data_i[10669] & sel_one_hot_i[83];
  assign data_masked[10668] = data_i[10668] & sel_one_hot_i[83];
  assign data_masked[10667] = data_i[10667] & sel_one_hot_i[83];
  assign data_masked[10666] = data_i[10666] & sel_one_hot_i[83];
  assign data_masked[10665] = data_i[10665] & sel_one_hot_i[83];
  assign data_masked[10664] = data_i[10664] & sel_one_hot_i[83];
  assign data_masked[10663] = data_i[10663] & sel_one_hot_i[83];
  assign data_masked[10662] = data_i[10662] & sel_one_hot_i[83];
  assign data_masked[10661] = data_i[10661] & sel_one_hot_i[83];
  assign data_masked[10660] = data_i[10660] & sel_one_hot_i[83];
  assign data_masked[10659] = data_i[10659] & sel_one_hot_i[83];
  assign data_masked[10658] = data_i[10658] & sel_one_hot_i[83];
  assign data_masked[10657] = data_i[10657] & sel_one_hot_i[83];
  assign data_masked[10656] = data_i[10656] & sel_one_hot_i[83];
  assign data_masked[10655] = data_i[10655] & sel_one_hot_i[83];
  assign data_masked[10654] = data_i[10654] & sel_one_hot_i[83];
  assign data_masked[10653] = data_i[10653] & sel_one_hot_i[83];
  assign data_masked[10652] = data_i[10652] & sel_one_hot_i[83];
  assign data_masked[10651] = data_i[10651] & sel_one_hot_i[83];
  assign data_masked[10650] = data_i[10650] & sel_one_hot_i[83];
  assign data_masked[10649] = data_i[10649] & sel_one_hot_i[83];
  assign data_masked[10648] = data_i[10648] & sel_one_hot_i[83];
  assign data_masked[10647] = data_i[10647] & sel_one_hot_i[83];
  assign data_masked[10646] = data_i[10646] & sel_one_hot_i[83];
  assign data_masked[10645] = data_i[10645] & sel_one_hot_i[83];
  assign data_masked[10644] = data_i[10644] & sel_one_hot_i[83];
  assign data_masked[10643] = data_i[10643] & sel_one_hot_i[83];
  assign data_masked[10642] = data_i[10642] & sel_one_hot_i[83];
  assign data_masked[10641] = data_i[10641] & sel_one_hot_i[83];
  assign data_masked[10640] = data_i[10640] & sel_one_hot_i[83];
  assign data_masked[10639] = data_i[10639] & sel_one_hot_i[83];
  assign data_masked[10638] = data_i[10638] & sel_one_hot_i[83];
  assign data_masked[10637] = data_i[10637] & sel_one_hot_i[83];
  assign data_masked[10636] = data_i[10636] & sel_one_hot_i[83];
  assign data_masked[10635] = data_i[10635] & sel_one_hot_i[83];
  assign data_masked[10634] = data_i[10634] & sel_one_hot_i[83];
  assign data_masked[10633] = data_i[10633] & sel_one_hot_i[83];
  assign data_masked[10632] = data_i[10632] & sel_one_hot_i[83];
  assign data_masked[10631] = data_i[10631] & sel_one_hot_i[83];
  assign data_masked[10630] = data_i[10630] & sel_one_hot_i[83];
  assign data_masked[10629] = data_i[10629] & sel_one_hot_i[83];
  assign data_masked[10628] = data_i[10628] & sel_one_hot_i[83];
  assign data_masked[10627] = data_i[10627] & sel_one_hot_i[83];
  assign data_masked[10626] = data_i[10626] & sel_one_hot_i[83];
  assign data_masked[10625] = data_i[10625] & sel_one_hot_i[83];
  assign data_masked[10624] = data_i[10624] & sel_one_hot_i[83];
  assign data_masked[10879] = data_i[10879] & sel_one_hot_i[84];
  assign data_masked[10878] = data_i[10878] & sel_one_hot_i[84];
  assign data_masked[10877] = data_i[10877] & sel_one_hot_i[84];
  assign data_masked[10876] = data_i[10876] & sel_one_hot_i[84];
  assign data_masked[10875] = data_i[10875] & sel_one_hot_i[84];
  assign data_masked[10874] = data_i[10874] & sel_one_hot_i[84];
  assign data_masked[10873] = data_i[10873] & sel_one_hot_i[84];
  assign data_masked[10872] = data_i[10872] & sel_one_hot_i[84];
  assign data_masked[10871] = data_i[10871] & sel_one_hot_i[84];
  assign data_masked[10870] = data_i[10870] & sel_one_hot_i[84];
  assign data_masked[10869] = data_i[10869] & sel_one_hot_i[84];
  assign data_masked[10868] = data_i[10868] & sel_one_hot_i[84];
  assign data_masked[10867] = data_i[10867] & sel_one_hot_i[84];
  assign data_masked[10866] = data_i[10866] & sel_one_hot_i[84];
  assign data_masked[10865] = data_i[10865] & sel_one_hot_i[84];
  assign data_masked[10864] = data_i[10864] & sel_one_hot_i[84];
  assign data_masked[10863] = data_i[10863] & sel_one_hot_i[84];
  assign data_masked[10862] = data_i[10862] & sel_one_hot_i[84];
  assign data_masked[10861] = data_i[10861] & sel_one_hot_i[84];
  assign data_masked[10860] = data_i[10860] & sel_one_hot_i[84];
  assign data_masked[10859] = data_i[10859] & sel_one_hot_i[84];
  assign data_masked[10858] = data_i[10858] & sel_one_hot_i[84];
  assign data_masked[10857] = data_i[10857] & sel_one_hot_i[84];
  assign data_masked[10856] = data_i[10856] & sel_one_hot_i[84];
  assign data_masked[10855] = data_i[10855] & sel_one_hot_i[84];
  assign data_masked[10854] = data_i[10854] & sel_one_hot_i[84];
  assign data_masked[10853] = data_i[10853] & sel_one_hot_i[84];
  assign data_masked[10852] = data_i[10852] & sel_one_hot_i[84];
  assign data_masked[10851] = data_i[10851] & sel_one_hot_i[84];
  assign data_masked[10850] = data_i[10850] & sel_one_hot_i[84];
  assign data_masked[10849] = data_i[10849] & sel_one_hot_i[84];
  assign data_masked[10848] = data_i[10848] & sel_one_hot_i[84];
  assign data_masked[10847] = data_i[10847] & sel_one_hot_i[84];
  assign data_masked[10846] = data_i[10846] & sel_one_hot_i[84];
  assign data_masked[10845] = data_i[10845] & sel_one_hot_i[84];
  assign data_masked[10844] = data_i[10844] & sel_one_hot_i[84];
  assign data_masked[10843] = data_i[10843] & sel_one_hot_i[84];
  assign data_masked[10842] = data_i[10842] & sel_one_hot_i[84];
  assign data_masked[10841] = data_i[10841] & sel_one_hot_i[84];
  assign data_masked[10840] = data_i[10840] & sel_one_hot_i[84];
  assign data_masked[10839] = data_i[10839] & sel_one_hot_i[84];
  assign data_masked[10838] = data_i[10838] & sel_one_hot_i[84];
  assign data_masked[10837] = data_i[10837] & sel_one_hot_i[84];
  assign data_masked[10836] = data_i[10836] & sel_one_hot_i[84];
  assign data_masked[10835] = data_i[10835] & sel_one_hot_i[84];
  assign data_masked[10834] = data_i[10834] & sel_one_hot_i[84];
  assign data_masked[10833] = data_i[10833] & sel_one_hot_i[84];
  assign data_masked[10832] = data_i[10832] & sel_one_hot_i[84];
  assign data_masked[10831] = data_i[10831] & sel_one_hot_i[84];
  assign data_masked[10830] = data_i[10830] & sel_one_hot_i[84];
  assign data_masked[10829] = data_i[10829] & sel_one_hot_i[84];
  assign data_masked[10828] = data_i[10828] & sel_one_hot_i[84];
  assign data_masked[10827] = data_i[10827] & sel_one_hot_i[84];
  assign data_masked[10826] = data_i[10826] & sel_one_hot_i[84];
  assign data_masked[10825] = data_i[10825] & sel_one_hot_i[84];
  assign data_masked[10824] = data_i[10824] & sel_one_hot_i[84];
  assign data_masked[10823] = data_i[10823] & sel_one_hot_i[84];
  assign data_masked[10822] = data_i[10822] & sel_one_hot_i[84];
  assign data_masked[10821] = data_i[10821] & sel_one_hot_i[84];
  assign data_masked[10820] = data_i[10820] & sel_one_hot_i[84];
  assign data_masked[10819] = data_i[10819] & sel_one_hot_i[84];
  assign data_masked[10818] = data_i[10818] & sel_one_hot_i[84];
  assign data_masked[10817] = data_i[10817] & sel_one_hot_i[84];
  assign data_masked[10816] = data_i[10816] & sel_one_hot_i[84];
  assign data_masked[10815] = data_i[10815] & sel_one_hot_i[84];
  assign data_masked[10814] = data_i[10814] & sel_one_hot_i[84];
  assign data_masked[10813] = data_i[10813] & sel_one_hot_i[84];
  assign data_masked[10812] = data_i[10812] & sel_one_hot_i[84];
  assign data_masked[10811] = data_i[10811] & sel_one_hot_i[84];
  assign data_masked[10810] = data_i[10810] & sel_one_hot_i[84];
  assign data_masked[10809] = data_i[10809] & sel_one_hot_i[84];
  assign data_masked[10808] = data_i[10808] & sel_one_hot_i[84];
  assign data_masked[10807] = data_i[10807] & sel_one_hot_i[84];
  assign data_masked[10806] = data_i[10806] & sel_one_hot_i[84];
  assign data_masked[10805] = data_i[10805] & sel_one_hot_i[84];
  assign data_masked[10804] = data_i[10804] & sel_one_hot_i[84];
  assign data_masked[10803] = data_i[10803] & sel_one_hot_i[84];
  assign data_masked[10802] = data_i[10802] & sel_one_hot_i[84];
  assign data_masked[10801] = data_i[10801] & sel_one_hot_i[84];
  assign data_masked[10800] = data_i[10800] & sel_one_hot_i[84];
  assign data_masked[10799] = data_i[10799] & sel_one_hot_i[84];
  assign data_masked[10798] = data_i[10798] & sel_one_hot_i[84];
  assign data_masked[10797] = data_i[10797] & sel_one_hot_i[84];
  assign data_masked[10796] = data_i[10796] & sel_one_hot_i[84];
  assign data_masked[10795] = data_i[10795] & sel_one_hot_i[84];
  assign data_masked[10794] = data_i[10794] & sel_one_hot_i[84];
  assign data_masked[10793] = data_i[10793] & sel_one_hot_i[84];
  assign data_masked[10792] = data_i[10792] & sel_one_hot_i[84];
  assign data_masked[10791] = data_i[10791] & sel_one_hot_i[84];
  assign data_masked[10790] = data_i[10790] & sel_one_hot_i[84];
  assign data_masked[10789] = data_i[10789] & sel_one_hot_i[84];
  assign data_masked[10788] = data_i[10788] & sel_one_hot_i[84];
  assign data_masked[10787] = data_i[10787] & sel_one_hot_i[84];
  assign data_masked[10786] = data_i[10786] & sel_one_hot_i[84];
  assign data_masked[10785] = data_i[10785] & sel_one_hot_i[84];
  assign data_masked[10784] = data_i[10784] & sel_one_hot_i[84];
  assign data_masked[10783] = data_i[10783] & sel_one_hot_i[84];
  assign data_masked[10782] = data_i[10782] & sel_one_hot_i[84];
  assign data_masked[10781] = data_i[10781] & sel_one_hot_i[84];
  assign data_masked[10780] = data_i[10780] & sel_one_hot_i[84];
  assign data_masked[10779] = data_i[10779] & sel_one_hot_i[84];
  assign data_masked[10778] = data_i[10778] & sel_one_hot_i[84];
  assign data_masked[10777] = data_i[10777] & sel_one_hot_i[84];
  assign data_masked[10776] = data_i[10776] & sel_one_hot_i[84];
  assign data_masked[10775] = data_i[10775] & sel_one_hot_i[84];
  assign data_masked[10774] = data_i[10774] & sel_one_hot_i[84];
  assign data_masked[10773] = data_i[10773] & sel_one_hot_i[84];
  assign data_masked[10772] = data_i[10772] & sel_one_hot_i[84];
  assign data_masked[10771] = data_i[10771] & sel_one_hot_i[84];
  assign data_masked[10770] = data_i[10770] & sel_one_hot_i[84];
  assign data_masked[10769] = data_i[10769] & sel_one_hot_i[84];
  assign data_masked[10768] = data_i[10768] & sel_one_hot_i[84];
  assign data_masked[10767] = data_i[10767] & sel_one_hot_i[84];
  assign data_masked[10766] = data_i[10766] & sel_one_hot_i[84];
  assign data_masked[10765] = data_i[10765] & sel_one_hot_i[84];
  assign data_masked[10764] = data_i[10764] & sel_one_hot_i[84];
  assign data_masked[10763] = data_i[10763] & sel_one_hot_i[84];
  assign data_masked[10762] = data_i[10762] & sel_one_hot_i[84];
  assign data_masked[10761] = data_i[10761] & sel_one_hot_i[84];
  assign data_masked[10760] = data_i[10760] & sel_one_hot_i[84];
  assign data_masked[10759] = data_i[10759] & sel_one_hot_i[84];
  assign data_masked[10758] = data_i[10758] & sel_one_hot_i[84];
  assign data_masked[10757] = data_i[10757] & sel_one_hot_i[84];
  assign data_masked[10756] = data_i[10756] & sel_one_hot_i[84];
  assign data_masked[10755] = data_i[10755] & sel_one_hot_i[84];
  assign data_masked[10754] = data_i[10754] & sel_one_hot_i[84];
  assign data_masked[10753] = data_i[10753] & sel_one_hot_i[84];
  assign data_masked[10752] = data_i[10752] & sel_one_hot_i[84];
  assign data_masked[11007] = data_i[11007] & sel_one_hot_i[85];
  assign data_masked[11006] = data_i[11006] & sel_one_hot_i[85];
  assign data_masked[11005] = data_i[11005] & sel_one_hot_i[85];
  assign data_masked[11004] = data_i[11004] & sel_one_hot_i[85];
  assign data_masked[11003] = data_i[11003] & sel_one_hot_i[85];
  assign data_masked[11002] = data_i[11002] & sel_one_hot_i[85];
  assign data_masked[11001] = data_i[11001] & sel_one_hot_i[85];
  assign data_masked[11000] = data_i[11000] & sel_one_hot_i[85];
  assign data_masked[10999] = data_i[10999] & sel_one_hot_i[85];
  assign data_masked[10998] = data_i[10998] & sel_one_hot_i[85];
  assign data_masked[10997] = data_i[10997] & sel_one_hot_i[85];
  assign data_masked[10996] = data_i[10996] & sel_one_hot_i[85];
  assign data_masked[10995] = data_i[10995] & sel_one_hot_i[85];
  assign data_masked[10994] = data_i[10994] & sel_one_hot_i[85];
  assign data_masked[10993] = data_i[10993] & sel_one_hot_i[85];
  assign data_masked[10992] = data_i[10992] & sel_one_hot_i[85];
  assign data_masked[10991] = data_i[10991] & sel_one_hot_i[85];
  assign data_masked[10990] = data_i[10990] & sel_one_hot_i[85];
  assign data_masked[10989] = data_i[10989] & sel_one_hot_i[85];
  assign data_masked[10988] = data_i[10988] & sel_one_hot_i[85];
  assign data_masked[10987] = data_i[10987] & sel_one_hot_i[85];
  assign data_masked[10986] = data_i[10986] & sel_one_hot_i[85];
  assign data_masked[10985] = data_i[10985] & sel_one_hot_i[85];
  assign data_masked[10984] = data_i[10984] & sel_one_hot_i[85];
  assign data_masked[10983] = data_i[10983] & sel_one_hot_i[85];
  assign data_masked[10982] = data_i[10982] & sel_one_hot_i[85];
  assign data_masked[10981] = data_i[10981] & sel_one_hot_i[85];
  assign data_masked[10980] = data_i[10980] & sel_one_hot_i[85];
  assign data_masked[10979] = data_i[10979] & sel_one_hot_i[85];
  assign data_masked[10978] = data_i[10978] & sel_one_hot_i[85];
  assign data_masked[10977] = data_i[10977] & sel_one_hot_i[85];
  assign data_masked[10976] = data_i[10976] & sel_one_hot_i[85];
  assign data_masked[10975] = data_i[10975] & sel_one_hot_i[85];
  assign data_masked[10974] = data_i[10974] & sel_one_hot_i[85];
  assign data_masked[10973] = data_i[10973] & sel_one_hot_i[85];
  assign data_masked[10972] = data_i[10972] & sel_one_hot_i[85];
  assign data_masked[10971] = data_i[10971] & sel_one_hot_i[85];
  assign data_masked[10970] = data_i[10970] & sel_one_hot_i[85];
  assign data_masked[10969] = data_i[10969] & sel_one_hot_i[85];
  assign data_masked[10968] = data_i[10968] & sel_one_hot_i[85];
  assign data_masked[10967] = data_i[10967] & sel_one_hot_i[85];
  assign data_masked[10966] = data_i[10966] & sel_one_hot_i[85];
  assign data_masked[10965] = data_i[10965] & sel_one_hot_i[85];
  assign data_masked[10964] = data_i[10964] & sel_one_hot_i[85];
  assign data_masked[10963] = data_i[10963] & sel_one_hot_i[85];
  assign data_masked[10962] = data_i[10962] & sel_one_hot_i[85];
  assign data_masked[10961] = data_i[10961] & sel_one_hot_i[85];
  assign data_masked[10960] = data_i[10960] & sel_one_hot_i[85];
  assign data_masked[10959] = data_i[10959] & sel_one_hot_i[85];
  assign data_masked[10958] = data_i[10958] & sel_one_hot_i[85];
  assign data_masked[10957] = data_i[10957] & sel_one_hot_i[85];
  assign data_masked[10956] = data_i[10956] & sel_one_hot_i[85];
  assign data_masked[10955] = data_i[10955] & sel_one_hot_i[85];
  assign data_masked[10954] = data_i[10954] & sel_one_hot_i[85];
  assign data_masked[10953] = data_i[10953] & sel_one_hot_i[85];
  assign data_masked[10952] = data_i[10952] & sel_one_hot_i[85];
  assign data_masked[10951] = data_i[10951] & sel_one_hot_i[85];
  assign data_masked[10950] = data_i[10950] & sel_one_hot_i[85];
  assign data_masked[10949] = data_i[10949] & sel_one_hot_i[85];
  assign data_masked[10948] = data_i[10948] & sel_one_hot_i[85];
  assign data_masked[10947] = data_i[10947] & sel_one_hot_i[85];
  assign data_masked[10946] = data_i[10946] & sel_one_hot_i[85];
  assign data_masked[10945] = data_i[10945] & sel_one_hot_i[85];
  assign data_masked[10944] = data_i[10944] & sel_one_hot_i[85];
  assign data_masked[10943] = data_i[10943] & sel_one_hot_i[85];
  assign data_masked[10942] = data_i[10942] & sel_one_hot_i[85];
  assign data_masked[10941] = data_i[10941] & sel_one_hot_i[85];
  assign data_masked[10940] = data_i[10940] & sel_one_hot_i[85];
  assign data_masked[10939] = data_i[10939] & sel_one_hot_i[85];
  assign data_masked[10938] = data_i[10938] & sel_one_hot_i[85];
  assign data_masked[10937] = data_i[10937] & sel_one_hot_i[85];
  assign data_masked[10936] = data_i[10936] & sel_one_hot_i[85];
  assign data_masked[10935] = data_i[10935] & sel_one_hot_i[85];
  assign data_masked[10934] = data_i[10934] & sel_one_hot_i[85];
  assign data_masked[10933] = data_i[10933] & sel_one_hot_i[85];
  assign data_masked[10932] = data_i[10932] & sel_one_hot_i[85];
  assign data_masked[10931] = data_i[10931] & sel_one_hot_i[85];
  assign data_masked[10930] = data_i[10930] & sel_one_hot_i[85];
  assign data_masked[10929] = data_i[10929] & sel_one_hot_i[85];
  assign data_masked[10928] = data_i[10928] & sel_one_hot_i[85];
  assign data_masked[10927] = data_i[10927] & sel_one_hot_i[85];
  assign data_masked[10926] = data_i[10926] & sel_one_hot_i[85];
  assign data_masked[10925] = data_i[10925] & sel_one_hot_i[85];
  assign data_masked[10924] = data_i[10924] & sel_one_hot_i[85];
  assign data_masked[10923] = data_i[10923] & sel_one_hot_i[85];
  assign data_masked[10922] = data_i[10922] & sel_one_hot_i[85];
  assign data_masked[10921] = data_i[10921] & sel_one_hot_i[85];
  assign data_masked[10920] = data_i[10920] & sel_one_hot_i[85];
  assign data_masked[10919] = data_i[10919] & sel_one_hot_i[85];
  assign data_masked[10918] = data_i[10918] & sel_one_hot_i[85];
  assign data_masked[10917] = data_i[10917] & sel_one_hot_i[85];
  assign data_masked[10916] = data_i[10916] & sel_one_hot_i[85];
  assign data_masked[10915] = data_i[10915] & sel_one_hot_i[85];
  assign data_masked[10914] = data_i[10914] & sel_one_hot_i[85];
  assign data_masked[10913] = data_i[10913] & sel_one_hot_i[85];
  assign data_masked[10912] = data_i[10912] & sel_one_hot_i[85];
  assign data_masked[10911] = data_i[10911] & sel_one_hot_i[85];
  assign data_masked[10910] = data_i[10910] & sel_one_hot_i[85];
  assign data_masked[10909] = data_i[10909] & sel_one_hot_i[85];
  assign data_masked[10908] = data_i[10908] & sel_one_hot_i[85];
  assign data_masked[10907] = data_i[10907] & sel_one_hot_i[85];
  assign data_masked[10906] = data_i[10906] & sel_one_hot_i[85];
  assign data_masked[10905] = data_i[10905] & sel_one_hot_i[85];
  assign data_masked[10904] = data_i[10904] & sel_one_hot_i[85];
  assign data_masked[10903] = data_i[10903] & sel_one_hot_i[85];
  assign data_masked[10902] = data_i[10902] & sel_one_hot_i[85];
  assign data_masked[10901] = data_i[10901] & sel_one_hot_i[85];
  assign data_masked[10900] = data_i[10900] & sel_one_hot_i[85];
  assign data_masked[10899] = data_i[10899] & sel_one_hot_i[85];
  assign data_masked[10898] = data_i[10898] & sel_one_hot_i[85];
  assign data_masked[10897] = data_i[10897] & sel_one_hot_i[85];
  assign data_masked[10896] = data_i[10896] & sel_one_hot_i[85];
  assign data_masked[10895] = data_i[10895] & sel_one_hot_i[85];
  assign data_masked[10894] = data_i[10894] & sel_one_hot_i[85];
  assign data_masked[10893] = data_i[10893] & sel_one_hot_i[85];
  assign data_masked[10892] = data_i[10892] & sel_one_hot_i[85];
  assign data_masked[10891] = data_i[10891] & sel_one_hot_i[85];
  assign data_masked[10890] = data_i[10890] & sel_one_hot_i[85];
  assign data_masked[10889] = data_i[10889] & sel_one_hot_i[85];
  assign data_masked[10888] = data_i[10888] & sel_one_hot_i[85];
  assign data_masked[10887] = data_i[10887] & sel_one_hot_i[85];
  assign data_masked[10886] = data_i[10886] & sel_one_hot_i[85];
  assign data_masked[10885] = data_i[10885] & sel_one_hot_i[85];
  assign data_masked[10884] = data_i[10884] & sel_one_hot_i[85];
  assign data_masked[10883] = data_i[10883] & sel_one_hot_i[85];
  assign data_masked[10882] = data_i[10882] & sel_one_hot_i[85];
  assign data_masked[10881] = data_i[10881] & sel_one_hot_i[85];
  assign data_masked[10880] = data_i[10880] & sel_one_hot_i[85];
  assign data_masked[11135] = data_i[11135] & sel_one_hot_i[86];
  assign data_masked[11134] = data_i[11134] & sel_one_hot_i[86];
  assign data_masked[11133] = data_i[11133] & sel_one_hot_i[86];
  assign data_masked[11132] = data_i[11132] & sel_one_hot_i[86];
  assign data_masked[11131] = data_i[11131] & sel_one_hot_i[86];
  assign data_masked[11130] = data_i[11130] & sel_one_hot_i[86];
  assign data_masked[11129] = data_i[11129] & sel_one_hot_i[86];
  assign data_masked[11128] = data_i[11128] & sel_one_hot_i[86];
  assign data_masked[11127] = data_i[11127] & sel_one_hot_i[86];
  assign data_masked[11126] = data_i[11126] & sel_one_hot_i[86];
  assign data_masked[11125] = data_i[11125] & sel_one_hot_i[86];
  assign data_masked[11124] = data_i[11124] & sel_one_hot_i[86];
  assign data_masked[11123] = data_i[11123] & sel_one_hot_i[86];
  assign data_masked[11122] = data_i[11122] & sel_one_hot_i[86];
  assign data_masked[11121] = data_i[11121] & sel_one_hot_i[86];
  assign data_masked[11120] = data_i[11120] & sel_one_hot_i[86];
  assign data_masked[11119] = data_i[11119] & sel_one_hot_i[86];
  assign data_masked[11118] = data_i[11118] & sel_one_hot_i[86];
  assign data_masked[11117] = data_i[11117] & sel_one_hot_i[86];
  assign data_masked[11116] = data_i[11116] & sel_one_hot_i[86];
  assign data_masked[11115] = data_i[11115] & sel_one_hot_i[86];
  assign data_masked[11114] = data_i[11114] & sel_one_hot_i[86];
  assign data_masked[11113] = data_i[11113] & sel_one_hot_i[86];
  assign data_masked[11112] = data_i[11112] & sel_one_hot_i[86];
  assign data_masked[11111] = data_i[11111] & sel_one_hot_i[86];
  assign data_masked[11110] = data_i[11110] & sel_one_hot_i[86];
  assign data_masked[11109] = data_i[11109] & sel_one_hot_i[86];
  assign data_masked[11108] = data_i[11108] & sel_one_hot_i[86];
  assign data_masked[11107] = data_i[11107] & sel_one_hot_i[86];
  assign data_masked[11106] = data_i[11106] & sel_one_hot_i[86];
  assign data_masked[11105] = data_i[11105] & sel_one_hot_i[86];
  assign data_masked[11104] = data_i[11104] & sel_one_hot_i[86];
  assign data_masked[11103] = data_i[11103] & sel_one_hot_i[86];
  assign data_masked[11102] = data_i[11102] & sel_one_hot_i[86];
  assign data_masked[11101] = data_i[11101] & sel_one_hot_i[86];
  assign data_masked[11100] = data_i[11100] & sel_one_hot_i[86];
  assign data_masked[11099] = data_i[11099] & sel_one_hot_i[86];
  assign data_masked[11098] = data_i[11098] & sel_one_hot_i[86];
  assign data_masked[11097] = data_i[11097] & sel_one_hot_i[86];
  assign data_masked[11096] = data_i[11096] & sel_one_hot_i[86];
  assign data_masked[11095] = data_i[11095] & sel_one_hot_i[86];
  assign data_masked[11094] = data_i[11094] & sel_one_hot_i[86];
  assign data_masked[11093] = data_i[11093] & sel_one_hot_i[86];
  assign data_masked[11092] = data_i[11092] & sel_one_hot_i[86];
  assign data_masked[11091] = data_i[11091] & sel_one_hot_i[86];
  assign data_masked[11090] = data_i[11090] & sel_one_hot_i[86];
  assign data_masked[11089] = data_i[11089] & sel_one_hot_i[86];
  assign data_masked[11088] = data_i[11088] & sel_one_hot_i[86];
  assign data_masked[11087] = data_i[11087] & sel_one_hot_i[86];
  assign data_masked[11086] = data_i[11086] & sel_one_hot_i[86];
  assign data_masked[11085] = data_i[11085] & sel_one_hot_i[86];
  assign data_masked[11084] = data_i[11084] & sel_one_hot_i[86];
  assign data_masked[11083] = data_i[11083] & sel_one_hot_i[86];
  assign data_masked[11082] = data_i[11082] & sel_one_hot_i[86];
  assign data_masked[11081] = data_i[11081] & sel_one_hot_i[86];
  assign data_masked[11080] = data_i[11080] & sel_one_hot_i[86];
  assign data_masked[11079] = data_i[11079] & sel_one_hot_i[86];
  assign data_masked[11078] = data_i[11078] & sel_one_hot_i[86];
  assign data_masked[11077] = data_i[11077] & sel_one_hot_i[86];
  assign data_masked[11076] = data_i[11076] & sel_one_hot_i[86];
  assign data_masked[11075] = data_i[11075] & sel_one_hot_i[86];
  assign data_masked[11074] = data_i[11074] & sel_one_hot_i[86];
  assign data_masked[11073] = data_i[11073] & sel_one_hot_i[86];
  assign data_masked[11072] = data_i[11072] & sel_one_hot_i[86];
  assign data_masked[11071] = data_i[11071] & sel_one_hot_i[86];
  assign data_masked[11070] = data_i[11070] & sel_one_hot_i[86];
  assign data_masked[11069] = data_i[11069] & sel_one_hot_i[86];
  assign data_masked[11068] = data_i[11068] & sel_one_hot_i[86];
  assign data_masked[11067] = data_i[11067] & sel_one_hot_i[86];
  assign data_masked[11066] = data_i[11066] & sel_one_hot_i[86];
  assign data_masked[11065] = data_i[11065] & sel_one_hot_i[86];
  assign data_masked[11064] = data_i[11064] & sel_one_hot_i[86];
  assign data_masked[11063] = data_i[11063] & sel_one_hot_i[86];
  assign data_masked[11062] = data_i[11062] & sel_one_hot_i[86];
  assign data_masked[11061] = data_i[11061] & sel_one_hot_i[86];
  assign data_masked[11060] = data_i[11060] & sel_one_hot_i[86];
  assign data_masked[11059] = data_i[11059] & sel_one_hot_i[86];
  assign data_masked[11058] = data_i[11058] & sel_one_hot_i[86];
  assign data_masked[11057] = data_i[11057] & sel_one_hot_i[86];
  assign data_masked[11056] = data_i[11056] & sel_one_hot_i[86];
  assign data_masked[11055] = data_i[11055] & sel_one_hot_i[86];
  assign data_masked[11054] = data_i[11054] & sel_one_hot_i[86];
  assign data_masked[11053] = data_i[11053] & sel_one_hot_i[86];
  assign data_masked[11052] = data_i[11052] & sel_one_hot_i[86];
  assign data_masked[11051] = data_i[11051] & sel_one_hot_i[86];
  assign data_masked[11050] = data_i[11050] & sel_one_hot_i[86];
  assign data_masked[11049] = data_i[11049] & sel_one_hot_i[86];
  assign data_masked[11048] = data_i[11048] & sel_one_hot_i[86];
  assign data_masked[11047] = data_i[11047] & sel_one_hot_i[86];
  assign data_masked[11046] = data_i[11046] & sel_one_hot_i[86];
  assign data_masked[11045] = data_i[11045] & sel_one_hot_i[86];
  assign data_masked[11044] = data_i[11044] & sel_one_hot_i[86];
  assign data_masked[11043] = data_i[11043] & sel_one_hot_i[86];
  assign data_masked[11042] = data_i[11042] & sel_one_hot_i[86];
  assign data_masked[11041] = data_i[11041] & sel_one_hot_i[86];
  assign data_masked[11040] = data_i[11040] & sel_one_hot_i[86];
  assign data_masked[11039] = data_i[11039] & sel_one_hot_i[86];
  assign data_masked[11038] = data_i[11038] & sel_one_hot_i[86];
  assign data_masked[11037] = data_i[11037] & sel_one_hot_i[86];
  assign data_masked[11036] = data_i[11036] & sel_one_hot_i[86];
  assign data_masked[11035] = data_i[11035] & sel_one_hot_i[86];
  assign data_masked[11034] = data_i[11034] & sel_one_hot_i[86];
  assign data_masked[11033] = data_i[11033] & sel_one_hot_i[86];
  assign data_masked[11032] = data_i[11032] & sel_one_hot_i[86];
  assign data_masked[11031] = data_i[11031] & sel_one_hot_i[86];
  assign data_masked[11030] = data_i[11030] & sel_one_hot_i[86];
  assign data_masked[11029] = data_i[11029] & sel_one_hot_i[86];
  assign data_masked[11028] = data_i[11028] & sel_one_hot_i[86];
  assign data_masked[11027] = data_i[11027] & sel_one_hot_i[86];
  assign data_masked[11026] = data_i[11026] & sel_one_hot_i[86];
  assign data_masked[11025] = data_i[11025] & sel_one_hot_i[86];
  assign data_masked[11024] = data_i[11024] & sel_one_hot_i[86];
  assign data_masked[11023] = data_i[11023] & sel_one_hot_i[86];
  assign data_masked[11022] = data_i[11022] & sel_one_hot_i[86];
  assign data_masked[11021] = data_i[11021] & sel_one_hot_i[86];
  assign data_masked[11020] = data_i[11020] & sel_one_hot_i[86];
  assign data_masked[11019] = data_i[11019] & sel_one_hot_i[86];
  assign data_masked[11018] = data_i[11018] & sel_one_hot_i[86];
  assign data_masked[11017] = data_i[11017] & sel_one_hot_i[86];
  assign data_masked[11016] = data_i[11016] & sel_one_hot_i[86];
  assign data_masked[11015] = data_i[11015] & sel_one_hot_i[86];
  assign data_masked[11014] = data_i[11014] & sel_one_hot_i[86];
  assign data_masked[11013] = data_i[11013] & sel_one_hot_i[86];
  assign data_masked[11012] = data_i[11012] & sel_one_hot_i[86];
  assign data_masked[11011] = data_i[11011] & sel_one_hot_i[86];
  assign data_masked[11010] = data_i[11010] & sel_one_hot_i[86];
  assign data_masked[11009] = data_i[11009] & sel_one_hot_i[86];
  assign data_masked[11008] = data_i[11008] & sel_one_hot_i[86];
  assign data_masked[11263] = data_i[11263] & sel_one_hot_i[87];
  assign data_masked[11262] = data_i[11262] & sel_one_hot_i[87];
  assign data_masked[11261] = data_i[11261] & sel_one_hot_i[87];
  assign data_masked[11260] = data_i[11260] & sel_one_hot_i[87];
  assign data_masked[11259] = data_i[11259] & sel_one_hot_i[87];
  assign data_masked[11258] = data_i[11258] & sel_one_hot_i[87];
  assign data_masked[11257] = data_i[11257] & sel_one_hot_i[87];
  assign data_masked[11256] = data_i[11256] & sel_one_hot_i[87];
  assign data_masked[11255] = data_i[11255] & sel_one_hot_i[87];
  assign data_masked[11254] = data_i[11254] & sel_one_hot_i[87];
  assign data_masked[11253] = data_i[11253] & sel_one_hot_i[87];
  assign data_masked[11252] = data_i[11252] & sel_one_hot_i[87];
  assign data_masked[11251] = data_i[11251] & sel_one_hot_i[87];
  assign data_masked[11250] = data_i[11250] & sel_one_hot_i[87];
  assign data_masked[11249] = data_i[11249] & sel_one_hot_i[87];
  assign data_masked[11248] = data_i[11248] & sel_one_hot_i[87];
  assign data_masked[11247] = data_i[11247] & sel_one_hot_i[87];
  assign data_masked[11246] = data_i[11246] & sel_one_hot_i[87];
  assign data_masked[11245] = data_i[11245] & sel_one_hot_i[87];
  assign data_masked[11244] = data_i[11244] & sel_one_hot_i[87];
  assign data_masked[11243] = data_i[11243] & sel_one_hot_i[87];
  assign data_masked[11242] = data_i[11242] & sel_one_hot_i[87];
  assign data_masked[11241] = data_i[11241] & sel_one_hot_i[87];
  assign data_masked[11240] = data_i[11240] & sel_one_hot_i[87];
  assign data_masked[11239] = data_i[11239] & sel_one_hot_i[87];
  assign data_masked[11238] = data_i[11238] & sel_one_hot_i[87];
  assign data_masked[11237] = data_i[11237] & sel_one_hot_i[87];
  assign data_masked[11236] = data_i[11236] & sel_one_hot_i[87];
  assign data_masked[11235] = data_i[11235] & sel_one_hot_i[87];
  assign data_masked[11234] = data_i[11234] & sel_one_hot_i[87];
  assign data_masked[11233] = data_i[11233] & sel_one_hot_i[87];
  assign data_masked[11232] = data_i[11232] & sel_one_hot_i[87];
  assign data_masked[11231] = data_i[11231] & sel_one_hot_i[87];
  assign data_masked[11230] = data_i[11230] & sel_one_hot_i[87];
  assign data_masked[11229] = data_i[11229] & sel_one_hot_i[87];
  assign data_masked[11228] = data_i[11228] & sel_one_hot_i[87];
  assign data_masked[11227] = data_i[11227] & sel_one_hot_i[87];
  assign data_masked[11226] = data_i[11226] & sel_one_hot_i[87];
  assign data_masked[11225] = data_i[11225] & sel_one_hot_i[87];
  assign data_masked[11224] = data_i[11224] & sel_one_hot_i[87];
  assign data_masked[11223] = data_i[11223] & sel_one_hot_i[87];
  assign data_masked[11222] = data_i[11222] & sel_one_hot_i[87];
  assign data_masked[11221] = data_i[11221] & sel_one_hot_i[87];
  assign data_masked[11220] = data_i[11220] & sel_one_hot_i[87];
  assign data_masked[11219] = data_i[11219] & sel_one_hot_i[87];
  assign data_masked[11218] = data_i[11218] & sel_one_hot_i[87];
  assign data_masked[11217] = data_i[11217] & sel_one_hot_i[87];
  assign data_masked[11216] = data_i[11216] & sel_one_hot_i[87];
  assign data_masked[11215] = data_i[11215] & sel_one_hot_i[87];
  assign data_masked[11214] = data_i[11214] & sel_one_hot_i[87];
  assign data_masked[11213] = data_i[11213] & sel_one_hot_i[87];
  assign data_masked[11212] = data_i[11212] & sel_one_hot_i[87];
  assign data_masked[11211] = data_i[11211] & sel_one_hot_i[87];
  assign data_masked[11210] = data_i[11210] & sel_one_hot_i[87];
  assign data_masked[11209] = data_i[11209] & sel_one_hot_i[87];
  assign data_masked[11208] = data_i[11208] & sel_one_hot_i[87];
  assign data_masked[11207] = data_i[11207] & sel_one_hot_i[87];
  assign data_masked[11206] = data_i[11206] & sel_one_hot_i[87];
  assign data_masked[11205] = data_i[11205] & sel_one_hot_i[87];
  assign data_masked[11204] = data_i[11204] & sel_one_hot_i[87];
  assign data_masked[11203] = data_i[11203] & sel_one_hot_i[87];
  assign data_masked[11202] = data_i[11202] & sel_one_hot_i[87];
  assign data_masked[11201] = data_i[11201] & sel_one_hot_i[87];
  assign data_masked[11200] = data_i[11200] & sel_one_hot_i[87];
  assign data_masked[11199] = data_i[11199] & sel_one_hot_i[87];
  assign data_masked[11198] = data_i[11198] & sel_one_hot_i[87];
  assign data_masked[11197] = data_i[11197] & sel_one_hot_i[87];
  assign data_masked[11196] = data_i[11196] & sel_one_hot_i[87];
  assign data_masked[11195] = data_i[11195] & sel_one_hot_i[87];
  assign data_masked[11194] = data_i[11194] & sel_one_hot_i[87];
  assign data_masked[11193] = data_i[11193] & sel_one_hot_i[87];
  assign data_masked[11192] = data_i[11192] & sel_one_hot_i[87];
  assign data_masked[11191] = data_i[11191] & sel_one_hot_i[87];
  assign data_masked[11190] = data_i[11190] & sel_one_hot_i[87];
  assign data_masked[11189] = data_i[11189] & sel_one_hot_i[87];
  assign data_masked[11188] = data_i[11188] & sel_one_hot_i[87];
  assign data_masked[11187] = data_i[11187] & sel_one_hot_i[87];
  assign data_masked[11186] = data_i[11186] & sel_one_hot_i[87];
  assign data_masked[11185] = data_i[11185] & sel_one_hot_i[87];
  assign data_masked[11184] = data_i[11184] & sel_one_hot_i[87];
  assign data_masked[11183] = data_i[11183] & sel_one_hot_i[87];
  assign data_masked[11182] = data_i[11182] & sel_one_hot_i[87];
  assign data_masked[11181] = data_i[11181] & sel_one_hot_i[87];
  assign data_masked[11180] = data_i[11180] & sel_one_hot_i[87];
  assign data_masked[11179] = data_i[11179] & sel_one_hot_i[87];
  assign data_masked[11178] = data_i[11178] & sel_one_hot_i[87];
  assign data_masked[11177] = data_i[11177] & sel_one_hot_i[87];
  assign data_masked[11176] = data_i[11176] & sel_one_hot_i[87];
  assign data_masked[11175] = data_i[11175] & sel_one_hot_i[87];
  assign data_masked[11174] = data_i[11174] & sel_one_hot_i[87];
  assign data_masked[11173] = data_i[11173] & sel_one_hot_i[87];
  assign data_masked[11172] = data_i[11172] & sel_one_hot_i[87];
  assign data_masked[11171] = data_i[11171] & sel_one_hot_i[87];
  assign data_masked[11170] = data_i[11170] & sel_one_hot_i[87];
  assign data_masked[11169] = data_i[11169] & sel_one_hot_i[87];
  assign data_masked[11168] = data_i[11168] & sel_one_hot_i[87];
  assign data_masked[11167] = data_i[11167] & sel_one_hot_i[87];
  assign data_masked[11166] = data_i[11166] & sel_one_hot_i[87];
  assign data_masked[11165] = data_i[11165] & sel_one_hot_i[87];
  assign data_masked[11164] = data_i[11164] & sel_one_hot_i[87];
  assign data_masked[11163] = data_i[11163] & sel_one_hot_i[87];
  assign data_masked[11162] = data_i[11162] & sel_one_hot_i[87];
  assign data_masked[11161] = data_i[11161] & sel_one_hot_i[87];
  assign data_masked[11160] = data_i[11160] & sel_one_hot_i[87];
  assign data_masked[11159] = data_i[11159] & sel_one_hot_i[87];
  assign data_masked[11158] = data_i[11158] & sel_one_hot_i[87];
  assign data_masked[11157] = data_i[11157] & sel_one_hot_i[87];
  assign data_masked[11156] = data_i[11156] & sel_one_hot_i[87];
  assign data_masked[11155] = data_i[11155] & sel_one_hot_i[87];
  assign data_masked[11154] = data_i[11154] & sel_one_hot_i[87];
  assign data_masked[11153] = data_i[11153] & sel_one_hot_i[87];
  assign data_masked[11152] = data_i[11152] & sel_one_hot_i[87];
  assign data_masked[11151] = data_i[11151] & sel_one_hot_i[87];
  assign data_masked[11150] = data_i[11150] & sel_one_hot_i[87];
  assign data_masked[11149] = data_i[11149] & sel_one_hot_i[87];
  assign data_masked[11148] = data_i[11148] & sel_one_hot_i[87];
  assign data_masked[11147] = data_i[11147] & sel_one_hot_i[87];
  assign data_masked[11146] = data_i[11146] & sel_one_hot_i[87];
  assign data_masked[11145] = data_i[11145] & sel_one_hot_i[87];
  assign data_masked[11144] = data_i[11144] & sel_one_hot_i[87];
  assign data_masked[11143] = data_i[11143] & sel_one_hot_i[87];
  assign data_masked[11142] = data_i[11142] & sel_one_hot_i[87];
  assign data_masked[11141] = data_i[11141] & sel_one_hot_i[87];
  assign data_masked[11140] = data_i[11140] & sel_one_hot_i[87];
  assign data_masked[11139] = data_i[11139] & sel_one_hot_i[87];
  assign data_masked[11138] = data_i[11138] & sel_one_hot_i[87];
  assign data_masked[11137] = data_i[11137] & sel_one_hot_i[87];
  assign data_masked[11136] = data_i[11136] & sel_one_hot_i[87];
  assign data_masked[11391] = data_i[11391] & sel_one_hot_i[88];
  assign data_masked[11390] = data_i[11390] & sel_one_hot_i[88];
  assign data_masked[11389] = data_i[11389] & sel_one_hot_i[88];
  assign data_masked[11388] = data_i[11388] & sel_one_hot_i[88];
  assign data_masked[11387] = data_i[11387] & sel_one_hot_i[88];
  assign data_masked[11386] = data_i[11386] & sel_one_hot_i[88];
  assign data_masked[11385] = data_i[11385] & sel_one_hot_i[88];
  assign data_masked[11384] = data_i[11384] & sel_one_hot_i[88];
  assign data_masked[11383] = data_i[11383] & sel_one_hot_i[88];
  assign data_masked[11382] = data_i[11382] & sel_one_hot_i[88];
  assign data_masked[11381] = data_i[11381] & sel_one_hot_i[88];
  assign data_masked[11380] = data_i[11380] & sel_one_hot_i[88];
  assign data_masked[11379] = data_i[11379] & sel_one_hot_i[88];
  assign data_masked[11378] = data_i[11378] & sel_one_hot_i[88];
  assign data_masked[11377] = data_i[11377] & sel_one_hot_i[88];
  assign data_masked[11376] = data_i[11376] & sel_one_hot_i[88];
  assign data_masked[11375] = data_i[11375] & sel_one_hot_i[88];
  assign data_masked[11374] = data_i[11374] & sel_one_hot_i[88];
  assign data_masked[11373] = data_i[11373] & sel_one_hot_i[88];
  assign data_masked[11372] = data_i[11372] & sel_one_hot_i[88];
  assign data_masked[11371] = data_i[11371] & sel_one_hot_i[88];
  assign data_masked[11370] = data_i[11370] & sel_one_hot_i[88];
  assign data_masked[11369] = data_i[11369] & sel_one_hot_i[88];
  assign data_masked[11368] = data_i[11368] & sel_one_hot_i[88];
  assign data_masked[11367] = data_i[11367] & sel_one_hot_i[88];
  assign data_masked[11366] = data_i[11366] & sel_one_hot_i[88];
  assign data_masked[11365] = data_i[11365] & sel_one_hot_i[88];
  assign data_masked[11364] = data_i[11364] & sel_one_hot_i[88];
  assign data_masked[11363] = data_i[11363] & sel_one_hot_i[88];
  assign data_masked[11362] = data_i[11362] & sel_one_hot_i[88];
  assign data_masked[11361] = data_i[11361] & sel_one_hot_i[88];
  assign data_masked[11360] = data_i[11360] & sel_one_hot_i[88];
  assign data_masked[11359] = data_i[11359] & sel_one_hot_i[88];
  assign data_masked[11358] = data_i[11358] & sel_one_hot_i[88];
  assign data_masked[11357] = data_i[11357] & sel_one_hot_i[88];
  assign data_masked[11356] = data_i[11356] & sel_one_hot_i[88];
  assign data_masked[11355] = data_i[11355] & sel_one_hot_i[88];
  assign data_masked[11354] = data_i[11354] & sel_one_hot_i[88];
  assign data_masked[11353] = data_i[11353] & sel_one_hot_i[88];
  assign data_masked[11352] = data_i[11352] & sel_one_hot_i[88];
  assign data_masked[11351] = data_i[11351] & sel_one_hot_i[88];
  assign data_masked[11350] = data_i[11350] & sel_one_hot_i[88];
  assign data_masked[11349] = data_i[11349] & sel_one_hot_i[88];
  assign data_masked[11348] = data_i[11348] & sel_one_hot_i[88];
  assign data_masked[11347] = data_i[11347] & sel_one_hot_i[88];
  assign data_masked[11346] = data_i[11346] & sel_one_hot_i[88];
  assign data_masked[11345] = data_i[11345] & sel_one_hot_i[88];
  assign data_masked[11344] = data_i[11344] & sel_one_hot_i[88];
  assign data_masked[11343] = data_i[11343] & sel_one_hot_i[88];
  assign data_masked[11342] = data_i[11342] & sel_one_hot_i[88];
  assign data_masked[11341] = data_i[11341] & sel_one_hot_i[88];
  assign data_masked[11340] = data_i[11340] & sel_one_hot_i[88];
  assign data_masked[11339] = data_i[11339] & sel_one_hot_i[88];
  assign data_masked[11338] = data_i[11338] & sel_one_hot_i[88];
  assign data_masked[11337] = data_i[11337] & sel_one_hot_i[88];
  assign data_masked[11336] = data_i[11336] & sel_one_hot_i[88];
  assign data_masked[11335] = data_i[11335] & sel_one_hot_i[88];
  assign data_masked[11334] = data_i[11334] & sel_one_hot_i[88];
  assign data_masked[11333] = data_i[11333] & sel_one_hot_i[88];
  assign data_masked[11332] = data_i[11332] & sel_one_hot_i[88];
  assign data_masked[11331] = data_i[11331] & sel_one_hot_i[88];
  assign data_masked[11330] = data_i[11330] & sel_one_hot_i[88];
  assign data_masked[11329] = data_i[11329] & sel_one_hot_i[88];
  assign data_masked[11328] = data_i[11328] & sel_one_hot_i[88];
  assign data_masked[11327] = data_i[11327] & sel_one_hot_i[88];
  assign data_masked[11326] = data_i[11326] & sel_one_hot_i[88];
  assign data_masked[11325] = data_i[11325] & sel_one_hot_i[88];
  assign data_masked[11324] = data_i[11324] & sel_one_hot_i[88];
  assign data_masked[11323] = data_i[11323] & sel_one_hot_i[88];
  assign data_masked[11322] = data_i[11322] & sel_one_hot_i[88];
  assign data_masked[11321] = data_i[11321] & sel_one_hot_i[88];
  assign data_masked[11320] = data_i[11320] & sel_one_hot_i[88];
  assign data_masked[11319] = data_i[11319] & sel_one_hot_i[88];
  assign data_masked[11318] = data_i[11318] & sel_one_hot_i[88];
  assign data_masked[11317] = data_i[11317] & sel_one_hot_i[88];
  assign data_masked[11316] = data_i[11316] & sel_one_hot_i[88];
  assign data_masked[11315] = data_i[11315] & sel_one_hot_i[88];
  assign data_masked[11314] = data_i[11314] & sel_one_hot_i[88];
  assign data_masked[11313] = data_i[11313] & sel_one_hot_i[88];
  assign data_masked[11312] = data_i[11312] & sel_one_hot_i[88];
  assign data_masked[11311] = data_i[11311] & sel_one_hot_i[88];
  assign data_masked[11310] = data_i[11310] & sel_one_hot_i[88];
  assign data_masked[11309] = data_i[11309] & sel_one_hot_i[88];
  assign data_masked[11308] = data_i[11308] & sel_one_hot_i[88];
  assign data_masked[11307] = data_i[11307] & sel_one_hot_i[88];
  assign data_masked[11306] = data_i[11306] & sel_one_hot_i[88];
  assign data_masked[11305] = data_i[11305] & sel_one_hot_i[88];
  assign data_masked[11304] = data_i[11304] & sel_one_hot_i[88];
  assign data_masked[11303] = data_i[11303] & sel_one_hot_i[88];
  assign data_masked[11302] = data_i[11302] & sel_one_hot_i[88];
  assign data_masked[11301] = data_i[11301] & sel_one_hot_i[88];
  assign data_masked[11300] = data_i[11300] & sel_one_hot_i[88];
  assign data_masked[11299] = data_i[11299] & sel_one_hot_i[88];
  assign data_masked[11298] = data_i[11298] & sel_one_hot_i[88];
  assign data_masked[11297] = data_i[11297] & sel_one_hot_i[88];
  assign data_masked[11296] = data_i[11296] & sel_one_hot_i[88];
  assign data_masked[11295] = data_i[11295] & sel_one_hot_i[88];
  assign data_masked[11294] = data_i[11294] & sel_one_hot_i[88];
  assign data_masked[11293] = data_i[11293] & sel_one_hot_i[88];
  assign data_masked[11292] = data_i[11292] & sel_one_hot_i[88];
  assign data_masked[11291] = data_i[11291] & sel_one_hot_i[88];
  assign data_masked[11290] = data_i[11290] & sel_one_hot_i[88];
  assign data_masked[11289] = data_i[11289] & sel_one_hot_i[88];
  assign data_masked[11288] = data_i[11288] & sel_one_hot_i[88];
  assign data_masked[11287] = data_i[11287] & sel_one_hot_i[88];
  assign data_masked[11286] = data_i[11286] & sel_one_hot_i[88];
  assign data_masked[11285] = data_i[11285] & sel_one_hot_i[88];
  assign data_masked[11284] = data_i[11284] & sel_one_hot_i[88];
  assign data_masked[11283] = data_i[11283] & sel_one_hot_i[88];
  assign data_masked[11282] = data_i[11282] & sel_one_hot_i[88];
  assign data_masked[11281] = data_i[11281] & sel_one_hot_i[88];
  assign data_masked[11280] = data_i[11280] & sel_one_hot_i[88];
  assign data_masked[11279] = data_i[11279] & sel_one_hot_i[88];
  assign data_masked[11278] = data_i[11278] & sel_one_hot_i[88];
  assign data_masked[11277] = data_i[11277] & sel_one_hot_i[88];
  assign data_masked[11276] = data_i[11276] & sel_one_hot_i[88];
  assign data_masked[11275] = data_i[11275] & sel_one_hot_i[88];
  assign data_masked[11274] = data_i[11274] & sel_one_hot_i[88];
  assign data_masked[11273] = data_i[11273] & sel_one_hot_i[88];
  assign data_masked[11272] = data_i[11272] & sel_one_hot_i[88];
  assign data_masked[11271] = data_i[11271] & sel_one_hot_i[88];
  assign data_masked[11270] = data_i[11270] & sel_one_hot_i[88];
  assign data_masked[11269] = data_i[11269] & sel_one_hot_i[88];
  assign data_masked[11268] = data_i[11268] & sel_one_hot_i[88];
  assign data_masked[11267] = data_i[11267] & sel_one_hot_i[88];
  assign data_masked[11266] = data_i[11266] & sel_one_hot_i[88];
  assign data_masked[11265] = data_i[11265] & sel_one_hot_i[88];
  assign data_masked[11264] = data_i[11264] & sel_one_hot_i[88];
  assign data_masked[11519] = data_i[11519] & sel_one_hot_i[89];
  assign data_masked[11518] = data_i[11518] & sel_one_hot_i[89];
  assign data_masked[11517] = data_i[11517] & sel_one_hot_i[89];
  assign data_masked[11516] = data_i[11516] & sel_one_hot_i[89];
  assign data_masked[11515] = data_i[11515] & sel_one_hot_i[89];
  assign data_masked[11514] = data_i[11514] & sel_one_hot_i[89];
  assign data_masked[11513] = data_i[11513] & sel_one_hot_i[89];
  assign data_masked[11512] = data_i[11512] & sel_one_hot_i[89];
  assign data_masked[11511] = data_i[11511] & sel_one_hot_i[89];
  assign data_masked[11510] = data_i[11510] & sel_one_hot_i[89];
  assign data_masked[11509] = data_i[11509] & sel_one_hot_i[89];
  assign data_masked[11508] = data_i[11508] & sel_one_hot_i[89];
  assign data_masked[11507] = data_i[11507] & sel_one_hot_i[89];
  assign data_masked[11506] = data_i[11506] & sel_one_hot_i[89];
  assign data_masked[11505] = data_i[11505] & sel_one_hot_i[89];
  assign data_masked[11504] = data_i[11504] & sel_one_hot_i[89];
  assign data_masked[11503] = data_i[11503] & sel_one_hot_i[89];
  assign data_masked[11502] = data_i[11502] & sel_one_hot_i[89];
  assign data_masked[11501] = data_i[11501] & sel_one_hot_i[89];
  assign data_masked[11500] = data_i[11500] & sel_one_hot_i[89];
  assign data_masked[11499] = data_i[11499] & sel_one_hot_i[89];
  assign data_masked[11498] = data_i[11498] & sel_one_hot_i[89];
  assign data_masked[11497] = data_i[11497] & sel_one_hot_i[89];
  assign data_masked[11496] = data_i[11496] & sel_one_hot_i[89];
  assign data_masked[11495] = data_i[11495] & sel_one_hot_i[89];
  assign data_masked[11494] = data_i[11494] & sel_one_hot_i[89];
  assign data_masked[11493] = data_i[11493] & sel_one_hot_i[89];
  assign data_masked[11492] = data_i[11492] & sel_one_hot_i[89];
  assign data_masked[11491] = data_i[11491] & sel_one_hot_i[89];
  assign data_masked[11490] = data_i[11490] & sel_one_hot_i[89];
  assign data_masked[11489] = data_i[11489] & sel_one_hot_i[89];
  assign data_masked[11488] = data_i[11488] & sel_one_hot_i[89];
  assign data_masked[11487] = data_i[11487] & sel_one_hot_i[89];
  assign data_masked[11486] = data_i[11486] & sel_one_hot_i[89];
  assign data_masked[11485] = data_i[11485] & sel_one_hot_i[89];
  assign data_masked[11484] = data_i[11484] & sel_one_hot_i[89];
  assign data_masked[11483] = data_i[11483] & sel_one_hot_i[89];
  assign data_masked[11482] = data_i[11482] & sel_one_hot_i[89];
  assign data_masked[11481] = data_i[11481] & sel_one_hot_i[89];
  assign data_masked[11480] = data_i[11480] & sel_one_hot_i[89];
  assign data_masked[11479] = data_i[11479] & sel_one_hot_i[89];
  assign data_masked[11478] = data_i[11478] & sel_one_hot_i[89];
  assign data_masked[11477] = data_i[11477] & sel_one_hot_i[89];
  assign data_masked[11476] = data_i[11476] & sel_one_hot_i[89];
  assign data_masked[11475] = data_i[11475] & sel_one_hot_i[89];
  assign data_masked[11474] = data_i[11474] & sel_one_hot_i[89];
  assign data_masked[11473] = data_i[11473] & sel_one_hot_i[89];
  assign data_masked[11472] = data_i[11472] & sel_one_hot_i[89];
  assign data_masked[11471] = data_i[11471] & sel_one_hot_i[89];
  assign data_masked[11470] = data_i[11470] & sel_one_hot_i[89];
  assign data_masked[11469] = data_i[11469] & sel_one_hot_i[89];
  assign data_masked[11468] = data_i[11468] & sel_one_hot_i[89];
  assign data_masked[11467] = data_i[11467] & sel_one_hot_i[89];
  assign data_masked[11466] = data_i[11466] & sel_one_hot_i[89];
  assign data_masked[11465] = data_i[11465] & sel_one_hot_i[89];
  assign data_masked[11464] = data_i[11464] & sel_one_hot_i[89];
  assign data_masked[11463] = data_i[11463] & sel_one_hot_i[89];
  assign data_masked[11462] = data_i[11462] & sel_one_hot_i[89];
  assign data_masked[11461] = data_i[11461] & sel_one_hot_i[89];
  assign data_masked[11460] = data_i[11460] & sel_one_hot_i[89];
  assign data_masked[11459] = data_i[11459] & sel_one_hot_i[89];
  assign data_masked[11458] = data_i[11458] & sel_one_hot_i[89];
  assign data_masked[11457] = data_i[11457] & sel_one_hot_i[89];
  assign data_masked[11456] = data_i[11456] & sel_one_hot_i[89];
  assign data_masked[11455] = data_i[11455] & sel_one_hot_i[89];
  assign data_masked[11454] = data_i[11454] & sel_one_hot_i[89];
  assign data_masked[11453] = data_i[11453] & sel_one_hot_i[89];
  assign data_masked[11452] = data_i[11452] & sel_one_hot_i[89];
  assign data_masked[11451] = data_i[11451] & sel_one_hot_i[89];
  assign data_masked[11450] = data_i[11450] & sel_one_hot_i[89];
  assign data_masked[11449] = data_i[11449] & sel_one_hot_i[89];
  assign data_masked[11448] = data_i[11448] & sel_one_hot_i[89];
  assign data_masked[11447] = data_i[11447] & sel_one_hot_i[89];
  assign data_masked[11446] = data_i[11446] & sel_one_hot_i[89];
  assign data_masked[11445] = data_i[11445] & sel_one_hot_i[89];
  assign data_masked[11444] = data_i[11444] & sel_one_hot_i[89];
  assign data_masked[11443] = data_i[11443] & sel_one_hot_i[89];
  assign data_masked[11442] = data_i[11442] & sel_one_hot_i[89];
  assign data_masked[11441] = data_i[11441] & sel_one_hot_i[89];
  assign data_masked[11440] = data_i[11440] & sel_one_hot_i[89];
  assign data_masked[11439] = data_i[11439] & sel_one_hot_i[89];
  assign data_masked[11438] = data_i[11438] & sel_one_hot_i[89];
  assign data_masked[11437] = data_i[11437] & sel_one_hot_i[89];
  assign data_masked[11436] = data_i[11436] & sel_one_hot_i[89];
  assign data_masked[11435] = data_i[11435] & sel_one_hot_i[89];
  assign data_masked[11434] = data_i[11434] & sel_one_hot_i[89];
  assign data_masked[11433] = data_i[11433] & sel_one_hot_i[89];
  assign data_masked[11432] = data_i[11432] & sel_one_hot_i[89];
  assign data_masked[11431] = data_i[11431] & sel_one_hot_i[89];
  assign data_masked[11430] = data_i[11430] & sel_one_hot_i[89];
  assign data_masked[11429] = data_i[11429] & sel_one_hot_i[89];
  assign data_masked[11428] = data_i[11428] & sel_one_hot_i[89];
  assign data_masked[11427] = data_i[11427] & sel_one_hot_i[89];
  assign data_masked[11426] = data_i[11426] & sel_one_hot_i[89];
  assign data_masked[11425] = data_i[11425] & sel_one_hot_i[89];
  assign data_masked[11424] = data_i[11424] & sel_one_hot_i[89];
  assign data_masked[11423] = data_i[11423] & sel_one_hot_i[89];
  assign data_masked[11422] = data_i[11422] & sel_one_hot_i[89];
  assign data_masked[11421] = data_i[11421] & sel_one_hot_i[89];
  assign data_masked[11420] = data_i[11420] & sel_one_hot_i[89];
  assign data_masked[11419] = data_i[11419] & sel_one_hot_i[89];
  assign data_masked[11418] = data_i[11418] & sel_one_hot_i[89];
  assign data_masked[11417] = data_i[11417] & sel_one_hot_i[89];
  assign data_masked[11416] = data_i[11416] & sel_one_hot_i[89];
  assign data_masked[11415] = data_i[11415] & sel_one_hot_i[89];
  assign data_masked[11414] = data_i[11414] & sel_one_hot_i[89];
  assign data_masked[11413] = data_i[11413] & sel_one_hot_i[89];
  assign data_masked[11412] = data_i[11412] & sel_one_hot_i[89];
  assign data_masked[11411] = data_i[11411] & sel_one_hot_i[89];
  assign data_masked[11410] = data_i[11410] & sel_one_hot_i[89];
  assign data_masked[11409] = data_i[11409] & sel_one_hot_i[89];
  assign data_masked[11408] = data_i[11408] & sel_one_hot_i[89];
  assign data_masked[11407] = data_i[11407] & sel_one_hot_i[89];
  assign data_masked[11406] = data_i[11406] & sel_one_hot_i[89];
  assign data_masked[11405] = data_i[11405] & sel_one_hot_i[89];
  assign data_masked[11404] = data_i[11404] & sel_one_hot_i[89];
  assign data_masked[11403] = data_i[11403] & sel_one_hot_i[89];
  assign data_masked[11402] = data_i[11402] & sel_one_hot_i[89];
  assign data_masked[11401] = data_i[11401] & sel_one_hot_i[89];
  assign data_masked[11400] = data_i[11400] & sel_one_hot_i[89];
  assign data_masked[11399] = data_i[11399] & sel_one_hot_i[89];
  assign data_masked[11398] = data_i[11398] & sel_one_hot_i[89];
  assign data_masked[11397] = data_i[11397] & sel_one_hot_i[89];
  assign data_masked[11396] = data_i[11396] & sel_one_hot_i[89];
  assign data_masked[11395] = data_i[11395] & sel_one_hot_i[89];
  assign data_masked[11394] = data_i[11394] & sel_one_hot_i[89];
  assign data_masked[11393] = data_i[11393] & sel_one_hot_i[89];
  assign data_masked[11392] = data_i[11392] & sel_one_hot_i[89];
  assign data_masked[11647] = data_i[11647] & sel_one_hot_i[90];
  assign data_masked[11646] = data_i[11646] & sel_one_hot_i[90];
  assign data_masked[11645] = data_i[11645] & sel_one_hot_i[90];
  assign data_masked[11644] = data_i[11644] & sel_one_hot_i[90];
  assign data_masked[11643] = data_i[11643] & sel_one_hot_i[90];
  assign data_masked[11642] = data_i[11642] & sel_one_hot_i[90];
  assign data_masked[11641] = data_i[11641] & sel_one_hot_i[90];
  assign data_masked[11640] = data_i[11640] & sel_one_hot_i[90];
  assign data_masked[11639] = data_i[11639] & sel_one_hot_i[90];
  assign data_masked[11638] = data_i[11638] & sel_one_hot_i[90];
  assign data_masked[11637] = data_i[11637] & sel_one_hot_i[90];
  assign data_masked[11636] = data_i[11636] & sel_one_hot_i[90];
  assign data_masked[11635] = data_i[11635] & sel_one_hot_i[90];
  assign data_masked[11634] = data_i[11634] & sel_one_hot_i[90];
  assign data_masked[11633] = data_i[11633] & sel_one_hot_i[90];
  assign data_masked[11632] = data_i[11632] & sel_one_hot_i[90];
  assign data_masked[11631] = data_i[11631] & sel_one_hot_i[90];
  assign data_masked[11630] = data_i[11630] & sel_one_hot_i[90];
  assign data_masked[11629] = data_i[11629] & sel_one_hot_i[90];
  assign data_masked[11628] = data_i[11628] & sel_one_hot_i[90];
  assign data_masked[11627] = data_i[11627] & sel_one_hot_i[90];
  assign data_masked[11626] = data_i[11626] & sel_one_hot_i[90];
  assign data_masked[11625] = data_i[11625] & sel_one_hot_i[90];
  assign data_masked[11624] = data_i[11624] & sel_one_hot_i[90];
  assign data_masked[11623] = data_i[11623] & sel_one_hot_i[90];
  assign data_masked[11622] = data_i[11622] & sel_one_hot_i[90];
  assign data_masked[11621] = data_i[11621] & sel_one_hot_i[90];
  assign data_masked[11620] = data_i[11620] & sel_one_hot_i[90];
  assign data_masked[11619] = data_i[11619] & sel_one_hot_i[90];
  assign data_masked[11618] = data_i[11618] & sel_one_hot_i[90];
  assign data_masked[11617] = data_i[11617] & sel_one_hot_i[90];
  assign data_masked[11616] = data_i[11616] & sel_one_hot_i[90];
  assign data_masked[11615] = data_i[11615] & sel_one_hot_i[90];
  assign data_masked[11614] = data_i[11614] & sel_one_hot_i[90];
  assign data_masked[11613] = data_i[11613] & sel_one_hot_i[90];
  assign data_masked[11612] = data_i[11612] & sel_one_hot_i[90];
  assign data_masked[11611] = data_i[11611] & sel_one_hot_i[90];
  assign data_masked[11610] = data_i[11610] & sel_one_hot_i[90];
  assign data_masked[11609] = data_i[11609] & sel_one_hot_i[90];
  assign data_masked[11608] = data_i[11608] & sel_one_hot_i[90];
  assign data_masked[11607] = data_i[11607] & sel_one_hot_i[90];
  assign data_masked[11606] = data_i[11606] & sel_one_hot_i[90];
  assign data_masked[11605] = data_i[11605] & sel_one_hot_i[90];
  assign data_masked[11604] = data_i[11604] & sel_one_hot_i[90];
  assign data_masked[11603] = data_i[11603] & sel_one_hot_i[90];
  assign data_masked[11602] = data_i[11602] & sel_one_hot_i[90];
  assign data_masked[11601] = data_i[11601] & sel_one_hot_i[90];
  assign data_masked[11600] = data_i[11600] & sel_one_hot_i[90];
  assign data_masked[11599] = data_i[11599] & sel_one_hot_i[90];
  assign data_masked[11598] = data_i[11598] & sel_one_hot_i[90];
  assign data_masked[11597] = data_i[11597] & sel_one_hot_i[90];
  assign data_masked[11596] = data_i[11596] & sel_one_hot_i[90];
  assign data_masked[11595] = data_i[11595] & sel_one_hot_i[90];
  assign data_masked[11594] = data_i[11594] & sel_one_hot_i[90];
  assign data_masked[11593] = data_i[11593] & sel_one_hot_i[90];
  assign data_masked[11592] = data_i[11592] & sel_one_hot_i[90];
  assign data_masked[11591] = data_i[11591] & sel_one_hot_i[90];
  assign data_masked[11590] = data_i[11590] & sel_one_hot_i[90];
  assign data_masked[11589] = data_i[11589] & sel_one_hot_i[90];
  assign data_masked[11588] = data_i[11588] & sel_one_hot_i[90];
  assign data_masked[11587] = data_i[11587] & sel_one_hot_i[90];
  assign data_masked[11586] = data_i[11586] & sel_one_hot_i[90];
  assign data_masked[11585] = data_i[11585] & sel_one_hot_i[90];
  assign data_masked[11584] = data_i[11584] & sel_one_hot_i[90];
  assign data_masked[11583] = data_i[11583] & sel_one_hot_i[90];
  assign data_masked[11582] = data_i[11582] & sel_one_hot_i[90];
  assign data_masked[11581] = data_i[11581] & sel_one_hot_i[90];
  assign data_masked[11580] = data_i[11580] & sel_one_hot_i[90];
  assign data_masked[11579] = data_i[11579] & sel_one_hot_i[90];
  assign data_masked[11578] = data_i[11578] & sel_one_hot_i[90];
  assign data_masked[11577] = data_i[11577] & sel_one_hot_i[90];
  assign data_masked[11576] = data_i[11576] & sel_one_hot_i[90];
  assign data_masked[11575] = data_i[11575] & sel_one_hot_i[90];
  assign data_masked[11574] = data_i[11574] & sel_one_hot_i[90];
  assign data_masked[11573] = data_i[11573] & sel_one_hot_i[90];
  assign data_masked[11572] = data_i[11572] & sel_one_hot_i[90];
  assign data_masked[11571] = data_i[11571] & sel_one_hot_i[90];
  assign data_masked[11570] = data_i[11570] & sel_one_hot_i[90];
  assign data_masked[11569] = data_i[11569] & sel_one_hot_i[90];
  assign data_masked[11568] = data_i[11568] & sel_one_hot_i[90];
  assign data_masked[11567] = data_i[11567] & sel_one_hot_i[90];
  assign data_masked[11566] = data_i[11566] & sel_one_hot_i[90];
  assign data_masked[11565] = data_i[11565] & sel_one_hot_i[90];
  assign data_masked[11564] = data_i[11564] & sel_one_hot_i[90];
  assign data_masked[11563] = data_i[11563] & sel_one_hot_i[90];
  assign data_masked[11562] = data_i[11562] & sel_one_hot_i[90];
  assign data_masked[11561] = data_i[11561] & sel_one_hot_i[90];
  assign data_masked[11560] = data_i[11560] & sel_one_hot_i[90];
  assign data_masked[11559] = data_i[11559] & sel_one_hot_i[90];
  assign data_masked[11558] = data_i[11558] & sel_one_hot_i[90];
  assign data_masked[11557] = data_i[11557] & sel_one_hot_i[90];
  assign data_masked[11556] = data_i[11556] & sel_one_hot_i[90];
  assign data_masked[11555] = data_i[11555] & sel_one_hot_i[90];
  assign data_masked[11554] = data_i[11554] & sel_one_hot_i[90];
  assign data_masked[11553] = data_i[11553] & sel_one_hot_i[90];
  assign data_masked[11552] = data_i[11552] & sel_one_hot_i[90];
  assign data_masked[11551] = data_i[11551] & sel_one_hot_i[90];
  assign data_masked[11550] = data_i[11550] & sel_one_hot_i[90];
  assign data_masked[11549] = data_i[11549] & sel_one_hot_i[90];
  assign data_masked[11548] = data_i[11548] & sel_one_hot_i[90];
  assign data_masked[11547] = data_i[11547] & sel_one_hot_i[90];
  assign data_masked[11546] = data_i[11546] & sel_one_hot_i[90];
  assign data_masked[11545] = data_i[11545] & sel_one_hot_i[90];
  assign data_masked[11544] = data_i[11544] & sel_one_hot_i[90];
  assign data_masked[11543] = data_i[11543] & sel_one_hot_i[90];
  assign data_masked[11542] = data_i[11542] & sel_one_hot_i[90];
  assign data_masked[11541] = data_i[11541] & sel_one_hot_i[90];
  assign data_masked[11540] = data_i[11540] & sel_one_hot_i[90];
  assign data_masked[11539] = data_i[11539] & sel_one_hot_i[90];
  assign data_masked[11538] = data_i[11538] & sel_one_hot_i[90];
  assign data_masked[11537] = data_i[11537] & sel_one_hot_i[90];
  assign data_masked[11536] = data_i[11536] & sel_one_hot_i[90];
  assign data_masked[11535] = data_i[11535] & sel_one_hot_i[90];
  assign data_masked[11534] = data_i[11534] & sel_one_hot_i[90];
  assign data_masked[11533] = data_i[11533] & sel_one_hot_i[90];
  assign data_masked[11532] = data_i[11532] & sel_one_hot_i[90];
  assign data_masked[11531] = data_i[11531] & sel_one_hot_i[90];
  assign data_masked[11530] = data_i[11530] & sel_one_hot_i[90];
  assign data_masked[11529] = data_i[11529] & sel_one_hot_i[90];
  assign data_masked[11528] = data_i[11528] & sel_one_hot_i[90];
  assign data_masked[11527] = data_i[11527] & sel_one_hot_i[90];
  assign data_masked[11526] = data_i[11526] & sel_one_hot_i[90];
  assign data_masked[11525] = data_i[11525] & sel_one_hot_i[90];
  assign data_masked[11524] = data_i[11524] & sel_one_hot_i[90];
  assign data_masked[11523] = data_i[11523] & sel_one_hot_i[90];
  assign data_masked[11522] = data_i[11522] & sel_one_hot_i[90];
  assign data_masked[11521] = data_i[11521] & sel_one_hot_i[90];
  assign data_masked[11520] = data_i[11520] & sel_one_hot_i[90];
  assign data_masked[11775] = data_i[11775] & sel_one_hot_i[91];
  assign data_masked[11774] = data_i[11774] & sel_one_hot_i[91];
  assign data_masked[11773] = data_i[11773] & sel_one_hot_i[91];
  assign data_masked[11772] = data_i[11772] & sel_one_hot_i[91];
  assign data_masked[11771] = data_i[11771] & sel_one_hot_i[91];
  assign data_masked[11770] = data_i[11770] & sel_one_hot_i[91];
  assign data_masked[11769] = data_i[11769] & sel_one_hot_i[91];
  assign data_masked[11768] = data_i[11768] & sel_one_hot_i[91];
  assign data_masked[11767] = data_i[11767] & sel_one_hot_i[91];
  assign data_masked[11766] = data_i[11766] & sel_one_hot_i[91];
  assign data_masked[11765] = data_i[11765] & sel_one_hot_i[91];
  assign data_masked[11764] = data_i[11764] & sel_one_hot_i[91];
  assign data_masked[11763] = data_i[11763] & sel_one_hot_i[91];
  assign data_masked[11762] = data_i[11762] & sel_one_hot_i[91];
  assign data_masked[11761] = data_i[11761] & sel_one_hot_i[91];
  assign data_masked[11760] = data_i[11760] & sel_one_hot_i[91];
  assign data_masked[11759] = data_i[11759] & sel_one_hot_i[91];
  assign data_masked[11758] = data_i[11758] & sel_one_hot_i[91];
  assign data_masked[11757] = data_i[11757] & sel_one_hot_i[91];
  assign data_masked[11756] = data_i[11756] & sel_one_hot_i[91];
  assign data_masked[11755] = data_i[11755] & sel_one_hot_i[91];
  assign data_masked[11754] = data_i[11754] & sel_one_hot_i[91];
  assign data_masked[11753] = data_i[11753] & sel_one_hot_i[91];
  assign data_masked[11752] = data_i[11752] & sel_one_hot_i[91];
  assign data_masked[11751] = data_i[11751] & sel_one_hot_i[91];
  assign data_masked[11750] = data_i[11750] & sel_one_hot_i[91];
  assign data_masked[11749] = data_i[11749] & sel_one_hot_i[91];
  assign data_masked[11748] = data_i[11748] & sel_one_hot_i[91];
  assign data_masked[11747] = data_i[11747] & sel_one_hot_i[91];
  assign data_masked[11746] = data_i[11746] & sel_one_hot_i[91];
  assign data_masked[11745] = data_i[11745] & sel_one_hot_i[91];
  assign data_masked[11744] = data_i[11744] & sel_one_hot_i[91];
  assign data_masked[11743] = data_i[11743] & sel_one_hot_i[91];
  assign data_masked[11742] = data_i[11742] & sel_one_hot_i[91];
  assign data_masked[11741] = data_i[11741] & sel_one_hot_i[91];
  assign data_masked[11740] = data_i[11740] & sel_one_hot_i[91];
  assign data_masked[11739] = data_i[11739] & sel_one_hot_i[91];
  assign data_masked[11738] = data_i[11738] & sel_one_hot_i[91];
  assign data_masked[11737] = data_i[11737] & sel_one_hot_i[91];
  assign data_masked[11736] = data_i[11736] & sel_one_hot_i[91];
  assign data_masked[11735] = data_i[11735] & sel_one_hot_i[91];
  assign data_masked[11734] = data_i[11734] & sel_one_hot_i[91];
  assign data_masked[11733] = data_i[11733] & sel_one_hot_i[91];
  assign data_masked[11732] = data_i[11732] & sel_one_hot_i[91];
  assign data_masked[11731] = data_i[11731] & sel_one_hot_i[91];
  assign data_masked[11730] = data_i[11730] & sel_one_hot_i[91];
  assign data_masked[11729] = data_i[11729] & sel_one_hot_i[91];
  assign data_masked[11728] = data_i[11728] & sel_one_hot_i[91];
  assign data_masked[11727] = data_i[11727] & sel_one_hot_i[91];
  assign data_masked[11726] = data_i[11726] & sel_one_hot_i[91];
  assign data_masked[11725] = data_i[11725] & sel_one_hot_i[91];
  assign data_masked[11724] = data_i[11724] & sel_one_hot_i[91];
  assign data_masked[11723] = data_i[11723] & sel_one_hot_i[91];
  assign data_masked[11722] = data_i[11722] & sel_one_hot_i[91];
  assign data_masked[11721] = data_i[11721] & sel_one_hot_i[91];
  assign data_masked[11720] = data_i[11720] & sel_one_hot_i[91];
  assign data_masked[11719] = data_i[11719] & sel_one_hot_i[91];
  assign data_masked[11718] = data_i[11718] & sel_one_hot_i[91];
  assign data_masked[11717] = data_i[11717] & sel_one_hot_i[91];
  assign data_masked[11716] = data_i[11716] & sel_one_hot_i[91];
  assign data_masked[11715] = data_i[11715] & sel_one_hot_i[91];
  assign data_masked[11714] = data_i[11714] & sel_one_hot_i[91];
  assign data_masked[11713] = data_i[11713] & sel_one_hot_i[91];
  assign data_masked[11712] = data_i[11712] & sel_one_hot_i[91];
  assign data_masked[11711] = data_i[11711] & sel_one_hot_i[91];
  assign data_masked[11710] = data_i[11710] & sel_one_hot_i[91];
  assign data_masked[11709] = data_i[11709] & sel_one_hot_i[91];
  assign data_masked[11708] = data_i[11708] & sel_one_hot_i[91];
  assign data_masked[11707] = data_i[11707] & sel_one_hot_i[91];
  assign data_masked[11706] = data_i[11706] & sel_one_hot_i[91];
  assign data_masked[11705] = data_i[11705] & sel_one_hot_i[91];
  assign data_masked[11704] = data_i[11704] & sel_one_hot_i[91];
  assign data_masked[11703] = data_i[11703] & sel_one_hot_i[91];
  assign data_masked[11702] = data_i[11702] & sel_one_hot_i[91];
  assign data_masked[11701] = data_i[11701] & sel_one_hot_i[91];
  assign data_masked[11700] = data_i[11700] & sel_one_hot_i[91];
  assign data_masked[11699] = data_i[11699] & sel_one_hot_i[91];
  assign data_masked[11698] = data_i[11698] & sel_one_hot_i[91];
  assign data_masked[11697] = data_i[11697] & sel_one_hot_i[91];
  assign data_masked[11696] = data_i[11696] & sel_one_hot_i[91];
  assign data_masked[11695] = data_i[11695] & sel_one_hot_i[91];
  assign data_masked[11694] = data_i[11694] & sel_one_hot_i[91];
  assign data_masked[11693] = data_i[11693] & sel_one_hot_i[91];
  assign data_masked[11692] = data_i[11692] & sel_one_hot_i[91];
  assign data_masked[11691] = data_i[11691] & sel_one_hot_i[91];
  assign data_masked[11690] = data_i[11690] & sel_one_hot_i[91];
  assign data_masked[11689] = data_i[11689] & sel_one_hot_i[91];
  assign data_masked[11688] = data_i[11688] & sel_one_hot_i[91];
  assign data_masked[11687] = data_i[11687] & sel_one_hot_i[91];
  assign data_masked[11686] = data_i[11686] & sel_one_hot_i[91];
  assign data_masked[11685] = data_i[11685] & sel_one_hot_i[91];
  assign data_masked[11684] = data_i[11684] & sel_one_hot_i[91];
  assign data_masked[11683] = data_i[11683] & sel_one_hot_i[91];
  assign data_masked[11682] = data_i[11682] & sel_one_hot_i[91];
  assign data_masked[11681] = data_i[11681] & sel_one_hot_i[91];
  assign data_masked[11680] = data_i[11680] & sel_one_hot_i[91];
  assign data_masked[11679] = data_i[11679] & sel_one_hot_i[91];
  assign data_masked[11678] = data_i[11678] & sel_one_hot_i[91];
  assign data_masked[11677] = data_i[11677] & sel_one_hot_i[91];
  assign data_masked[11676] = data_i[11676] & sel_one_hot_i[91];
  assign data_masked[11675] = data_i[11675] & sel_one_hot_i[91];
  assign data_masked[11674] = data_i[11674] & sel_one_hot_i[91];
  assign data_masked[11673] = data_i[11673] & sel_one_hot_i[91];
  assign data_masked[11672] = data_i[11672] & sel_one_hot_i[91];
  assign data_masked[11671] = data_i[11671] & sel_one_hot_i[91];
  assign data_masked[11670] = data_i[11670] & sel_one_hot_i[91];
  assign data_masked[11669] = data_i[11669] & sel_one_hot_i[91];
  assign data_masked[11668] = data_i[11668] & sel_one_hot_i[91];
  assign data_masked[11667] = data_i[11667] & sel_one_hot_i[91];
  assign data_masked[11666] = data_i[11666] & sel_one_hot_i[91];
  assign data_masked[11665] = data_i[11665] & sel_one_hot_i[91];
  assign data_masked[11664] = data_i[11664] & sel_one_hot_i[91];
  assign data_masked[11663] = data_i[11663] & sel_one_hot_i[91];
  assign data_masked[11662] = data_i[11662] & sel_one_hot_i[91];
  assign data_masked[11661] = data_i[11661] & sel_one_hot_i[91];
  assign data_masked[11660] = data_i[11660] & sel_one_hot_i[91];
  assign data_masked[11659] = data_i[11659] & sel_one_hot_i[91];
  assign data_masked[11658] = data_i[11658] & sel_one_hot_i[91];
  assign data_masked[11657] = data_i[11657] & sel_one_hot_i[91];
  assign data_masked[11656] = data_i[11656] & sel_one_hot_i[91];
  assign data_masked[11655] = data_i[11655] & sel_one_hot_i[91];
  assign data_masked[11654] = data_i[11654] & sel_one_hot_i[91];
  assign data_masked[11653] = data_i[11653] & sel_one_hot_i[91];
  assign data_masked[11652] = data_i[11652] & sel_one_hot_i[91];
  assign data_masked[11651] = data_i[11651] & sel_one_hot_i[91];
  assign data_masked[11650] = data_i[11650] & sel_one_hot_i[91];
  assign data_masked[11649] = data_i[11649] & sel_one_hot_i[91];
  assign data_masked[11648] = data_i[11648] & sel_one_hot_i[91];
  assign data_masked[11903] = data_i[11903] & sel_one_hot_i[92];
  assign data_masked[11902] = data_i[11902] & sel_one_hot_i[92];
  assign data_masked[11901] = data_i[11901] & sel_one_hot_i[92];
  assign data_masked[11900] = data_i[11900] & sel_one_hot_i[92];
  assign data_masked[11899] = data_i[11899] & sel_one_hot_i[92];
  assign data_masked[11898] = data_i[11898] & sel_one_hot_i[92];
  assign data_masked[11897] = data_i[11897] & sel_one_hot_i[92];
  assign data_masked[11896] = data_i[11896] & sel_one_hot_i[92];
  assign data_masked[11895] = data_i[11895] & sel_one_hot_i[92];
  assign data_masked[11894] = data_i[11894] & sel_one_hot_i[92];
  assign data_masked[11893] = data_i[11893] & sel_one_hot_i[92];
  assign data_masked[11892] = data_i[11892] & sel_one_hot_i[92];
  assign data_masked[11891] = data_i[11891] & sel_one_hot_i[92];
  assign data_masked[11890] = data_i[11890] & sel_one_hot_i[92];
  assign data_masked[11889] = data_i[11889] & sel_one_hot_i[92];
  assign data_masked[11888] = data_i[11888] & sel_one_hot_i[92];
  assign data_masked[11887] = data_i[11887] & sel_one_hot_i[92];
  assign data_masked[11886] = data_i[11886] & sel_one_hot_i[92];
  assign data_masked[11885] = data_i[11885] & sel_one_hot_i[92];
  assign data_masked[11884] = data_i[11884] & sel_one_hot_i[92];
  assign data_masked[11883] = data_i[11883] & sel_one_hot_i[92];
  assign data_masked[11882] = data_i[11882] & sel_one_hot_i[92];
  assign data_masked[11881] = data_i[11881] & sel_one_hot_i[92];
  assign data_masked[11880] = data_i[11880] & sel_one_hot_i[92];
  assign data_masked[11879] = data_i[11879] & sel_one_hot_i[92];
  assign data_masked[11878] = data_i[11878] & sel_one_hot_i[92];
  assign data_masked[11877] = data_i[11877] & sel_one_hot_i[92];
  assign data_masked[11876] = data_i[11876] & sel_one_hot_i[92];
  assign data_masked[11875] = data_i[11875] & sel_one_hot_i[92];
  assign data_masked[11874] = data_i[11874] & sel_one_hot_i[92];
  assign data_masked[11873] = data_i[11873] & sel_one_hot_i[92];
  assign data_masked[11872] = data_i[11872] & sel_one_hot_i[92];
  assign data_masked[11871] = data_i[11871] & sel_one_hot_i[92];
  assign data_masked[11870] = data_i[11870] & sel_one_hot_i[92];
  assign data_masked[11869] = data_i[11869] & sel_one_hot_i[92];
  assign data_masked[11868] = data_i[11868] & sel_one_hot_i[92];
  assign data_masked[11867] = data_i[11867] & sel_one_hot_i[92];
  assign data_masked[11866] = data_i[11866] & sel_one_hot_i[92];
  assign data_masked[11865] = data_i[11865] & sel_one_hot_i[92];
  assign data_masked[11864] = data_i[11864] & sel_one_hot_i[92];
  assign data_masked[11863] = data_i[11863] & sel_one_hot_i[92];
  assign data_masked[11862] = data_i[11862] & sel_one_hot_i[92];
  assign data_masked[11861] = data_i[11861] & sel_one_hot_i[92];
  assign data_masked[11860] = data_i[11860] & sel_one_hot_i[92];
  assign data_masked[11859] = data_i[11859] & sel_one_hot_i[92];
  assign data_masked[11858] = data_i[11858] & sel_one_hot_i[92];
  assign data_masked[11857] = data_i[11857] & sel_one_hot_i[92];
  assign data_masked[11856] = data_i[11856] & sel_one_hot_i[92];
  assign data_masked[11855] = data_i[11855] & sel_one_hot_i[92];
  assign data_masked[11854] = data_i[11854] & sel_one_hot_i[92];
  assign data_masked[11853] = data_i[11853] & sel_one_hot_i[92];
  assign data_masked[11852] = data_i[11852] & sel_one_hot_i[92];
  assign data_masked[11851] = data_i[11851] & sel_one_hot_i[92];
  assign data_masked[11850] = data_i[11850] & sel_one_hot_i[92];
  assign data_masked[11849] = data_i[11849] & sel_one_hot_i[92];
  assign data_masked[11848] = data_i[11848] & sel_one_hot_i[92];
  assign data_masked[11847] = data_i[11847] & sel_one_hot_i[92];
  assign data_masked[11846] = data_i[11846] & sel_one_hot_i[92];
  assign data_masked[11845] = data_i[11845] & sel_one_hot_i[92];
  assign data_masked[11844] = data_i[11844] & sel_one_hot_i[92];
  assign data_masked[11843] = data_i[11843] & sel_one_hot_i[92];
  assign data_masked[11842] = data_i[11842] & sel_one_hot_i[92];
  assign data_masked[11841] = data_i[11841] & sel_one_hot_i[92];
  assign data_masked[11840] = data_i[11840] & sel_one_hot_i[92];
  assign data_masked[11839] = data_i[11839] & sel_one_hot_i[92];
  assign data_masked[11838] = data_i[11838] & sel_one_hot_i[92];
  assign data_masked[11837] = data_i[11837] & sel_one_hot_i[92];
  assign data_masked[11836] = data_i[11836] & sel_one_hot_i[92];
  assign data_masked[11835] = data_i[11835] & sel_one_hot_i[92];
  assign data_masked[11834] = data_i[11834] & sel_one_hot_i[92];
  assign data_masked[11833] = data_i[11833] & sel_one_hot_i[92];
  assign data_masked[11832] = data_i[11832] & sel_one_hot_i[92];
  assign data_masked[11831] = data_i[11831] & sel_one_hot_i[92];
  assign data_masked[11830] = data_i[11830] & sel_one_hot_i[92];
  assign data_masked[11829] = data_i[11829] & sel_one_hot_i[92];
  assign data_masked[11828] = data_i[11828] & sel_one_hot_i[92];
  assign data_masked[11827] = data_i[11827] & sel_one_hot_i[92];
  assign data_masked[11826] = data_i[11826] & sel_one_hot_i[92];
  assign data_masked[11825] = data_i[11825] & sel_one_hot_i[92];
  assign data_masked[11824] = data_i[11824] & sel_one_hot_i[92];
  assign data_masked[11823] = data_i[11823] & sel_one_hot_i[92];
  assign data_masked[11822] = data_i[11822] & sel_one_hot_i[92];
  assign data_masked[11821] = data_i[11821] & sel_one_hot_i[92];
  assign data_masked[11820] = data_i[11820] & sel_one_hot_i[92];
  assign data_masked[11819] = data_i[11819] & sel_one_hot_i[92];
  assign data_masked[11818] = data_i[11818] & sel_one_hot_i[92];
  assign data_masked[11817] = data_i[11817] & sel_one_hot_i[92];
  assign data_masked[11816] = data_i[11816] & sel_one_hot_i[92];
  assign data_masked[11815] = data_i[11815] & sel_one_hot_i[92];
  assign data_masked[11814] = data_i[11814] & sel_one_hot_i[92];
  assign data_masked[11813] = data_i[11813] & sel_one_hot_i[92];
  assign data_masked[11812] = data_i[11812] & sel_one_hot_i[92];
  assign data_masked[11811] = data_i[11811] & sel_one_hot_i[92];
  assign data_masked[11810] = data_i[11810] & sel_one_hot_i[92];
  assign data_masked[11809] = data_i[11809] & sel_one_hot_i[92];
  assign data_masked[11808] = data_i[11808] & sel_one_hot_i[92];
  assign data_masked[11807] = data_i[11807] & sel_one_hot_i[92];
  assign data_masked[11806] = data_i[11806] & sel_one_hot_i[92];
  assign data_masked[11805] = data_i[11805] & sel_one_hot_i[92];
  assign data_masked[11804] = data_i[11804] & sel_one_hot_i[92];
  assign data_masked[11803] = data_i[11803] & sel_one_hot_i[92];
  assign data_masked[11802] = data_i[11802] & sel_one_hot_i[92];
  assign data_masked[11801] = data_i[11801] & sel_one_hot_i[92];
  assign data_masked[11800] = data_i[11800] & sel_one_hot_i[92];
  assign data_masked[11799] = data_i[11799] & sel_one_hot_i[92];
  assign data_masked[11798] = data_i[11798] & sel_one_hot_i[92];
  assign data_masked[11797] = data_i[11797] & sel_one_hot_i[92];
  assign data_masked[11796] = data_i[11796] & sel_one_hot_i[92];
  assign data_masked[11795] = data_i[11795] & sel_one_hot_i[92];
  assign data_masked[11794] = data_i[11794] & sel_one_hot_i[92];
  assign data_masked[11793] = data_i[11793] & sel_one_hot_i[92];
  assign data_masked[11792] = data_i[11792] & sel_one_hot_i[92];
  assign data_masked[11791] = data_i[11791] & sel_one_hot_i[92];
  assign data_masked[11790] = data_i[11790] & sel_one_hot_i[92];
  assign data_masked[11789] = data_i[11789] & sel_one_hot_i[92];
  assign data_masked[11788] = data_i[11788] & sel_one_hot_i[92];
  assign data_masked[11787] = data_i[11787] & sel_one_hot_i[92];
  assign data_masked[11786] = data_i[11786] & sel_one_hot_i[92];
  assign data_masked[11785] = data_i[11785] & sel_one_hot_i[92];
  assign data_masked[11784] = data_i[11784] & sel_one_hot_i[92];
  assign data_masked[11783] = data_i[11783] & sel_one_hot_i[92];
  assign data_masked[11782] = data_i[11782] & sel_one_hot_i[92];
  assign data_masked[11781] = data_i[11781] & sel_one_hot_i[92];
  assign data_masked[11780] = data_i[11780] & sel_one_hot_i[92];
  assign data_masked[11779] = data_i[11779] & sel_one_hot_i[92];
  assign data_masked[11778] = data_i[11778] & sel_one_hot_i[92];
  assign data_masked[11777] = data_i[11777] & sel_one_hot_i[92];
  assign data_masked[11776] = data_i[11776] & sel_one_hot_i[92];
  assign data_masked[12031] = data_i[12031] & sel_one_hot_i[93];
  assign data_masked[12030] = data_i[12030] & sel_one_hot_i[93];
  assign data_masked[12029] = data_i[12029] & sel_one_hot_i[93];
  assign data_masked[12028] = data_i[12028] & sel_one_hot_i[93];
  assign data_masked[12027] = data_i[12027] & sel_one_hot_i[93];
  assign data_masked[12026] = data_i[12026] & sel_one_hot_i[93];
  assign data_masked[12025] = data_i[12025] & sel_one_hot_i[93];
  assign data_masked[12024] = data_i[12024] & sel_one_hot_i[93];
  assign data_masked[12023] = data_i[12023] & sel_one_hot_i[93];
  assign data_masked[12022] = data_i[12022] & sel_one_hot_i[93];
  assign data_masked[12021] = data_i[12021] & sel_one_hot_i[93];
  assign data_masked[12020] = data_i[12020] & sel_one_hot_i[93];
  assign data_masked[12019] = data_i[12019] & sel_one_hot_i[93];
  assign data_masked[12018] = data_i[12018] & sel_one_hot_i[93];
  assign data_masked[12017] = data_i[12017] & sel_one_hot_i[93];
  assign data_masked[12016] = data_i[12016] & sel_one_hot_i[93];
  assign data_masked[12015] = data_i[12015] & sel_one_hot_i[93];
  assign data_masked[12014] = data_i[12014] & sel_one_hot_i[93];
  assign data_masked[12013] = data_i[12013] & sel_one_hot_i[93];
  assign data_masked[12012] = data_i[12012] & sel_one_hot_i[93];
  assign data_masked[12011] = data_i[12011] & sel_one_hot_i[93];
  assign data_masked[12010] = data_i[12010] & sel_one_hot_i[93];
  assign data_masked[12009] = data_i[12009] & sel_one_hot_i[93];
  assign data_masked[12008] = data_i[12008] & sel_one_hot_i[93];
  assign data_masked[12007] = data_i[12007] & sel_one_hot_i[93];
  assign data_masked[12006] = data_i[12006] & sel_one_hot_i[93];
  assign data_masked[12005] = data_i[12005] & sel_one_hot_i[93];
  assign data_masked[12004] = data_i[12004] & sel_one_hot_i[93];
  assign data_masked[12003] = data_i[12003] & sel_one_hot_i[93];
  assign data_masked[12002] = data_i[12002] & sel_one_hot_i[93];
  assign data_masked[12001] = data_i[12001] & sel_one_hot_i[93];
  assign data_masked[12000] = data_i[12000] & sel_one_hot_i[93];
  assign data_masked[11999] = data_i[11999] & sel_one_hot_i[93];
  assign data_masked[11998] = data_i[11998] & sel_one_hot_i[93];
  assign data_masked[11997] = data_i[11997] & sel_one_hot_i[93];
  assign data_masked[11996] = data_i[11996] & sel_one_hot_i[93];
  assign data_masked[11995] = data_i[11995] & sel_one_hot_i[93];
  assign data_masked[11994] = data_i[11994] & sel_one_hot_i[93];
  assign data_masked[11993] = data_i[11993] & sel_one_hot_i[93];
  assign data_masked[11992] = data_i[11992] & sel_one_hot_i[93];
  assign data_masked[11991] = data_i[11991] & sel_one_hot_i[93];
  assign data_masked[11990] = data_i[11990] & sel_one_hot_i[93];
  assign data_masked[11989] = data_i[11989] & sel_one_hot_i[93];
  assign data_masked[11988] = data_i[11988] & sel_one_hot_i[93];
  assign data_masked[11987] = data_i[11987] & sel_one_hot_i[93];
  assign data_masked[11986] = data_i[11986] & sel_one_hot_i[93];
  assign data_masked[11985] = data_i[11985] & sel_one_hot_i[93];
  assign data_masked[11984] = data_i[11984] & sel_one_hot_i[93];
  assign data_masked[11983] = data_i[11983] & sel_one_hot_i[93];
  assign data_masked[11982] = data_i[11982] & sel_one_hot_i[93];
  assign data_masked[11981] = data_i[11981] & sel_one_hot_i[93];
  assign data_masked[11980] = data_i[11980] & sel_one_hot_i[93];
  assign data_masked[11979] = data_i[11979] & sel_one_hot_i[93];
  assign data_masked[11978] = data_i[11978] & sel_one_hot_i[93];
  assign data_masked[11977] = data_i[11977] & sel_one_hot_i[93];
  assign data_masked[11976] = data_i[11976] & sel_one_hot_i[93];
  assign data_masked[11975] = data_i[11975] & sel_one_hot_i[93];
  assign data_masked[11974] = data_i[11974] & sel_one_hot_i[93];
  assign data_masked[11973] = data_i[11973] & sel_one_hot_i[93];
  assign data_masked[11972] = data_i[11972] & sel_one_hot_i[93];
  assign data_masked[11971] = data_i[11971] & sel_one_hot_i[93];
  assign data_masked[11970] = data_i[11970] & sel_one_hot_i[93];
  assign data_masked[11969] = data_i[11969] & sel_one_hot_i[93];
  assign data_masked[11968] = data_i[11968] & sel_one_hot_i[93];
  assign data_masked[11967] = data_i[11967] & sel_one_hot_i[93];
  assign data_masked[11966] = data_i[11966] & sel_one_hot_i[93];
  assign data_masked[11965] = data_i[11965] & sel_one_hot_i[93];
  assign data_masked[11964] = data_i[11964] & sel_one_hot_i[93];
  assign data_masked[11963] = data_i[11963] & sel_one_hot_i[93];
  assign data_masked[11962] = data_i[11962] & sel_one_hot_i[93];
  assign data_masked[11961] = data_i[11961] & sel_one_hot_i[93];
  assign data_masked[11960] = data_i[11960] & sel_one_hot_i[93];
  assign data_masked[11959] = data_i[11959] & sel_one_hot_i[93];
  assign data_masked[11958] = data_i[11958] & sel_one_hot_i[93];
  assign data_masked[11957] = data_i[11957] & sel_one_hot_i[93];
  assign data_masked[11956] = data_i[11956] & sel_one_hot_i[93];
  assign data_masked[11955] = data_i[11955] & sel_one_hot_i[93];
  assign data_masked[11954] = data_i[11954] & sel_one_hot_i[93];
  assign data_masked[11953] = data_i[11953] & sel_one_hot_i[93];
  assign data_masked[11952] = data_i[11952] & sel_one_hot_i[93];
  assign data_masked[11951] = data_i[11951] & sel_one_hot_i[93];
  assign data_masked[11950] = data_i[11950] & sel_one_hot_i[93];
  assign data_masked[11949] = data_i[11949] & sel_one_hot_i[93];
  assign data_masked[11948] = data_i[11948] & sel_one_hot_i[93];
  assign data_masked[11947] = data_i[11947] & sel_one_hot_i[93];
  assign data_masked[11946] = data_i[11946] & sel_one_hot_i[93];
  assign data_masked[11945] = data_i[11945] & sel_one_hot_i[93];
  assign data_masked[11944] = data_i[11944] & sel_one_hot_i[93];
  assign data_masked[11943] = data_i[11943] & sel_one_hot_i[93];
  assign data_masked[11942] = data_i[11942] & sel_one_hot_i[93];
  assign data_masked[11941] = data_i[11941] & sel_one_hot_i[93];
  assign data_masked[11940] = data_i[11940] & sel_one_hot_i[93];
  assign data_masked[11939] = data_i[11939] & sel_one_hot_i[93];
  assign data_masked[11938] = data_i[11938] & sel_one_hot_i[93];
  assign data_masked[11937] = data_i[11937] & sel_one_hot_i[93];
  assign data_masked[11936] = data_i[11936] & sel_one_hot_i[93];
  assign data_masked[11935] = data_i[11935] & sel_one_hot_i[93];
  assign data_masked[11934] = data_i[11934] & sel_one_hot_i[93];
  assign data_masked[11933] = data_i[11933] & sel_one_hot_i[93];
  assign data_masked[11932] = data_i[11932] & sel_one_hot_i[93];
  assign data_masked[11931] = data_i[11931] & sel_one_hot_i[93];
  assign data_masked[11930] = data_i[11930] & sel_one_hot_i[93];
  assign data_masked[11929] = data_i[11929] & sel_one_hot_i[93];
  assign data_masked[11928] = data_i[11928] & sel_one_hot_i[93];
  assign data_masked[11927] = data_i[11927] & sel_one_hot_i[93];
  assign data_masked[11926] = data_i[11926] & sel_one_hot_i[93];
  assign data_masked[11925] = data_i[11925] & sel_one_hot_i[93];
  assign data_masked[11924] = data_i[11924] & sel_one_hot_i[93];
  assign data_masked[11923] = data_i[11923] & sel_one_hot_i[93];
  assign data_masked[11922] = data_i[11922] & sel_one_hot_i[93];
  assign data_masked[11921] = data_i[11921] & sel_one_hot_i[93];
  assign data_masked[11920] = data_i[11920] & sel_one_hot_i[93];
  assign data_masked[11919] = data_i[11919] & sel_one_hot_i[93];
  assign data_masked[11918] = data_i[11918] & sel_one_hot_i[93];
  assign data_masked[11917] = data_i[11917] & sel_one_hot_i[93];
  assign data_masked[11916] = data_i[11916] & sel_one_hot_i[93];
  assign data_masked[11915] = data_i[11915] & sel_one_hot_i[93];
  assign data_masked[11914] = data_i[11914] & sel_one_hot_i[93];
  assign data_masked[11913] = data_i[11913] & sel_one_hot_i[93];
  assign data_masked[11912] = data_i[11912] & sel_one_hot_i[93];
  assign data_masked[11911] = data_i[11911] & sel_one_hot_i[93];
  assign data_masked[11910] = data_i[11910] & sel_one_hot_i[93];
  assign data_masked[11909] = data_i[11909] & sel_one_hot_i[93];
  assign data_masked[11908] = data_i[11908] & sel_one_hot_i[93];
  assign data_masked[11907] = data_i[11907] & sel_one_hot_i[93];
  assign data_masked[11906] = data_i[11906] & sel_one_hot_i[93];
  assign data_masked[11905] = data_i[11905] & sel_one_hot_i[93];
  assign data_masked[11904] = data_i[11904] & sel_one_hot_i[93];
  assign data_masked[12159] = data_i[12159] & sel_one_hot_i[94];
  assign data_masked[12158] = data_i[12158] & sel_one_hot_i[94];
  assign data_masked[12157] = data_i[12157] & sel_one_hot_i[94];
  assign data_masked[12156] = data_i[12156] & sel_one_hot_i[94];
  assign data_masked[12155] = data_i[12155] & sel_one_hot_i[94];
  assign data_masked[12154] = data_i[12154] & sel_one_hot_i[94];
  assign data_masked[12153] = data_i[12153] & sel_one_hot_i[94];
  assign data_masked[12152] = data_i[12152] & sel_one_hot_i[94];
  assign data_masked[12151] = data_i[12151] & sel_one_hot_i[94];
  assign data_masked[12150] = data_i[12150] & sel_one_hot_i[94];
  assign data_masked[12149] = data_i[12149] & sel_one_hot_i[94];
  assign data_masked[12148] = data_i[12148] & sel_one_hot_i[94];
  assign data_masked[12147] = data_i[12147] & sel_one_hot_i[94];
  assign data_masked[12146] = data_i[12146] & sel_one_hot_i[94];
  assign data_masked[12145] = data_i[12145] & sel_one_hot_i[94];
  assign data_masked[12144] = data_i[12144] & sel_one_hot_i[94];
  assign data_masked[12143] = data_i[12143] & sel_one_hot_i[94];
  assign data_masked[12142] = data_i[12142] & sel_one_hot_i[94];
  assign data_masked[12141] = data_i[12141] & sel_one_hot_i[94];
  assign data_masked[12140] = data_i[12140] & sel_one_hot_i[94];
  assign data_masked[12139] = data_i[12139] & sel_one_hot_i[94];
  assign data_masked[12138] = data_i[12138] & sel_one_hot_i[94];
  assign data_masked[12137] = data_i[12137] & sel_one_hot_i[94];
  assign data_masked[12136] = data_i[12136] & sel_one_hot_i[94];
  assign data_masked[12135] = data_i[12135] & sel_one_hot_i[94];
  assign data_masked[12134] = data_i[12134] & sel_one_hot_i[94];
  assign data_masked[12133] = data_i[12133] & sel_one_hot_i[94];
  assign data_masked[12132] = data_i[12132] & sel_one_hot_i[94];
  assign data_masked[12131] = data_i[12131] & sel_one_hot_i[94];
  assign data_masked[12130] = data_i[12130] & sel_one_hot_i[94];
  assign data_masked[12129] = data_i[12129] & sel_one_hot_i[94];
  assign data_masked[12128] = data_i[12128] & sel_one_hot_i[94];
  assign data_masked[12127] = data_i[12127] & sel_one_hot_i[94];
  assign data_masked[12126] = data_i[12126] & sel_one_hot_i[94];
  assign data_masked[12125] = data_i[12125] & sel_one_hot_i[94];
  assign data_masked[12124] = data_i[12124] & sel_one_hot_i[94];
  assign data_masked[12123] = data_i[12123] & sel_one_hot_i[94];
  assign data_masked[12122] = data_i[12122] & sel_one_hot_i[94];
  assign data_masked[12121] = data_i[12121] & sel_one_hot_i[94];
  assign data_masked[12120] = data_i[12120] & sel_one_hot_i[94];
  assign data_masked[12119] = data_i[12119] & sel_one_hot_i[94];
  assign data_masked[12118] = data_i[12118] & sel_one_hot_i[94];
  assign data_masked[12117] = data_i[12117] & sel_one_hot_i[94];
  assign data_masked[12116] = data_i[12116] & sel_one_hot_i[94];
  assign data_masked[12115] = data_i[12115] & sel_one_hot_i[94];
  assign data_masked[12114] = data_i[12114] & sel_one_hot_i[94];
  assign data_masked[12113] = data_i[12113] & sel_one_hot_i[94];
  assign data_masked[12112] = data_i[12112] & sel_one_hot_i[94];
  assign data_masked[12111] = data_i[12111] & sel_one_hot_i[94];
  assign data_masked[12110] = data_i[12110] & sel_one_hot_i[94];
  assign data_masked[12109] = data_i[12109] & sel_one_hot_i[94];
  assign data_masked[12108] = data_i[12108] & sel_one_hot_i[94];
  assign data_masked[12107] = data_i[12107] & sel_one_hot_i[94];
  assign data_masked[12106] = data_i[12106] & sel_one_hot_i[94];
  assign data_masked[12105] = data_i[12105] & sel_one_hot_i[94];
  assign data_masked[12104] = data_i[12104] & sel_one_hot_i[94];
  assign data_masked[12103] = data_i[12103] & sel_one_hot_i[94];
  assign data_masked[12102] = data_i[12102] & sel_one_hot_i[94];
  assign data_masked[12101] = data_i[12101] & sel_one_hot_i[94];
  assign data_masked[12100] = data_i[12100] & sel_one_hot_i[94];
  assign data_masked[12099] = data_i[12099] & sel_one_hot_i[94];
  assign data_masked[12098] = data_i[12098] & sel_one_hot_i[94];
  assign data_masked[12097] = data_i[12097] & sel_one_hot_i[94];
  assign data_masked[12096] = data_i[12096] & sel_one_hot_i[94];
  assign data_masked[12095] = data_i[12095] & sel_one_hot_i[94];
  assign data_masked[12094] = data_i[12094] & sel_one_hot_i[94];
  assign data_masked[12093] = data_i[12093] & sel_one_hot_i[94];
  assign data_masked[12092] = data_i[12092] & sel_one_hot_i[94];
  assign data_masked[12091] = data_i[12091] & sel_one_hot_i[94];
  assign data_masked[12090] = data_i[12090] & sel_one_hot_i[94];
  assign data_masked[12089] = data_i[12089] & sel_one_hot_i[94];
  assign data_masked[12088] = data_i[12088] & sel_one_hot_i[94];
  assign data_masked[12087] = data_i[12087] & sel_one_hot_i[94];
  assign data_masked[12086] = data_i[12086] & sel_one_hot_i[94];
  assign data_masked[12085] = data_i[12085] & sel_one_hot_i[94];
  assign data_masked[12084] = data_i[12084] & sel_one_hot_i[94];
  assign data_masked[12083] = data_i[12083] & sel_one_hot_i[94];
  assign data_masked[12082] = data_i[12082] & sel_one_hot_i[94];
  assign data_masked[12081] = data_i[12081] & sel_one_hot_i[94];
  assign data_masked[12080] = data_i[12080] & sel_one_hot_i[94];
  assign data_masked[12079] = data_i[12079] & sel_one_hot_i[94];
  assign data_masked[12078] = data_i[12078] & sel_one_hot_i[94];
  assign data_masked[12077] = data_i[12077] & sel_one_hot_i[94];
  assign data_masked[12076] = data_i[12076] & sel_one_hot_i[94];
  assign data_masked[12075] = data_i[12075] & sel_one_hot_i[94];
  assign data_masked[12074] = data_i[12074] & sel_one_hot_i[94];
  assign data_masked[12073] = data_i[12073] & sel_one_hot_i[94];
  assign data_masked[12072] = data_i[12072] & sel_one_hot_i[94];
  assign data_masked[12071] = data_i[12071] & sel_one_hot_i[94];
  assign data_masked[12070] = data_i[12070] & sel_one_hot_i[94];
  assign data_masked[12069] = data_i[12069] & sel_one_hot_i[94];
  assign data_masked[12068] = data_i[12068] & sel_one_hot_i[94];
  assign data_masked[12067] = data_i[12067] & sel_one_hot_i[94];
  assign data_masked[12066] = data_i[12066] & sel_one_hot_i[94];
  assign data_masked[12065] = data_i[12065] & sel_one_hot_i[94];
  assign data_masked[12064] = data_i[12064] & sel_one_hot_i[94];
  assign data_masked[12063] = data_i[12063] & sel_one_hot_i[94];
  assign data_masked[12062] = data_i[12062] & sel_one_hot_i[94];
  assign data_masked[12061] = data_i[12061] & sel_one_hot_i[94];
  assign data_masked[12060] = data_i[12060] & sel_one_hot_i[94];
  assign data_masked[12059] = data_i[12059] & sel_one_hot_i[94];
  assign data_masked[12058] = data_i[12058] & sel_one_hot_i[94];
  assign data_masked[12057] = data_i[12057] & sel_one_hot_i[94];
  assign data_masked[12056] = data_i[12056] & sel_one_hot_i[94];
  assign data_masked[12055] = data_i[12055] & sel_one_hot_i[94];
  assign data_masked[12054] = data_i[12054] & sel_one_hot_i[94];
  assign data_masked[12053] = data_i[12053] & sel_one_hot_i[94];
  assign data_masked[12052] = data_i[12052] & sel_one_hot_i[94];
  assign data_masked[12051] = data_i[12051] & sel_one_hot_i[94];
  assign data_masked[12050] = data_i[12050] & sel_one_hot_i[94];
  assign data_masked[12049] = data_i[12049] & sel_one_hot_i[94];
  assign data_masked[12048] = data_i[12048] & sel_one_hot_i[94];
  assign data_masked[12047] = data_i[12047] & sel_one_hot_i[94];
  assign data_masked[12046] = data_i[12046] & sel_one_hot_i[94];
  assign data_masked[12045] = data_i[12045] & sel_one_hot_i[94];
  assign data_masked[12044] = data_i[12044] & sel_one_hot_i[94];
  assign data_masked[12043] = data_i[12043] & sel_one_hot_i[94];
  assign data_masked[12042] = data_i[12042] & sel_one_hot_i[94];
  assign data_masked[12041] = data_i[12041] & sel_one_hot_i[94];
  assign data_masked[12040] = data_i[12040] & sel_one_hot_i[94];
  assign data_masked[12039] = data_i[12039] & sel_one_hot_i[94];
  assign data_masked[12038] = data_i[12038] & sel_one_hot_i[94];
  assign data_masked[12037] = data_i[12037] & sel_one_hot_i[94];
  assign data_masked[12036] = data_i[12036] & sel_one_hot_i[94];
  assign data_masked[12035] = data_i[12035] & sel_one_hot_i[94];
  assign data_masked[12034] = data_i[12034] & sel_one_hot_i[94];
  assign data_masked[12033] = data_i[12033] & sel_one_hot_i[94];
  assign data_masked[12032] = data_i[12032] & sel_one_hot_i[94];
  assign data_masked[12287] = data_i[12287] & sel_one_hot_i[95];
  assign data_masked[12286] = data_i[12286] & sel_one_hot_i[95];
  assign data_masked[12285] = data_i[12285] & sel_one_hot_i[95];
  assign data_masked[12284] = data_i[12284] & sel_one_hot_i[95];
  assign data_masked[12283] = data_i[12283] & sel_one_hot_i[95];
  assign data_masked[12282] = data_i[12282] & sel_one_hot_i[95];
  assign data_masked[12281] = data_i[12281] & sel_one_hot_i[95];
  assign data_masked[12280] = data_i[12280] & sel_one_hot_i[95];
  assign data_masked[12279] = data_i[12279] & sel_one_hot_i[95];
  assign data_masked[12278] = data_i[12278] & sel_one_hot_i[95];
  assign data_masked[12277] = data_i[12277] & sel_one_hot_i[95];
  assign data_masked[12276] = data_i[12276] & sel_one_hot_i[95];
  assign data_masked[12275] = data_i[12275] & sel_one_hot_i[95];
  assign data_masked[12274] = data_i[12274] & sel_one_hot_i[95];
  assign data_masked[12273] = data_i[12273] & sel_one_hot_i[95];
  assign data_masked[12272] = data_i[12272] & sel_one_hot_i[95];
  assign data_masked[12271] = data_i[12271] & sel_one_hot_i[95];
  assign data_masked[12270] = data_i[12270] & sel_one_hot_i[95];
  assign data_masked[12269] = data_i[12269] & sel_one_hot_i[95];
  assign data_masked[12268] = data_i[12268] & sel_one_hot_i[95];
  assign data_masked[12267] = data_i[12267] & sel_one_hot_i[95];
  assign data_masked[12266] = data_i[12266] & sel_one_hot_i[95];
  assign data_masked[12265] = data_i[12265] & sel_one_hot_i[95];
  assign data_masked[12264] = data_i[12264] & sel_one_hot_i[95];
  assign data_masked[12263] = data_i[12263] & sel_one_hot_i[95];
  assign data_masked[12262] = data_i[12262] & sel_one_hot_i[95];
  assign data_masked[12261] = data_i[12261] & sel_one_hot_i[95];
  assign data_masked[12260] = data_i[12260] & sel_one_hot_i[95];
  assign data_masked[12259] = data_i[12259] & sel_one_hot_i[95];
  assign data_masked[12258] = data_i[12258] & sel_one_hot_i[95];
  assign data_masked[12257] = data_i[12257] & sel_one_hot_i[95];
  assign data_masked[12256] = data_i[12256] & sel_one_hot_i[95];
  assign data_masked[12255] = data_i[12255] & sel_one_hot_i[95];
  assign data_masked[12254] = data_i[12254] & sel_one_hot_i[95];
  assign data_masked[12253] = data_i[12253] & sel_one_hot_i[95];
  assign data_masked[12252] = data_i[12252] & sel_one_hot_i[95];
  assign data_masked[12251] = data_i[12251] & sel_one_hot_i[95];
  assign data_masked[12250] = data_i[12250] & sel_one_hot_i[95];
  assign data_masked[12249] = data_i[12249] & sel_one_hot_i[95];
  assign data_masked[12248] = data_i[12248] & sel_one_hot_i[95];
  assign data_masked[12247] = data_i[12247] & sel_one_hot_i[95];
  assign data_masked[12246] = data_i[12246] & sel_one_hot_i[95];
  assign data_masked[12245] = data_i[12245] & sel_one_hot_i[95];
  assign data_masked[12244] = data_i[12244] & sel_one_hot_i[95];
  assign data_masked[12243] = data_i[12243] & sel_one_hot_i[95];
  assign data_masked[12242] = data_i[12242] & sel_one_hot_i[95];
  assign data_masked[12241] = data_i[12241] & sel_one_hot_i[95];
  assign data_masked[12240] = data_i[12240] & sel_one_hot_i[95];
  assign data_masked[12239] = data_i[12239] & sel_one_hot_i[95];
  assign data_masked[12238] = data_i[12238] & sel_one_hot_i[95];
  assign data_masked[12237] = data_i[12237] & sel_one_hot_i[95];
  assign data_masked[12236] = data_i[12236] & sel_one_hot_i[95];
  assign data_masked[12235] = data_i[12235] & sel_one_hot_i[95];
  assign data_masked[12234] = data_i[12234] & sel_one_hot_i[95];
  assign data_masked[12233] = data_i[12233] & sel_one_hot_i[95];
  assign data_masked[12232] = data_i[12232] & sel_one_hot_i[95];
  assign data_masked[12231] = data_i[12231] & sel_one_hot_i[95];
  assign data_masked[12230] = data_i[12230] & sel_one_hot_i[95];
  assign data_masked[12229] = data_i[12229] & sel_one_hot_i[95];
  assign data_masked[12228] = data_i[12228] & sel_one_hot_i[95];
  assign data_masked[12227] = data_i[12227] & sel_one_hot_i[95];
  assign data_masked[12226] = data_i[12226] & sel_one_hot_i[95];
  assign data_masked[12225] = data_i[12225] & sel_one_hot_i[95];
  assign data_masked[12224] = data_i[12224] & sel_one_hot_i[95];
  assign data_masked[12223] = data_i[12223] & sel_one_hot_i[95];
  assign data_masked[12222] = data_i[12222] & sel_one_hot_i[95];
  assign data_masked[12221] = data_i[12221] & sel_one_hot_i[95];
  assign data_masked[12220] = data_i[12220] & sel_one_hot_i[95];
  assign data_masked[12219] = data_i[12219] & sel_one_hot_i[95];
  assign data_masked[12218] = data_i[12218] & sel_one_hot_i[95];
  assign data_masked[12217] = data_i[12217] & sel_one_hot_i[95];
  assign data_masked[12216] = data_i[12216] & sel_one_hot_i[95];
  assign data_masked[12215] = data_i[12215] & sel_one_hot_i[95];
  assign data_masked[12214] = data_i[12214] & sel_one_hot_i[95];
  assign data_masked[12213] = data_i[12213] & sel_one_hot_i[95];
  assign data_masked[12212] = data_i[12212] & sel_one_hot_i[95];
  assign data_masked[12211] = data_i[12211] & sel_one_hot_i[95];
  assign data_masked[12210] = data_i[12210] & sel_one_hot_i[95];
  assign data_masked[12209] = data_i[12209] & sel_one_hot_i[95];
  assign data_masked[12208] = data_i[12208] & sel_one_hot_i[95];
  assign data_masked[12207] = data_i[12207] & sel_one_hot_i[95];
  assign data_masked[12206] = data_i[12206] & sel_one_hot_i[95];
  assign data_masked[12205] = data_i[12205] & sel_one_hot_i[95];
  assign data_masked[12204] = data_i[12204] & sel_one_hot_i[95];
  assign data_masked[12203] = data_i[12203] & sel_one_hot_i[95];
  assign data_masked[12202] = data_i[12202] & sel_one_hot_i[95];
  assign data_masked[12201] = data_i[12201] & sel_one_hot_i[95];
  assign data_masked[12200] = data_i[12200] & sel_one_hot_i[95];
  assign data_masked[12199] = data_i[12199] & sel_one_hot_i[95];
  assign data_masked[12198] = data_i[12198] & sel_one_hot_i[95];
  assign data_masked[12197] = data_i[12197] & sel_one_hot_i[95];
  assign data_masked[12196] = data_i[12196] & sel_one_hot_i[95];
  assign data_masked[12195] = data_i[12195] & sel_one_hot_i[95];
  assign data_masked[12194] = data_i[12194] & sel_one_hot_i[95];
  assign data_masked[12193] = data_i[12193] & sel_one_hot_i[95];
  assign data_masked[12192] = data_i[12192] & sel_one_hot_i[95];
  assign data_masked[12191] = data_i[12191] & sel_one_hot_i[95];
  assign data_masked[12190] = data_i[12190] & sel_one_hot_i[95];
  assign data_masked[12189] = data_i[12189] & sel_one_hot_i[95];
  assign data_masked[12188] = data_i[12188] & sel_one_hot_i[95];
  assign data_masked[12187] = data_i[12187] & sel_one_hot_i[95];
  assign data_masked[12186] = data_i[12186] & sel_one_hot_i[95];
  assign data_masked[12185] = data_i[12185] & sel_one_hot_i[95];
  assign data_masked[12184] = data_i[12184] & sel_one_hot_i[95];
  assign data_masked[12183] = data_i[12183] & sel_one_hot_i[95];
  assign data_masked[12182] = data_i[12182] & sel_one_hot_i[95];
  assign data_masked[12181] = data_i[12181] & sel_one_hot_i[95];
  assign data_masked[12180] = data_i[12180] & sel_one_hot_i[95];
  assign data_masked[12179] = data_i[12179] & sel_one_hot_i[95];
  assign data_masked[12178] = data_i[12178] & sel_one_hot_i[95];
  assign data_masked[12177] = data_i[12177] & sel_one_hot_i[95];
  assign data_masked[12176] = data_i[12176] & sel_one_hot_i[95];
  assign data_masked[12175] = data_i[12175] & sel_one_hot_i[95];
  assign data_masked[12174] = data_i[12174] & sel_one_hot_i[95];
  assign data_masked[12173] = data_i[12173] & sel_one_hot_i[95];
  assign data_masked[12172] = data_i[12172] & sel_one_hot_i[95];
  assign data_masked[12171] = data_i[12171] & sel_one_hot_i[95];
  assign data_masked[12170] = data_i[12170] & sel_one_hot_i[95];
  assign data_masked[12169] = data_i[12169] & sel_one_hot_i[95];
  assign data_masked[12168] = data_i[12168] & sel_one_hot_i[95];
  assign data_masked[12167] = data_i[12167] & sel_one_hot_i[95];
  assign data_masked[12166] = data_i[12166] & sel_one_hot_i[95];
  assign data_masked[12165] = data_i[12165] & sel_one_hot_i[95];
  assign data_masked[12164] = data_i[12164] & sel_one_hot_i[95];
  assign data_masked[12163] = data_i[12163] & sel_one_hot_i[95];
  assign data_masked[12162] = data_i[12162] & sel_one_hot_i[95];
  assign data_masked[12161] = data_i[12161] & sel_one_hot_i[95];
  assign data_masked[12160] = data_i[12160] & sel_one_hot_i[95];
  assign data_masked[12415] = data_i[12415] & sel_one_hot_i[96];
  assign data_masked[12414] = data_i[12414] & sel_one_hot_i[96];
  assign data_masked[12413] = data_i[12413] & sel_one_hot_i[96];
  assign data_masked[12412] = data_i[12412] & sel_one_hot_i[96];
  assign data_masked[12411] = data_i[12411] & sel_one_hot_i[96];
  assign data_masked[12410] = data_i[12410] & sel_one_hot_i[96];
  assign data_masked[12409] = data_i[12409] & sel_one_hot_i[96];
  assign data_masked[12408] = data_i[12408] & sel_one_hot_i[96];
  assign data_masked[12407] = data_i[12407] & sel_one_hot_i[96];
  assign data_masked[12406] = data_i[12406] & sel_one_hot_i[96];
  assign data_masked[12405] = data_i[12405] & sel_one_hot_i[96];
  assign data_masked[12404] = data_i[12404] & sel_one_hot_i[96];
  assign data_masked[12403] = data_i[12403] & sel_one_hot_i[96];
  assign data_masked[12402] = data_i[12402] & sel_one_hot_i[96];
  assign data_masked[12401] = data_i[12401] & sel_one_hot_i[96];
  assign data_masked[12400] = data_i[12400] & sel_one_hot_i[96];
  assign data_masked[12399] = data_i[12399] & sel_one_hot_i[96];
  assign data_masked[12398] = data_i[12398] & sel_one_hot_i[96];
  assign data_masked[12397] = data_i[12397] & sel_one_hot_i[96];
  assign data_masked[12396] = data_i[12396] & sel_one_hot_i[96];
  assign data_masked[12395] = data_i[12395] & sel_one_hot_i[96];
  assign data_masked[12394] = data_i[12394] & sel_one_hot_i[96];
  assign data_masked[12393] = data_i[12393] & sel_one_hot_i[96];
  assign data_masked[12392] = data_i[12392] & sel_one_hot_i[96];
  assign data_masked[12391] = data_i[12391] & sel_one_hot_i[96];
  assign data_masked[12390] = data_i[12390] & sel_one_hot_i[96];
  assign data_masked[12389] = data_i[12389] & sel_one_hot_i[96];
  assign data_masked[12388] = data_i[12388] & sel_one_hot_i[96];
  assign data_masked[12387] = data_i[12387] & sel_one_hot_i[96];
  assign data_masked[12386] = data_i[12386] & sel_one_hot_i[96];
  assign data_masked[12385] = data_i[12385] & sel_one_hot_i[96];
  assign data_masked[12384] = data_i[12384] & sel_one_hot_i[96];
  assign data_masked[12383] = data_i[12383] & sel_one_hot_i[96];
  assign data_masked[12382] = data_i[12382] & sel_one_hot_i[96];
  assign data_masked[12381] = data_i[12381] & sel_one_hot_i[96];
  assign data_masked[12380] = data_i[12380] & sel_one_hot_i[96];
  assign data_masked[12379] = data_i[12379] & sel_one_hot_i[96];
  assign data_masked[12378] = data_i[12378] & sel_one_hot_i[96];
  assign data_masked[12377] = data_i[12377] & sel_one_hot_i[96];
  assign data_masked[12376] = data_i[12376] & sel_one_hot_i[96];
  assign data_masked[12375] = data_i[12375] & sel_one_hot_i[96];
  assign data_masked[12374] = data_i[12374] & sel_one_hot_i[96];
  assign data_masked[12373] = data_i[12373] & sel_one_hot_i[96];
  assign data_masked[12372] = data_i[12372] & sel_one_hot_i[96];
  assign data_masked[12371] = data_i[12371] & sel_one_hot_i[96];
  assign data_masked[12370] = data_i[12370] & sel_one_hot_i[96];
  assign data_masked[12369] = data_i[12369] & sel_one_hot_i[96];
  assign data_masked[12368] = data_i[12368] & sel_one_hot_i[96];
  assign data_masked[12367] = data_i[12367] & sel_one_hot_i[96];
  assign data_masked[12366] = data_i[12366] & sel_one_hot_i[96];
  assign data_masked[12365] = data_i[12365] & sel_one_hot_i[96];
  assign data_masked[12364] = data_i[12364] & sel_one_hot_i[96];
  assign data_masked[12363] = data_i[12363] & sel_one_hot_i[96];
  assign data_masked[12362] = data_i[12362] & sel_one_hot_i[96];
  assign data_masked[12361] = data_i[12361] & sel_one_hot_i[96];
  assign data_masked[12360] = data_i[12360] & sel_one_hot_i[96];
  assign data_masked[12359] = data_i[12359] & sel_one_hot_i[96];
  assign data_masked[12358] = data_i[12358] & sel_one_hot_i[96];
  assign data_masked[12357] = data_i[12357] & sel_one_hot_i[96];
  assign data_masked[12356] = data_i[12356] & sel_one_hot_i[96];
  assign data_masked[12355] = data_i[12355] & sel_one_hot_i[96];
  assign data_masked[12354] = data_i[12354] & sel_one_hot_i[96];
  assign data_masked[12353] = data_i[12353] & sel_one_hot_i[96];
  assign data_masked[12352] = data_i[12352] & sel_one_hot_i[96];
  assign data_masked[12351] = data_i[12351] & sel_one_hot_i[96];
  assign data_masked[12350] = data_i[12350] & sel_one_hot_i[96];
  assign data_masked[12349] = data_i[12349] & sel_one_hot_i[96];
  assign data_masked[12348] = data_i[12348] & sel_one_hot_i[96];
  assign data_masked[12347] = data_i[12347] & sel_one_hot_i[96];
  assign data_masked[12346] = data_i[12346] & sel_one_hot_i[96];
  assign data_masked[12345] = data_i[12345] & sel_one_hot_i[96];
  assign data_masked[12344] = data_i[12344] & sel_one_hot_i[96];
  assign data_masked[12343] = data_i[12343] & sel_one_hot_i[96];
  assign data_masked[12342] = data_i[12342] & sel_one_hot_i[96];
  assign data_masked[12341] = data_i[12341] & sel_one_hot_i[96];
  assign data_masked[12340] = data_i[12340] & sel_one_hot_i[96];
  assign data_masked[12339] = data_i[12339] & sel_one_hot_i[96];
  assign data_masked[12338] = data_i[12338] & sel_one_hot_i[96];
  assign data_masked[12337] = data_i[12337] & sel_one_hot_i[96];
  assign data_masked[12336] = data_i[12336] & sel_one_hot_i[96];
  assign data_masked[12335] = data_i[12335] & sel_one_hot_i[96];
  assign data_masked[12334] = data_i[12334] & sel_one_hot_i[96];
  assign data_masked[12333] = data_i[12333] & sel_one_hot_i[96];
  assign data_masked[12332] = data_i[12332] & sel_one_hot_i[96];
  assign data_masked[12331] = data_i[12331] & sel_one_hot_i[96];
  assign data_masked[12330] = data_i[12330] & sel_one_hot_i[96];
  assign data_masked[12329] = data_i[12329] & sel_one_hot_i[96];
  assign data_masked[12328] = data_i[12328] & sel_one_hot_i[96];
  assign data_masked[12327] = data_i[12327] & sel_one_hot_i[96];
  assign data_masked[12326] = data_i[12326] & sel_one_hot_i[96];
  assign data_masked[12325] = data_i[12325] & sel_one_hot_i[96];
  assign data_masked[12324] = data_i[12324] & sel_one_hot_i[96];
  assign data_masked[12323] = data_i[12323] & sel_one_hot_i[96];
  assign data_masked[12322] = data_i[12322] & sel_one_hot_i[96];
  assign data_masked[12321] = data_i[12321] & sel_one_hot_i[96];
  assign data_masked[12320] = data_i[12320] & sel_one_hot_i[96];
  assign data_masked[12319] = data_i[12319] & sel_one_hot_i[96];
  assign data_masked[12318] = data_i[12318] & sel_one_hot_i[96];
  assign data_masked[12317] = data_i[12317] & sel_one_hot_i[96];
  assign data_masked[12316] = data_i[12316] & sel_one_hot_i[96];
  assign data_masked[12315] = data_i[12315] & sel_one_hot_i[96];
  assign data_masked[12314] = data_i[12314] & sel_one_hot_i[96];
  assign data_masked[12313] = data_i[12313] & sel_one_hot_i[96];
  assign data_masked[12312] = data_i[12312] & sel_one_hot_i[96];
  assign data_masked[12311] = data_i[12311] & sel_one_hot_i[96];
  assign data_masked[12310] = data_i[12310] & sel_one_hot_i[96];
  assign data_masked[12309] = data_i[12309] & sel_one_hot_i[96];
  assign data_masked[12308] = data_i[12308] & sel_one_hot_i[96];
  assign data_masked[12307] = data_i[12307] & sel_one_hot_i[96];
  assign data_masked[12306] = data_i[12306] & sel_one_hot_i[96];
  assign data_masked[12305] = data_i[12305] & sel_one_hot_i[96];
  assign data_masked[12304] = data_i[12304] & sel_one_hot_i[96];
  assign data_masked[12303] = data_i[12303] & sel_one_hot_i[96];
  assign data_masked[12302] = data_i[12302] & sel_one_hot_i[96];
  assign data_masked[12301] = data_i[12301] & sel_one_hot_i[96];
  assign data_masked[12300] = data_i[12300] & sel_one_hot_i[96];
  assign data_masked[12299] = data_i[12299] & sel_one_hot_i[96];
  assign data_masked[12298] = data_i[12298] & sel_one_hot_i[96];
  assign data_masked[12297] = data_i[12297] & sel_one_hot_i[96];
  assign data_masked[12296] = data_i[12296] & sel_one_hot_i[96];
  assign data_masked[12295] = data_i[12295] & sel_one_hot_i[96];
  assign data_masked[12294] = data_i[12294] & sel_one_hot_i[96];
  assign data_masked[12293] = data_i[12293] & sel_one_hot_i[96];
  assign data_masked[12292] = data_i[12292] & sel_one_hot_i[96];
  assign data_masked[12291] = data_i[12291] & sel_one_hot_i[96];
  assign data_masked[12290] = data_i[12290] & sel_one_hot_i[96];
  assign data_masked[12289] = data_i[12289] & sel_one_hot_i[96];
  assign data_masked[12288] = data_i[12288] & sel_one_hot_i[96];
  assign data_masked[12543] = data_i[12543] & sel_one_hot_i[97];
  assign data_masked[12542] = data_i[12542] & sel_one_hot_i[97];
  assign data_masked[12541] = data_i[12541] & sel_one_hot_i[97];
  assign data_masked[12540] = data_i[12540] & sel_one_hot_i[97];
  assign data_masked[12539] = data_i[12539] & sel_one_hot_i[97];
  assign data_masked[12538] = data_i[12538] & sel_one_hot_i[97];
  assign data_masked[12537] = data_i[12537] & sel_one_hot_i[97];
  assign data_masked[12536] = data_i[12536] & sel_one_hot_i[97];
  assign data_masked[12535] = data_i[12535] & sel_one_hot_i[97];
  assign data_masked[12534] = data_i[12534] & sel_one_hot_i[97];
  assign data_masked[12533] = data_i[12533] & sel_one_hot_i[97];
  assign data_masked[12532] = data_i[12532] & sel_one_hot_i[97];
  assign data_masked[12531] = data_i[12531] & sel_one_hot_i[97];
  assign data_masked[12530] = data_i[12530] & sel_one_hot_i[97];
  assign data_masked[12529] = data_i[12529] & sel_one_hot_i[97];
  assign data_masked[12528] = data_i[12528] & sel_one_hot_i[97];
  assign data_masked[12527] = data_i[12527] & sel_one_hot_i[97];
  assign data_masked[12526] = data_i[12526] & sel_one_hot_i[97];
  assign data_masked[12525] = data_i[12525] & sel_one_hot_i[97];
  assign data_masked[12524] = data_i[12524] & sel_one_hot_i[97];
  assign data_masked[12523] = data_i[12523] & sel_one_hot_i[97];
  assign data_masked[12522] = data_i[12522] & sel_one_hot_i[97];
  assign data_masked[12521] = data_i[12521] & sel_one_hot_i[97];
  assign data_masked[12520] = data_i[12520] & sel_one_hot_i[97];
  assign data_masked[12519] = data_i[12519] & sel_one_hot_i[97];
  assign data_masked[12518] = data_i[12518] & sel_one_hot_i[97];
  assign data_masked[12517] = data_i[12517] & sel_one_hot_i[97];
  assign data_masked[12516] = data_i[12516] & sel_one_hot_i[97];
  assign data_masked[12515] = data_i[12515] & sel_one_hot_i[97];
  assign data_masked[12514] = data_i[12514] & sel_one_hot_i[97];
  assign data_masked[12513] = data_i[12513] & sel_one_hot_i[97];
  assign data_masked[12512] = data_i[12512] & sel_one_hot_i[97];
  assign data_masked[12511] = data_i[12511] & sel_one_hot_i[97];
  assign data_masked[12510] = data_i[12510] & sel_one_hot_i[97];
  assign data_masked[12509] = data_i[12509] & sel_one_hot_i[97];
  assign data_masked[12508] = data_i[12508] & sel_one_hot_i[97];
  assign data_masked[12507] = data_i[12507] & sel_one_hot_i[97];
  assign data_masked[12506] = data_i[12506] & sel_one_hot_i[97];
  assign data_masked[12505] = data_i[12505] & sel_one_hot_i[97];
  assign data_masked[12504] = data_i[12504] & sel_one_hot_i[97];
  assign data_masked[12503] = data_i[12503] & sel_one_hot_i[97];
  assign data_masked[12502] = data_i[12502] & sel_one_hot_i[97];
  assign data_masked[12501] = data_i[12501] & sel_one_hot_i[97];
  assign data_masked[12500] = data_i[12500] & sel_one_hot_i[97];
  assign data_masked[12499] = data_i[12499] & sel_one_hot_i[97];
  assign data_masked[12498] = data_i[12498] & sel_one_hot_i[97];
  assign data_masked[12497] = data_i[12497] & sel_one_hot_i[97];
  assign data_masked[12496] = data_i[12496] & sel_one_hot_i[97];
  assign data_masked[12495] = data_i[12495] & sel_one_hot_i[97];
  assign data_masked[12494] = data_i[12494] & sel_one_hot_i[97];
  assign data_masked[12493] = data_i[12493] & sel_one_hot_i[97];
  assign data_masked[12492] = data_i[12492] & sel_one_hot_i[97];
  assign data_masked[12491] = data_i[12491] & sel_one_hot_i[97];
  assign data_masked[12490] = data_i[12490] & sel_one_hot_i[97];
  assign data_masked[12489] = data_i[12489] & sel_one_hot_i[97];
  assign data_masked[12488] = data_i[12488] & sel_one_hot_i[97];
  assign data_masked[12487] = data_i[12487] & sel_one_hot_i[97];
  assign data_masked[12486] = data_i[12486] & sel_one_hot_i[97];
  assign data_masked[12485] = data_i[12485] & sel_one_hot_i[97];
  assign data_masked[12484] = data_i[12484] & sel_one_hot_i[97];
  assign data_masked[12483] = data_i[12483] & sel_one_hot_i[97];
  assign data_masked[12482] = data_i[12482] & sel_one_hot_i[97];
  assign data_masked[12481] = data_i[12481] & sel_one_hot_i[97];
  assign data_masked[12480] = data_i[12480] & sel_one_hot_i[97];
  assign data_masked[12479] = data_i[12479] & sel_one_hot_i[97];
  assign data_masked[12478] = data_i[12478] & sel_one_hot_i[97];
  assign data_masked[12477] = data_i[12477] & sel_one_hot_i[97];
  assign data_masked[12476] = data_i[12476] & sel_one_hot_i[97];
  assign data_masked[12475] = data_i[12475] & sel_one_hot_i[97];
  assign data_masked[12474] = data_i[12474] & sel_one_hot_i[97];
  assign data_masked[12473] = data_i[12473] & sel_one_hot_i[97];
  assign data_masked[12472] = data_i[12472] & sel_one_hot_i[97];
  assign data_masked[12471] = data_i[12471] & sel_one_hot_i[97];
  assign data_masked[12470] = data_i[12470] & sel_one_hot_i[97];
  assign data_masked[12469] = data_i[12469] & sel_one_hot_i[97];
  assign data_masked[12468] = data_i[12468] & sel_one_hot_i[97];
  assign data_masked[12467] = data_i[12467] & sel_one_hot_i[97];
  assign data_masked[12466] = data_i[12466] & sel_one_hot_i[97];
  assign data_masked[12465] = data_i[12465] & sel_one_hot_i[97];
  assign data_masked[12464] = data_i[12464] & sel_one_hot_i[97];
  assign data_masked[12463] = data_i[12463] & sel_one_hot_i[97];
  assign data_masked[12462] = data_i[12462] & sel_one_hot_i[97];
  assign data_masked[12461] = data_i[12461] & sel_one_hot_i[97];
  assign data_masked[12460] = data_i[12460] & sel_one_hot_i[97];
  assign data_masked[12459] = data_i[12459] & sel_one_hot_i[97];
  assign data_masked[12458] = data_i[12458] & sel_one_hot_i[97];
  assign data_masked[12457] = data_i[12457] & sel_one_hot_i[97];
  assign data_masked[12456] = data_i[12456] & sel_one_hot_i[97];
  assign data_masked[12455] = data_i[12455] & sel_one_hot_i[97];
  assign data_masked[12454] = data_i[12454] & sel_one_hot_i[97];
  assign data_masked[12453] = data_i[12453] & sel_one_hot_i[97];
  assign data_masked[12452] = data_i[12452] & sel_one_hot_i[97];
  assign data_masked[12451] = data_i[12451] & sel_one_hot_i[97];
  assign data_masked[12450] = data_i[12450] & sel_one_hot_i[97];
  assign data_masked[12449] = data_i[12449] & sel_one_hot_i[97];
  assign data_masked[12448] = data_i[12448] & sel_one_hot_i[97];
  assign data_masked[12447] = data_i[12447] & sel_one_hot_i[97];
  assign data_masked[12446] = data_i[12446] & sel_one_hot_i[97];
  assign data_masked[12445] = data_i[12445] & sel_one_hot_i[97];
  assign data_masked[12444] = data_i[12444] & sel_one_hot_i[97];
  assign data_masked[12443] = data_i[12443] & sel_one_hot_i[97];
  assign data_masked[12442] = data_i[12442] & sel_one_hot_i[97];
  assign data_masked[12441] = data_i[12441] & sel_one_hot_i[97];
  assign data_masked[12440] = data_i[12440] & sel_one_hot_i[97];
  assign data_masked[12439] = data_i[12439] & sel_one_hot_i[97];
  assign data_masked[12438] = data_i[12438] & sel_one_hot_i[97];
  assign data_masked[12437] = data_i[12437] & sel_one_hot_i[97];
  assign data_masked[12436] = data_i[12436] & sel_one_hot_i[97];
  assign data_masked[12435] = data_i[12435] & sel_one_hot_i[97];
  assign data_masked[12434] = data_i[12434] & sel_one_hot_i[97];
  assign data_masked[12433] = data_i[12433] & sel_one_hot_i[97];
  assign data_masked[12432] = data_i[12432] & sel_one_hot_i[97];
  assign data_masked[12431] = data_i[12431] & sel_one_hot_i[97];
  assign data_masked[12430] = data_i[12430] & sel_one_hot_i[97];
  assign data_masked[12429] = data_i[12429] & sel_one_hot_i[97];
  assign data_masked[12428] = data_i[12428] & sel_one_hot_i[97];
  assign data_masked[12427] = data_i[12427] & sel_one_hot_i[97];
  assign data_masked[12426] = data_i[12426] & sel_one_hot_i[97];
  assign data_masked[12425] = data_i[12425] & sel_one_hot_i[97];
  assign data_masked[12424] = data_i[12424] & sel_one_hot_i[97];
  assign data_masked[12423] = data_i[12423] & sel_one_hot_i[97];
  assign data_masked[12422] = data_i[12422] & sel_one_hot_i[97];
  assign data_masked[12421] = data_i[12421] & sel_one_hot_i[97];
  assign data_masked[12420] = data_i[12420] & sel_one_hot_i[97];
  assign data_masked[12419] = data_i[12419] & sel_one_hot_i[97];
  assign data_masked[12418] = data_i[12418] & sel_one_hot_i[97];
  assign data_masked[12417] = data_i[12417] & sel_one_hot_i[97];
  assign data_masked[12416] = data_i[12416] & sel_one_hot_i[97];
  assign data_masked[12671] = data_i[12671] & sel_one_hot_i[98];
  assign data_masked[12670] = data_i[12670] & sel_one_hot_i[98];
  assign data_masked[12669] = data_i[12669] & sel_one_hot_i[98];
  assign data_masked[12668] = data_i[12668] & sel_one_hot_i[98];
  assign data_masked[12667] = data_i[12667] & sel_one_hot_i[98];
  assign data_masked[12666] = data_i[12666] & sel_one_hot_i[98];
  assign data_masked[12665] = data_i[12665] & sel_one_hot_i[98];
  assign data_masked[12664] = data_i[12664] & sel_one_hot_i[98];
  assign data_masked[12663] = data_i[12663] & sel_one_hot_i[98];
  assign data_masked[12662] = data_i[12662] & sel_one_hot_i[98];
  assign data_masked[12661] = data_i[12661] & sel_one_hot_i[98];
  assign data_masked[12660] = data_i[12660] & sel_one_hot_i[98];
  assign data_masked[12659] = data_i[12659] & sel_one_hot_i[98];
  assign data_masked[12658] = data_i[12658] & sel_one_hot_i[98];
  assign data_masked[12657] = data_i[12657] & sel_one_hot_i[98];
  assign data_masked[12656] = data_i[12656] & sel_one_hot_i[98];
  assign data_masked[12655] = data_i[12655] & sel_one_hot_i[98];
  assign data_masked[12654] = data_i[12654] & sel_one_hot_i[98];
  assign data_masked[12653] = data_i[12653] & sel_one_hot_i[98];
  assign data_masked[12652] = data_i[12652] & sel_one_hot_i[98];
  assign data_masked[12651] = data_i[12651] & sel_one_hot_i[98];
  assign data_masked[12650] = data_i[12650] & sel_one_hot_i[98];
  assign data_masked[12649] = data_i[12649] & sel_one_hot_i[98];
  assign data_masked[12648] = data_i[12648] & sel_one_hot_i[98];
  assign data_masked[12647] = data_i[12647] & sel_one_hot_i[98];
  assign data_masked[12646] = data_i[12646] & sel_one_hot_i[98];
  assign data_masked[12645] = data_i[12645] & sel_one_hot_i[98];
  assign data_masked[12644] = data_i[12644] & sel_one_hot_i[98];
  assign data_masked[12643] = data_i[12643] & sel_one_hot_i[98];
  assign data_masked[12642] = data_i[12642] & sel_one_hot_i[98];
  assign data_masked[12641] = data_i[12641] & sel_one_hot_i[98];
  assign data_masked[12640] = data_i[12640] & sel_one_hot_i[98];
  assign data_masked[12639] = data_i[12639] & sel_one_hot_i[98];
  assign data_masked[12638] = data_i[12638] & sel_one_hot_i[98];
  assign data_masked[12637] = data_i[12637] & sel_one_hot_i[98];
  assign data_masked[12636] = data_i[12636] & sel_one_hot_i[98];
  assign data_masked[12635] = data_i[12635] & sel_one_hot_i[98];
  assign data_masked[12634] = data_i[12634] & sel_one_hot_i[98];
  assign data_masked[12633] = data_i[12633] & sel_one_hot_i[98];
  assign data_masked[12632] = data_i[12632] & sel_one_hot_i[98];
  assign data_masked[12631] = data_i[12631] & sel_one_hot_i[98];
  assign data_masked[12630] = data_i[12630] & sel_one_hot_i[98];
  assign data_masked[12629] = data_i[12629] & sel_one_hot_i[98];
  assign data_masked[12628] = data_i[12628] & sel_one_hot_i[98];
  assign data_masked[12627] = data_i[12627] & sel_one_hot_i[98];
  assign data_masked[12626] = data_i[12626] & sel_one_hot_i[98];
  assign data_masked[12625] = data_i[12625] & sel_one_hot_i[98];
  assign data_masked[12624] = data_i[12624] & sel_one_hot_i[98];
  assign data_masked[12623] = data_i[12623] & sel_one_hot_i[98];
  assign data_masked[12622] = data_i[12622] & sel_one_hot_i[98];
  assign data_masked[12621] = data_i[12621] & sel_one_hot_i[98];
  assign data_masked[12620] = data_i[12620] & sel_one_hot_i[98];
  assign data_masked[12619] = data_i[12619] & sel_one_hot_i[98];
  assign data_masked[12618] = data_i[12618] & sel_one_hot_i[98];
  assign data_masked[12617] = data_i[12617] & sel_one_hot_i[98];
  assign data_masked[12616] = data_i[12616] & sel_one_hot_i[98];
  assign data_masked[12615] = data_i[12615] & sel_one_hot_i[98];
  assign data_masked[12614] = data_i[12614] & sel_one_hot_i[98];
  assign data_masked[12613] = data_i[12613] & sel_one_hot_i[98];
  assign data_masked[12612] = data_i[12612] & sel_one_hot_i[98];
  assign data_masked[12611] = data_i[12611] & sel_one_hot_i[98];
  assign data_masked[12610] = data_i[12610] & sel_one_hot_i[98];
  assign data_masked[12609] = data_i[12609] & sel_one_hot_i[98];
  assign data_masked[12608] = data_i[12608] & sel_one_hot_i[98];
  assign data_masked[12607] = data_i[12607] & sel_one_hot_i[98];
  assign data_masked[12606] = data_i[12606] & sel_one_hot_i[98];
  assign data_masked[12605] = data_i[12605] & sel_one_hot_i[98];
  assign data_masked[12604] = data_i[12604] & sel_one_hot_i[98];
  assign data_masked[12603] = data_i[12603] & sel_one_hot_i[98];
  assign data_masked[12602] = data_i[12602] & sel_one_hot_i[98];
  assign data_masked[12601] = data_i[12601] & sel_one_hot_i[98];
  assign data_masked[12600] = data_i[12600] & sel_one_hot_i[98];
  assign data_masked[12599] = data_i[12599] & sel_one_hot_i[98];
  assign data_masked[12598] = data_i[12598] & sel_one_hot_i[98];
  assign data_masked[12597] = data_i[12597] & sel_one_hot_i[98];
  assign data_masked[12596] = data_i[12596] & sel_one_hot_i[98];
  assign data_masked[12595] = data_i[12595] & sel_one_hot_i[98];
  assign data_masked[12594] = data_i[12594] & sel_one_hot_i[98];
  assign data_masked[12593] = data_i[12593] & sel_one_hot_i[98];
  assign data_masked[12592] = data_i[12592] & sel_one_hot_i[98];
  assign data_masked[12591] = data_i[12591] & sel_one_hot_i[98];
  assign data_masked[12590] = data_i[12590] & sel_one_hot_i[98];
  assign data_masked[12589] = data_i[12589] & sel_one_hot_i[98];
  assign data_masked[12588] = data_i[12588] & sel_one_hot_i[98];
  assign data_masked[12587] = data_i[12587] & sel_one_hot_i[98];
  assign data_masked[12586] = data_i[12586] & sel_one_hot_i[98];
  assign data_masked[12585] = data_i[12585] & sel_one_hot_i[98];
  assign data_masked[12584] = data_i[12584] & sel_one_hot_i[98];
  assign data_masked[12583] = data_i[12583] & sel_one_hot_i[98];
  assign data_masked[12582] = data_i[12582] & sel_one_hot_i[98];
  assign data_masked[12581] = data_i[12581] & sel_one_hot_i[98];
  assign data_masked[12580] = data_i[12580] & sel_one_hot_i[98];
  assign data_masked[12579] = data_i[12579] & sel_one_hot_i[98];
  assign data_masked[12578] = data_i[12578] & sel_one_hot_i[98];
  assign data_masked[12577] = data_i[12577] & sel_one_hot_i[98];
  assign data_masked[12576] = data_i[12576] & sel_one_hot_i[98];
  assign data_masked[12575] = data_i[12575] & sel_one_hot_i[98];
  assign data_masked[12574] = data_i[12574] & sel_one_hot_i[98];
  assign data_masked[12573] = data_i[12573] & sel_one_hot_i[98];
  assign data_masked[12572] = data_i[12572] & sel_one_hot_i[98];
  assign data_masked[12571] = data_i[12571] & sel_one_hot_i[98];
  assign data_masked[12570] = data_i[12570] & sel_one_hot_i[98];
  assign data_masked[12569] = data_i[12569] & sel_one_hot_i[98];
  assign data_masked[12568] = data_i[12568] & sel_one_hot_i[98];
  assign data_masked[12567] = data_i[12567] & sel_one_hot_i[98];
  assign data_masked[12566] = data_i[12566] & sel_one_hot_i[98];
  assign data_masked[12565] = data_i[12565] & sel_one_hot_i[98];
  assign data_masked[12564] = data_i[12564] & sel_one_hot_i[98];
  assign data_masked[12563] = data_i[12563] & sel_one_hot_i[98];
  assign data_masked[12562] = data_i[12562] & sel_one_hot_i[98];
  assign data_masked[12561] = data_i[12561] & sel_one_hot_i[98];
  assign data_masked[12560] = data_i[12560] & sel_one_hot_i[98];
  assign data_masked[12559] = data_i[12559] & sel_one_hot_i[98];
  assign data_masked[12558] = data_i[12558] & sel_one_hot_i[98];
  assign data_masked[12557] = data_i[12557] & sel_one_hot_i[98];
  assign data_masked[12556] = data_i[12556] & sel_one_hot_i[98];
  assign data_masked[12555] = data_i[12555] & sel_one_hot_i[98];
  assign data_masked[12554] = data_i[12554] & sel_one_hot_i[98];
  assign data_masked[12553] = data_i[12553] & sel_one_hot_i[98];
  assign data_masked[12552] = data_i[12552] & sel_one_hot_i[98];
  assign data_masked[12551] = data_i[12551] & sel_one_hot_i[98];
  assign data_masked[12550] = data_i[12550] & sel_one_hot_i[98];
  assign data_masked[12549] = data_i[12549] & sel_one_hot_i[98];
  assign data_masked[12548] = data_i[12548] & sel_one_hot_i[98];
  assign data_masked[12547] = data_i[12547] & sel_one_hot_i[98];
  assign data_masked[12546] = data_i[12546] & sel_one_hot_i[98];
  assign data_masked[12545] = data_i[12545] & sel_one_hot_i[98];
  assign data_masked[12544] = data_i[12544] & sel_one_hot_i[98];
  assign data_masked[12799] = data_i[12799] & sel_one_hot_i[99];
  assign data_masked[12798] = data_i[12798] & sel_one_hot_i[99];
  assign data_masked[12797] = data_i[12797] & sel_one_hot_i[99];
  assign data_masked[12796] = data_i[12796] & sel_one_hot_i[99];
  assign data_masked[12795] = data_i[12795] & sel_one_hot_i[99];
  assign data_masked[12794] = data_i[12794] & sel_one_hot_i[99];
  assign data_masked[12793] = data_i[12793] & sel_one_hot_i[99];
  assign data_masked[12792] = data_i[12792] & sel_one_hot_i[99];
  assign data_masked[12791] = data_i[12791] & sel_one_hot_i[99];
  assign data_masked[12790] = data_i[12790] & sel_one_hot_i[99];
  assign data_masked[12789] = data_i[12789] & sel_one_hot_i[99];
  assign data_masked[12788] = data_i[12788] & sel_one_hot_i[99];
  assign data_masked[12787] = data_i[12787] & sel_one_hot_i[99];
  assign data_masked[12786] = data_i[12786] & sel_one_hot_i[99];
  assign data_masked[12785] = data_i[12785] & sel_one_hot_i[99];
  assign data_masked[12784] = data_i[12784] & sel_one_hot_i[99];
  assign data_masked[12783] = data_i[12783] & sel_one_hot_i[99];
  assign data_masked[12782] = data_i[12782] & sel_one_hot_i[99];
  assign data_masked[12781] = data_i[12781] & sel_one_hot_i[99];
  assign data_masked[12780] = data_i[12780] & sel_one_hot_i[99];
  assign data_masked[12779] = data_i[12779] & sel_one_hot_i[99];
  assign data_masked[12778] = data_i[12778] & sel_one_hot_i[99];
  assign data_masked[12777] = data_i[12777] & sel_one_hot_i[99];
  assign data_masked[12776] = data_i[12776] & sel_one_hot_i[99];
  assign data_masked[12775] = data_i[12775] & sel_one_hot_i[99];
  assign data_masked[12774] = data_i[12774] & sel_one_hot_i[99];
  assign data_masked[12773] = data_i[12773] & sel_one_hot_i[99];
  assign data_masked[12772] = data_i[12772] & sel_one_hot_i[99];
  assign data_masked[12771] = data_i[12771] & sel_one_hot_i[99];
  assign data_masked[12770] = data_i[12770] & sel_one_hot_i[99];
  assign data_masked[12769] = data_i[12769] & sel_one_hot_i[99];
  assign data_masked[12768] = data_i[12768] & sel_one_hot_i[99];
  assign data_masked[12767] = data_i[12767] & sel_one_hot_i[99];
  assign data_masked[12766] = data_i[12766] & sel_one_hot_i[99];
  assign data_masked[12765] = data_i[12765] & sel_one_hot_i[99];
  assign data_masked[12764] = data_i[12764] & sel_one_hot_i[99];
  assign data_masked[12763] = data_i[12763] & sel_one_hot_i[99];
  assign data_masked[12762] = data_i[12762] & sel_one_hot_i[99];
  assign data_masked[12761] = data_i[12761] & sel_one_hot_i[99];
  assign data_masked[12760] = data_i[12760] & sel_one_hot_i[99];
  assign data_masked[12759] = data_i[12759] & sel_one_hot_i[99];
  assign data_masked[12758] = data_i[12758] & sel_one_hot_i[99];
  assign data_masked[12757] = data_i[12757] & sel_one_hot_i[99];
  assign data_masked[12756] = data_i[12756] & sel_one_hot_i[99];
  assign data_masked[12755] = data_i[12755] & sel_one_hot_i[99];
  assign data_masked[12754] = data_i[12754] & sel_one_hot_i[99];
  assign data_masked[12753] = data_i[12753] & sel_one_hot_i[99];
  assign data_masked[12752] = data_i[12752] & sel_one_hot_i[99];
  assign data_masked[12751] = data_i[12751] & sel_one_hot_i[99];
  assign data_masked[12750] = data_i[12750] & sel_one_hot_i[99];
  assign data_masked[12749] = data_i[12749] & sel_one_hot_i[99];
  assign data_masked[12748] = data_i[12748] & sel_one_hot_i[99];
  assign data_masked[12747] = data_i[12747] & sel_one_hot_i[99];
  assign data_masked[12746] = data_i[12746] & sel_one_hot_i[99];
  assign data_masked[12745] = data_i[12745] & sel_one_hot_i[99];
  assign data_masked[12744] = data_i[12744] & sel_one_hot_i[99];
  assign data_masked[12743] = data_i[12743] & sel_one_hot_i[99];
  assign data_masked[12742] = data_i[12742] & sel_one_hot_i[99];
  assign data_masked[12741] = data_i[12741] & sel_one_hot_i[99];
  assign data_masked[12740] = data_i[12740] & sel_one_hot_i[99];
  assign data_masked[12739] = data_i[12739] & sel_one_hot_i[99];
  assign data_masked[12738] = data_i[12738] & sel_one_hot_i[99];
  assign data_masked[12737] = data_i[12737] & sel_one_hot_i[99];
  assign data_masked[12736] = data_i[12736] & sel_one_hot_i[99];
  assign data_masked[12735] = data_i[12735] & sel_one_hot_i[99];
  assign data_masked[12734] = data_i[12734] & sel_one_hot_i[99];
  assign data_masked[12733] = data_i[12733] & sel_one_hot_i[99];
  assign data_masked[12732] = data_i[12732] & sel_one_hot_i[99];
  assign data_masked[12731] = data_i[12731] & sel_one_hot_i[99];
  assign data_masked[12730] = data_i[12730] & sel_one_hot_i[99];
  assign data_masked[12729] = data_i[12729] & sel_one_hot_i[99];
  assign data_masked[12728] = data_i[12728] & sel_one_hot_i[99];
  assign data_masked[12727] = data_i[12727] & sel_one_hot_i[99];
  assign data_masked[12726] = data_i[12726] & sel_one_hot_i[99];
  assign data_masked[12725] = data_i[12725] & sel_one_hot_i[99];
  assign data_masked[12724] = data_i[12724] & sel_one_hot_i[99];
  assign data_masked[12723] = data_i[12723] & sel_one_hot_i[99];
  assign data_masked[12722] = data_i[12722] & sel_one_hot_i[99];
  assign data_masked[12721] = data_i[12721] & sel_one_hot_i[99];
  assign data_masked[12720] = data_i[12720] & sel_one_hot_i[99];
  assign data_masked[12719] = data_i[12719] & sel_one_hot_i[99];
  assign data_masked[12718] = data_i[12718] & sel_one_hot_i[99];
  assign data_masked[12717] = data_i[12717] & sel_one_hot_i[99];
  assign data_masked[12716] = data_i[12716] & sel_one_hot_i[99];
  assign data_masked[12715] = data_i[12715] & sel_one_hot_i[99];
  assign data_masked[12714] = data_i[12714] & sel_one_hot_i[99];
  assign data_masked[12713] = data_i[12713] & sel_one_hot_i[99];
  assign data_masked[12712] = data_i[12712] & sel_one_hot_i[99];
  assign data_masked[12711] = data_i[12711] & sel_one_hot_i[99];
  assign data_masked[12710] = data_i[12710] & sel_one_hot_i[99];
  assign data_masked[12709] = data_i[12709] & sel_one_hot_i[99];
  assign data_masked[12708] = data_i[12708] & sel_one_hot_i[99];
  assign data_masked[12707] = data_i[12707] & sel_one_hot_i[99];
  assign data_masked[12706] = data_i[12706] & sel_one_hot_i[99];
  assign data_masked[12705] = data_i[12705] & sel_one_hot_i[99];
  assign data_masked[12704] = data_i[12704] & sel_one_hot_i[99];
  assign data_masked[12703] = data_i[12703] & sel_one_hot_i[99];
  assign data_masked[12702] = data_i[12702] & sel_one_hot_i[99];
  assign data_masked[12701] = data_i[12701] & sel_one_hot_i[99];
  assign data_masked[12700] = data_i[12700] & sel_one_hot_i[99];
  assign data_masked[12699] = data_i[12699] & sel_one_hot_i[99];
  assign data_masked[12698] = data_i[12698] & sel_one_hot_i[99];
  assign data_masked[12697] = data_i[12697] & sel_one_hot_i[99];
  assign data_masked[12696] = data_i[12696] & sel_one_hot_i[99];
  assign data_masked[12695] = data_i[12695] & sel_one_hot_i[99];
  assign data_masked[12694] = data_i[12694] & sel_one_hot_i[99];
  assign data_masked[12693] = data_i[12693] & sel_one_hot_i[99];
  assign data_masked[12692] = data_i[12692] & sel_one_hot_i[99];
  assign data_masked[12691] = data_i[12691] & sel_one_hot_i[99];
  assign data_masked[12690] = data_i[12690] & sel_one_hot_i[99];
  assign data_masked[12689] = data_i[12689] & sel_one_hot_i[99];
  assign data_masked[12688] = data_i[12688] & sel_one_hot_i[99];
  assign data_masked[12687] = data_i[12687] & sel_one_hot_i[99];
  assign data_masked[12686] = data_i[12686] & sel_one_hot_i[99];
  assign data_masked[12685] = data_i[12685] & sel_one_hot_i[99];
  assign data_masked[12684] = data_i[12684] & sel_one_hot_i[99];
  assign data_masked[12683] = data_i[12683] & sel_one_hot_i[99];
  assign data_masked[12682] = data_i[12682] & sel_one_hot_i[99];
  assign data_masked[12681] = data_i[12681] & sel_one_hot_i[99];
  assign data_masked[12680] = data_i[12680] & sel_one_hot_i[99];
  assign data_masked[12679] = data_i[12679] & sel_one_hot_i[99];
  assign data_masked[12678] = data_i[12678] & sel_one_hot_i[99];
  assign data_masked[12677] = data_i[12677] & sel_one_hot_i[99];
  assign data_masked[12676] = data_i[12676] & sel_one_hot_i[99];
  assign data_masked[12675] = data_i[12675] & sel_one_hot_i[99];
  assign data_masked[12674] = data_i[12674] & sel_one_hot_i[99];
  assign data_masked[12673] = data_i[12673] & sel_one_hot_i[99];
  assign data_masked[12672] = data_i[12672] & sel_one_hot_i[99];
  assign data_masked[12927] = data_i[12927] & sel_one_hot_i[100];
  assign data_masked[12926] = data_i[12926] & sel_one_hot_i[100];
  assign data_masked[12925] = data_i[12925] & sel_one_hot_i[100];
  assign data_masked[12924] = data_i[12924] & sel_one_hot_i[100];
  assign data_masked[12923] = data_i[12923] & sel_one_hot_i[100];
  assign data_masked[12922] = data_i[12922] & sel_one_hot_i[100];
  assign data_masked[12921] = data_i[12921] & sel_one_hot_i[100];
  assign data_masked[12920] = data_i[12920] & sel_one_hot_i[100];
  assign data_masked[12919] = data_i[12919] & sel_one_hot_i[100];
  assign data_masked[12918] = data_i[12918] & sel_one_hot_i[100];
  assign data_masked[12917] = data_i[12917] & sel_one_hot_i[100];
  assign data_masked[12916] = data_i[12916] & sel_one_hot_i[100];
  assign data_masked[12915] = data_i[12915] & sel_one_hot_i[100];
  assign data_masked[12914] = data_i[12914] & sel_one_hot_i[100];
  assign data_masked[12913] = data_i[12913] & sel_one_hot_i[100];
  assign data_masked[12912] = data_i[12912] & sel_one_hot_i[100];
  assign data_masked[12911] = data_i[12911] & sel_one_hot_i[100];
  assign data_masked[12910] = data_i[12910] & sel_one_hot_i[100];
  assign data_masked[12909] = data_i[12909] & sel_one_hot_i[100];
  assign data_masked[12908] = data_i[12908] & sel_one_hot_i[100];
  assign data_masked[12907] = data_i[12907] & sel_one_hot_i[100];
  assign data_masked[12906] = data_i[12906] & sel_one_hot_i[100];
  assign data_masked[12905] = data_i[12905] & sel_one_hot_i[100];
  assign data_masked[12904] = data_i[12904] & sel_one_hot_i[100];
  assign data_masked[12903] = data_i[12903] & sel_one_hot_i[100];
  assign data_masked[12902] = data_i[12902] & sel_one_hot_i[100];
  assign data_masked[12901] = data_i[12901] & sel_one_hot_i[100];
  assign data_masked[12900] = data_i[12900] & sel_one_hot_i[100];
  assign data_masked[12899] = data_i[12899] & sel_one_hot_i[100];
  assign data_masked[12898] = data_i[12898] & sel_one_hot_i[100];
  assign data_masked[12897] = data_i[12897] & sel_one_hot_i[100];
  assign data_masked[12896] = data_i[12896] & sel_one_hot_i[100];
  assign data_masked[12895] = data_i[12895] & sel_one_hot_i[100];
  assign data_masked[12894] = data_i[12894] & sel_one_hot_i[100];
  assign data_masked[12893] = data_i[12893] & sel_one_hot_i[100];
  assign data_masked[12892] = data_i[12892] & sel_one_hot_i[100];
  assign data_masked[12891] = data_i[12891] & sel_one_hot_i[100];
  assign data_masked[12890] = data_i[12890] & sel_one_hot_i[100];
  assign data_masked[12889] = data_i[12889] & sel_one_hot_i[100];
  assign data_masked[12888] = data_i[12888] & sel_one_hot_i[100];
  assign data_masked[12887] = data_i[12887] & sel_one_hot_i[100];
  assign data_masked[12886] = data_i[12886] & sel_one_hot_i[100];
  assign data_masked[12885] = data_i[12885] & sel_one_hot_i[100];
  assign data_masked[12884] = data_i[12884] & sel_one_hot_i[100];
  assign data_masked[12883] = data_i[12883] & sel_one_hot_i[100];
  assign data_masked[12882] = data_i[12882] & sel_one_hot_i[100];
  assign data_masked[12881] = data_i[12881] & sel_one_hot_i[100];
  assign data_masked[12880] = data_i[12880] & sel_one_hot_i[100];
  assign data_masked[12879] = data_i[12879] & sel_one_hot_i[100];
  assign data_masked[12878] = data_i[12878] & sel_one_hot_i[100];
  assign data_masked[12877] = data_i[12877] & sel_one_hot_i[100];
  assign data_masked[12876] = data_i[12876] & sel_one_hot_i[100];
  assign data_masked[12875] = data_i[12875] & sel_one_hot_i[100];
  assign data_masked[12874] = data_i[12874] & sel_one_hot_i[100];
  assign data_masked[12873] = data_i[12873] & sel_one_hot_i[100];
  assign data_masked[12872] = data_i[12872] & sel_one_hot_i[100];
  assign data_masked[12871] = data_i[12871] & sel_one_hot_i[100];
  assign data_masked[12870] = data_i[12870] & sel_one_hot_i[100];
  assign data_masked[12869] = data_i[12869] & sel_one_hot_i[100];
  assign data_masked[12868] = data_i[12868] & sel_one_hot_i[100];
  assign data_masked[12867] = data_i[12867] & sel_one_hot_i[100];
  assign data_masked[12866] = data_i[12866] & sel_one_hot_i[100];
  assign data_masked[12865] = data_i[12865] & sel_one_hot_i[100];
  assign data_masked[12864] = data_i[12864] & sel_one_hot_i[100];
  assign data_masked[12863] = data_i[12863] & sel_one_hot_i[100];
  assign data_masked[12862] = data_i[12862] & sel_one_hot_i[100];
  assign data_masked[12861] = data_i[12861] & sel_one_hot_i[100];
  assign data_masked[12860] = data_i[12860] & sel_one_hot_i[100];
  assign data_masked[12859] = data_i[12859] & sel_one_hot_i[100];
  assign data_masked[12858] = data_i[12858] & sel_one_hot_i[100];
  assign data_masked[12857] = data_i[12857] & sel_one_hot_i[100];
  assign data_masked[12856] = data_i[12856] & sel_one_hot_i[100];
  assign data_masked[12855] = data_i[12855] & sel_one_hot_i[100];
  assign data_masked[12854] = data_i[12854] & sel_one_hot_i[100];
  assign data_masked[12853] = data_i[12853] & sel_one_hot_i[100];
  assign data_masked[12852] = data_i[12852] & sel_one_hot_i[100];
  assign data_masked[12851] = data_i[12851] & sel_one_hot_i[100];
  assign data_masked[12850] = data_i[12850] & sel_one_hot_i[100];
  assign data_masked[12849] = data_i[12849] & sel_one_hot_i[100];
  assign data_masked[12848] = data_i[12848] & sel_one_hot_i[100];
  assign data_masked[12847] = data_i[12847] & sel_one_hot_i[100];
  assign data_masked[12846] = data_i[12846] & sel_one_hot_i[100];
  assign data_masked[12845] = data_i[12845] & sel_one_hot_i[100];
  assign data_masked[12844] = data_i[12844] & sel_one_hot_i[100];
  assign data_masked[12843] = data_i[12843] & sel_one_hot_i[100];
  assign data_masked[12842] = data_i[12842] & sel_one_hot_i[100];
  assign data_masked[12841] = data_i[12841] & sel_one_hot_i[100];
  assign data_masked[12840] = data_i[12840] & sel_one_hot_i[100];
  assign data_masked[12839] = data_i[12839] & sel_one_hot_i[100];
  assign data_masked[12838] = data_i[12838] & sel_one_hot_i[100];
  assign data_masked[12837] = data_i[12837] & sel_one_hot_i[100];
  assign data_masked[12836] = data_i[12836] & sel_one_hot_i[100];
  assign data_masked[12835] = data_i[12835] & sel_one_hot_i[100];
  assign data_masked[12834] = data_i[12834] & sel_one_hot_i[100];
  assign data_masked[12833] = data_i[12833] & sel_one_hot_i[100];
  assign data_masked[12832] = data_i[12832] & sel_one_hot_i[100];
  assign data_masked[12831] = data_i[12831] & sel_one_hot_i[100];
  assign data_masked[12830] = data_i[12830] & sel_one_hot_i[100];
  assign data_masked[12829] = data_i[12829] & sel_one_hot_i[100];
  assign data_masked[12828] = data_i[12828] & sel_one_hot_i[100];
  assign data_masked[12827] = data_i[12827] & sel_one_hot_i[100];
  assign data_masked[12826] = data_i[12826] & sel_one_hot_i[100];
  assign data_masked[12825] = data_i[12825] & sel_one_hot_i[100];
  assign data_masked[12824] = data_i[12824] & sel_one_hot_i[100];
  assign data_masked[12823] = data_i[12823] & sel_one_hot_i[100];
  assign data_masked[12822] = data_i[12822] & sel_one_hot_i[100];
  assign data_masked[12821] = data_i[12821] & sel_one_hot_i[100];
  assign data_masked[12820] = data_i[12820] & sel_one_hot_i[100];
  assign data_masked[12819] = data_i[12819] & sel_one_hot_i[100];
  assign data_masked[12818] = data_i[12818] & sel_one_hot_i[100];
  assign data_masked[12817] = data_i[12817] & sel_one_hot_i[100];
  assign data_masked[12816] = data_i[12816] & sel_one_hot_i[100];
  assign data_masked[12815] = data_i[12815] & sel_one_hot_i[100];
  assign data_masked[12814] = data_i[12814] & sel_one_hot_i[100];
  assign data_masked[12813] = data_i[12813] & sel_one_hot_i[100];
  assign data_masked[12812] = data_i[12812] & sel_one_hot_i[100];
  assign data_masked[12811] = data_i[12811] & sel_one_hot_i[100];
  assign data_masked[12810] = data_i[12810] & sel_one_hot_i[100];
  assign data_masked[12809] = data_i[12809] & sel_one_hot_i[100];
  assign data_masked[12808] = data_i[12808] & sel_one_hot_i[100];
  assign data_masked[12807] = data_i[12807] & sel_one_hot_i[100];
  assign data_masked[12806] = data_i[12806] & sel_one_hot_i[100];
  assign data_masked[12805] = data_i[12805] & sel_one_hot_i[100];
  assign data_masked[12804] = data_i[12804] & sel_one_hot_i[100];
  assign data_masked[12803] = data_i[12803] & sel_one_hot_i[100];
  assign data_masked[12802] = data_i[12802] & sel_one_hot_i[100];
  assign data_masked[12801] = data_i[12801] & sel_one_hot_i[100];
  assign data_masked[12800] = data_i[12800] & sel_one_hot_i[100];
  assign data_masked[13055] = data_i[13055] & sel_one_hot_i[101];
  assign data_masked[13054] = data_i[13054] & sel_one_hot_i[101];
  assign data_masked[13053] = data_i[13053] & sel_one_hot_i[101];
  assign data_masked[13052] = data_i[13052] & sel_one_hot_i[101];
  assign data_masked[13051] = data_i[13051] & sel_one_hot_i[101];
  assign data_masked[13050] = data_i[13050] & sel_one_hot_i[101];
  assign data_masked[13049] = data_i[13049] & sel_one_hot_i[101];
  assign data_masked[13048] = data_i[13048] & sel_one_hot_i[101];
  assign data_masked[13047] = data_i[13047] & sel_one_hot_i[101];
  assign data_masked[13046] = data_i[13046] & sel_one_hot_i[101];
  assign data_masked[13045] = data_i[13045] & sel_one_hot_i[101];
  assign data_masked[13044] = data_i[13044] & sel_one_hot_i[101];
  assign data_masked[13043] = data_i[13043] & sel_one_hot_i[101];
  assign data_masked[13042] = data_i[13042] & sel_one_hot_i[101];
  assign data_masked[13041] = data_i[13041] & sel_one_hot_i[101];
  assign data_masked[13040] = data_i[13040] & sel_one_hot_i[101];
  assign data_masked[13039] = data_i[13039] & sel_one_hot_i[101];
  assign data_masked[13038] = data_i[13038] & sel_one_hot_i[101];
  assign data_masked[13037] = data_i[13037] & sel_one_hot_i[101];
  assign data_masked[13036] = data_i[13036] & sel_one_hot_i[101];
  assign data_masked[13035] = data_i[13035] & sel_one_hot_i[101];
  assign data_masked[13034] = data_i[13034] & sel_one_hot_i[101];
  assign data_masked[13033] = data_i[13033] & sel_one_hot_i[101];
  assign data_masked[13032] = data_i[13032] & sel_one_hot_i[101];
  assign data_masked[13031] = data_i[13031] & sel_one_hot_i[101];
  assign data_masked[13030] = data_i[13030] & sel_one_hot_i[101];
  assign data_masked[13029] = data_i[13029] & sel_one_hot_i[101];
  assign data_masked[13028] = data_i[13028] & sel_one_hot_i[101];
  assign data_masked[13027] = data_i[13027] & sel_one_hot_i[101];
  assign data_masked[13026] = data_i[13026] & sel_one_hot_i[101];
  assign data_masked[13025] = data_i[13025] & sel_one_hot_i[101];
  assign data_masked[13024] = data_i[13024] & sel_one_hot_i[101];
  assign data_masked[13023] = data_i[13023] & sel_one_hot_i[101];
  assign data_masked[13022] = data_i[13022] & sel_one_hot_i[101];
  assign data_masked[13021] = data_i[13021] & sel_one_hot_i[101];
  assign data_masked[13020] = data_i[13020] & sel_one_hot_i[101];
  assign data_masked[13019] = data_i[13019] & sel_one_hot_i[101];
  assign data_masked[13018] = data_i[13018] & sel_one_hot_i[101];
  assign data_masked[13017] = data_i[13017] & sel_one_hot_i[101];
  assign data_masked[13016] = data_i[13016] & sel_one_hot_i[101];
  assign data_masked[13015] = data_i[13015] & sel_one_hot_i[101];
  assign data_masked[13014] = data_i[13014] & sel_one_hot_i[101];
  assign data_masked[13013] = data_i[13013] & sel_one_hot_i[101];
  assign data_masked[13012] = data_i[13012] & sel_one_hot_i[101];
  assign data_masked[13011] = data_i[13011] & sel_one_hot_i[101];
  assign data_masked[13010] = data_i[13010] & sel_one_hot_i[101];
  assign data_masked[13009] = data_i[13009] & sel_one_hot_i[101];
  assign data_masked[13008] = data_i[13008] & sel_one_hot_i[101];
  assign data_masked[13007] = data_i[13007] & sel_one_hot_i[101];
  assign data_masked[13006] = data_i[13006] & sel_one_hot_i[101];
  assign data_masked[13005] = data_i[13005] & sel_one_hot_i[101];
  assign data_masked[13004] = data_i[13004] & sel_one_hot_i[101];
  assign data_masked[13003] = data_i[13003] & sel_one_hot_i[101];
  assign data_masked[13002] = data_i[13002] & sel_one_hot_i[101];
  assign data_masked[13001] = data_i[13001] & sel_one_hot_i[101];
  assign data_masked[13000] = data_i[13000] & sel_one_hot_i[101];
  assign data_masked[12999] = data_i[12999] & sel_one_hot_i[101];
  assign data_masked[12998] = data_i[12998] & sel_one_hot_i[101];
  assign data_masked[12997] = data_i[12997] & sel_one_hot_i[101];
  assign data_masked[12996] = data_i[12996] & sel_one_hot_i[101];
  assign data_masked[12995] = data_i[12995] & sel_one_hot_i[101];
  assign data_masked[12994] = data_i[12994] & sel_one_hot_i[101];
  assign data_masked[12993] = data_i[12993] & sel_one_hot_i[101];
  assign data_masked[12992] = data_i[12992] & sel_one_hot_i[101];
  assign data_masked[12991] = data_i[12991] & sel_one_hot_i[101];
  assign data_masked[12990] = data_i[12990] & sel_one_hot_i[101];
  assign data_masked[12989] = data_i[12989] & sel_one_hot_i[101];
  assign data_masked[12988] = data_i[12988] & sel_one_hot_i[101];
  assign data_masked[12987] = data_i[12987] & sel_one_hot_i[101];
  assign data_masked[12986] = data_i[12986] & sel_one_hot_i[101];
  assign data_masked[12985] = data_i[12985] & sel_one_hot_i[101];
  assign data_masked[12984] = data_i[12984] & sel_one_hot_i[101];
  assign data_masked[12983] = data_i[12983] & sel_one_hot_i[101];
  assign data_masked[12982] = data_i[12982] & sel_one_hot_i[101];
  assign data_masked[12981] = data_i[12981] & sel_one_hot_i[101];
  assign data_masked[12980] = data_i[12980] & sel_one_hot_i[101];
  assign data_masked[12979] = data_i[12979] & sel_one_hot_i[101];
  assign data_masked[12978] = data_i[12978] & sel_one_hot_i[101];
  assign data_masked[12977] = data_i[12977] & sel_one_hot_i[101];
  assign data_masked[12976] = data_i[12976] & sel_one_hot_i[101];
  assign data_masked[12975] = data_i[12975] & sel_one_hot_i[101];
  assign data_masked[12974] = data_i[12974] & sel_one_hot_i[101];
  assign data_masked[12973] = data_i[12973] & sel_one_hot_i[101];
  assign data_masked[12972] = data_i[12972] & sel_one_hot_i[101];
  assign data_masked[12971] = data_i[12971] & sel_one_hot_i[101];
  assign data_masked[12970] = data_i[12970] & sel_one_hot_i[101];
  assign data_masked[12969] = data_i[12969] & sel_one_hot_i[101];
  assign data_masked[12968] = data_i[12968] & sel_one_hot_i[101];
  assign data_masked[12967] = data_i[12967] & sel_one_hot_i[101];
  assign data_masked[12966] = data_i[12966] & sel_one_hot_i[101];
  assign data_masked[12965] = data_i[12965] & sel_one_hot_i[101];
  assign data_masked[12964] = data_i[12964] & sel_one_hot_i[101];
  assign data_masked[12963] = data_i[12963] & sel_one_hot_i[101];
  assign data_masked[12962] = data_i[12962] & sel_one_hot_i[101];
  assign data_masked[12961] = data_i[12961] & sel_one_hot_i[101];
  assign data_masked[12960] = data_i[12960] & sel_one_hot_i[101];
  assign data_masked[12959] = data_i[12959] & sel_one_hot_i[101];
  assign data_masked[12958] = data_i[12958] & sel_one_hot_i[101];
  assign data_masked[12957] = data_i[12957] & sel_one_hot_i[101];
  assign data_masked[12956] = data_i[12956] & sel_one_hot_i[101];
  assign data_masked[12955] = data_i[12955] & sel_one_hot_i[101];
  assign data_masked[12954] = data_i[12954] & sel_one_hot_i[101];
  assign data_masked[12953] = data_i[12953] & sel_one_hot_i[101];
  assign data_masked[12952] = data_i[12952] & sel_one_hot_i[101];
  assign data_masked[12951] = data_i[12951] & sel_one_hot_i[101];
  assign data_masked[12950] = data_i[12950] & sel_one_hot_i[101];
  assign data_masked[12949] = data_i[12949] & sel_one_hot_i[101];
  assign data_masked[12948] = data_i[12948] & sel_one_hot_i[101];
  assign data_masked[12947] = data_i[12947] & sel_one_hot_i[101];
  assign data_masked[12946] = data_i[12946] & sel_one_hot_i[101];
  assign data_masked[12945] = data_i[12945] & sel_one_hot_i[101];
  assign data_masked[12944] = data_i[12944] & sel_one_hot_i[101];
  assign data_masked[12943] = data_i[12943] & sel_one_hot_i[101];
  assign data_masked[12942] = data_i[12942] & sel_one_hot_i[101];
  assign data_masked[12941] = data_i[12941] & sel_one_hot_i[101];
  assign data_masked[12940] = data_i[12940] & sel_one_hot_i[101];
  assign data_masked[12939] = data_i[12939] & sel_one_hot_i[101];
  assign data_masked[12938] = data_i[12938] & sel_one_hot_i[101];
  assign data_masked[12937] = data_i[12937] & sel_one_hot_i[101];
  assign data_masked[12936] = data_i[12936] & sel_one_hot_i[101];
  assign data_masked[12935] = data_i[12935] & sel_one_hot_i[101];
  assign data_masked[12934] = data_i[12934] & sel_one_hot_i[101];
  assign data_masked[12933] = data_i[12933] & sel_one_hot_i[101];
  assign data_masked[12932] = data_i[12932] & sel_one_hot_i[101];
  assign data_masked[12931] = data_i[12931] & sel_one_hot_i[101];
  assign data_masked[12930] = data_i[12930] & sel_one_hot_i[101];
  assign data_masked[12929] = data_i[12929] & sel_one_hot_i[101];
  assign data_masked[12928] = data_i[12928] & sel_one_hot_i[101];
  assign data_masked[13183] = data_i[13183] & sel_one_hot_i[102];
  assign data_masked[13182] = data_i[13182] & sel_one_hot_i[102];
  assign data_masked[13181] = data_i[13181] & sel_one_hot_i[102];
  assign data_masked[13180] = data_i[13180] & sel_one_hot_i[102];
  assign data_masked[13179] = data_i[13179] & sel_one_hot_i[102];
  assign data_masked[13178] = data_i[13178] & sel_one_hot_i[102];
  assign data_masked[13177] = data_i[13177] & sel_one_hot_i[102];
  assign data_masked[13176] = data_i[13176] & sel_one_hot_i[102];
  assign data_masked[13175] = data_i[13175] & sel_one_hot_i[102];
  assign data_masked[13174] = data_i[13174] & sel_one_hot_i[102];
  assign data_masked[13173] = data_i[13173] & sel_one_hot_i[102];
  assign data_masked[13172] = data_i[13172] & sel_one_hot_i[102];
  assign data_masked[13171] = data_i[13171] & sel_one_hot_i[102];
  assign data_masked[13170] = data_i[13170] & sel_one_hot_i[102];
  assign data_masked[13169] = data_i[13169] & sel_one_hot_i[102];
  assign data_masked[13168] = data_i[13168] & sel_one_hot_i[102];
  assign data_masked[13167] = data_i[13167] & sel_one_hot_i[102];
  assign data_masked[13166] = data_i[13166] & sel_one_hot_i[102];
  assign data_masked[13165] = data_i[13165] & sel_one_hot_i[102];
  assign data_masked[13164] = data_i[13164] & sel_one_hot_i[102];
  assign data_masked[13163] = data_i[13163] & sel_one_hot_i[102];
  assign data_masked[13162] = data_i[13162] & sel_one_hot_i[102];
  assign data_masked[13161] = data_i[13161] & sel_one_hot_i[102];
  assign data_masked[13160] = data_i[13160] & sel_one_hot_i[102];
  assign data_masked[13159] = data_i[13159] & sel_one_hot_i[102];
  assign data_masked[13158] = data_i[13158] & sel_one_hot_i[102];
  assign data_masked[13157] = data_i[13157] & sel_one_hot_i[102];
  assign data_masked[13156] = data_i[13156] & sel_one_hot_i[102];
  assign data_masked[13155] = data_i[13155] & sel_one_hot_i[102];
  assign data_masked[13154] = data_i[13154] & sel_one_hot_i[102];
  assign data_masked[13153] = data_i[13153] & sel_one_hot_i[102];
  assign data_masked[13152] = data_i[13152] & sel_one_hot_i[102];
  assign data_masked[13151] = data_i[13151] & sel_one_hot_i[102];
  assign data_masked[13150] = data_i[13150] & sel_one_hot_i[102];
  assign data_masked[13149] = data_i[13149] & sel_one_hot_i[102];
  assign data_masked[13148] = data_i[13148] & sel_one_hot_i[102];
  assign data_masked[13147] = data_i[13147] & sel_one_hot_i[102];
  assign data_masked[13146] = data_i[13146] & sel_one_hot_i[102];
  assign data_masked[13145] = data_i[13145] & sel_one_hot_i[102];
  assign data_masked[13144] = data_i[13144] & sel_one_hot_i[102];
  assign data_masked[13143] = data_i[13143] & sel_one_hot_i[102];
  assign data_masked[13142] = data_i[13142] & sel_one_hot_i[102];
  assign data_masked[13141] = data_i[13141] & sel_one_hot_i[102];
  assign data_masked[13140] = data_i[13140] & sel_one_hot_i[102];
  assign data_masked[13139] = data_i[13139] & sel_one_hot_i[102];
  assign data_masked[13138] = data_i[13138] & sel_one_hot_i[102];
  assign data_masked[13137] = data_i[13137] & sel_one_hot_i[102];
  assign data_masked[13136] = data_i[13136] & sel_one_hot_i[102];
  assign data_masked[13135] = data_i[13135] & sel_one_hot_i[102];
  assign data_masked[13134] = data_i[13134] & sel_one_hot_i[102];
  assign data_masked[13133] = data_i[13133] & sel_one_hot_i[102];
  assign data_masked[13132] = data_i[13132] & sel_one_hot_i[102];
  assign data_masked[13131] = data_i[13131] & sel_one_hot_i[102];
  assign data_masked[13130] = data_i[13130] & sel_one_hot_i[102];
  assign data_masked[13129] = data_i[13129] & sel_one_hot_i[102];
  assign data_masked[13128] = data_i[13128] & sel_one_hot_i[102];
  assign data_masked[13127] = data_i[13127] & sel_one_hot_i[102];
  assign data_masked[13126] = data_i[13126] & sel_one_hot_i[102];
  assign data_masked[13125] = data_i[13125] & sel_one_hot_i[102];
  assign data_masked[13124] = data_i[13124] & sel_one_hot_i[102];
  assign data_masked[13123] = data_i[13123] & sel_one_hot_i[102];
  assign data_masked[13122] = data_i[13122] & sel_one_hot_i[102];
  assign data_masked[13121] = data_i[13121] & sel_one_hot_i[102];
  assign data_masked[13120] = data_i[13120] & sel_one_hot_i[102];
  assign data_masked[13119] = data_i[13119] & sel_one_hot_i[102];
  assign data_masked[13118] = data_i[13118] & sel_one_hot_i[102];
  assign data_masked[13117] = data_i[13117] & sel_one_hot_i[102];
  assign data_masked[13116] = data_i[13116] & sel_one_hot_i[102];
  assign data_masked[13115] = data_i[13115] & sel_one_hot_i[102];
  assign data_masked[13114] = data_i[13114] & sel_one_hot_i[102];
  assign data_masked[13113] = data_i[13113] & sel_one_hot_i[102];
  assign data_masked[13112] = data_i[13112] & sel_one_hot_i[102];
  assign data_masked[13111] = data_i[13111] & sel_one_hot_i[102];
  assign data_masked[13110] = data_i[13110] & sel_one_hot_i[102];
  assign data_masked[13109] = data_i[13109] & sel_one_hot_i[102];
  assign data_masked[13108] = data_i[13108] & sel_one_hot_i[102];
  assign data_masked[13107] = data_i[13107] & sel_one_hot_i[102];
  assign data_masked[13106] = data_i[13106] & sel_one_hot_i[102];
  assign data_masked[13105] = data_i[13105] & sel_one_hot_i[102];
  assign data_masked[13104] = data_i[13104] & sel_one_hot_i[102];
  assign data_masked[13103] = data_i[13103] & sel_one_hot_i[102];
  assign data_masked[13102] = data_i[13102] & sel_one_hot_i[102];
  assign data_masked[13101] = data_i[13101] & sel_one_hot_i[102];
  assign data_masked[13100] = data_i[13100] & sel_one_hot_i[102];
  assign data_masked[13099] = data_i[13099] & sel_one_hot_i[102];
  assign data_masked[13098] = data_i[13098] & sel_one_hot_i[102];
  assign data_masked[13097] = data_i[13097] & sel_one_hot_i[102];
  assign data_masked[13096] = data_i[13096] & sel_one_hot_i[102];
  assign data_masked[13095] = data_i[13095] & sel_one_hot_i[102];
  assign data_masked[13094] = data_i[13094] & sel_one_hot_i[102];
  assign data_masked[13093] = data_i[13093] & sel_one_hot_i[102];
  assign data_masked[13092] = data_i[13092] & sel_one_hot_i[102];
  assign data_masked[13091] = data_i[13091] & sel_one_hot_i[102];
  assign data_masked[13090] = data_i[13090] & sel_one_hot_i[102];
  assign data_masked[13089] = data_i[13089] & sel_one_hot_i[102];
  assign data_masked[13088] = data_i[13088] & sel_one_hot_i[102];
  assign data_masked[13087] = data_i[13087] & sel_one_hot_i[102];
  assign data_masked[13086] = data_i[13086] & sel_one_hot_i[102];
  assign data_masked[13085] = data_i[13085] & sel_one_hot_i[102];
  assign data_masked[13084] = data_i[13084] & sel_one_hot_i[102];
  assign data_masked[13083] = data_i[13083] & sel_one_hot_i[102];
  assign data_masked[13082] = data_i[13082] & sel_one_hot_i[102];
  assign data_masked[13081] = data_i[13081] & sel_one_hot_i[102];
  assign data_masked[13080] = data_i[13080] & sel_one_hot_i[102];
  assign data_masked[13079] = data_i[13079] & sel_one_hot_i[102];
  assign data_masked[13078] = data_i[13078] & sel_one_hot_i[102];
  assign data_masked[13077] = data_i[13077] & sel_one_hot_i[102];
  assign data_masked[13076] = data_i[13076] & sel_one_hot_i[102];
  assign data_masked[13075] = data_i[13075] & sel_one_hot_i[102];
  assign data_masked[13074] = data_i[13074] & sel_one_hot_i[102];
  assign data_masked[13073] = data_i[13073] & sel_one_hot_i[102];
  assign data_masked[13072] = data_i[13072] & sel_one_hot_i[102];
  assign data_masked[13071] = data_i[13071] & sel_one_hot_i[102];
  assign data_masked[13070] = data_i[13070] & sel_one_hot_i[102];
  assign data_masked[13069] = data_i[13069] & sel_one_hot_i[102];
  assign data_masked[13068] = data_i[13068] & sel_one_hot_i[102];
  assign data_masked[13067] = data_i[13067] & sel_one_hot_i[102];
  assign data_masked[13066] = data_i[13066] & sel_one_hot_i[102];
  assign data_masked[13065] = data_i[13065] & sel_one_hot_i[102];
  assign data_masked[13064] = data_i[13064] & sel_one_hot_i[102];
  assign data_masked[13063] = data_i[13063] & sel_one_hot_i[102];
  assign data_masked[13062] = data_i[13062] & sel_one_hot_i[102];
  assign data_masked[13061] = data_i[13061] & sel_one_hot_i[102];
  assign data_masked[13060] = data_i[13060] & sel_one_hot_i[102];
  assign data_masked[13059] = data_i[13059] & sel_one_hot_i[102];
  assign data_masked[13058] = data_i[13058] & sel_one_hot_i[102];
  assign data_masked[13057] = data_i[13057] & sel_one_hot_i[102];
  assign data_masked[13056] = data_i[13056] & sel_one_hot_i[102];
  assign data_masked[13311] = data_i[13311] & sel_one_hot_i[103];
  assign data_masked[13310] = data_i[13310] & sel_one_hot_i[103];
  assign data_masked[13309] = data_i[13309] & sel_one_hot_i[103];
  assign data_masked[13308] = data_i[13308] & sel_one_hot_i[103];
  assign data_masked[13307] = data_i[13307] & sel_one_hot_i[103];
  assign data_masked[13306] = data_i[13306] & sel_one_hot_i[103];
  assign data_masked[13305] = data_i[13305] & sel_one_hot_i[103];
  assign data_masked[13304] = data_i[13304] & sel_one_hot_i[103];
  assign data_masked[13303] = data_i[13303] & sel_one_hot_i[103];
  assign data_masked[13302] = data_i[13302] & sel_one_hot_i[103];
  assign data_masked[13301] = data_i[13301] & sel_one_hot_i[103];
  assign data_masked[13300] = data_i[13300] & sel_one_hot_i[103];
  assign data_masked[13299] = data_i[13299] & sel_one_hot_i[103];
  assign data_masked[13298] = data_i[13298] & sel_one_hot_i[103];
  assign data_masked[13297] = data_i[13297] & sel_one_hot_i[103];
  assign data_masked[13296] = data_i[13296] & sel_one_hot_i[103];
  assign data_masked[13295] = data_i[13295] & sel_one_hot_i[103];
  assign data_masked[13294] = data_i[13294] & sel_one_hot_i[103];
  assign data_masked[13293] = data_i[13293] & sel_one_hot_i[103];
  assign data_masked[13292] = data_i[13292] & sel_one_hot_i[103];
  assign data_masked[13291] = data_i[13291] & sel_one_hot_i[103];
  assign data_masked[13290] = data_i[13290] & sel_one_hot_i[103];
  assign data_masked[13289] = data_i[13289] & sel_one_hot_i[103];
  assign data_masked[13288] = data_i[13288] & sel_one_hot_i[103];
  assign data_masked[13287] = data_i[13287] & sel_one_hot_i[103];
  assign data_masked[13286] = data_i[13286] & sel_one_hot_i[103];
  assign data_masked[13285] = data_i[13285] & sel_one_hot_i[103];
  assign data_masked[13284] = data_i[13284] & sel_one_hot_i[103];
  assign data_masked[13283] = data_i[13283] & sel_one_hot_i[103];
  assign data_masked[13282] = data_i[13282] & sel_one_hot_i[103];
  assign data_masked[13281] = data_i[13281] & sel_one_hot_i[103];
  assign data_masked[13280] = data_i[13280] & sel_one_hot_i[103];
  assign data_masked[13279] = data_i[13279] & sel_one_hot_i[103];
  assign data_masked[13278] = data_i[13278] & sel_one_hot_i[103];
  assign data_masked[13277] = data_i[13277] & sel_one_hot_i[103];
  assign data_masked[13276] = data_i[13276] & sel_one_hot_i[103];
  assign data_masked[13275] = data_i[13275] & sel_one_hot_i[103];
  assign data_masked[13274] = data_i[13274] & sel_one_hot_i[103];
  assign data_masked[13273] = data_i[13273] & sel_one_hot_i[103];
  assign data_masked[13272] = data_i[13272] & sel_one_hot_i[103];
  assign data_masked[13271] = data_i[13271] & sel_one_hot_i[103];
  assign data_masked[13270] = data_i[13270] & sel_one_hot_i[103];
  assign data_masked[13269] = data_i[13269] & sel_one_hot_i[103];
  assign data_masked[13268] = data_i[13268] & sel_one_hot_i[103];
  assign data_masked[13267] = data_i[13267] & sel_one_hot_i[103];
  assign data_masked[13266] = data_i[13266] & sel_one_hot_i[103];
  assign data_masked[13265] = data_i[13265] & sel_one_hot_i[103];
  assign data_masked[13264] = data_i[13264] & sel_one_hot_i[103];
  assign data_masked[13263] = data_i[13263] & sel_one_hot_i[103];
  assign data_masked[13262] = data_i[13262] & sel_one_hot_i[103];
  assign data_masked[13261] = data_i[13261] & sel_one_hot_i[103];
  assign data_masked[13260] = data_i[13260] & sel_one_hot_i[103];
  assign data_masked[13259] = data_i[13259] & sel_one_hot_i[103];
  assign data_masked[13258] = data_i[13258] & sel_one_hot_i[103];
  assign data_masked[13257] = data_i[13257] & sel_one_hot_i[103];
  assign data_masked[13256] = data_i[13256] & sel_one_hot_i[103];
  assign data_masked[13255] = data_i[13255] & sel_one_hot_i[103];
  assign data_masked[13254] = data_i[13254] & sel_one_hot_i[103];
  assign data_masked[13253] = data_i[13253] & sel_one_hot_i[103];
  assign data_masked[13252] = data_i[13252] & sel_one_hot_i[103];
  assign data_masked[13251] = data_i[13251] & sel_one_hot_i[103];
  assign data_masked[13250] = data_i[13250] & sel_one_hot_i[103];
  assign data_masked[13249] = data_i[13249] & sel_one_hot_i[103];
  assign data_masked[13248] = data_i[13248] & sel_one_hot_i[103];
  assign data_masked[13247] = data_i[13247] & sel_one_hot_i[103];
  assign data_masked[13246] = data_i[13246] & sel_one_hot_i[103];
  assign data_masked[13245] = data_i[13245] & sel_one_hot_i[103];
  assign data_masked[13244] = data_i[13244] & sel_one_hot_i[103];
  assign data_masked[13243] = data_i[13243] & sel_one_hot_i[103];
  assign data_masked[13242] = data_i[13242] & sel_one_hot_i[103];
  assign data_masked[13241] = data_i[13241] & sel_one_hot_i[103];
  assign data_masked[13240] = data_i[13240] & sel_one_hot_i[103];
  assign data_masked[13239] = data_i[13239] & sel_one_hot_i[103];
  assign data_masked[13238] = data_i[13238] & sel_one_hot_i[103];
  assign data_masked[13237] = data_i[13237] & sel_one_hot_i[103];
  assign data_masked[13236] = data_i[13236] & sel_one_hot_i[103];
  assign data_masked[13235] = data_i[13235] & sel_one_hot_i[103];
  assign data_masked[13234] = data_i[13234] & sel_one_hot_i[103];
  assign data_masked[13233] = data_i[13233] & sel_one_hot_i[103];
  assign data_masked[13232] = data_i[13232] & sel_one_hot_i[103];
  assign data_masked[13231] = data_i[13231] & sel_one_hot_i[103];
  assign data_masked[13230] = data_i[13230] & sel_one_hot_i[103];
  assign data_masked[13229] = data_i[13229] & sel_one_hot_i[103];
  assign data_masked[13228] = data_i[13228] & sel_one_hot_i[103];
  assign data_masked[13227] = data_i[13227] & sel_one_hot_i[103];
  assign data_masked[13226] = data_i[13226] & sel_one_hot_i[103];
  assign data_masked[13225] = data_i[13225] & sel_one_hot_i[103];
  assign data_masked[13224] = data_i[13224] & sel_one_hot_i[103];
  assign data_masked[13223] = data_i[13223] & sel_one_hot_i[103];
  assign data_masked[13222] = data_i[13222] & sel_one_hot_i[103];
  assign data_masked[13221] = data_i[13221] & sel_one_hot_i[103];
  assign data_masked[13220] = data_i[13220] & sel_one_hot_i[103];
  assign data_masked[13219] = data_i[13219] & sel_one_hot_i[103];
  assign data_masked[13218] = data_i[13218] & sel_one_hot_i[103];
  assign data_masked[13217] = data_i[13217] & sel_one_hot_i[103];
  assign data_masked[13216] = data_i[13216] & sel_one_hot_i[103];
  assign data_masked[13215] = data_i[13215] & sel_one_hot_i[103];
  assign data_masked[13214] = data_i[13214] & sel_one_hot_i[103];
  assign data_masked[13213] = data_i[13213] & sel_one_hot_i[103];
  assign data_masked[13212] = data_i[13212] & sel_one_hot_i[103];
  assign data_masked[13211] = data_i[13211] & sel_one_hot_i[103];
  assign data_masked[13210] = data_i[13210] & sel_one_hot_i[103];
  assign data_masked[13209] = data_i[13209] & sel_one_hot_i[103];
  assign data_masked[13208] = data_i[13208] & sel_one_hot_i[103];
  assign data_masked[13207] = data_i[13207] & sel_one_hot_i[103];
  assign data_masked[13206] = data_i[13206] & sel_one_hot_i[103];
  assign data_masked[13205] = data_i[13205] & sel_one_hot_i[103];
  assign data_masked[13204] = data_i[13204] & sel_one_hot_i[103];
  assign data_masked[13203] = data_i[13203] & sel_one_hot_i[103];
  assign data_masked[13202] = data_i[13202] & sel_one_hot_i[103];
  assign data_masked[13201] = data_i[13201] & sel_one_hot_i[103];
  assign data_masked[13200] = data_i[13200] & sel_one_hot_i[103];
  assign data_masked[13199] = data_i[13199] & sel_one_hot_i[103];
  assign data_masked[13198] = data_i[13198] & sel_one_hot_i[103];
  assign data_masked[13197] = data_i[13197] & sel_one_hot_i[103];
  assign data_masked[13196] = data_i[13196] & sel_one_hot_i[103];
  assign data_masked[13195] = data_i[13195] & sel_one_hot_i[103];
  assign data_masked[13194] = data_i[13194] & sel_one_hot_i[103];
  assign data_masked[13193] = data_i[13193] & sel_one_hot_i[103];
  assign data_masked[13192] = data_i[13192] & sel_one_hot_i[103];
  assign data_masked[13191] = data_i[13191] & sel_one_hot_i[103];
  assign data_masked[13190] = data_i[13190] & sel_one_hot_i[103];
  assign data_masked[13189] = data_i[13189] & sel_one_hot_i[103];
  assign data_masked[13188] = data_i[13188] & sel_one_hot_i[103];
  assign data_masked[13187] = data_i[13187] & sel_one_hot_i[103];
  assign data_masked[13186] = data_i[13186] & sel_one_hot_i[103];
  assign data_masked[13185] = data_i[13185] & sel_one_hot_i[103];
  assign data_masked[13184] = data_i[13184] & sel_one_hot_i[103];
  assign data_masked[13439] = data_i[13439] & sel_one_hot_i[104];
  assign data_masked[13438] = data_i[13438] & sel_one_hot_i[104];
  assign data_masked[13437] = data_i[13437] & sel_one_hot_i[104];
  assign data_masked[13436] = data_i[13436] & sel_one_hot_i[104];
  assign data_masked[13435] = data_i[13435] & sel_one_hot_i[104];
  assign data_masked[13434] = data_i[13434] & sel_one_hot_i[104];
  assign data_masked[13433] = data_i[13433] & sel_one_hot_i[104];
  assign data_masked[13432] = data_i[13432] & sel_one_hot_i[104];
  assign data_masked[13431] = data_i[13431] & sel_one_hot_i[104];
  assign data_masked[13430] = data_i[13430] & sel_one_hot_i[104];
  assign data_masked[13429] = data_i[13429] & sel_one_hot_i[104];
  assign data_masked[13428] = data_i[13428] & sel_one_hot_i[104];
  assign data_masked[13427] = data_i[13427] & sel_one_hot_i[104];
  assign data_masked[13426] = data_i[13426] & sel_one_hot_i[104];
  assign data_masked[13425] = data_i[13425] & sel_one_hot_i[104];
  assign data_masked[13424] = data_i[13424] & sel_one_hot_i[104];
  assign data_masked[13423] = data_i[13423] & sel_one_hot_i[104];
  assign data_masked[13422] = data_i[13422] & sel_one_hot_i[104];
  assign data_masked[13421] = data_i[13421] & sel_one_hot_i[104];
  assign data_masked[13420] = data_i[13420] & sel_one_hot_i[104];
  assign data_masked[13419] = data_i[13419] & sel_one_hot_i[104];
  assign data_masked[13418] = data_i[13418] & sel_one_hot_i[104];
  assign data_masked[13417] = data_i[13417] & sel_one_hot_i[104];
  assign data_masked[13416] = data_i[13416] & sel_one_hot_i[104];
  assign data_masked[13415] = data_i[13415] & sel_one_hot_i[104];
  assign data_masked[13414] = data_i[13414] & sel_one_hot_i[104];
  assign data_masked[13413] = data_i[13413] & sel_one_hot_i[104];
  assign data_masked[13412] = data_i[13412] & sel_one_hot_i[104];
  assign data_masked[13411] = data_i[13411] & sel_one_hot_i[104];
  assign data_masked[13410] = data_i[13410] & sel_one_hot_i[104];
  assign data_masked[13409] = data_i[13409] & sel_one_hot_i[104];
  assign data_masked[13408] = data_i[13408] & sel_one_hot_i[104];
  assign data_masked[13407] = data_i[13407] & sel_one_hot_i[104];
  assign data_masked[13406] = data_i[13406] & sel_one_hot_i[104];
  assign data_masked[13405] = data_i[13405] & sel_one_hot_i[104];
  assign data_masked[13404] = data_i[13404] & sel_one_hot_i[104];
  assign data_masked[13403] = data_i[13403] & sel_one_hot_i[104];
  assign data_masked[13402] = data_i[13402] & sel_one_hot_i[104];
  assign data_masked[13401] = data_i[13401] & sel_one_hot_i[104];
  assign data_masked[13400] = data_i[13400] & sel_one_hot_i[104];
  assign data_masked[13399] = data_i[13399] & sel_one_hot_i[104];
  assign data_masked[13398] = data_i[13398] & sel_one_hot_i[104];
  assign data_masked[13397] = data_i[13397] & sel_one_hot_i[104];
  assign data_masked[13396] = data_i[13396] & sel_one_hot_i[104];
  assign data_masked[13395] = data_i[13395] & sel_one_hot_i[104];
  assign data_masked[13394] = data_i[13394] & sel_one_hot_i[104];
  assign data_masked[13393] = data_i[13393] & sel_one_hot_i[104];
  assign data_masked[13392] = data_i[13392] & sel_one_hot_i[104];
  assign data_masked[13391] = data_i[13391] & sel_one_hot_i[104];
  assign data_masked[13390] = data_i[13390] & sel_one_hot_i[104];
  assign data_masked[13389] = data_i[13389] & sel_one_hot_i[104];
  assign data_masked[13388] = data_i[13388] & sel_one_hot_i[104];
  assign data_masked[13387] = data_i[13387] & sel_one_hot_i[104];
  assign data_masked[13386] = data_i[13386] & sel_one_hot_i[104];
  assign data_masked[13385] = data_i[13385] & sel_one_hot_i[104];
  assign data_masked[13384] = data_i[13384] & sel_one_hot_i[104];
  assign data_masked[13383] = data_i[13383] & sel_one_hot_i[104];
  assign data_masked[13382] = data_i[13382] & sel_one_hot_i[104];
  assign data_masked[13381] = data_i[13381] & sel_one_hot_i[104];
  assign data_masked[13380] = data_i[13380] & sel_one_hot_i[104];
  assign data_masked[13379] = data_i[13379] & sel_one_hot_i[104];
  assign data_masked[13378] = data_i[13378] & sel_one_hot_i[104];
  assign data_masked[13377] = data_i[13377] & sel_one_hot_i[104];
  assign data_masked[13376] = data_i[13376] & sel_one_hot_i[104];
  assign data_masked[13375] = data_i[13375] & sel_one_hot_i[104];
  assign data_masked[13374] = data_i[13374] & sel_one_hot_i[104];
  assign data_masked[13373] = data_i[13373] & sel_one_hot_i[104];
  assign data_masked[13372] = data_i[13372] & sel_one_hot_i[104];
  assign data_masked[13371] = data_i[13371] & sel_one_hot_i[104];
  assign data_masked[13370] = data_i[13370] & sel_one_hot_i[104];
  assign data_masked[13369] = data_i[13369] & sel_one_hot_i[104];
  assign data_masked[13368] = data_i[13368] & sel_one_hot_i[104];
  assign data_masked[13367] = data_i[13367] & sel_one_hot_i[104];
  assign data_masked[13366] = data_i[13366] & sel_one_hot_i[104];
  assign data_masked[13365] = data_i[13365] & sel_one_hot_i[104];
  assign data_masked[13364] = data_i[13364] & sel_one_hot_i[104];
  assign data_masked[13363] = data_i[13363] & sel_one_hot_i[104];
  assign data_masked[13362] = data_i[13362] & sel_one_hot_i[104];
  assign data_masked[13361] = data_i[13361] & sel_one_hot_i[104];
  assign data_masked[13360] = data_i[13360] & sel_one_hot_i[104];
  assign data_masked[13359] = data_i[13359] & sel_one_hot_i[104];
  assign data_masked[13358] = data_i[13358] & sel_one_hot_i[104];
  assign data_masked[13357] = data_i[13357] & sel_one_hot_i[104];
  assign data_masked[13356] = data_i[13356] & sel_one_hot_i[104];
  assign data_masked[13355] = data_i[13355] & sel_one_hot_i[104];
  assign data_masked[13354] = data_i[13354] & sel_one_hot_i[104];
  assign data_masked[13353] = data_i[13353] & sel_one_hot_i[104];
  assign data_masked[13352] = data_i[13352] & sel_one_hot_i[104];
  assign data_masked[13351] = data_i[13351] & sel_one_hot_i[104];
  assign data_masked[13350] = data_i[13350] & sel_one_hot_i[104];
  assign data_masked[13349] = data_i[13349] & sel_one_hot_i[104];
  assign data_masked[13348] = data_i[13348] & sel_one_hot_i[104];
  assign data_masked[13347] = data_i[13347] & sel_one_hot_i[104];
  assign data_masked[13346] = data_i[13346] & sel_one_hot_i[104];
  assign data_masked[13345] = data_i[13345] & sel_one_hot_i[104];
  assign data_masked[13344] = data_i[13344] & sel_one_hot_i[104];
  assign data_masked[13343] = data_i[13343] & sel_one_hot_i[104];
  assign data_masked[13342] = data_i[13342] & sel_one_hot_i[104];
  assign data_masked[13341] = data_i[13341] & sel_one_hot_i[104];
  assign data_masked[13340] = data_i[13340] & sel_one_hot_i[104];
  assign data_masked[13339] = data_i[13339] & sel_one_hot_i[104];
  assign data_masked[13338] = data_i[13338] & sel_one_hot_i[104];
  assign data_masked[13337] = data_i[13337] & sel_one_hot_i[104];
  assign data_masked[13336] = data_i[13336] & sel_one_hot_i[104];
  assign data_masked[13335] = data_i[13335] & sel_one_hot_i[104];
  assign data_masked[13334] = data_i[13334] & sel_one_hot_i[104];
  assign data_masked[13333] = data_i[13333] & sel_one_hot_i[104];
  assign data_masked[13332] = data_i[13332] & sel_one_hot_i[104];
  assign data_masked[13331] = data_i[13331] & sel_one_hot_i[104];
  assign data_masked[13330] = data_i[13330] & sel_one_hot_i[104];
  assign data_masked[13329] = data_i[13329] & sel_one_hot_i[104];
  assign data_masked[13328] = data_i[13328] & sel_one_hot_i[104];
  assign data_masked[13327] = data_i[13327] & sel_one_hot_i[104];
  assign data_masked[13326] = data_i[13326] & sel_one_hot_i[104];
  assign data_masked[13325] = data_i[13325] & sel_one_hot_i[104];
  assign data_masked[13324] = data_i[13324] & sel_one_hot_i[104];
  assign data_masked[13323] = data_i[13323] & sel_one_hot_i[104];
  assign data_masked[13322] = data_i[13322] & sel_one_hot_i[104];
  assign data_masked[13321] = data_i[13321] & sel_one_hot_i[104];
  assign data_masked[13320] = data_i[13320] & sel_one_hot_i[104];
  assign data_masked[13319] = data_i[13319] & sel_one_hot_i[104];
  assign data_masked[13318] = data_i[13318] & sel_one_hot_i[104];
  assign data_masked[13317] = data_i[13317] & sel_one_hot_i[104];
  assign data_masked[13316] = data_i[13316] & sel_one_hot_i[104];
  assign data_masked[13315] = data_i[13315] & sel_one_hot_i[104];
  assign data_masked[13314] = data_i[13314] & sel_one_hot_i[104];
  assign data_masked[13313] = data_i[13313] & sel_one_hot_i[104];
  assign data_masked[13312] = data_i[13312] & sel_one_hot_i[104];
  assign data_masked[13567] = data_i[13567] & sel_one_hot_i[105];
  assign data_masked[13566] = data_i[13566] & sel_one_hot_i[105];
  assign data_masked[13565] = data_i[13565] & sel_one_hot_i[105];
  assign data_masked[13564] = data_i[13564] & sel_one_hot_i[105];
  assign data_masked[13563] = data_i[13563] & sel_one_hot_i[105];
  assign data_masked[13562] = data_i[13562] & sel_one_hot_i[105];
  assign data_masked[13561] = data_i[13561] & sel_one_hot_i[105];
  assign data_masked[13560] = data_i[13560] & sel_one_hot_i[105];
  assign data_masked[13559] = data_i[13559] & sel_one_hot_i[105];
  assign data_masked[13558] = data_i[13558] & sel_one_hot_i[105];
  assign data_masked[13557] = data_i[13557] & sel_one_hot_i[105];
  assign data_masked[13556] = data_i[13556] & sel_one_hot_i[105];
  assign data_masked[13555] = data_i[13555] & sel_one_hot_i[105];
  assign data_masked[13554] = data_i[13554] & sel_one_hot_i[105];
  assign data_masked[13553] = data_i[13553] & sel_one_hot_i[105];
  assign data_masked[13552] = data_i[13552] & sel_one_hot_i[105];
  assign data_masked[13551] = data_i[13551] & sel_one_hot_i[105];
  assign data_masked[13550] = data_i[13550] & sel_one_hot_i[105];
  assign data_masked[13549] = data_i[13549] & sel_one_hot_i[105];
  assign data_masked[13548] = data_i[13548] & sel_one_hot_i[105];
  assign data_masked[13547] = data_i[13547] & sel_one_hot_i[105];
  assign data_masked[13546] = data_i[13546] & sel_one_hot_i[105];
  assign data_masked[13545] = data_i[13545] & sel_one_hot_i[105];
  assign data_masked[13544] = data_i[13544] & sel_one_hot_i[105];
  assign data_masked[13543] = data_i[13543] & sel_one_hot_i[105];
  assign data_masked[13542] = data_i[13542] & sel_one_hot_i[105];
  assign data_masked[13541] = data_i[13541] & sel_one_hot_i[105];
  assign data_masked[13540] = data_i[13540] & sel_one_hot_i[105];
  assign data_masked[13539] = data_i[13539] & sel_one_hot_i[105];
  assign data_masked[13538] = data_i[13538] & sel_one_hot_i[105];
  assign data_masked[13537] = data_i[13537] & sel_one_hot_i[105];
  assign data_masked[13536] = data_i[13536] & sel_one_hot_i[105];
  assign data_masked[13535] = data_i[13535] & sel_one_hot_i[105];
  assign data_masked[13534] = data_i[13534] & sel_one_hot_i[105];
  assign data_masked[13533] = data_i[13533] & sel_one_hot_i[105];
  assign data_masked[13532] = data_i[13532] & sel_one_hot_i[105];
  assign data_masked[13531] = data_i[13531] & sel_one_hot_i[105];
  assign data_masked[13530] = data_i[13530] & sel_one_hot_i[105];
  assign data_masked[13529] = data_i[13529] & sel_one_hot_i[105];
  assign data_masked[13528] = data_i[13528] & sel_one_hot_i[105];
  assign data_masked[13527] = data_i[13527] & sel_one_hot_i[105];
  assign data_masked[13526] = data_i[13526] & sel_one_hot_i[105];
  assign data_masked[13525] = data_i[13525] & sel_one_hot_i[105];
  assign data_masked[13524] = data_i[13524] & sel_one_hot_i[105];
  assign data_masked[13523] = data_i[13523] & sel_one_hot_i[105];
  assign data_masked[13522] = data_i[13522] & sel_one_hot_i[105];
  assign data_masked[13521] = data_i[13521] & sel_one_hot_i[105];
  assign data_masked[13520] = data_i[13520] & sel_one_hot_i[105];
  assign data_masked[13519] = data_i[13519] & sel_one_hot_i[105];
  assign data_masked[13518] = data_i[13518] & sel_one_hot_i[105];
  assign data_masked[13517] = data_i[13517] & sel_one_hot_i[105];
  assign data_masked[13516] = data_i[13516] & sel_one_hot_i[105];
  assign data_masked[13515] = data_i[13515] & sel_one_hot_i[105];
  assign data_masked[13514] = data_i[13514] & sel_one_hot_i[105];
  assign data_masked[13513] = data_i[13513] & sel_one_hot_i[105];
  assign data_masked[13512] = data_i[13512] & sel_one_hot_i[105];
  assign data_masked[13511] = data_i[13511] & sel_one_hot_i[105];
  assign data_masked[13510] = data_i[13510] & sel_one_hot_i[105];
  assign data_masked[13509] = data_i[13509] & sel_one_hot_i[105];
  assign data_masked[13508] = data_i[13508] & sel_one_hot_i[105];
  assign data_masked[13507] = data_i[13507] & sel_one_hot_i[105];
  assign data_masked[13506] = data_i[13506] & sel_one_hot_i[105];
  assign data_masked[13505] = data_i[13505] & sel_one_hot_i[105];
  assign data_masked[13504] = data_i[13504] & sel_one_hot_i[105];
  assign data_masked[13503] = data_i[13503] & sel_one_hot_i[105];
  assign data_masked[13502] = data_i[13502] & sel_one_hot_i[105];
  assign data_masked[13501] = data_i[13501] & sel_one_hot_i[105];
  assign data_masked[13500] = data_i[13500] & sel_one_hot_i[105];
  assign data_masked[13499] = data_i[13499] & sel_one_hot_i[105];
  assign data_masked[13498] = data_i[13498] & sel_one_hot_i[105];
  assign data_masked[13497] = data_i[13497] & sel_one_hot_i[105];
  assign data_masked[13496] = data_i[13496] & sel_one_hot_i[105];
  assign data_masked[13495] = data_i[13495] & sel_one_hot_i[105];
  assign data_masked[13494] = data_i[13494] & sel_one_hot_i[105];
  assign data_masked[13493] = data_i[13493] & sel_one_hot_i[105];
  assign data_masked[13492] = data_i[13492] & sel_one_hot_i[105];
  assign data_masked[13491] = data_i[13491] & sel_one_hot_i[105];
  assign data_masked[13490] = data_i[13490] & sel_one_hot_i[105];
  assign data_masked[13489] = data_i[13489] & sel_one_hot_i[105];
  assign data_masked[13488] = data_i[13488] & sel_one_hot_i[105];
  assign data_masked[13487] = data_i[13487] & sel_one_hot_i[105];
  assign data_masked[13486] = data_i[13486] & sel_one_hot_i[105];
  assign data_masked[13485] = data_i[13485] & sel_one_hot_i[105];
  assign data_masked[13484] = data_i[13484] & sel_one_hot_i[105];
  assign data_masked[13483] = data_i[13483] & sel_one_hot_i[105];
  assign data_masked[13482] = data_i[13482] & sel_one_hot_i[105];
  assign data_masked[13481] = data_i[13481] & sel_one_hot_i[105];
  assign data_masked[13480] = data_i[13480] & sel_one_hot_i[105];
  assign data_masked[13479] = data_i[13479] & sel_one_hot_i[105];
  assign data_masked[13478] = data_i[13478] & sel_one_hot_i[105];
  assign data_masked[13477] = data_i[13477] & sel_one_hot_i[105];
  assign data_masked[13476] = data_i[13476] & sel_one_hot_i[105];
  assign data_masked[13475] = data_i[13475] & sel_one_hot_i[105];
  assign data_masked[13474] = data_i[13474] & sel_one_hot_i[105];
  assign data_masked[13473] = data_i[13473] & sel_one_hot_i[105];
  assign data_masked[13472] = data_i[13472] & sel_one_hot_i[105];
  assign data_masked[13471] = data_i[13471] & sel_one_hot_i[105];
  assign data_masked[13470] = data_i[13470] & sel_one_hot_i[105];
  assign data_masked[13469] = data_i[13469] & sel_one_hot_i[105];
  assign data_masked[13468] = data_i[13468] & sel_one_hot_i[105];
  assign data_masked[13467] = data_i[13467] & sel_one_hot_i[105];
  assign data_masked[13466] = data_i[13466] & sel_one_hot_i[105];
  assign data_masked[13465] = data_i[13465] & sel_one_hot_i[105];
  assign data_masked[13464] = data_i[13464] & sel_one_hot_i[105];
  assign data_masked[13463] = data_i[13463] & sel_one_hot_i[105];
  assign data_masked[13462] = data_i[13462] & sel_one_hot_i[105];
  assign data_masked[13461] = data_i[13461] & sel_one_hot_i[105];
  assign data_masked[13460] = data_i[13460] & sel_one_hot_i[105];
  assign data_masked[13459] = data_i[13459] & sel_one_hot_i[105];
  assign data_masked[13458] = data_i[13458] & sel_one_hot_i[105];
  assign data_masked[13457] = data_i[13457] & sel_one_hot_i[105];
  assign data_masked[13456] = data_i[13456] & sel_one_hot_i[105];
  assign data_masked[13455] = data_i[13455] & sel_one_hot_i[105];
  assign data_masked[13454] = data_i[13454] & sel_one_hot_i[105];
  assign data_masked[13453] = data_i[13453] & sel_one_hot_i[105];
  assign data_masked[13452] = data_i[13452] & sel_one_hot_i[105];
  assign data_masked[13451] = data_i[13451] & sel_one_hot_i[105];
  assign data_masked[13450] = data_i[13450] & sel_one_hot_i[105];
  assign data_masked[13449] = data_i[13449] & sel_one_hot_i[105];
  assign data_masked[13448] = data_i[13448] & sel_one_hot_i[105];
  assign data_masked[13447] = data_i[13447] & sel_one_hot_i[105];
  assign data_masked[13446] = data_i[13446] & sel_one_hot_i[105];
  assign data_masked[13445] = data_i[13445] & sel_one_hot_i[105];
  assign data_masked[13444] = data_i[13444] & sel_one_hot_i[105];
  assign data_masked[13443] = data_i[13443] & sel_one_hot_i[105];
  assign data_masked[13442] = data_i[13442] & sel_one_hot_i[105];
  assign data_masked[13441] = data_i[13441] & sel_one_hot_i[105];
  assign data_masked[13440] = data_i[13440] & sel_one_hot_i[105];
  assign data_masked[13695] = data_i[13695] & sel_one_hot_i[106];
  assign data_masked[13694] = data_i[13694] & sel_one_hot_i[106];
  assign data_masked[13693] = data_i[13693] & sel_one_hot_i[106];
  assign data_masked[13692] = data_i[13692] & sel_one_hot_i[106];
  assign data_masked[13691] = data_i[13691] & sel_one_hot_i[106];
  assign data_masked[13690] = data_i[13690] & sel_one_hot_i[106];
  assign data_masked[13689] = data_i[13689] & sel_one_hot_i[106];
  assign data_masked[13688] = data_i[13688] & sel_one_hot_i[106];
  assign data_masked[13687] = data_i[13687] & sel_one_hot_i[106];
  assign data_masked[13686] = data_i[13686] & sel_one_hot_i[106];
  assign data_masked[13685] = data_i[13685] & sel_one_hot_i[106];
  assign data_masked[13684] = data_i[13684] & sel_one_hot_i[106];
  assign data_masked[13683] = data_i[13683] & sel_one_hot_i[106];
  assign data_masked[13682] = data_i[13682] & sel_one_hot_i[106];
  assign data_masked[13681] = data_i[13681] & sel_one_hot_i[106];
  assign data_masked[13680] = data_i[13680] & sel_one_hot_i[106];
  assign data_masked[13679] = data_i[13679] & sel_one_hot_i[106];
  assign data_masked[13678] = data_i[13678] & sel_one_hot_i[106];
  assign data_masked[13677] = data_i[13677] & sel_one_hot_i[106];
  assign data_masked[13676] = data_i[13676] & sel_one_hot_i[106];
  assign data_masked[13675] = data_i[13675] & sel_one_hot_i[106];
  assign data_masked[13674] = data_i[13674] & sel_one_hot_i[106];
  assign data_masked[13673] = data_i[13673] & sel_one_hot_i[106];
  assign data_masked[13672] = data_i[13672] & sel_one_hot_i[106];
  assign data_masked[13671] = data_i[13671] & sel_one_hot_i[106];
  assign data_masked[13670] = data_i[13670] & sel_one_hot_i[106];
  assign data_masked[13669] = data_i[13669] & sel_one_hot_i[106];
  assign data_masked[13668] = data_i[13668] & sel_one_hot_i[106];
  assign data_masked[13667] = data_i[13667] & sel_one_hot_i[106];
  assign data_masked[13666] = data_i[13666] & sel_one_hot_i[106];
  assign data_masked[13665] = data_i[13665] & sel_one_hot_i[106];
  assign data_masked[13664] = data_i[13664] & sel_one_hot_i[106];
  assign data_masked[13663] = data_i[13663] & sel_one_hot_i[106];
  assign data_masked[13662] = data_i[13662] & sel_one_hot_i[106];
  assign data_masked[13661] = data_i[13661] & sel_one_hot_i[106];
  assign data_masked[13660] = data_i[13660] & sel_one_hot_i[106];
  assign data_masked[13659] = data_i[13659] & sel_one_hot_i[106];
  assign data_masked[13658] = data_i[13658] & sel_one_hot_i[106];
  assign data_masked[13657] = data_i[13657] & sel_one_hot_i[106];
  assign data_masked[13656] = data_i[13656] & sel_one_hot_i[106];
  assign data_masked[13655] = data_i[13655] & sel_one_hot_i[106];
  assign data_masked[13654] = data_i[13654] & sel_one_hot_i[106];
  assign data_masked[13653] = data_i[13653] & sel_one_hot_i[106];
  assign data_masked[13652] = data_i[13652] & sel_one_hot_i[106];
  assign data_masked[13651] = data_i[13651] & sel_one_hot_i[106];
  assign data_masked[13650] = data_i[13650] & sel_one_hot_i[106];
  assign data_masked[13649] = data_i[13649] & sel_one_hot_i[106];
  assign data_masked[13648] = data_i[13648] & sel_one_hot_i[106];
  assign data_masked[13647] = data_i[13647] & sel_one_hot_i[106];
  assign data_masked[13646] = data_i[13646] & sel_one_hot_i[106];
  assign data_masked[13645] = data_i[13645] & sel_one_hot_i[106];
  assign data_masked[13644] = data_i[13644] & sel_one_hot_i[106];
  assign data_masked[13643] = data_i[13643] & sel_one_hot_i[106];
  assign data_masked[13642] = data_i[13642] & sel_one_hot_i[106];
  assign data_masked[13641] = data_i[13641] & sel_one_hot_i[106];
  assign data_masked[13640] = data_i[13640] & sel_one_hot_i[106];
  assign data_masked[13639] = data_i[13639] & sel_one_hot_i[106];
  assign data_masked[13638] = data_i[13638] & sel_one_hot_i[106];
  assign data_masked[13637] = data_i[13637] & sel_one_hot_i[106];
  assign data_masked[13636] = data_i[13636] & sel_one_hot_i[106];
  assign data_masked[13635] = data_i[13635] & sel_one_hot_i[106];
  assign data_masked[13634] = data_i[13634] & sel_one_hot_i[106];
  assign data_masked[13633] = data_i[13633] & sel_one_hot_i[106];
  assign data_masked[13632] = data_i[13632] & sel_one_hot_i[106];
  assign data_masked[13631] = data_i[13631] & sel_one_hot_i[106];
  assign data_masked[13630] = data_i[13630] & sel_one_hot_i[106];
  assign data_masked[13629] = data_i[13629] & sel_one_hot_i[106];
  assign data_masked[13628] = data_i[13628] & sel_one_hot_i[106];
  assign data_masked[13627] = data_i[13627] & sel_one_hot_i[106];
  assign data_masked[13626] = data_i[13626] & sel_one_hot_i[106];
  assign data_masked[13625] = data_i[13625] & sel_one_hot_i[106];
  assign data_masked[13624] = data_i[13624] & sel_one_hot_i[106];
  assign data_masked[13623] = data_i[13623] & sel_one_hot_i[106];
  assign data_masked[13622] = data_i[13622] & sel_one_hot_i[106];
  assign data_masked[13621] = data_i[13621] & sel_one_hot_i[106];
  assign data_masked[13620] = data_i[13620] & sel_one_hot_i[106];
  assign data_masked[13619] = data_i[13619] & sel_one_hot_i[106];
  assign data_masked[13618] = data_i[13618] & sel_one_hot_i[106];
  assign data_masked[13617] = data_i[13617] & sel_one_hot_i[106];
  assign data_masked[13616] = data_i[13616] & sel_one_hot_i[106];
  assign data_masked[13615] = data_i[13615] & sel_one_hot_i[106];
  assign data_masked[13614] = data_i[13614] & sel_one_hot_i[106];
  assign data_masked[13613] = data_i[13613] & sel_one_hot_i[106];
  assign data_masked[13612] = data_i[13612] & sel_one_hot_i[106];
  assign data_masked[13611] = data_i[13611] & sel_one_hot_i[106];
  assign data_masked[13610] = data_i[13610] & sel_one_hot_i[106];
  assign data_masked[13609] = data_i[13609] & sel_one_hot_i[106];
  assign data_masked[13608] = data_i[13608] & sel_one_hot_i[106];
  assign data_masked[13607] = data_i[13607] & sel_one_hot_i[106];
  assign data_masked[13606] = data_i[13606] & sel_one_hot_i[106];
  assign data_masked[13605] = data_i[13605] & sel_one_hot_i[106];
  assign data_masked[13604] = data_i[13604] & sel_one_hot_i[106];
  assign data_masked[13603] = data_i[13603] & sel_one_hot_i[106];
  assign data_masked[13602] = data_i[13602] & sel_one_hot_i[106];
  assign data_masked[13601] = data_i[13601] & sel_one_hot_i[106];
  assign data_masked[13600] = data_i[13600] & sel_one_hot_i[106];
  assign data_masked[13599] = data_i[13599] & sel_one_hot_i[106];
  assign data_masked[13598] = data_i[13598] & sel_one_hot_i[106];
  assign data_masked[13597] = data_i[13597] & sel_one_hot_i[106];
  assign data_masked[13596] = data_i[13596] & sel_one_hot_i[106];
  assign data_masked[13595] = data_i[13595] & sel_one_hot_i[106];
  assign data_masked[13594] = data_i[13594] & sel_one_hot_i[106];
  assign data_masked[13593] = data_i[13593] & sel_one_hot_i[106];
  assign data_masked[13592] = data_i[13592] & sel_one_hot_i[106];
  assign data_masked[13591] = data_i[13591] & sel_one_hot_i[106];
  assign data_masked[13590] = data_i[13590] & sel_one_hot_i[106];
  assign data_masked[13589] = data_i[13589] & sel_one_hot_i[106];
  assign data_masked[13588] = data_i[13588] & sel_one_hot_i[106];
  assign data_masked[13587] = data_i[13587] & sel_one_hot_i[106];
  assign data_masked[13586] = data_i[13586] & sel_one_hot_i[106];
  assign data_masked[13585] = data_i[13585] & sel_one_hot_i[106];
  assign data_masked[13584] = data_i[13584] & sel_one_hot_i[106];
  assign data_masked[13583] = data_i[13583] & sel_one_hot_i[106];
  assign data_masked[13582] = data_i[13582] & sel_one_hot_i[106];
  assign data_masked[13581] = data_i[13581] & sel_one_hot_i[106];
  assign data_masked[13580] = data_i[13580] & sel_one_hot_i[106];
  assign data_masked[13579] = data_i[13579] & sel_one_hot_i[106];
  assign data_masked[13578] = data_i[13578] & sel_one_hot_i[106];
  assign data_masked[13577] = data_i[13577] & sel_one_hot_i[106];
  assign data_masked[13576] = data_i[13576] & sel_one_hot_i[106];
  assign data_masked[13575] = data_i[13575] & sel_one_hot_i[106];
  assign data_masked[13574] = data_i[13574] & sel_one_hot_i[106];
  assign data_masked[13573] = data_i[13573] & sel_one_hot_i[106];
  assign data_masked[13572] = data_i[13572] & sel_one_hot_i[106];
  assign data_masked[13571] = data_i[13571] & sel_one_hot_i[106];
  assign data_masked[13570] = data_i[13570] & sel_one_hot_i[106];
  assign data_masked[13569] = data_i[13569] & sel_one_hot_i[106];
  assign data_masked[13568] = data_i[13568] & sel_one_hot_i[106];
  assign data_masked[13823] = data_i[13823] & sel_one_hot_i[107];
  assign data_masked[13822] = data_i[13822] & sel_one_hot_i[107];
  assign data_masked[13821] = data_i[13821] & sel_one_hot_i[107];
  assign data_masked[13820] = data_i[13820] & sel_one_hot_i[107];
  assign data_masked[13819] = data_i[13819] & sel_one_hot_i[107];
  assign data_masked[13818] = data_i[13818] & sel_one_hot_i[107];
  assign data_masked[13817] = data_i[13817] & sel_one_hot_i[107];
  assign data_masked[13816] = data_i[13816] & sel_one_hot_i[107];
  assign data_masked[13815] = data_i[13815] & sel_one_hot_i[107];
  assign data_masked[13814] = data_i[13814] & sel_one_hot_i[107];
  assign data_masked[13813] = data_i[13813] & sel_one_hot_i[107];
  assign data_masked[13812] = data_i[13812] & sel_one_hot_i[107];
  assign data_masked[13811] = data_i[13811] & sel_one_hot_i[107];
  assign data_masked[13810] = data_i[13810] & sel_one_hot_i[107];
  assign data_masked[13809] = data_i[13809] & sel_one_hot_i[107];
  assign data_masked[13808] = data_i[13808] & sel_one_hot_i[107];
  assign data_masked[13807] = data_i[13807] & sel_one_hot_i[107];
  assign data_masked[13806] = data_i[13806] & sel_one_hot_i[107];
  assign data_masked[13805] = data_i[13805] & sel_one_hot_i[107];
  assign data_masked[13804] = data_i[13804] & sel_one_hot_i[107];
  assign data_masked[13803] = data_i[13803] & sel_one_hot_i[107];
  assign data_masked[13802] = data_i[13802] & sel_one_hot_i[107];
  assign data_masked[13801] = data_i[13801] & sel_one_hot_i[107];
  assign data_masked[13800] = data_i[13800] & sel_one_hot_i[107];
  assign data_masked[13799] = data_i[13799] & sel_one_hot_i[107];
  assign data_masked[13798] = data_i[13798] & sel_one_hot_i[107];
  assign data_masked[13797] = data_i[13797] & sel_one_hot_i[107];
  assign data_masked[13796] = data_i[13796] & sel_one_hot_i[107];
  assign data_masked[13795] = data_i[13795] & sel_one_hot_i[107];
  assign data_masked[13794] = data_i[13794] & sel_one_hot_i[107];
  assign data_masked[13793] = data_i[13793] & sel_one_hot_i[107];
  assign data_masked[13792] = data_i[13792] & sel_one_hot_i[107];
  assign data_masked[13791] = data_i[13791] & sel_one_hot_i[107];
  assign data_masked[13790] = data_i[13790] & sel_one_hot_i[107];
  assign data_masked[13789] = data_i[13789] & sel_one_hot_i[107];
  assign data_masked[13788] = data_i[13788] & sel_one_hot_i[107];
  assign data_masked[13787] = data_i[13787] & sel_one_hot_i[107];
  assign data_masked[13786] = data_i[13786] & sel_one_hot_i[107];
  assign data_masked[13785] = data_i[13785] & sel_one_hot_i[107];
  assign data_masked[13784] = data_i[13784] & sel_one_hot_i[107];
  assign data_masked[13783] = data_i[13783] & sel_one_hot_i[107];
  assign data_masked[13782] = data_i[13782] & sel_one_hot_i[107];
  assign data_masked[13781] = data_i[13781] & sel_one_hot_i[107];
  assign data_masked[13780] = data_i[13780] & sel_one_hot_i[107];
  assign data_masked[13779] = data_i[13779] & sel_one_hot_i[107];
  assign data_masked[13778] = data_i[13778] & sel_one_hot_i[107];
  assign data_masked[13777] = data_i[13777] & sel_one_hot_i[107];
  assign data_masked[13776] = data_i[13776] & sel_one_hot_i[107];
  assign data_masked[13775] = data_i[13775] & sel_one_hot_i[107];
  assign data_masked[13774] = data_i[13774] & sel_one_hot_i[107];
  assign data_masked[13773] = data_i[13773] & sel_one_hot_i[107];
  assign data_masked[13772] = data_i[13772] & sel_one_hot_i[107];
  assign data_masked[13771] = data_i[13771] & sel_one_hot_i[107];
  assign data_masked[13770] = data_i[13770] & sel_one_hot_i[107];
  assign data_masked[13769] = data_i[13769] & sel_one_hot_i[107];
  assign data_masked[13768] = data_i[13768] & sel_one_hot_i[107];
  assign data_masked[13767] = data_i[13767] & sel_one_hot_i[107];
  assign data_masked[13766] = data_i[13766] & sel_one_hot_i[107];
  assign data_masked[13765] = data_i[13765] & sel_one_hot_i[107];
  assign data_masked[13764] = data_i[13764] & sel_one_hot_i[107];
  assign data_masked[13763] = data_i[13763] & sel_one_hot_i[107];
  assign data_masked[13762] = data_i[13762] & sel_one_hot_i[107];
  assign data_masked[13761] = data_i[13761] & sel_one_hot_i[107];
  assign data_masked[13760] = data_i[13760] & sel_one_hot_i[107];
  assign data_masked[13759] = data_i[13759] & sel_one_hot_i[107];
  assign data_masked[13758] = data_i[13758] & sel_one_hot_i[107];
  assign data_masked[13757] = data_i[13757] & sel_one_hot_i[107];
  assign data_masked[13756] = data_i[13756] & sel_one_hot_i[107];
  assign data_masked[13755] = data_i[13755] & sel_one_hot_i[107];
  assign data_masked[13754] = data_i[13754] & sel_one_hot_i[107];
  assign data_masked[13753] = data_i[13753] & sel_one_hot_i[107];
  assign data_masked[13752] = data_i[13752] & sel_one_hot_i[107];
  assign data_masked[13751] = data_i[13751] & sel_one_hot_i[107];
  assign data_masked[13750] = data_i[13750] & sel_one_hot_i[107];
  assign data_masked[13749] = data_i[13749] & sel_one_hot_i[107];
  assign data_masked[13748] = data_i[13748] & sel_one_hot_i[107];
  assign data_masked[13747] = data_i[13747] & sel_one_hot_i[107];
  assign data_masked[13746] = data_i[13746] & sel_one_hot_i[107];
  assign data_masked[13745] = data_i[13745] & sel_one_hot_i[107];
  assign data_masked[13744] = data_i[13744] & sel_one_hot_i[107];
  assign data_masked[13743] = data_i[13743] & sel_one_hot_i[107];
  assign data_masked[13742] = data_i[13742] & sel_one_hot_i[107];
  assign data_masked[13741] = data_i[13741] & sel_one_hot_i[107];
  assign data_masked[13740] = data_i[13740] & sel_one_hot_i[107];
  assign data_masked[13739] = data_i[13739] & sel_one_hot_i[107];
  assign data_masked[13738] = data_i[13738] & sel_one_hot_i[107];
  assign data_masked[13737] = data_i[13737] & sel_one_hot_i[107];
  assign data_masked[13736] = data_i[13736] & sel_one_hot_i[107];
  assign data_masked[13735] = data_i[13735] & sel_one_hot_i[107];
  assign data_masked[13734] = data_i[13734] & sel_one_hot_i[107];
  assign data_masked[13733] = data_i[13733] & sel_one_hot_i[107];
  assign data_masked[13732] = data_i[13732] & sel_one_hot_i[107];
  assign data_masked[13731] = data_i[13731] & sel_one_hot_i[107];
  assign data_masked[13730] = data_i[13730] & sel_one_hot_i[107];
  assign data_masked[13729] = data_i[13729] & sel_one_hot_i[107];
  assign data_masked[13728] = data_i[13728] & sel_one_hot_i[107];
  assign data_masked[13727] = data_i[13727] & sel_one_hot_i[107];
  assign data_masked[13726] = data_i[13726] & sel_one_hot_i[107];
  assign data_masked[13725] = data_i[13725] & sel_one_hot_i[107];
  assign data_masked[13724] = data_i[13724] & sel_one_hot_i[107];
  assign data_masked[13723] = data_i[13723] & sel_one_hot_i[107];
  assign data_masked[13722] = data_i[13722] & sel_one_hot_i[107];
  assign data_masked[13721] = data_i[13721] & sel_one_hot_i[107];
  assign data_masked[13720] = data_i[13720] & sel_one_hot_i[107];
  assign data_masked[13719] = data_i[13719] & sel_one_hot_i[107];
  assign data_masked[13718] = data_i[13718] & sel_one_hot_i[107];
  assign data_masked[13717] = data_i[13717] & sel_one_hot_i[107];
  assign data_masked[13716] = data_i[13716] & sel_one_hot_i[107];
  assign data_masked[13715] = data_i[13715] & sel_one_hot_i[107];
  assign data_masked[13714] = data_i[13714] & sel_one_hot_i[107];
  assign data_masked[13713] = data_i[13713] & sel_one_hot_i[107];
  assign data_masked[13712] = data_i[13712] & sel_one_hot_i[107];
  assign data_masked[13711] = data_i[13711] & sel_one_hot_i[107];
  assign data_masked[13710] = data_i[13710] & sel_one_hot_i[107];
  assign data_masked[13709] = data_i[13709] & sel_one_hot_i[107];
  assign data_masked[13708] = data_i[13708] & sel_one_hot_i[107];
  assign data_masked[13707] = data_i[13707] & sel_one_hot_i[107];
  assign data_masked[13706] = data_i[13706] & sel_one_hot_i[107];
  assign data_masked[13705] = data_i[13705] & sel_one_hot_i[107];
  assign data_masked[13704] = data_i[13704] & sel_one_hot_i[107];
  assign data_masked[13703] = data_i[13703] & sel_one_hot_i[107];
  assign data_masked[13702] = data_i[13702] & sel_one_hot_i[107];
  assign data_masked[13701] = data_i[13701] & sel_one_hot_i[107];
  assign data_masked[13700] = data_i[13700] & sel_one_hot_i[107];
  assign data_masked[13699] = data_i[13699] & sel_one_hot_i[107];
  assign data_masked[13698] = data_i[13698] & sel_one_hot_i[107];
  assign data_masked[13697] = data_i[13697] & sel_one_hot_i[107];
  assign data_masked[13696] = data_i[13696] & sel_one_hot_i[107];
  assign data_masked[13951] = data_i[13951] & sel_one_hot_i[108];
  assign data_masked[13950] = data_i[13950] & sel_one_hot_i[108];
  assign data_masked[13949] = data_i[13949] & sel_one_hot_i[108];
  assign data_masked[13948] = data_i[13948] & sel_one_hot_i[108];
  assign data_masked[13947] = data_i[13947] & sel_one_hot_i[108];
  assign data_masked[13946] = data_i[13946] & sel_one_hot_i[108];
  assign data_masked[13945] = data_i[13945] & sel_one_hot_i[108];
  assign data_masked[13944] = data_i[13944] & sel_one_hot_i[108];
  assign data_masked[13943] = data_i[13943] & sel_one_hot_i[108];
  assign data_masked[13942] = data_i[13942] & sel_one_hot_i[108];
  assign data_masked[13941] = data_i[13941] & sel_one_hot_i[108];
  assign data_masked[13940] = data_i[13940] & sel_one_hot_i[108];
  assign data_masked[13939] = data_i[13939] & sel_one_hot_i[108];
  assign data_masked[13938] = data_i[13938] & sel_one_hot_i[108];
  assign data_masked[13937] = data_i[13937] & sel_one_hot_i[108];
  assign data_masked[13936] = data_i[13936] & sel_one_hot_i[108];
  assign data_masked[13935] = data_i[13935] & sel_one_hot_i[108];
  assign data_masked[13934] = data_i[13934] & sel_one_hot_i[108];
  assign data_masked[13933] = data_i[13933] & sel_one_hot_i[108];
  assign data_masked[13932] = data_i[13932] & sel_one_hot_i[108];
  assign data_masked[13931] = data_i[13931] & sel_one_hot_i[108];
  assign data_masked[13930] = data_i[13930] & sel_one_hot_i[108];
  assign data_masked[13929] = data_i[13929] & sel_one_hot_i[108];
  assign data_masked[13928] = data_i[13928] & sel_one_hot_i[108];
  assign data_masked[13927] = data_i[13927] & sel_one_hot_i[108];
  assign data_masked[13926] = data_i[13926] & sel_one_hot_i[108];
  assign data_masked[13925] = data_i[13925] & sel_one_hot_i[108];
  assign data_masked[13924] = data_i[13924] & sel_one_hot_i[108];
  assign data_masked[13923] = data_i[13923] & sel_one_hot_i[108];
  assign data_masked[13922] = data_i[13922] & sel_one_hot_i[108];
  assign data_masked[13921] = data_i[13921] & sel_one_hot_i[108];
  assign data_masked[13920] = data_i[13920] & sel_one_hot_i[108];
  assign data_masked[13919] = data_i[13919] & sel_one_hot_i[108];
  assign data_masked[13918] = data_i[13918] & sel_one_hot_i[108];
  assign data_masked[13917] = data_i[13917] & sel_one_hot_i[108];
  assign data_masked[13916] = data_i[13916] & sel_one_hot_i[108];
  assign data_masked[13915] = data_i[13915] & sel_one_hot_i[108];
  assign data_masked[13914] = data_i[13914] & sel_one_hot_i[108];
  assign data_masked[13913] = data_i[13913] & sel_one_hot_i[108];
  assign data_masked[13912] = data_i[13912] & sel_one_hot_i[108];
  assign data_masked[13911] = data_i[13911] & sel_one_hot_i[108];
  assign data_masked[13910] = data_i[13910] & sel_one_hot_i[108];
  assign data_masked[13909] = data_i[13909] & sel_one_hot_i[108];
  assign data_masked[13908] = data_i[13908] & sel_one_hot_i[108];
  assign data_masked[13907] = data_i[13907] & sel_one_hot_i[108];
  assign data_masked[13906] = data_i[13906] & sel_one_hot_i[108];
  assign data_masked[13905] = data_i[13905] & sel_one_hot_i[108];
  assign data_masked[13904] = data_i[13904] & sel_one_hot_i[108];
  assign data_masked[13903] = data_i[13903] & sel_one_hot_i[108];
  assign data_masked[13902] = data_i[13902] & sel_one_hot_i[108];
  assign data_masked[13901] = data_i[13901] & sel_one_hot_i[108];
  assign data_masked[13900] = data_i[13900] & sel_one_hot_i[108];
  assign data_masked[13899] = data_i[13899] & sel_one_hot_i[108];
  assign data_masked[13898] = data_i[13898] & sel_one_hot_i[108];
  assign data_masked[13897] = data_i[13897] & sel_one_hot_i[108];
  assign data_masked[13896] = data_i[13896] & sel_one_hot_i[108];
  assign data_masked[13895] = data_i[13895] & sel_one_hot_i[108];
  assign data_masked[13894] = data_i[13894] & sel_one_hot_i[108];
  assign data_masked[13893] = data_i[13893] & sel_one_hot_i[108];
  assign data_masked[13892] = data_i[13892] & sel_one_hot_i[108];
  assign data_masked[13891] = data_i[13891] & sel_one_hot_i[108];
  assign data_masked[13890] = data_i[13890] & sel_one_hot_i[108];
  assign data_masked[13889] = data_i[13889] & sel_one_hot_i[108];
  assign data_masked[13888] = data_i[13888] & sel_one_hot_i[108];
  assign data_masked[13887] = data_i[13887] & sel_one_hot_i[108];
  assign data_masked[13886] = data_i[13886] & sel_one_hot_i[108];
  assign data_masked[13885] = data_i[13885] & sel_one_hot_i[108];
  assign data_masked[13884] = data_i[13884] & sel_one_hot_i[108];
  assign data_masked[13883] = data_i[13883] & sel_one_hot_i[108];
  assign data_masked[13882] = data_i[13882] & sel_one_hot_i[108];
  assign data_masked[13881] = data_i[13881] & sel_one_hot_i[108];
  assign data_masked[13880] = data_i[13880] & sel_one_hot_i[108];
  assign data_masked[13879] = data_i[13879] & sel_one_hot_i[108];
  assign data_masked[13878] = data_i[13878] & sel_one_hot_i[108];
  assign data_masked[13877] = data_i[13877] & sel_one_hot_i[108];
  assign data_masked[13876] = data_i[13876] & sel_one_hot_i[108];
  assign data_masked[13875] = data_i[13875] & sel_one_hot_i[108];
  assign data_masked[13874] = data_i[13874] & sel_one_hot_i[108];
  assign data_masked[13873] = data_i[13873] & sel_one_hot_i[108];
  assign data_masked[13872] = data_i[13872] & sel_one_hot_i[108];
  assign data_masked[13871] = data_i[13871] & sel_one_hot_i[108];
  assign data_masked[13870] = data_i[13870] & sel_one_hot_i[108];
  assign data_masked[13869] = data_i[13869] & sel_one_hot_i[108];
  assign data_masked[13868] = data_i[13868] & sel_one_hot_i[108];
  assign data_masked[13867] = data_i[13867] & sel_one_hot_i[108];
  assign data_masked[13866] = data_i[13866] & sel_one_hot_i[108];
  assign data_masked[13865] = data_i[13865] & sel_one_hot_i[108];
  assign data_masked[13864] = data_i[13864] & sel_one_hot_i[108];
  assign data_masked[13863] = data_i[13863] & sel_one_hot_i[108];
  assign data_masked[13862] = data_i[13862] & sel_one_hot_i[108];
  assign data_masked[13861] = data_i[13861] & sel_one_hot_i[108];
  assign data_masked[13860] = data_i[13860] & sel_one_hot_i[108];
  assign data_masked[13859] = data_i[13859] & sel_one_hot_i[108];
  assign data_masked[13858] = data_i[13858] & sel_one_hot_i[108];
  assign data_masked[13857] = data_i[13857] & sel_one_hot_i[108];
  assign data_masked[13856] = data_i[13856] & sel_one_hot_i[108];
  assign data_masked[13855] = data_i[13855] & sel_one_hot_i[108];
  assign data_masked[13854] = data_i[13854] & sel_one_hot_i[108];
  assign data_masked[13853] = data_i[13853] & sel_one_hot_i[108];
  assign data_masked[13852] = data_i[13852] & sel_one_hot_i[108];
  assign data_masked[13851] = data_i[13851] & sel_one_hot_i[108];
  assign data_masked[13850] = data_i[13850] & sel_one_hot_i[108];
  assign data_masked[13849] = data_i[13849] & sel_one_hot_i[108];
  assign data_masked[13848] = data_i[13848] & sel_one_hot_i[108];
  assign data_masked[13847] = data_i[13847] & sel_one_hot_i[108];
  assign data_masked[13846] = data_i[13846] & sel_one_hot_i[108];
  assign data_masked[13845] = data_i[13845] & sel_one_hot_i[108];
  assign data_masked[13844] = data_i[13844] & sel_one_hot_i[108];
  assign data_masked[13843] = data_i[13843] & sel_one_hot_i[108];
  assign data_masked[13842] = data_i[13842] & sel_one_hot_i[108];
  assign data_masked[13841] = data_i[13841] & sel_one_hot_i[108];
  assign data_masked[13840] = data_i[13840] & sel_one_hot_i[108];
  assign data_masked[13839] = data_i[13839] & sel_one_hot_i[108];
  assign data_masked[13838] = data_i[13838] & sel_one_hot_i[108];
  assign data_masked[13837] = data_i[13837] & sel_one_hot_i[108];
  assign data_masked[13836] = data_i[13836] & sel_one_hot_i[108];
  assign data_masked[13835] = data_i[13835] & sel_one_hot_i[108];
  assign data_masked[13834] = data_i[13834] & sel_one_hot_i[108];
  assign data_masked[13833] = data_i[13833] & sel_one_hot_i[108];
  assign data_masked[13832] = data_i[13832] & sel_one_hot_i[108];
  assign data_masked[13831] = data_i[13831] & sel_one_hot_i[108];
  assign data_masked[13830] = data_i[13830] & sel_one_hot_i[108];
  assign data_masked[13829] = data_i[13829] & sel_one_hot_i[108];
  assign data_masked[13828] = data_i[13828] & sel_one_hot_i[108];
  assign data_masked[13827] = data_i[13827] & sel_one_hot_i[108];
  assign data_masked[13826] = data_i[13826] & sel_one_hot_i[108];
  assign data_masked[13825] = data_i[13825] & sel_one_hot_i[108];
  assign data_masked[13824] = data_i[13824] & sel_one_hot_i[108];
  assign data_masked[14079] = data_i[14079] & sel_one_hot_i[109];
  assign data_masked[14078] = data_i[14078] & sel_one_hot_i[109];
  assign data_masked[14077] = data_i[14077] & sel_one_hot_i[109];
  assign data_masked[14076] = data_i[14076] & sel_one_hot_i[109];
  assign data_masked[14075] = data_i[14075] & sel_one_hot_i[109];
  assign data_masked[14074] = data_i[14074] & sel_one_hot_i[109];
  assign data_masked[14073] = data_i[14073] & sel_one_hot_i[109];
  assign data_masked[14072] = data_i[14072] & sel_one_hot_i[109];
  assign data_masked[14071] = data_i[14071] & sel_one_hot_i[109];
  assign data_masked[14070] = data_i[14070] & sel_one_hot_i[109];
  assign data_masked[14069] = data_i[14069] & sel_one_hot_i[109];
  assign data_masked[14068] = data_i[14068] & sel_one_hot_i[109];
  assign data_masked[14067] = data_i[14067] & sel_one_hot_i[109];
  assign data_masked[14066] = data_i[14066] & sel_one_hot_i[109];
  assign data_masked[14065] = data_i[14065] & sel_one_hot_i[109];
  assign data_masked[14064] = data_i[14064] & sel_one_hot_i[109];
  assign data_masked[14063] = data_i[14063] & sel_one_hot_i[109];
  assign data_masked[14062] = data_i[14062] & sel_one_hot_i[109];
  assign data_masked[14061] = data_i[14061] & sel_one_hot_i[109];
  assign data_masked[14060] = data_i[14060] & sel_one_hot_i[109];
  assign data_masked[14059] = data_i[14059] & sel_one_hot_i[109];
  assign data_masked[14058] = data_i[14058] & sel_one_hot_i[109];
  assign data_masked[14057] = data_i[14057] & sel_one_hot_i[109];
  assign data_masked[14056] = data_i[14056] & sel_one_hot_i[109];
  assign data_masked[14055] = data_i[14055] & sel_one_hot_i[109];
  assign data_masked[14054] = data_i[14054] & sel_one_hot_i[109];
  assign data_masked[14053] = data_i[14053] & sel_one_hot_i[109];
  assign data_masked[14052] = data_i[14052] & sel_one_hot_i[109];
  assign data_masked[14051] = data_i[14051] & sel_one_hot_i[109];
  assign data_masked[14050] = data_i[14050] & sel_one_hot_i[109];
  assign data_masked[14049] = data_i[14049] & sel_one_hot_i[109];
  assign data_masked[14048] = data_i[14048] & sel_one_hot_i[109];
  assign data_masked[14047] = data_i[14047] & sel_one_hot_i[109];
  assign data_masked[14046] = data_i[14046] & sel_one_hot_i[109];
  assign data_masked[14045] = data_i[14045] & sel_one_hot_i[109];
  assign data_masked[14044] = data_i[14044] & sel_one_hot_i[109];
  assign data_masked[14043] = data_i[14043] & sel_one_hot_i[109];
  assign data_masked[14042] = data_i[14042] & sel_one_hot_i[109];
  assign data_masked[14041] = data_i[14041] & sel_one_hot_i[109];
  assign data_masked[14040] = data_i[14040] & sel_one_hot_i[109];
  assign data_masked[14039] = data_i[14039] & sel_one_hot_i[109];
  assign data_masked[14038] = data_i[14038] & sel_one_hot_i[109];
  assign data_masked[14037] = data_i[14037] & sel_one_hot_i[109];
  assign data_masked[14036] = data_i[14036] & sel_one_hot_i[109];
  assign data_masked[14035] = data_i[14035] & sel_one_hot_i[109];
  assign data_masked[14034] = data_i[14034] & sel_one_hot_i[109];
  assign data_masked[14033] = data_i[14033] & sel_one_hot_i[109];
  assign data_masked[14032] = data_i[14032] & sel_one_hot_i[109];
  assign data_masked[14031] = data_i[14031] & sel_one_hot_i[109];
  assign data_masked[14030] = data_i[14030] & sel_one_hot_i[109];
  assign data_masked[14029] = data_i[14029] & sel_one_hot_i[109];
  assign data_masked[14028] = data_i[14028] & sel_one_hot_i[109];
  assign data_masked[14027] = data_i[14027] & sel_one_hot_i[109];
  assign data_masked[14026] = data_i[14026] & sel_one_hot_i[109];
  assign data_masked[14025] = data_i[14025] & sel_one_hot_i[109];
  assign data_masked[14024] = data_i[14024] & sel_one_hot_i[109];
  assign data_masked[14023] = data_i[14023] & sel_one_hot_i[109];
  assign data_masked[14022] = data_i[14022] & sel_one_hot_i[109];
  assign data_masked[14021] = data_i[14021] & sel_one_hot_i[109];
  assign data_masked[14020] = data_i[14020] & sel_one_hot_i[109];
  assign data_masked[14019] = data_i[14019] & sel_one_hot_i[109];
  assign data_masked[14018] = data_i[14018] & sel_one_hot_i[109];
  assign data_masked[14017] = data_i[14017] & sel_one_hot_i[109];
  assign data_masked[14016] = data_i[14016] & sel_one_hot_i[109];
  assign data_masked[14015] = data_i[14015] & sel_one_hot_i[109];
  assign data_masked[14014] = data_i[14014] & sel_one_hot_i[109];
  assign data_masked[14013] = data_i[14013] & sel_one_hot_i[109];
  assign data_masked[14012] = data_i[14012] & sel_one_hot_i[109];
  assign data_masked[14011] = data_i[14011] & sel_one_hot_i[109];
  assign data_masked[14010] = data_i[14010] & sel_one_hot_i[109];
  assign data_masked[14009] = data_i[14009] & sel_one_hot_i[109];
  assign data_masked[14008] = data_i[14008] & sel_one_hot_i[109];
  assign data_masked[14007] = data_i[14007] & sel_one_hot_i[109];
  assign data_masked[14006] = data_i[14006] & sel_one_hot_i[109];
  assign data_masked[14005] = data_i[14005] & sel_one_hot_i[109];
  assign data_masked[14004] = data_i[14004] & sel_one_hot_i[109];
  assign data_masked[14003] = data_i[14003] & sel_one_hot_i[109];
  assign data_masked[14002] = data_i[14002] & sel_one_hot_i[109];
  assign data_masked[14001] = data_i[14001] & sel_one_hot_i[109];
  assign data_masked[14000] = data_i[14000] & sel_one_hot_i[109];
  assign data_masked[13999] = data_i[13999] & sel_one_hot_i[109];
  assign data_masked[13998] = data_i[13998] & sel_one_hot_i[109];
  assign data_masked[13997] = data_i[13997] & sel_one_hot_i[109];
  assign data_masked[13996] = data_i[13996] & sel_one_hot_i[109];
  assign data_masked[13995] = data_i[13995] & sel_one_hot_i[109];
  assign data_masked[13994] = data_i[13994] & sel_one_hot_i[109];
  assign data_masked[13993] = data_i[13993] & sel_one_hot_i[109];
  assign data_masked[13992] = data_i[13992] & sel_one_hot_i[109];
  assign data_masked[13991] = data_i[13991] & sel_one_hot_i[109];
  assign data_masked[13990] = data_i[13990] & sel_one_hot_i[109];
  assign data_masked[13989] = data_i[13989] & sel_one_hot_i[109];
  assign data_masked[13988] = data_i[13988] & sel_one_hot_i[109];
  assign data_masked[13987] = data_i[13987] & sel_one_hot_i[109];
  assign data_masked[13986] = data_i[13986] & sel_one_hot_i[109];
  assign data_masked[13985] = data_i[13985] & sel_one_hot_i[109];
  assign data_masked[13984] = data_i[13984] & sel_one_hot_i[109];
  assign data_masked[13983] = data_i[13983] & sel_one_hot_i[109];
  assign data_masked[13982] = data_i[13982] & sel_one_hot_i[109];
  assign data_masked[13981] = data_i[13981] & sel_one_hot_i[109];
  assign data_masked[13980] = data_i[13980] & sel_one_hot_i[109];
  assign data_masked[13979] = data_i[13979] & sel_one_hot_i[109];
  assign data_masked[13978] = data_i[13978] & sel_one_hot_i[109];
  assign data_masked[13977] = data_i[13977] & sel_one_hot_i[109];
  assign data_masked[13976] = data_i[13976] & sel_one_hot_i[109];
  assign data_masked[13975] = data_i[13975] & sel_one_hot_i[109];
  assign data_masked[13974] = data_i[13974] & sel_one_hot_i[109];
  assign data_masked[13973] = data_i[13973] & sel_one_hot_i[109];
  assign data_masked[13972] = data_i[13972] & sel_one_hot_i[109];
  assign data_masked[13971] = data_i[13971] & sel_one_hot_i[109];
  assign data_masked[13970] = data_i[13970] & sel_one_hot_i[109];
  assign data_masked[13969] = data_i[13969] & sel_one_hot_i[109];
  assign data_masked[13968] = data_i[13968] & sel_one_hot_i[109];
  assign data_masked[13967] = data_i[13967] & sel_one_hot_i[109];
  assign data_masked[13966] = data_i[13966] & sel_one_hot_i[109];
  assign data_masked[13965] = data_i[13965] & sel_one_hot_i[109];
  assign data_masked[13964] = data_i[13964] & sel_one_hot_i[109];
  assign data_masked[13963] = data_i[13963] & sel_one_hot_i[109];
  assign data_masked[13962] = data_i[13962] & sel_one_hot_i[109];
  assign data_masked[13961] = data_i[13961] & sel_one_hot_i[109];
  assign data_masked[13960] = data_i[13960] & sel_one_hot_i[109];
  assign data_masked[13959] = data_i[13959] & sel_one_hot_i[109];
  assign data_masked[13958] = data_i[13958] & sel_one_hot_i[109];
  assign data_masked[13957] = data_i[13957] & sel_one_hot_i[109];
  assign data_masked[13956] = data_i[13956] & sel_one_hot_i[109];
  assign data_masked[13955] = data_i[13955] & sel_one_hot_i[109];
  assign data_masked[13954] = data_i[13954] & sel_one_hot_i[109];
  assign data_masked[13953] = data_i[13953] & sel_one_hot_i[109];
  assign data_masked[13952] = data_i[13952] & sel_one_hot_i[109];
  assign data_masked[14207] = data_i[14207] & sel_one_hot_i[110];
  assign data_masked[14206] = data_i[14206] & sel_one_hot_i[110];
  assign data_masked[14205] = data_i[14205] & sel_one_hot_i[110];
  assign data_masked[14204] = data_i[14204] & sel_one_hot_i[110];
  assign data_masked[14203] = data_i[14203] & sel_one_hot_i[110];
  assign data_masked[14202] = data_i[14202] & sel_one_hot_i[110];
  assign data_masked[14201] = data_i[14201] & sel_one_hot_i[110];
  assign data_masked[14200] = data_i[14200] & sel_one_hot_i[110];
  assign data_masked[14199] = data_i[14199] & sel_one_hot_i[110];
  assign data_masked[14198] = data_i[14198] & sel_one_hot_i[110];
  assign data_masked[14197] = data_i[14197] & sel_one_hot_i[110];
  assign data_masked[14196] = data_i[14196] & sel_one_hot_i[110];
  assign data_masked[14195] = data_i[14195] & sel_one_hot_i[110];
  assign data_masked[14194] = data_i[14194] & sel_one_hot_i[110];
  assign data_masked[14193] = data_i[14193] & sel_one_hot_i[110];
  assign data_masked[14192] = data_i[14192] & sel_one_hot_i[110];
  assign data_masked[14191] = data_i[14191] & sel_one_hot_i[110];
  assign data_masked[14190] = data_i[14190] & sel_one_hot_i[110];
  assign data_masked[14189] = data_i[14189] & sel_one_hot_i[110];
  assign data_masked[14188] = data_i[14188] & sel_one_hot_i[110];
  assign data_masked[14187] = data_i[14187] & sel_one_hot_i[110];
  assign data_masked[14186] = data_i[14186] & sel_one_hot_i[110];
  assign data_masked[14185] = data_i[14185] & sel_one_hot_i[110];
  assign data_masked[14184] = data_i[14184] & sel_one_hot_i[110];
  assign data_masked[14183] = data_i[14183] & sel_one_hot_i[110];
  assign data_masked[14182] = data_i[14182] & sel_one_hot_i[110];
  assign data_masked[14181] = data_i[14181] & sel_one_hot_i[110];
  assign data_masked[14180] = data_i[14180] & sel_one_hot_i[110];
  assign data_masked[14179] = data_i[14179] & sel_one_hot_i[110];
  assign data_masked[14178] = data_i[14178] & sel_one_hot_i[110];
  assign data_masked[14177] = data_i[14177] & sel_one_hot_i[110];
  assign data_masked[14176] = data_i[14176] & sel_one_hot_i[110];
  assign data_masked[14175] = data_i[14175] & sel_one_hot_i[110];
  assign data_masked[14174] = data_i[14174] & sel_one_hot_i[110];
  assign data_masked[14173] = data_i[14173] & sel_one_hot_i[110];
  assign data_masked[14172] = data_i[14172] & sel_one_hot_i[110];
  assign data_masked[14171] = data_i[14171] & sel_one_hot_i[110];
  assign data_masked[14170] = data_i[14170] & sel_one_hot_i[110];
  assign data_masked[14169] = data_i[14169] & sel_one_hot_i[110];
  assign data_masked[14168] = data_i[14168] & sel_one_hot_i[110];
  assign data_masked[14167] = data_i[14167] & sel_one_hot_i[110];
  assign data_masked[14166] = data_i[14166] & sel_one_hot_i[110];
  assign data_masked[14165] = data_i[14165] & sel_one_hot_i[110];
  assign data_masked[14164] = data_i[14164] & sel_one_hot_i[110];
  assign data_masked[14163] = data_i[14163] & sel_one_hot_i[110];
  assign data_masked[14162] = data_i[14162] & sel_one_hot_i[110];
  assign data_masked[14161] = data_i[14161] & sel_one_hot_i[110];
  assign data_masked[14160] = data_i[14160] & sel_one_hot_i[110];
  assign data_masked[14159] = data_i[14159] & sel_one_hot_i[110];
  assign data_masked[14158] = data_i[14158] & sel_one_hot_i[110];
  assign data_masked[14157] = data_i[14157] & sel_one_hot_i[110];
  assign data_masked[14156] = data_i[14156] & sel_one_hot_i[110];
  assign data_masked[14155] = data_i[14155] & sel_one_hot_i[110];
  assign data_masked[14154] = data_i[14154] & sel_one_hot_i[110];
  assign data_masked[14153] = data_i[14153] & sel_one_hot_i[110];
  assign data_masked[14152] = data_i[14152] & sel_one_hot_i[110];
  assign data_masked[14151] = data_i[14151] & sel_one_hot_i[110];
  assign data_masked[14150] = data_i[14150] & sel_one_hot_i[110];
  assign data_masked[14149] = data_i[14149] & sel_one_hot_i[110];
  assign data_masked[14148] = data_i[14148] & sel_one_hot_i[110];
  assign data_masked[14147] = data_i[14147] & sel_one_hot_i[110];
  assign data_masked[14146] = data_i[14146] & sel_one_hot_i[110];
  assign data_masked[14145] = data_i[14145] & sel_one_hot_i[110];
  assign data_masked[14144] = data_i[14144] & sel_one_hot_i[110];
  assign data_masked[14143] = data_i[14143] & sel_one_hot_i[110];
  assign data_masked[14142] = data_i[14142] & sel_one_hot_i[110];
  assign data_masked[14141] = data_i[14141] & sel_one_hot_i[110];
  assign data_masked[14140] = data_i[14140] & sel_one_hot_i[110];
  assign data_masked[14139] = data_i[14139] & sel_one_hot_i[110];
  assign data_masked[14138] = data_i[14138] & sel_one_hot_i[110];
  assign data_masked[14137] = data_i[14137] & sel_one_hot_i[110];
  assign data_masked[14136] = data_i[14136] & sel_one_hot_i[110];
  assign data_masked[14135] = data_i[14135] & sel_one_hot_i[110];
  assign data_masked[14134] = data_i[14134] & sel_one_hot_i[110];
  assign data_masked[14133] = data_i[14133] & sel_one_hot_i[110];
  assign data_masked[14132] = data_i[14132] & sel_one_hot_i[110];
  assign data_masked[14131] = data_i[14131] & sel_one_hot_i[110];
  assign data_masked[14130] = data_i[14130] & sel_one_hot_i[110];
  assign data_masked[14129] = data_i[14129] & sel_one_hot_i[110];
  assign data_masked[14128] = data_i[14128] & sel_one_hot_i[110];
  assign data_masked[14127] = data_i[14127] & sel_one_hot_i[110];
  assign data_masked[14126] = data_i[14126] & sel_one_hot_i[110];
  assign data_masked[14125] = data_i[14125] & sel_one_hot_i[110];
  assign data_masked[14124] = data_i[14124] & sel_one_hot_i[110];
  assign data_masked[14123] = data_i[14123] & sel_one_hot_i[110];
  assign data_masked[14122] = data_i[14122] & sel_one_hot_i[110];
  assign data_masked[14121] = data_i[14121] & sel_one_hot_i[110];
  assign data_masked[14120] = data_i[14120] & sel_one_hot_i[110];
  assign data_masked[14119] = data_i[14119] & sel_one_hot_i[110];
  assign data_masked[14118] = data_i[14118] & sel_one_hot_i[110];
  assign data_masked[14117] = data_i[14117] & sel_one_hot_i[110];
  assign data_masked[14116] = data_i[14116] & sel_one_hot_i[110];
  assign data_masked[14115] = data_i[14115] & sel_one_hot_i[110];
  assign data_masked[14114] = data_i[14114] & sel_one_hot_i[110];
  assign data_masked[14113] = data_i[14113] & sel_one_hot_i[110];
  assign data_masked[14112] = data_i[14112] & sel_one_hot_i[110];
  assign data_masked[14111] = data_i[14111] & sel_one_hot_i[110];
  assign data_masked[14110] = data_i[14110] & sel_one_hot_i[110];
  assign data_masked[14109] = data_i[14109] & sel_one_hot_i[110];
  assign data_masked[14108] = data_i[14108] & sel_one_hot_i[110];
  assign data_masked[14107] = data_i[14107] & sel_one_hot_i[110];
  assign data_masked[14106] = data_i[14106] & sel_one_hot_i[110];
  assign data_masked[14105] = data_i[14105] & sel_one_hot_i[110];
  assign data_masked[14104] = data_i[14104] & sel_one_hot_i[110];
  assign data_masked[14103] = data_i[14103] & sel_one_hot_i[110];
  assign data_masked[14102] = data_i[14102] & sel_one_hot_i[110];
  assign data_masked[14101] = data_i[14101] & sel_one_hot_i[110];
  assign data_masked[14100] = data_i[14100] & sel_one_hot_i[110];
  assign data_masked[14099] = data_i[14099] & sel_one_hot_i[110];
  assign data_masked[14098] = data_i[14098] & sel_one_hot_i[110];
  assign data_masked[14097] = data_i[14097] & sel_one_hot_i[110];
  assign data_masked[14096] = data_i[14096] & sel_one_hot_i[110];
  assign data_masked[14095] = data_i[14095] & sel_one_hot_i[110];
  assign data_masked[14094] = data_i[14094] & sel_one_hot_i[110];
  assign data_masked[14093] = data_i[14093] & sel_one_hot_i[110];
  assign data_masked[14092] = data_i[14092] & sel_one_hot_i[110];
  assign data_masked[14091] = data_i[14091] & sel_one_hot_i[110];
  assign data_masked[14090] = data_i[14090] & sel_one_hot_i[110];
  assign data_masked[14089] = data_i[14089] & sel_one_hot_i[110];
  assign data_masked[14088] = data_i[14088] & sel_one_hot_i[110];
  assign data_masked[14087] = data_i[14087] & sel_one_hot_i[110];
  assign data_masked[14086] = data_i[14086] & sel_one_hot_i[110];
  assign data_masked[14085] = data_i[14085] & sel_one_hot_i[110];
  assign data_masked[14084] = data_i[14084] & sel_one_hot_i[110];
  assign data_masked[14083] = data_i[14083] & sel_one_hot_i[110];
  assign data_masked[14082] = data_i[14082] & sel_one_hot_i[110];
  assign data_masked[14081] = data_i[14081] & sel_one_hot_i[110];
  assign data_masked[14080] = data_i[14080] & sel_one_hot_i[110];
  assign data_masked[14335] = data_i[14335] & sel_one_hot_i[111];
  assign data_masked[14334] = data_i[14334] & sel_one_hot_i[111];
  assign data_masked[14333] = data_i[14333] & sel_one_hot_i[111];
  assign data_masked[14332] = data_i[14332] & sel_one_hot_i[111];
  assign data_masked[14331] = data_i[14331] & sel_one_hot_i[111];
  assign data_masked[14330] = data_i[14330] & sel_one_hot_i[111];
  assign data_masked[14329] = data_i[14329] & sel_one_hot_i[111];
  assign data_masked[14328] = data_i[14328] & sel_one_hot_i[111];
  assign data_masked[14327] = data_i[14327] & sel_one_hot_i[111];
  assign data_masked[14326] = data_i[14326] & sel_one_hot_i[111];
  assign data_masked[14325] = data_i[14325] & sel_one_hot_i[111];
  assign data_masked[14324] = data_i[14324] & sel_one_hot_i[111];
  assign data_masked[14323] = data_i[14323] & sel_one_hot_i[111];
  assign data_masked[14322] = data_i[14322] & sel_one_hot_i[111];
  assign data_masked[14321] = data_i[14321] & sel_one_hot_i[111];
  assign data_masked[14320] = data_i[14320] & sel_one_hot_i[111];
  assign data_masked[14319] = data_i[14319] & sel_one_hot_i[111];
  assign data_masked[14318] = data_i[14318] & sel_one_hot_i[111];
  assign data_masked[14317] = data_i[14317] & sel_one_hot_i[111];
  assign data_masked[14316] = data_i[14316] & sel_one_hot_i[111];
  assign data_masked[14315] = data_i[14315] & sel_one_hot_i[111];
  assign data_masked[14314] = data_i[14314] & sel_one_hot_i[111];
  assign data_masked[14313] = data_i[14313] & sel_one_hot_i[111];
  assign data_masked[14312] = data_i[14312] & sel_one_hot_i[111];
  assign data_masked[14311] = data_i[14311] & sel_one_hot_i[111];
  assign data_masked[14310] = data_i[14310] & sel_one_hot_i[111];
  assign data_masked[14309] = data_i[14309] & sel_one_hot_i[111];
  assign data_masked[14308] = data_i[14308] & sel_one_hot_i[111];
  assign data_masked[14307] = data_i[14307] & sel_one_hot_i[111];
  assign data_masked[14306] = data_i[14306] & sel_one_hot_i[111];
  assign data_masked[14305] = data_i[14305] & sel_one_hot_i[111];
  assign data_masked[14304] = data_i[14304] & sel_one_hot_i[111];
  assign data_masked[14303] = data_i[14303] & sel_one_hot_i[111];
  assign data_masked[14302] = data_i[14302] & sel_one_hot_i[111];
  assign data_masked[14301] = data_i[14301] & sel_one_hot_i[111];
  assign data_masked[14300] = data_i[14300] & sel_one_hot_i[111];
  assign data_masked[14299] = data_i[14299] & sel_one_hot_i[111];
  assign data_masked[14298] = data_i[14298] & sel_one_hot_i[111];
  assign data_masked[14297] = data_i[14297] & sel_one_hot_i[111];
  assign data_masked[14296] = data_i[14296] & sel_one_hot_i[111];
  assign data_masked[14295] = data_i[14295] & sel_one_hot_i[111];
  assign data_masked[14294] = data_i[14294] & sel_one_hot_i[111];
  assign data_masked[14293] = data_i[14293] & sel_one_hot_i[111];
  assign data_masked[14292] = data_i[14292] & sel_one_hot_i[111];
  assign data_masked[14291] = data_i[14291] & sel_one_hot_i[111];
  assign data_masked[14290] = data_i[14290] & sel_one_hot_i[111];
  assign data_masked[14289] = data_i[14289] & sel_one_hot_i[111];
  assign data_masked[14288] = data_i[14288] & sel_one_hot_i[111];
  assign data_masked[14287] = data_i[14287] & sel_one_hot_i[111];
  assign data_masked[14286] = data_i[14286] & sel_one_hot_i[111];
  assign data_masked[14285] = data_i[14285] & sel_one_hot_i[111];
  assign data_masked[14284] = data_i[14284] & sel_one_hot_i[111];
  assign data_masked[14283] = data_i[14283] & sel_one_hot_i[111];
  assign data_masked[14282] = data_i[14282] & sel_one_hot_i[111];
  assign data_masked[14281] = data_i[14281] & sel_one_hot_i[111];
  assign data_masked[14280] = data_i[14280] & sel_one_hot_i[111];
  assign data_masked[14279] = data_i[14279] & sel_one_hot_i[111];
  assign data_masked[14278] = data_i[14278] & sel_one_hot_i[111];
  assign data_masked[14277] = data_i[14277] & sel_one_hot_i[111];
  assign data_masked[14276] = data_i[14276] & sel_one_hot_i[111];
  assign data_masked[14275] = data_i[14275] & sel_one_hot_i[111];
  assign data_masked[14274] = data_i[14274] & sel_one_hot_i[111];
  assign data_masked[14273] = data_i[14273] & sel_one_hot_i[111];
  assign data_masked[14272] = data_i[14272] & sel_one_hot_i[111];
  assign data_masked[14271] = data_i[14271] & sel_one_hot_i[111];
  assign data_masked[14270] = data_i[14270] & sel_one_hot_i[111];
  assign data_masked[14269] = data_i[14269] & sel_one_hot_i[111];
  assign data_masked[14268] = data_i[14268] & sel_one_hot_i[111];
  assign data_masked[14267] = data_i[14267] & sel_one_hot_i[111];
  assign data_masked[14266] = data_i[14266] & sel_one_hot_i[111];
  assign data_masked[14265] = data_i[14265] & sel_one_hot_i[111];
  assign data_masked[14264] = data_i[14264] & sel_one_hot_i[111];
  assign data_masked[14263] = data_i[14263] & sel_one_hot_i[111];
  assign data_masked[14262] = data_i[14262] & sel_one_hot_i[111];
  assign data_masked[14261] = data_i[14261] & sel_one_hot_i[111];
  assign data_masked[14260] = data_i[14260] & sel_one_hot_i[111];
  assign data_masked[14259] = data_i[14259] & sel_one_hot_i[111];
  assign data_masked[14258] = data_i[14258] & sel_one_hot_i[111];
  assign data_masked[14257] = data_i[14257] & sel_one_hot_i[111];
  assign data_masked[14256] = data_i[14256] & sel_one_hot_i[111];
  assign data_masked[14255] = data_i[14255] & sel_one_hot_i[111];
  assign data_masked[14254] = data_i[14254] & sel_one_hot_i[111];
  assign data_masked[14253] = data_i[14253] & sel_one_hot_i[111];
  assign data_masked[14252] = data_i[14252] & sel_one_hot_i[111];
  assign data_masked[14251] = data_i[14251] & sel_one_hot_i[111];
  assign data_masked[14250] = data_i[14250] & sel_one_hot_i[111];
  assign data_masked[14249] = data_i[14249] & sel_one_hot_i[111];
  assign data_masked[14248] = data_i[14248] & sel_one_hot_i[111];
  assign data_masked[14247] = data_i[14247] & sel_one_hot_i[111];
  assign data_masked[14246] = data_i[14246] & sel_one_hot_i[111];
  assign data_masked[14245] = data_i[14245] & sel_one_hot_i[111];
  assign data_masked[14244] = data_i[14244] & sel_one_hot_i[111];
  assign data_masked[14243] = data_i[14243] & sel_one_hot_i[111];
  assign data_masked[14242] = data_i[14242] & sel_one_hot_i[111];
  assign data_masked[14241] = data_i[14241] & sel_one_hot_i[111];
  assign data_masked[14240] = data_i[14240] & sel_one_hot_i[111];
  assign data_masked[14239] = data_i[14239] & sel_one_hot_i[111];
  assign data_masked[14238] = data_i[14238] & sel_one_hot_i[111];
  assign data_masked[14237] = data_i[14237] & sel_one_hot_i[111];
  assign data_masked[14236] = data_i[14236] & sel_one_hot_i[111];
  assign data_masked[14235] = data_i[14235] & sel_one_hot_i[111];
  assign data_masked[14234] = data_i[14234] & sel_one_hot_i[111];
  assign data_masked[14233] = data_i[14233] & sel_one_hot_i[111];
  assign data_masked[14232] = data_i[14232] & sel_one_hot_i[111];
  assign data_masked[14231] = data_i[14231] & sel_one_hot_i[111];
  assign data_masked[14230] = data_i[14230] & sel_one_hot_i[111];
  assign data_masked[14229] = data_i[14229] & sel_one_hot_i[111];
  assign data_masked[14228] = data_i[14228] & sel_one_hot_i[111];
  assign data_masked[14227] = data_i[14227] & sel_one_hot_i[111];
  assign data_masked[14226] = data_i[14226] & sel_one_hot_i[111];
  assign data_masked[14225] = data_i[14225] & sel_one_hot_i[111];
  assign data_masked[14224] = data_i[14224] & sel_one_hot_i[111];
  assign data_masked[14223] = data_i[14223] & sel_one_hot_i[111];
  assign data_masked[14222] = data_i[14222] & sel_one_hot_i[111];
  assign data_masked[14221] = data_i[14221] & sel_one_hot_i[111];
  assign data_masked[14220] = data_i[14220] & sel_one_hot_i[111];
  assign data_masked[14219] = data_i[14219] & sel_one_hot_i[111];
  assign data_masked[14218] = data_i[14218] & sel_one_hot_i[111];
  assign data_masked[14217] = data_i[14217] & sel_one_hot_i[111];
  assign data_masked[14216] = data_i[14216] & sel_one_hot_i[111];
  assign data_masked[14215] = data_i[14215] & sel_one_hot_i[111];
  assign data_masked[14214] = data_i[14214] & sel_one_hot_i[111];
  assign data_masked[14213] = data_i[14213] & sel_one_hot_i[111];
  assign data_masked[14212] = data_i[14212] & sel_one_hot_i[111];
  assign data_masked[14211] = data_i[14211] & sel_one_hot_i[111];
  assign data_masked[14210] = data_i[14210] & sel_one_hot_i[111];
  assign data_masked[14209] = data_i[14209] & sel_one_hot_i[111];
  assign data_masked[14208] = data_i[14208] & sel_one_hot_i[111];
  assign data_masked[14463] = data_i[14463] & sel_one_hot_i[112];
  assign data_masked[14462] = data_i[14462] & sel_one_hot_i[112];
  assign data_masked[14461] = data_i[14461] & sel_one_hot_i[112];
  assign data_masked[14460] = data_i[14460] & sel_one_hot_i[112];
  assign data_masked[14459] = data_i[14459] & sel_one_hot_i[112];
  assign data_masked[14458] = data_i[14458] & sel_one_hot_i[112];
  assign data_masked[14457] = data_i[14457] & sel_one_hot_i[112];
  assign data_masked[14456] = data_i[14456] & sel_one_hot_i[112];
  assign data_masked[14455] = data_i[14455] & sel_one_hot_i[112];
  assign data_masked[14454] = data_i[14454] & sel_one_hot_i[112];
  assign data_masked[14453] = data_i[14453] & sel_one_hot_i[112];
  assign data_masked[14452] = data_i[14452] & sel_one_hot_i[112];
  assign data_masked[14451] = data_i[14451] & sel_one_hot_i[112];
  assign data_masked[14450] = data_i[14450] & sel_one_hot_i[112];
  assign data_masked[14449] = data_i[14449] & sel_one_hot_i[112];
  assign data_masked[14448] = data_i[14448] & sel_one_hot_i[112];
  assign data_masked[14447] = data_i[14447] & sel_one_hot_i[112];
  assign data_masked[14446] = data_i[14446] & sel_one_hot_i[112];
  assign data_masked[14445] = data_i[14445] & sel_one_hot_i[112];
  assign data_masked[14444] = data_i[14444] & sel_one_hot_i[112];
  assign data_masked[14443] = data_i[14443] & sel_one_hot_i[112];
  assign data_masked[14442] = data_i[14442] & sel_one_hot_i[112];
  assign data_masked[14441] = data_i[14441] & sel_one_hot_i[112];
  assign data_masked[14440] = data_i[14440] & sel_one_hot_i[112];
  assign data_masked[14439] = data_i[14439] & sel_one_hot_i[112];
  assign data_masked[14438] = data_i[14438] & sel_one_hot_i[112];
  assign data_masked[14437] = data_i[14437] & sel_one_hot_i[112];
  assign data_masked[14436] = data_i[14436] & sel_one_hot_i[112];
  assign data_masked[14435] = data_i[14435] & sel_one_hot_i[112];
  assign data_masked[14434] = data_i[14434] & sel_one_hot_i[112];
  assign data_masked[14433] = data_i[14433] & sel_one_hot_i[112];
  assign data_masked[14432] = data_i[14432] & sel_one_hot_i[112];
  assign data_masked[14431] = data_i[14431] & sel_one_hot_i[112];
  assign data_masked[14430] = data_i[14430] & sel_one_hot_i[112];
  assign data_masked[14429] = data_i[14429] & sel_one_hot_i[112];
  assign data_masked[14428] = data_i[14428] & sel_one_hot_i[112];
  assign data_masked[14427] = data_i[14427] & sel_one_hot_i[112];
  assign data_masked[14426] = data_i[14426] & sel_one_hot_i[112];
  assign data_masked[14425] = data_i[14425] & sel_one_hot_i[112];
  assign data_masked[14424] = data_i[14424] & sel_one_hot_i[112];
  assign data_masked[14423] = data_i[14423] & sel_one_hot_i[112];
  assign data_masked[14422] = data_i[14422] & sel_one_hot_i[112];
  assign data_masked[14421] = data_i[14421] & sel_one_hot_i[112];
  assign data_masked[14420] = data_i[14420] & sel_one_hot_i[112];
  assign data_masked[14419] = data_i[14419] & sel_one_hot_i[112];
  assign data_masked[14418] = data_i[14418] & sel_one_hot_i[112];
  assign data_masked[14417] = data_i[14417] & sel_one_hot_i[112];
  assign data_masked[14416] = data_i[14416] & sel_one_hot_i[112];
  assign data_masked[14415] = data_i[14415] & sel_one_hot_i[112];
  assign data_masked[14414] = data_i[14414] & sel_one_hot_i[112];
  assign data_masked[14413] = data_i[14413] & sel_one_hot_i[112];
  assign data_masked[14412] = data_i[14412] & sel_one_hot_i[112];
  assign data_masked[14411] = data_i[14411] & sel_one_hot_i[112];
  assign data_masked[14410] = data_i[14410] & sel_one_hot_i[112];
  assign data_masked[14409] = data_i[14409] & sel_one_hot_i[112];
  assign data_masked[14408] = data_i[14408] & sel_one_hot_i[112];
  assign data_masked[14407] = data_i[14407] & sel_one_hot_i[112];
  assign data_masked[14406] = data_i[14406] & sel_one_hot_i[112];
  assign data_masked[14405] = data_i[14405] & sel_one_hot_i[112];
  assign data_masked[14404] = data_i[14404] & sel_one_hot_i[112];
  assign data_masked[14403] = data_i[14403] & sel_one_hot_i[112];
  assign data_masked[14402] = data_i[14402] & sel_one_hot_i[112];
  assign data_masked[14401] = data_i[14401] & sel_one_hot_i[112];
  assign data_masked[14400] = data_i[14400] & sel_one_hot_i[112];
  assign data_masked[14399] = data_i[14399] & sel_one_hot_i[112];
  assign data_masked[14398] = data_i[14398] & sel_one_hot_i[112];
  assign data_masked[14397] = data_i[14397] & sel_one_hot_i[112];
  assign data_masked[14396] = data_i[14396] & sel_one_hot_i[112];
  assign data_masked[14395] = data_i[14395] & sel_one_hot_i[112];
  assign data_masked[14394] = data_i[14394] & sel_one_hot_i[112];
  assign data_masked[14393] = data_i[14393] & sel_one_hot_i[112];
  assign data_masked[14392] = data_i[14392] & sel_one_hot_i[112];
  assign data_masked[14391] = data_i[14391] & sel_one_hot_i[112];
  assign data_masked[14390] = data_i[14390] & sel_one_hot_i[112];
  assign data_masked[14389] = data_i[14389] & sel_one_hot_i[112];
  assign data_masked[14388] = data_i[14388] & sel_one_hot_i[112];
  assign data_masked[14387] = data_i[14387] & sel_one_hot_i[112];
  assign data_masked[14386] = data_i[14386] & sel_one_hot_i[112];
  assign data_masked[14385] = data_i[14385] & sel_one_hot_i[112];
  assign data_masked[14384] = data_i[14384] & sel_one_hot_i[112];
  assign data_masked[14383] = data_i[14383] & sel_one_hot_i[112];
  assign data_masked[14382] = data_i[14382] & sel_one_hot_i[112];
  assign data_masked[14381] = data_i[14381] & sel_one_hot_i[112];
  assign data_masked[14380] = data_i[14380] & sel_one_hot_i[112];
  assign data_masked[14379] = data_i[14379] & sel_one_hot_i[112];
  assign data_masked[14378] = data_i[14378] & sel_one_hot_i[112];
  assign data_masked[14377] = data_i[14377] & sel_one_hot_i[112];
  assign data_masked[14376] = data_i[14376] & sel_one_hot_i[112];
  assign data_masked[14375] = data_i[14375] & sel_one_hot_i[112];
  assign data_masked[14374] = data_i[14374] & sel_one_hot_i[112];
  assign data_masked[14373] = data_i[14373] & sel_one_hot_i[112];
  assign data_masked[14372] = data_i[14372] & sel_one_hot_i[112];
  assign data_masked[14371] = data_i[14371] & sel_one_hot_i[112];
  assign data_masked[14370] = data_i[14370] & sel_one_hot_i[112];
  assign data_masked[14369] = data_i[14369] & sel_one_hot_i[112];
  assign data_masked[14368] = data_i[14368] & sel_one_hot_i[112];
  assign data_masked[14367] = data_i[14367] & sel_one_hot_i[112];
  assign data_masked[14366] = data_i[14366] & sel_one_hot_i[112];
  assign data_masked[14365] = data_i[14365] & sel_one_hot_i[112];
  assign data_masked[14364] = data_i[14364] & sel_one_hot_i[112];
  assign data_masked[14363] = data_i[14363] & sel_one_hot_i[112];
  assign data_masked[14362] = data_i[14362] & sel_one_hot_i[112];
  assign data_masked[14361] = data_i[14361] & sel_one_hot_i[112];
  assign data_masked[14360] = data_i[14360] & sel_one_hot_i[112];
  assign data_masked[14359] = data_i[14359] & sel_one_hot_i[112];
  assign data_masked[14358] = data_i[14358] & sel_one_hot_i[112];
  assign data_masked[14357] = data_i[14357] & sel_one_hot_i[112];
  assign data_masked[14356] = data_i[14356] & sel_one_hot_i[112];
  assign data_masked[14355] = data_i[14355] & sel_one_hot_i[112];
  assign data_masked[14354] = data_i[14354] & sel_one_hot_i[112];
  assign data_masked[14353] = data_i[14353] & sel_one_hot_i[112];
  assign data_masked[14352] = data_i[14352] & sel_one_hot_i[112];
  assign data_masked[14351] = data_i[14351] & sel_one_hot_i[112];
  assign data_masked[14350] = data_i[14350] & sel_one_hot_i[112];
  assign data_masked[14349] = data_i[14349] & sel_one_hot_i[112];
  assign data_masked[14348] = data_i[14348] & sel_one_hot_i[112];
  assign data_masked[14347] = data_i[14347] & sel_one_hot_i[112];
  assign data_masked[14346] = data_i[14346] & sel_one_hot_i[112];
  assign data_masked[14345] = data_i[14345] & sel_one_hot_i[112];
  assign data_masked[14344] = data_i[14344] & sel_one_hot_i[112];
  assign data_masked[14343] = data_i[14343] & sel_one_hot_i[112];
  assign data_masked[14342] = data_i[14342] & sel_one_hot_i[112];
  assign data_masked[14341] = data_i[14341] & sel_one_hot_i[112];
  assign data_masked[14340] = data_i[14340] & sel_one_hot_i[112];
  assign data_masked[14339] = data_i[14339] & sel_one_hot_i[112];
  assign data_masked[14338] = data_i[14338] & sel_one_hot_i[112];
  assign data_masked[14337] = data_i[14337] & sel_one_hot_i[112];
  assign data_masked[14336] = data_i[14336] & sel_one_hot_i[112];
  assign data_masked[14591] = data_i[14591] & sel_one_hot_i[113];
  assign data_masked[14590] = data_i[14590] & sel_one_hot_i[113];
  assign data_masked[14589] = data_i[14589] & sel_one_hot_i[113];
  assign data_masked[14588] = data_i[14588] & sel_one_hot_i[113];
  assign data_masked[14587] = data_i[14587] & sel_one_hot_i[113];
  assign data_masked[14586] = data_i[14586] & sel_one_hot_i[113];
  assign data_masked[14585] = data_i[14585] & sel_one_hot_i[113];
  assign data_masked[14584] = data_i[14584] & sel_one_hot_i[113];
  assign data_masked[14583] = data_i[14583] & sel_one_hot_i[113];
  assign data_masked[14582] = data_i[14582] & sel_one_hot_i[113];
  assign data_masked[14581] = data_i[14581] & sel_one_hot_i[113];
  assign data_masked[14580] = data_i[14580] & sel_one_hot_i[113];
  assign data_masked[14579] = data_i[14579] & sel_one_hot_i[113];
  assign data_masked[14578] = data_i[14578] & sel_one_hot_i[113];
  assign data_masked[14577] = data_i[14577] & sel_one_hot_i[113];
  assign data_masked[14576] = data_i[14576] & sel_one_hot_i[113];
  assign data_masked[14575] = data_i[14575] & sel_one_hot_i[113];
  assign data_masked[14574] = data_i[14574] & sel_one_hot_i[113];
  assign data_masked[14573] = data_i[14573] & sel_one_hot_i[113];
  assign data_masked[14572] = data_i[14572] & sel_one_hot_i[113];
  assign data_masked[14571] = data_i[14571] & sel_one_hot_i[113];
  assign data_masked[14570] = data_i[14570] & sel_one_hot_i[113];
  assign data_masked[14569] = data_i[14569] & sel_one_hot_i[113];
  assign data_masked[14568] = data_i[14568] & sel_one_hot_i[113];
  assign data_masked[14567] = data_i[14567] & sel_one_hot_i[113];
  assign data_masked[14566] = data_i[14566] & sel_one_hot_i[113];
  assign data_masked[14565] = data_i[14565] & sel_one_hot_i[113];
  assign data_masked[14564] = data_i[14564] & sel_one_hot_i[113];
  assign data_masked[14563] = data_i[14563] & sel_one_hot_i[113];
  assign data_masked[14562] = data_i[14562] & sel_one_hot_i[113];
  assign data_masked[14561] = data_i[14561] & sel_one_hot_i[113];
  assign data_masked[14560] = data_i[14560] & sel_one_hot_i[113];
  assign data_masked[14559] = data_i[14559] & sel_one_hot_i[113];
  assign data_masked[14558] = data_i[14558] & sel_one_hot_i[113];
  assign data_masked[14557] = data_i[14557] & sel_one_hot_i[113];
  assign data_masked[14556] = data_i[14556] & sel_one_hot_i[113];
  assign data_masked[14555] = data_i[14555] & sel_one_hot_i[113];
  assign data_masked[14554] = data_i[14554] & sel_one_hot_i[113];
  assign data_masked[14553] = data_i[14553] & sel_one_hot_i[113];
  assign data_masked[14552] = data_i[14552] & sel_one_hot_i[113];
  assign data_masked[14551] = data_i[14551] & sel_one_hot_i[113];
  assign data_masked[14550] = data_i[14550] & sel_one_hot_i[113];
  assign data_masked[14549] = data_i[14549] & sel_one_hot_i[113];
  assign data_masked[14548] = data_i[14548] & sel_one_hot_i[113];
  assign data_masked[14547] = data_i[14547] & sel_one_hot_i[113];
  assign data_masked[14546] = data_i[14546] & sel_one_hot_i[113];
  assign data_masked[14545] = data_i[14545] & sel_one_hot_i[113];
  assign data_masked[14544] = data_i[14544] & sel_one_hot_i[113];
  assign data_masked[14543] = data_i[14543] & sel_one_hot_i[113];
  assign data_masked[14542] = data_i[14542] & sel_one_hot_i[113];
  assign data_masked[14541] = data_i[14541] & sel_one_hot_i[113];
  assign data_masked[14540] = data_i[14540] & sel_one_hot_i[113];
  assign data_masked[14539] = data_i[14539] & sel_one_hot_i[113];
  assign data_masked[14538] = data_i[14538] & sel_one_hot_i[113];
  assign data_masked[14537] = data_i[14537] & sel_one_hot_i[113];
  assign data_masked[14536] = data_i[14536] & sel_one_hot_i[113];
  assign data_masked[14535] = data_i[14535] & sel_one_hot_i[113];
  assign data_masked[14534] = data_i[14534] & sel_one_hot_i[113];
  assign data_masked[14533] = data_i[14533] & sel_one_hot_i[113];
  assign data_masked[14532] = data_i[14532] & sel_one_hot_i[113];
  assign data_masked[14531] = data_i[14531] & sel_one_hot_i[113];
  assign data_masked[14530] = data_i[14530] & sel_one_hot_i[113];
  assign data_masked[14529] = data_i[14529] & sel_one_hot_i[113];
  assign data_masked[14528] = data_i[14528] & sel_one_hot_i[113];
  assign data_masked[14527] = data_i[14527] & sel_one_hot_i[113];
  assign data_masked[14526] = data_i[14526] & sel_one_hot_i[113];
  assign data_masked[14525] = data_i[14525] & sel_one_hot_i[113];
  assign data_masked[14524] = data_i[14524] & sel_one_hot_i[113];
  assign data_masked[14523] = data_i[14523] & sel_one_hot_i[113];
  assign data_masked[14522] = data_i[14522] & sel_one_hot_i[113];
  assign data_masked[14521] = data_i[14521] & sel_one_hot_i[113];
  assign data_masked[14520] = data_i[14520] & sel_one_hot_i[113];
  assign data_masked[14519] = data_i[14519] & sel_one_hot_i[113];
  assign data_masked[14518] = data_i[14518] & sel_one_hot_i[113];
  assign data_masked[14517] = data_i[14517] & sel_one_hot_i[113];
  assign data_masked[14516] = data_i[14516] & sel_one_hot_i[113];
  assign data_masked[14515] = data_i[14515] & sel_one_hot_i[113];
  assign data_masked[14514] = data_i[14514] & sel_one_hot_i[113];
  assign data_masked[14513] = data_i[14513] & sel_one_hot_i[113];
  assign data_masked[14512] = data_i[14512] & sel_one_hot_i[113];
  assign data_masked[14511] = data_i[14511] & sel_one_hot_i[113];
  assign data_masked[14510] = data_i[14510] & sel_one_hot_i[113];
  assign data_masked[14509] = data_i[14509] & sel_one_hot_i[113];
  assign data_masked[14508] = data_i[14508] & sel_one_hot_i[113];
  assign data_masked[14507] = data_i[14507] & sel_one_hot_i[113];
  assign data_masked[14506] = data_i[14506] & sel_one_hot_i[113];
  assign data_masked[14505] = data_i[14505] & sel_one_hot_i[113];
  assign data_masked[14504] = data_i[14504] & sel_one_hot_i[113];
  assign data_masked[14503] = data_i[14503] & sel_one_hot_i[113];
  assign data_masked[14502] = data_i[14502] & sel_one_hot_i[113];
  assign data_masked[14501] = data_i[14501] & sel_one_hot_i[113];
  assign data_masked[14500] = data_i[14500] & sel_one_hot_i[113];
  assign data_masked[14499] = data_i[14499] & sel_one_hot_i[113];
  assign data_masked[14498] = data_i[14498] & sel_one_hot_i[113];
  assign data_masked[14497] = data_i[14497] & sel_one_hot_i[113];
  assign data_masked[14496] = data_i[14496] & sel_one_hot_i[113];
  assign data_masked[14495] = data_i[14495] & sel_one_hot_i[113];
  assign data_masked[14494] = data_i[14494] & sel_one_hot_i[113];
  assign data_masked[14493] = data_i[14493] & sel_one_hot_i[113];
  assign data_masked[14492] = data_i[14492] & sel_one_hot_i[113];
  assign data_masked[14491] = data_i[14491] & sel_one_hot_i[113];
  assign data_masked[14490] = data_i[14490] & sel_one_hot_i[113];
  assign data_masked[14489] = data_i[14489] & sel_one_hot_i[113];
  assign data_masked[14488] = data_i[14488] & sel_one_hot_i[113];
  assign data_masked[14487] = data_i[14487] & sel_one_hot_i[113];
  assign data_masked[14486] = data_i[14486] & sel_one_hot_i[113];
  assign data_masked[14485] = data_i[14485] & sel_one_hot_i[113];
  assign data_masked[14484] = data_i[14484] & sel_one_hot_i[113];
  assign data_masked[14483] = data_i[14483] & sel_one_hot_i[113];
  assign data_masked[14482] = data_i[14482] & sel_one_hot_i[113];
  assign data_masked[14481] = data_i[14481] & sel_one_hot_i[113];
  assign data_masked[14480] = data_i[14480] & sel_one_hot_i[113];
  assign data_masked[14479] = data_i[14479] & sel_one_hot_i[113];
  assign data_masked[14478] = data_i[14478] & sel_one_hot_i[113];
  assign data_masked[14477] = data_i[14477] & sel_one_hot_i[113];
  assign data_masked[14476] = data_i[14476] & sel_one_hot_i[113];
  assign data_masked[14475] = data_i[14475] & sel_one_hot_i[113];
  assign data_masked[14474] = data_i[14474] & sel_one_hot_i[113];
  assign data_masked[14473] = data_i[14473] & sel_one_hot_i[113];
  assign data_masked[14472] = data_i[14472] & sel_one_hot_i[113];
  assign data_masked[14471] = data_i[14471] & sel_one_hot_i[113];
  assign data_masked[14470] = data_i[14470] & sel_one_hot_i[113];
  assign data_masked[14469] = data_i[14469] & sel_one_hot_i[113];
  assign data_masked[14468] = data_i[14468] & sel_one_hot_i[113];
  assign data_masked[14467] = data_i[14467] & sel_one_hot_i[113];
  assign data_masked[14466] = data_i[14466] & sel_one_hot_i[113];
  assign data_masked[14465] = data_i[14465] & sel_one_hot_i[113];
  assign data_masked[14464] = data_i[14464] & sel_one_hot_i[113];
  assign data_masked[14719] = data_i[14719] & sel_one_hot_i[114];
  assign data_masked[14718] = data_i[14718] & sel_one_hot_i[114];
  assign data_masked[14717] = data_i[14717] & sel_one_hot_i[114];
  assign data_masked[14716] = data_i[14716] & sel_one_hot_i[114];
  assign data_masked[14715] = data_i[14715] & sel_one_hot_i[114];
  assign data_masked[14714] = data_i[14714] & sel_one_hot_i[114];
  assign data_masked[14713] = data_i[14713] & sel_one_hot_i[114];
  assign data_masked[14712] = data_i[14712] & sel_one_hot_i[114];
  assign data_masked[14711] = data_i[14711] & sel_one_hot_i[114];
  assign data_masked[14710] = data_i[14710] & sel_one_hot_i[114];
  assign data_masked[14709] = data_i[14709] & sel_one_hot_i[114];
  assign data_masked[14708] = data_i[14708] & sel_one_hot_i[114];
  assign data_masked[14707] = data_i[14707] & sel_one_hot_i[114];
  assign data_masked[14706] = data_i[14706] & sel_one_hot_i[114];
  assign data_masked[14705] = data_i[14705] & sel_one_hot_i[114];
  assign data_masked[14704] = data_i[14704] & sel_one_hot_i[114];
  assign data_masked[14703] = data_i[14703] & sel_one_hot_i[114];
  assign data_masked[14702] = data_i[14702] & sel_one_hot_i[114];
  assign data_masked[14701] = data_i[14701] & sel_one_hot_i[114];
  assign data_masked[14700] = data_i[14700] & sel_one_hot_i[114];
  assign data_masked[14699] = data_i[14699] & sel_one_hot_i[114];
  assign data_masked[14698] = data_i[14698] & sel_one_hot_i[114];
  assign data_masked[14697] = data_i[14697] & sel_one_hot_i[114];
  assign data_masked[14696] = data_i[14696] & sel_one_hot_i[114];
  assign data_masked[14695] = data_i[14695] & sel_one_hot_i[114];
  assign data_masked[14694] = data_i[14694] & sel_one_hot_i[114];
  assign data_masked[14693] = data_i[14693] & sel_one_hot_i[114];
  assign data_masked[14692] = data_i[14692] & sel_one_hot_i[114];
  assign data_masked[14691] = data_i[14691] & sel_one_hot_i[114];
  assign data_masked[14690] = data_i[14690] & sel_one_hot_i[114];
  assign data_masked[14689] = data_i[14689] & sel_one_hot_i[114];
  assign data_masked[14688] = data_i[14688] & sel_one_hot_i[114];
  assign data_masked[14687] = data_i[14687] & sel_one_hot_i[114];
  assign data_masked[14686] = data_i[14686] & sel_one_hot_i[114];
  assign data_masked[14685] = data_i[14685] & sel_one_hot_i[114];
  assign data_masked[14684] = data_i[14684] & sel_one_hot_i[114];
  assign data_masked[14683] = data_i[14683] & sel_one_hot_i[114];
  assign data_masked[14682] = data_i[14682] & sel_one_hot_i[114];
  assign data_masked[14681] = data_i[14681] & sel_one_hot_i[114];
  assign data_masked[14680] = data_i[14680] & sel_one_hot_i[114];
  assign data_masked[14679] = data_i[14679] & sel_one_hot_i[114];
  assign data_masked[14678] = data_i[14678] & sel_one_hot_i[114];
  assign data_masked[14677] = data_i[14677] & sel_one_hot_i[114];
  assign data_masked[14676] = data_i[14676] & sel_one_hot_i[114];
  assign data_masked[14675] = data_i[14675] & sel_one_hot_i[114];
  assign data_masked[14674] = data_i[14674] & sel_one_hot_i[114];
  assign data_masked[14673] = data_i[14673] & sel_one_hot_i[114];
  assign data_masked[14672] = data_i[14672] & sel_one_hot_i[114];
  assign data_masked[14671] = data_i[14671] & sel_one_hot_i[114];
  assign data_masked[14670] = data_i[14670] & sel_one_hot_i[114];
  assign data_masked[14669] = data_i[14669] & sel_one_hot_i[114];
  assign data_masked[14668] = data_i[14668] & sel_one_hot_i[114];
  assign data_masked[14667] = data_i[14667] & sel_one_hot_i[114];
  assign data_masked[14666] = data_i[14666] & sel_one_hot_i[114];
  assign data_masked[14665] = data_i[14665] & sel_one_hot_i[114];
  assign data_masked[14664] = data_i[14664] & sel_one_hot_i[114];
  assign data_masked[14663] = data_i[14663] & sel_one_hot_i[114];
  assign data_masked[14662] = data_i[14662] & sel_one_hot_i[114];
  assign data_masked[14661] = data_i[14661] & sel_one_hot_i[114];
  assign data_masked[14660] = data_i[14660] & sel_one_hot_i[114];
  assign data_masked[14659] = data_i[14659] & sel_one_hot_i[114];
  assign data_masked[14658] = data_i[14658] & sel_one_hot_i[114];
  assign data_masked[14657] = data_i[14657] & sel_one_hot_i[114];
  assign data_masked[14656] = data_i[14656] & sel_one_hot_i[114];
  assign data_masked[14655] = data_i[14655] & sel_one_hot_i[114];
  assign data_masked[14654] = data_i[14654] & sel_one_hot_i[114];
  assign data_masked[14653] = data_i[14653] & sel_one_hot_i[114];
  assign data_masked[14652] = data_i[14652] & sel_one_hot_i[114];
  assign data_masked[14651] = data_i[14651] & sel_one_hot_i[114];
  assign data_masked[14650] = data_i[14650] & sel_one_hot_i[114];
  assign data_masked[14649] = data_i[14649] & sel_one_hot_i[114];
  assign data_masked[14648] = data_i[14648] & sel_one_hot_i[114];
  assign data_masked[14647] = data_i[14647] & sel_one_hot_i[114];
  assign data_masked[14646] = data_i[14646] & sel_one_hot_i[114];
  assign data_masked[14645] = data_i[14645] & sel_one_hot_i[114];
  assign data_masked[14644] = data_i[14644] & sel_one_hot_i[114];
  assign data_masked[14643] = data_i[14643] & sel_one_hot_i[114];
  assign data_masked[14642] = data_i[14642] & sel_one_hot_i[114];
  assign data_masked[14641] = data_i[14641] & sel_one_hot_i[114];
  assign data_masked[14640] = data_i[14640] & sel_one_hot_i[114];
  assign data_masked[14639] = data_i[14639] & sel_one_hot_i[114];
  assign data_masked[14638] = data_i[14638] & sel_one_hot_i[114];
  assign data_masked[14637] = data_i[14637] & sel_one_hot_i[114];
  assign data_masked[14636] = data_i[14636] & sel_one_hot_i[114];
  assign data_masked[14635] = data_i[14635] & sel_one_hot_i[114];
  assign data_masked[14634] = data_i[14634] & sel_one_hot_i[114];
  assign data_masked[14633] = data_i[14633] & sel_one_hot_i[114];
  assign data_masked[14632] = data_i[14632] & sel_one_hot_i[114];
  assign data_masked[14631] = data_i[14631] & sel_one_hot_i[114];
  assign data_masked[14630] = data_i[14630] & sel_one_hot_i[114];
  assign data_masked[14629] = data_i[14629] & sel_one_hot_i[114];
  assign data_masked[14628] = data_i[14628] & sel_one_hot_i[114];
  assign data_masked[14627] = data_i[14627] & sel_one_hot_i[114];
  assign data_masked[14626] = data_i[14626] & sel_one_hot_i[114];
  assign data_masked[14625] = data_i[14625] & sel_one_hot_i[114];
  assign data_masked[14624] = data_i[14624] & sel_one_hot_i[114];
  assign data_masked[14623] = data_i[14623] & sel_one_hot_i[114];
  assign data_masked[14622] = data_i[14622] & sel_one_hot_i[114];
  assign data_masked[14621] = data_i[14621] & sel_one_hot_i[114];
  assign data_masked[14620] = data_i[14620] & sel_one_hot_i[114];
  assign data_masked[14619] = data_i[14619] & sel_one_hot_i[114];
  assign data_masked[14618] = data_i[14618] & sel_one_hot_i[114];
  assign data_masked[14617] = data_i[14617] & sel_one_hot_i[114];
  assign data_masked[14616] = data_i[14616] & sel_one_hot_i[114];
  assign data_masked[14615] = data_i[14615] & sel_one_hot_i[114];
  assign data_masked[14614] = data_i[14614] & sel_one_hot_i[114];
  assign data_masked[14613] = data_i[14613] & sel_one_hot_i[114];
  assign data_masked[14612] = data_i[14612] & sel_one_hot_i[114];
  assign data_masked[14611] = data_i[14611] & sel_one_hot_i[114];
  assign data_masked[14610] = data_i[14610] & sel_one_hot_i[114];
  assign data_masked[14609] = data_i[14609] & sel_one_hot_i[114];
  assign data_masked[14608] = data_i[14608] & sel_one_hot_i[114];
  assign data_masked[14607] = data_i[14607] & sel_one_hot_i[114];
  assign data_masked[14606] = data_i[14606] & sel_one_hot_i[114];
  assign data_masked[14605] = data_i[14605] & sel_one_hot_i[114];
  assign data_masked[14604] = data_i[14604] & sel_one_hot_i[114];
  assign data_masked[14603] = data_i[14603] & sel_one_hot_i[114];
  assign data_masked[14602] = data_i[14602] & sel_one_hot_i[114];
  assign data_masked[14601] = data_i[14601] & sel_one_hot_i[114];
  assign data_masked[14600] = data_i[14600] & sel_one_hot_i[114];
  assign data_masked[14599] = data_i[14599] & sel_one_hot_i[114];
  assign data_masked[14598] = data_i[14598] & sel_one_hot_i[114];
  assign data_masked[14597] = data_i[14597] & sel_one_hot_i[114];
  assign data_masked[14596] = data_i[14596] & sel_one_hot_i[114];
  assign data_masked[14595] = data_i[14595] & sel_one_hot_i[114];
  assign data_masked[14594] = data_i[14594] & sel_one_hot_i[114];
  assign data_masked[14593] = data_i[14593] & sel_one_hot_i[114];
  assign data_masked[14592] = data_i[14592] & sel_one_hot_i[114];
  assign data_masked[14847] = data_i[14847] & sel_one_hot_i[115];
  assign data_masked[14846] = data_i[14846] & sel_one_hot_i[115];
  assign data_masked[14845] = data_i[14845] & sel_one_hot_i[115];
  assign data_masked[14844] = data_i[14844] & sel_one_hot_i[115];
  assign data_masked[14843] = data_i[14843] & sel_one_hot_i[115];
  assign data_masked[14842] = data_i[14842] & sel_one_hot_i[115];
  assign data_masked[14841] = data_i[14841] & sel_one_hot_i[115];
  assign data_masked[14840] = data_i[14840] & sel_one_hot_i[115];
  assign data_masked[14839] = data_i[14839] & sel_one_hot_i[115];
  assign data_masked[14838] = data_i[14838] & sel_one_hot_i[115];
  assign data_masked[14837] = data_i[14837] & sel_one_hot_i[115];
  assign data_masked[14836] = data_i[14836] & sel_one_hot_i[115];
  assign data_masked[14835] = data_i[14835] & sel_one_hot_i[115];
  assign data_masked[14834] = data_i[14834] & sel_one_hot_i[115];
  assign data_masked[14833] = data_i[14833] & sel_one_hot_i[115];
  assign data_masked[14832] = data_i[14832] & sel_one_hot_i[115];
  assign data_masked[14831] = data_i[14831] & sel_one_hot_i[115];
  assign data_masked[14830] = data_i[14830] & sel_one_hot_i[115];
  assign data_masked[14829] = data_i[14829] & sel_one_hot_i[115];
  assign data_masked[14828] = data_i[14828] & sel_one_hot_i[115];
  assign data_masked[14827] = data_i[14827] & sel_one_hot_i[115];
  assign data_masked[14826] = data_i[14826] & sel_one_hot_i[115];
  assign data_masked[14825] = data_i[14825] & sel_one_hot_i[115];
  assign data_masked[14824] = data_i[14824] & sel_one_hot_i[115];
  assign data_masked[14823] = data_i[14823] & sel_one_hot_i[115];
  assign data_masked[14822] = data_i[14822] & sel_one_hot_i[115];
  assign data_masked[14821] = data_i[14821] & sel_one_hot_i[115];
  assign data_masked[14820] = data_i[14820] & sel_one_hot_i[115];
  assign data_masked[14819] = data_i[14819] & sel_one_hot_i[115];
  assign data_masked[14818] = data_i[14818] & sel_one_hot_i[115];
  assign data_masked[14817] = data_i[14817] & sel_one_hot_i[115];
  assign data_masked[14816] = data_i[14816] & sel_one_hot_i[115];
  assign data_masked[14815] = data_i[14815] & sel_one_hot_i[115];
  assign data_masked[14814] = data_i[14814] & sel_one_hot_i[115];
  assign data_masked[14813] = data_i[14813] & sel_one_hot_i[115];
  assign data_masked[14812] = data_i[14812] & sel_one_hot_i[115];
  assign data_masked[14811] = data_i[14811] & sel_one_hot_i[115];
  assign data_masked[14810] = data_i[14810] & sel_one_hot_i[115];
  assign data_masked[14809] = data_i[14809] & sel_one_hot_i[115];
  assign data_masked[14808] = data_i[14808] & sel_one_hot_i[115];
  assign data_masked[14807] = data_i[14807] & sel_one_hot_i[115];
  assign data_masked[14806] = data_i[14806] & sel_one_hot_i[115];
  assign data_masked[14805] = data_i[14805] & sel_one_hot_i[115];
  assign data_masked[14804] = data_i[14804] & sel_one_hot_i[115];
  assign data_masked[14803] = data_i[14803] & sel_one_hot_i[115];
  assign data_masked[14802] = data_i[14802] & sel_one_hot_i[115];
  assign data_masked[14801] = data_i[14801] & sel_one_hot_i[115];
  assign data_masked[14800] = data_i[14800] & sel_one_hot_i[115];
  assign data_masked[14799] = data_i[14799] & sel_one_hot_i[115];
  assign data_masked[14798] = data_i[14798] & sel_one_hot_i[115];
  assign data_masked[14797] = data_i[14797] & sel_one_hot_i[115];
  assign data_masked[14796] = data_i[14796] & sel_one_hot_i[115];
  assign data_masked[14795] = data_i[14795] & sel_one_hot_i[115];
  assign data_masked[14794] = data_i[14794] & sel_one_hot_i[115];
  assign data_masked[14793] = data_i[14793] & sel_one_hot_i[115];
  assign data_masked[14792] = data_i[14792] & sel_one_hot_i[115];
  assign data_masked[14791] = data_i[14791] & sel_one_hot_i[115];
  assign data_masked[14790] = data_i[14790] & sel_one_hot_i[115];
  assign data_masked[14789] = data_i[14789] & sel_one_hot_i[115];
  assign data_masked[14788] = data_i[14788] & sel_one_hot_i[115];
  assign data_masked[14787] = data_i[14787] & sel_one_hot_i[115];
  assign data_masked[14786] = data_i[14786] & sel_one_hot_i[115];
  assign data_masked[14785] = data_i[14785] & sel_one_hot_i[115];
  assign data_masked[14784] = data_i[14784] & sel_one_hot_i[115];
  assign data_masked[14783] = data_i[14783] & sel_one_hot_i[115];
  assign data_masked[14782] = data_i[14782] & sel_one_hot_i[115];
  assign data_masked[14781] = data_i[14781] & sel_one_hot_i[115];
  assign data_masked[14780] = data_i[14780] & sel_one_hot_i[115];
  assign data_masked[14779] = data_i[14779] & sel_one_hot_i[115];
  assign data_masked[14778] = data_i[14778] & sel_one_hot_i[115];
  assign data_masked[14777] = data_i[14777] & sel_one_hot_i[115];
  assign data_masked[14776] = data_i[14776] & sel_one_hot_i[115];
  assign data_masked[14775] = data_i[14775] & sel_one_hot_i[115];
  assign data_masked[14774] = data_i[14774] & sel_one_hot_i[115];
  assign data_masked[14773] = data_i[14773] & sel_one_hot_i[115];
  assign data_masked[14772] = data_i[14772] & sel_one_hot_i[115];
  assign data_masked[14771] = data_i[14771] & sel_one_hot_i[115];
  assign data_masked[14770] = data_i[14770] & sel_one_hot_i[115];
  assign data_masked[14769] = data_i[14769] & sel_one_hot_i[115];
  assign data_masked[14768] = data_i[14768] & sel_one_hot_i[115];
  assign data_masked[14767] = data_i[14767] & sel_one_hot_i[115];
  assign data_masked[14766] = data_i[14766] & sel_one_hot_i[115];
  assign data_masked[14765] = data_i[14765] & sel_one_hot_i[115];
  assign data_masked[14764] = data_i[14764] & sel_one_hot_i[115];
  assign data_masked[14763] = data_i[14763] & sel_one_hot_i[115];
  assign data_masked[14762] = data_i[14762] & sel_one_hot_i[115];
  assign data_masked[14761] = data_i[14761] & sel_one_hot_i[115];
  assign data_masked[14760] = data_i[14760] & sel_one_hot_i[115];
  assign data_masked[14759] = data_i[14759] & sel_one_hot_i[115];
  assign data_masked[14758] = data_i[14758] & sel_one_hot_i[115];
  assign data_masked[14757] = data_i[14757] & sel_one_hot_i[115];
  assign data_masked[14756] = data_i[14756] & sel_one_hot_i[115];
  assign data_masked[14755] = data_i[14755] & sel_one_hot_i[115];
  assign data_masked[14754] = data_i[14754] & sel_one_hot_i[115];
  assign data_masked[14753] = data_i[14753] & sel_one_hot_i[115];
  assign data_masked[14752] = data_i[14752] & sel_one_hot_i[115];
  assign data_masked[14751] = data_i[14751] & sel_one_hot_i[115];
  assign data_masked[14750] = data_i[14750] & sel_one_hot_i[115];
  assign data_masked[14749] = data_i[14749] & sel_one_hot_i[115];
  assign data_masked[14748] = data_i[14748] & sel_one_hot_i[115];
  assign data_masked[14747] = data_i[14747] & sel_one_hot_i[115];
  assign data_masked[14746] = data_i[14746] & sel_one_hot_i[115];
  assign data_masked[14745] = data_i[14745] & sel_one_hot_i[115];
  assign data_masked[14744] = data_i[14744] & sel_one_hot_i[115];
  assign data_masked[14743] = data_i[14743] & sel_one_hot_i[115];
  assign data_masked[14742] = data_i[14742] & sel_one_hot_i[115];
  assign data_masked[14741] = data_i[14741] & sel_one_hot_i[115];
  assign data_masked[14740] = data_i[14740] & sel_one_hot_i[115];
  assign data_masked[14739] = data_i[14739] & sel_one_hot_i[115];
  assign data_masked[14738] = data_i[14738] & sel_one_hot_i[115];
  assign data_masked[14737] = data_i[14737] & sel_one_hot_i[115];
  assign data_masked[14736] = data_i[14736] & sel_one_hot_i[115];
  assign data_masked[14735] = data_i[14735] & sel_one_hot_i[115];
  assign data_masked[14734] = data_i[14734] & sel_one_hot_i[115];
  assign data_masked[14733] = data_i[14733] & sel_one_hot_i[115];
  assign data_masked[14732] = data_i[14732] & sel_one_hot_i[115];
  assign data_masked[14731] = data_i[14731] & sel_one_hot_i[115];
  assign data_masked[14730] = data_i[14730] & sel_one_hot_i[115];
  assign data_masked[14729] = data_i[14729] & sel_one_hot_i[115];
  assign data_masked[14728] = data_i[14728] & sel_one_hot_i[115];
  assign data_masked[14727] = data_i[14727] & sel_one_hot_i[115];
  assign data_masked[14726] = data_i[14726] & sel_one_hot_i[115];
  assign data_masked[14725] = data_i[14725] & sel_one_hot_i[115];
  assign data_masked[14724] = data_i[14724] & sel_one_hot_i[115];
  assign data_masked[14723] = data_i[14723] & sel_one_hot_i[115];
  assign data_masked[14722] = data_i[14722] & sel_one_hot_i[115];
  assign data_masked[14721] = data_i[14721] & sel_one_hot_i[115];
  assign data_masked[14720] = data_i[14720] & sel_one_hot_i[115];
  assign data_masked[14975] = data_i[14975] & sel_one_hot_i[116];
  assign data_masked[14974] = data_i[14974] & sel_one_hot_i[116];
  assign data_masked[14973] = data_i[14973] & sel_one_hot_i[116];
  assign data_masked[14972] = data_i[14972] & sel_one_hot_i[116];
  assign data_masked[14971] = data_i[14971] & sel_one_hot_i[116];
  assign data_masked[14970] = data_i[14970] & sel_one_hot_i[116];
  assign data_masked[14969] = data_i[14969] & sel_one_hot_i[116];
  assign data_masked[14968] = data_i[14968] & sel_one_hot_i[116];
  assign data_masked[14967] = data_i[14967] & sel_one_hot_i[116];
  assign data_masked[14966] = data_i[14966] & sel_one_hot_i[116];
  assign data_masked[14965] = data_i[14965] & sel_one_hot_i[116];
  assign data_masked[14964] = data_i[14964] & sel_one_hot_i[116];
  assign data_masked[14963] = data_i[14963] & sel_one_hot_i[116];
  assign data_masked[14962] = data_i[14962] & sel_one_hot_i[116];
  assign data_masked[14961] = data_i[14961] & sel_one_hot_i[116];
  assign data_masked[14960] = data_i[14960] & sel_one_hot_i[116];
  assign data_masked[14959] = data_i[14959] & sel_one_hot_i[116];
  assign data_masked[14958] = data_i[14958] & sel_one_hot_i[116];
  assign data_masked[14957] = data_i[14957] & sel_one_hot_i[116];
  assign data_masked[14956] = data_i[14956] & sel_one_hot_i[116];
  assign data_masked[14955] = data_i[14955] & sel_one_hot_i[116];
  assign data_masked[14954] = data_i[14954] & sel_one_hot_i[116];
  assign data_masked[14953] = data_i[14953] & sel_one_hot_i[116];
  assign data_masked[14952] = data_i[14952] & sel_one_hot_i[116];
  assign data_masked[14951] = data_i[14951] & sel_one_hot_i[116];
  assign data_masked[14950] = data_i[14950] & sel_one_hot_i[116];
  assign data_masked[14949] = data_i[14949] & sel_one_hot_i[116];
  assign data_masked[14948] = data_i[14948] & sel_one_hot_i[116];
  assign data_masked[14947] = data_i[14947] & sel_one_hot_i[116];
  assign data_masked[14946] = data_i[14946] & sel_one_hot_i[116];
  assign data_masked[14945] = data_i[14945] & sel_one_hot_i[116];
  assign data_masked[14944] = data_i[14944] & sel_one_hot_i[116];
  assign data_masked[14943] = data_i[14943] & sel_one_hot_i[116];
  assign data_masked[14942] = data_i[14942] & sel_one_hot_i[116];
  assign data_masked[14941] = data_i[14941] & sel_one_hot_i[116];
  assign data_masked[14940] = data_i[14940] & sel_one_hot_i[116];
  assign data_masked[14939] = data_i[14939] & sel_one_hot_i[116];
  assign data_masked[14938] = data_i[14938] & sel_one_hot_i[116];
  assign data_masked[14937] = data_i[14937] & sel_one_hot_i[116];
  assign data_masked[14936] = data_i[14936] & sel_one_hot_i[116];
  assign data_masked[14935] = data_i[14935] & sel_one_hot_i[116];
  assign data_masked[14934] = data_i[14934] & sel_one_hot_i[116];
  assign data_masked[14933] = data_i[14933] & sel_one_hot_i[116];
  assign data_masked[14932] = data_i[14932] & sel_one_hot_i[116];
  assign data_masked[14931] = data_i[14931] & sel_one_hot_i[116];
  assign data_masked[14930] = data_i[14930] & sel_one_hot_i[116];
  assign data_masked[14929] = data_i[14929] & sel_one_hot_i[116];
  assign data_masked[14928] = data_i[14928] & sel_one_hot_i[116];
  assign data_masked[14927] = data_i[14927] & sel_one_hot_i[116];
  assign data_masked[14926] = data_i[14926] & sel_one_hot_i[116];
  assign data_masked[14925] = data_i[14925] & sel_one_hot_i[116];
  assign data_masked[14924] = data_i[14924] & sel_one_hot_i[116];
  assign data_masked[14923] = data_i[14923] & sel_one_hot_i[116];
  assign data_masked[14922] = data_i[14922] & sel_one_hot_i[116];
  assign data_masked[14921] = data_i[14921] & sel_one_hot_i[116];
  assign data_masked[14920] = data_i[14920] & sel_one_hot_i[116];
  assign data_masked[14919] = data_i[14919] & sel_one_hot_i[116];
  assign data_masked[14918] = data_i[14918] & sel_one_hot_i[116];
  assign data_masked[14917] = data_i[14917] & sel_one_hot_i[116];
  assign data_masked[14916] = data_i[14916] & sel_one_hot_i[116];
  assign data_masked[14915] = data_i[14915] & sel_one_hot_i[116];
  assign data_masked[14914] = data_i[14914] & sel_one_hot_i[116];
  assign data_masked[14913] = data_i[14913] & sel_one_hot_i[116];
  assign data_masked[14912] = data_i[14912] & sel_one_hot_i[116];
  assign data_masked[14911] = data_i[14911] & sel_one_hot_i[116];
  assign data_masked[14910] = data_i[14910] & sel_one_hot_i[116];
  assign data_masked[14909] = data_i[14909] & sel_one_hot_i[116];
  assign data_masked[14908] = data_i[14908] & sel_one_hot_i[116];
  assign data_masked[14907] = data_i[14907] & sel_one_hot_i[116];
  assign data_masked[14906] = data_i[14906] & sel_one_hot_i[116];
  assign data_masked[14905] = data_i[14905] & sel_one_hot_i[116];
  assign data_masked[14904] = data_i[14904] & sel_one_hot_i[116];
  assign data_masked[14903] = data_i[14903] & sel_one_hot_i[116];
  assign data_masked[14902] = data_i[14902] & sel_one_hot_i[116];
  assign data_masked[14901] = data_i[14901] & sel_one_hot_i[116];
  assign data_masked[14900] = data_i[14900] & sel_one_hot_i[116];
  assign data_masked[14899] = data_i[14899] & sel_one_hot_i[116];
  assign data_masked[14898] = data_i[14898] & sel_one_hot_i[116];
  assign data_masked[14897] = data_i[14897] & sel_one_hot_i[116];
  assign data_masked[14896] = data_i[14896] & sel_one_hot_i[116];
  assign data_masked[14895] = data_i[14895] & sel_one_hot_i[116];
  assign data_masked[14894] = data_i[14894] & sel_one_hot_i[116];
  assign data_masked[14893] = data_i[14893] & sel_one_hot_i[116];
  assign data_masked[14892] = data_i[14892] & sel_one_hot_i[116];
  assign data_masked[14891] = data_i[14891] & sel_one_hot_i[116];
  assign data_masked[14890] = data_i[14890] & sel_one_hot_i[116];
  assign data_masked[14889] = data_i[14889] & sel_one_hot_i[116];
  assign data_masked[14888] = data_i[14888] & sel_one_hot_i[116];
  assign data_masked[14887] = data_i[14887] & sel_one_hot_i[116];
  assign data_masked[14886] = data_i[14886] & sel_one_hot_i[116];
  assign data_masked[14885] = data_i[14885] & sel_one_hot_i[116];
  assign data_masked[14884] = data_i[14884] & sel_one_hot_i[116];
  assign data_masked[14883] = data_i[14883] & sel_one_hot_i[116];
  assign data_masked[14882] = data_i[14882] & sel_one_hot_i[116];
  assign data_masked[14881] = data_i[14881] & sel_one_hot_i[116];
  assign data_masked[14880] = data_i[14880] & sel_one_hot_i[116];
  assign data_masked[14879] = data_i[14879] & sel_one_hot_i[116];
  assign data_masked[14878] = data_i[14878] & sel_one_hot_i[116];
  assign data_masked[14877] = data_i[14877] & sel_one_hot_i[116];
  assign data_masked[14876] = data_i[14876] & sel_one_hot_i[116];
  assign data_masked[14875] = data_i[14875] & sel_one_hot_i[116];
  assign data_masked[14874] = data_i[14874] & sel_one_hot_i[116];
  assign data_masked[14873] = data_i[14873] & sel_one_hot_i[116];
  assign data_masked[14872] = data_i[14872] & sel_one_hot_i[116];
  assign data_masked[14871] = data_i[14871] & sel_one_hot_i[116];
  assign data_masked[14870] = data_i[14870] & sel_one_hot_i[116];
  assign data_masked[14869] = data_i[14869] & sel_one_hot_i[116];
  assign data_masked[14868] = data_i[14868] & sel_one_hot_i[116];
  assign data_masked[14867] = data_i[14867] & sel_one_hot_i[116];
  assign data_masked[14866] = data_i[14866] & sel_one_hot_i[116];
  assign data_masked[14865] = data_i[14865] & sel_one_hot_i[116];
  assign data_masked[14864] = data_i[14864] & sel_one_hot_i[116];
  assign data_masked[14863] = data_i[14863] & sel_one_hot_i[116];
  assign data_masked[14862] = data_i[14862] & sel_one_hot_i[116];
  assign data_masked[14861] = data_i[14861] & sel_one_hot_i[116];
  assign data_masked[14860] = data_i[14860] & sel_one_hot_i[116];
  assign data_masked[14859] = data_i[14859] & sel_one_hot_i[116];
  assign data_masked[14858] = data_i[14858] & sel_one_hot_i[116];
  assign data_masked[14857] = data_i[14857] & sel_one_hot_i[116];
  assign data_masked[14856] = data_i[14856] & sel_one_hot_i[116];
  assign data_masked[14855] = data_i[14855] & sel_one_hot_i[116];
  assign data_masked[14854] = data_i[14854] & sel_one_hot_i[116];
  assign data_masked[14853] = data_i[14853] & sel_one_hot_i[116];
  assign data_masked[14852] = data_i[14852] & sel_one_hot_i[116];
  assign data_masked[14851] = data_i[14851] & sel_one_hot_i[116];
  assign data_masked[14850] = data_i[14850] & sel_one_hot_i[116];
  assign data_masked[14849] = data_i[14849] & sel_one_hot_i[116];
  assign data_masked[14848] = data_i[14848] & sel_one_hot_i[116];
  assign data_masked[15103] = data_i[15103] & sel_one_hot_i[117];
  assign data_masked[15102] = data_i[15102] & sel_one_hot_i[117];
  assign data_masked[15101] = data_i[15101] & sel_one_hot_i[117];
  assign data_masked[15100] = data_i[15100] & sel_one_hot_i[117];
  assign data_masked[15099] = data_i[15099] & sel_one_hot_i[117];
  assign data_masked[15098] = data_i[15098] & sel_one_hot_i[117];
  assign data_masked[15097] = data_i[15097] & sel_one_hot_i[117];
  assign data_masked[15096] = data_i[15096] & sel_one_hot_i[117];
  assign data_masked[15095] = data_i[15095] & sel_one_hot_i[117];
  assign data_masked[15094] = data_i[15094] & sel_one_hot_i[117];
  assign data_masked[15093] = data_i[15093] & sel_one_hot_i[117];
  assign data_masked[15092] = data_i[15092] & sel_one_hot_i[117];
  assign data_masked[15091] = data_i[15091] & sel_one_hot_i[117];
  assign data_masked[15090] = data_i[15090] & sel_one_hot_i[117];
  assign data_masked[15089] = data_i[15089] & sel_one_hot_i[117];
  assign data_masked[15088] = data_i[15088] & sel_one_hot_i[117];
  assign data_masked[15087] = data_i[15087] & sel_one_hot_i[117];
  assign data_masked[15086] = data_i[15086] & sel_one_hot_i[117];
  assign data_masked[15085] = data_i[15085] & sel_one_hot_i[117];
  assign data_masked[15084] = data_i[15084] & sel_one_hot_i[117];
  assign data_masked[15083] = data_i[15083] & sel_one_hot_i[117];
  assign data_masked[15082] = data_i[15082] & sel_one_hot_i[117];
  assign data_masked[15081] = data_i[15081] & sel_one_hot_i[117];
  assign data_masked[15080] = data_i[15080] & sel_one_hot_i[117];
  assign data_masked[15079] = data_i[15079] & sel_one_hot_i[117];
  assign data_masked[15078] = data_i[15078] & sel_one_hot_i[117];
  assign data_masked[15077] = data_i[15077] & sel_one_hot_i[117];
  assign data_masked[15076] = data_i[15076] & sel_one_hot_i[117];
  assign data_masked[15075] = data_i[15075] & sel_one_hot_i[117];
  assign data_masked[15074] = data_i[15074] & sel_one_hot_i[117];
  assign data_masked[15073] = data_i[15073] & sel_one_hot_i[117];
  assign data_masked[15072] = data_i[15072] & sel_one_hot_i[117];
  assign data_masked[15071] = data_i[15071] & sel_one_hot_i[117];
  assign data_masked[15070] = data_i[15070] & sel_one_hot_i[117];
  assign data_masked[15069] = data_i[15069] & sel_one_hot_i[117];
  assign data_masked[15068] = data_i[15068] & sel_one_hot_i[117];
  assign data_masked[15067] = data_i[15067] & sel_one_hot_i[117];
  assign data_masked[15066] = data_i[15066] & sel_one_hot_i[117];
  assign data_masked[15065] = data_i[15065] & sel_one_hot_i[117];
  assign data_masked[15064] = data_i[15064] & sel_one_hot_i[117];
  assign data_masked[15063] = data_i[15063] & sel_one_hot_i[117];
  assign data_masked[15062] = data_i[15062] & sel_one_hot_i[117];
  assign data_masked[15061] = data_i[15061] & sel_one_hot_i[117];
  assign data_masked[15060] = data_i[15060] & sel_one_hot_i[117];
  assign data_masked[15059] = data_i[15059] & sel_one_hot_i[117];
  assign data_masked[15058] = data_i[15058] & sel_one_hot_i[117];
  assign data_masked[15057] = data_i[15057] & sel_one_hot_i[117];
  assign data_masked[15056] = data_i[15056] & sel_one_hot_i[117];
  assign data_masked[15055] = data_i[15055] & sel_one_hot_i[117];
  assign data_masked[15054] = data_i[15054] & sel_one_hot_i[117];
  assign data_masked[15053] = data_i[15053] & sel_one_hot_i[117];
  assign data_masked[15052] = data_i[15052] & sel_one_hot_i[117];
  assign data_masked[15051] = data_i[15051] & sel_one_hot_i[117];
  assign data_masked[15050] = data_i[15050] & sel_one_hot_i[117];
  assign data_masked[15049] = data_i[15049] & sel_one_hot_i[117];
  assign data_masked[15048] = data_i[15048] & sel_one_hot_i[117];
  assign data_masked[15047] = data_i[15047] & sel_one_hot_i[117];
  assign data_masked[15046] = data_i[15046] & sel_one_hot_i[117];
  assign data_masked[15045] = data_i[15045] & sel_one_hot_i[117];
  assign data_masked[15044] = data_i[15044] & sel_one_hot_i[117];
  assign data_masked[15043] = data_i[15043] & sel_one_hot_i[117];
  assign data_masked[15042] = data_i[15042] & sel_one_hot_i[117];
  assign data_masked[15041] = data_i[15041] & sel_one_hot_i[117];
  assign data_masked[15040] = data_i[15040] & sel_one_hot_i[117];
  assign data_masked[15039] = data_i[15039] & sel_one_hot_i[117];
  assign data_masked[15038] = data_i[15038] & sel_one_hot_i[117];
  assign data_masked[15037] = data_i[15037] & sel_one_hot_i[117];
  assign data_masked[15036] = data_i[15036] & sel_one_hot_i[117];
  assign data_masked[15035] = data_i[15035] & sel_one_hot_i[117];
  assign data_masked[15034] = data_i[15034] & sel_one_hot_i[117];
  assign data_masked[15033] = data_i[15033] & sel_one_hot_i[117];
  assign data_masked[15032] = data_i[15032] & sel_one_hot_i[117];
  assign data_masked[15031] = data_i[15031] & sel_one_hot_i[117];
  assign data_masked[15030] = data_i[15030] & sel_one_hot_i[117];
  assign data_masked[15029] = data_i[15029] & sel_one_hot_i[117];
  assign data_masked[15028] = data_i[15028] & sel_one_hot_i[117];
  assign data_masked[15027] = data_i[15027] & sel_one_hot_i[117];
  assign data_masked[15026] = data_i[15026] & sel_one_hot_i[117];
  assign data_masked[15025] = data_i[15025] & sel_one_hot_i[117];
  assign data_masked[15024] = data_i[15024] & sel_one_hot_i[117];
  assign data_masked[15023] = data_i[15023] & sel_one_hot_i[117];
  assign data_masked[15022] = data_i[15022] & sel_one_hot_i[117];
  assign data_masked[15021] = data_i[15021] & sel_one_hot_i[117];
  assign data_masked[15020] = data_i[15020] & sel_one_hot_i[117];
  assign data_masked[15019] = data_i[15019] & sel_one_hot_i[117];
  assign data_masked[15018] = data_i[15018] & sel_one_hot_i[117];
  assign data_masked[15017] = data_i[15017] & sel_one_hot_i[117];
  assign data_masked[15016] = data_i[15016] & sel_one_hot_i[117];
  assign data_masked[15015] = data_i[15015] & sel_one_hot_i[117];
  assign data_masked[15014] = data_i[15014] & sel_one_hot_i[117];
  assign data_masked[15013] = data_i[15013] & sel_one_hot_i[117];
  assign data_masked[15012] = data_i[15012] & sel_one_hot_i[117];
  assign data_masked[15011] = data_i[15011] & sel_one_hot_i[117];
  assign data_masked[15010] = data_i[15010] & sel_one_hot_i[117];
  assign data_masked[15009] = data_i[15009] & sel_one_hot_i[117];
  assign data_masked[15008] = data_i[15008] & sel_one_hot_i[117];
  assign data_masked[15007] = data_i[15007] & sel_one_hot_i[117];
  assign data_masked[15006] = data_i[15006] & sel_one_hot_i[117];
  assign data_masked[15005] = data_i[15005] & sel_one_hot_i[117];
  assign data_masked[15004] = data_i[15004] & sel_one_hot_i[117];
  assign data_masked[15003] = data_i[15003] & sel_one_hot_i[117];
  assign data_masked[15002] = data_i[15002] & sel_one_hot_i[117];
  assign data_masked[15001] = data_i[15001] & sel_one_hot_i[117];
  assign data_masked[15000] = data_i[15000] & sel_one_hot_i[117];
  assign data_masked[14999] = data_i[14999] & sel_one_hot_i[117];
  assign data_masked[14998] = data_i[14998] & sel_one_hot_i[117];
  assign data_masked[14997] = data_i[14997] & sel_one_hot_i[117];
  assign data_masked[14996] = data_i[14996] & sel_one_hot_i[117];
  assign data_masked[14995] = data_i[14995] & sel_one_hot_i[117];
  assign data_masked[14994] = data_i[14994] & sel_one_hot_i[117];
  assign data_masked[14993] = data_i[14993] & sel_one_hot_i[117];
  assign data_masked[14992] = data_i[14992] & sel_one_hot_i[117];
  assign data_masked[14991] = data_i[14991] & sel_one_hot_i[117];
  assign data_masked[14990] = data_i[14990] & sel_one_hot_i[117];
  assign data_masked[14989] = data_i[14989] & sel_one_hot_i[117];
  assign data_masked[14988] = data_i[14988] & sel_one_hot_i[117];
  assign data_masked[14987] = data_i[14987] & sel_one_hot_i[117];
  assign data_masked[14986] = data_i[14986] & sel_one_hot_i[117];
  assign data_masked[14985] = data_i[14985] & sel_one_hot_i[117];
  assign data_masked[14984] = data_i[14984] & sel_one_hot_i[117];
  assign data_masked[14983] = data_i[14983] & sel_one_hot_i[117];
  assign data_masked[14982] = data_i[14982] & sel_one_hot_i[117];
  assign data_masked[14981] = data_i[14981] & sel_one_hot_i[117];
  assign data_masked[14980] = data_i[14980] & sel_one_hot_i[117];
  assign data_masked[14979] = data_i[14979] & sel_one_hot_i[117];
  assign data_masked[14978] = data_i[14978] & sel_one_hot_i[117];
  assign data_masked[14977] = data_i[14977] & sel_one_hot_i[117];
  assign data_masked[14976] = data_i[14976] & sel_one_hot_i[117];
  assign data_masked[15231] = data_i[15231] & sel_one_hot_i[118];
  assign data_masked[15230] = data_i[15230] & sel_one_hot_i[118];
  assign data_masked[15229] = data_i[15229] & sel_one_hot_i[118];
  assign data_masked[15228] = data_i[15228] & sel_one_hot_i[118];
  assign data_masked[15227] = data_i[15227] & sel_one_hot_i[118];
  assign data_masked[15226] = data_i[15226] & sel_one_hot_i[118];
  assign data_masked[15225] = data_i[15225] & sel_one_hot_i[118];
  assign data_masked[15224] = data_i[15224] & sel_one_hot_i[118];
  assign data_masked[15223] = data_i[15223] & sel_one_hot_i[118];
  assign data_masked[15222] = data_i[15222] & sel_one_hot_i[118];
  assign data_masked[15221] = data_i[15221] & sel_one_hot_i[118];
  assign data_masked[15220] = data_i[15220] & sel_one_hot_i[118];
  assign data_masked[15219] = data_i[15219] & sel_one_hot_i[118];
  assign data_masked[15218] = data_i[15218] & sel_one_hot_i[118];
  assign data_masked[15217] = data_i[15217] & sel_one_hot_i[118];
  assign data_masked[15216] = data_i[15216] & sel_one_hot_i[118];
  assign data_masked[15215] = data_i[15215] & sel_one_hot_i[118];
  assign data_masked[15214] = data_i[15214] & sel_one_hot_i[118];
  assign data_masked[15213] = data_i[15213] & sel_one_hot_i[118];
  assign data_masked[15212] = data_i[15212] & sel_one_hot_i[118];
  assign data_masked[15211] = data_i[15211] & sel_one_hot_i[118];
  assign data_masked[15210] = data_i[15210] & sel_one_hot_i[118];
  assign data_masked[15209] = data_i[15209] & sel_one_hot_i[118];
  assign data_masked[15208] = data_i[15208] & sel_one_hot_i[118];
  assign data_masked[15207] = data_i[15207] & sel_one_hot_i[118];
  assign data_masked[15206] = data_i[15206] & sel_one_hot_i[118];
  assign data_masked[15205] = data_i[15205] & sel_one_hot_i[118];
  assign data_masked[15204] = data_i[15204] & sel_one_hot_i[118];
  assign data_masked[15203] = data_i[15203] & sel_one_hot_i[118];
  assign data_masked[15202] = data_i[15202] & sel_one_hot_i[118];
  assign data_masked[15201] = data_i[15201] & sel_one_hot_i[118];
  assign data_masked[15200] = data_i[15200] & sel_one_hot_i[118];
  assign data_masked[15199] = data_i[15199] & sel_one_hot_i[118];
  assign data_masked[15198] = data_i[15198] & sel_one_hot_i[118];
  assign data_masked[15197] = data_i[15197] & sel_one_hot_i[118];
  assign data_masked[15196] = data_i[15196] & sel_one_hot_i[118];
  assign data_masked[15195] = data_i[15195] & sel_one_hot_i[118];
  assign data_masked[15194] = data_i[15194] & sel_one_hot_i[118];
  assign data_masked[15193] = data_i[15193] & sel_one_hot_i[118];
  assign data_masked[15192] = data_i[15192] & sel_one_hot_i[118];
  assign data_masked[15191] = data_i[15191] & sel_one_hot_i[118];
  assign data_masked[15190] = data_i[15190] & sel_one_hot_i[118];
  assign data_masked[15189] = data_i[15189] & sel_one_hot_i[118];
  assign data_masked[15188] = data_i[15188] & sel_one_hot_i[118];
  assign data_masked[15187] = data_i[15187] & sel_one_hot_i[118];
  assign data_masked[15186] = data_i[15186] & sel_one_hot_i[118];
  assign data_masked[15185] = data_i[15185] & sel_one_hot_i[118];
  assign data_masked[15184] = data_i[15184] & sel_one_hot_i[118];
  assign data_masked[15183] = data_i[15183] & sel_one_hot_i[118];
  assign data_masked[15182] = data_i[15182] & sel_one_hot_i[118];
  assign data_masked[15181] = data_i[15181] & sel_one_hot_i[118];
  assign data_masked[15180] = data_i[15180] & sel_one_hot_i[118];
  assign data_masked[15179] = data_i[15179] & sel_one_hot_i[118];
  assign data_masked[15178] = data_i[15178] & sel_one_hot_i[118];
  assign data_masked[15177] = data_i[15177] & sel_one_hot_i[118];
  assign data_masked[15176] = data_i[15176] & sel_one_hot_i[118];
  assign data_masked[15175] = data_i[15175] & sel_one_hot_i[118];
  assign data_masked[15174] = data_i[15174] & sel_one_hot_i[118];
  assign data_masked[15173] = data_i[15173] & sel_one_hot_i[118];
  assign data_masked[15172] = data_i[15172] & sel_one_hot_i[118];
  assign data_masked[15171] = data_i[15171] & sel_one_hot_i[118];
  assign data_masked[15170] = data_i[15170] & sel_one_hot_i[118];
  assign data_masked[15169] = data_i[15169] & sel_one_hot_i[118];
  assign data_masked[15168] = data_i[15168] & sel_one_hot_i[118];
  assign data_masked[15167] = data_i[15167] & sel_one_hot_i[118];
  assign data_masked[15166] = data_i[15166] & sel_one_hot_i[118];
  assign data_masked[15165] = data_i[15165] & sel_one_hot_i[118];
  assign data_masked[15164] = data_i[15164] & sel_one_hot_i[118];
  assign data_masked[15163] = data_i[15163] & sel_one_hot_i[118];
  assign data_masked[15162] = data_i[15162] & sel_one_hot_i[118];
  assign data_masked[15161] = data_i[15161] & sel_one_hot_i[118];
  assign data_masked[15160] = data_i[15160] & sel_one_hot_i[118];
  assign data_masked[15159] = data_i[15159] & sel_one_hot_i[118];
  assign data_masked[15158] = data_i[15158] & sel_one_hot_i[118];
  assign data_masked[15157] = data_i[15157] & sel_one_hot_i[118];
  assign data_masked[15156] = data_i[15156] & sel_one_hot_i[118];
  assign data_masked[15155] = data_i[15155] & sel_one_hot_i[118];
  assign data_masked[15154] = data_i[15154] & sel_one_hot_i[118];
  assign data_masked[15153] = data_i[15153] & sel_one_hot_i[118];
  assign data_masked[15152] = data_i[15152] & sel_one_hot_i[118];
  assign data_masked[15151] = data_i[15151] & sel_one_hot_i[118];
  assign data_masked[15150] = data_i[15150] & sel_one_hot_i[118];
  assign data_masked[15149] = data_i[15149] & sel_one_hot_i[118];
  assign data_masked[15148] = data_i[15148] & sel_one_hot_i[118];
  assign data_masked[15147] = data_i[15147] & sel_one_hot_i[118];
  assign data_masked[15146] = data_i[15146] & sel_one_hot_i[118];
  assign data_masked[15145] = data_i[15145] & sel_one_hot_i[118];
  assign data_masked[15144] = data_i[15144] & sel_one_hot_i[118];
  assign data_masked[15143] = data_i[15143] & sel_one_hot_i[118];
  assign data_masked[15142] = data_i[15142] & sel_one_hot_i[118];
  assign data_masked[15141] = data_i[15141] & sel_one_hot_i[118];
  assign data_masked[15140] = data_i[15140] & sel_one_hot_i[118];
  assign data_masked[15139] = data_i[15139] & sel_one_hot_i[118];
  assign data_masked[15138] = data_i[15138] & sel_one_hot_i[118];
  assign data_masked[15137] = data_i[15137] & sel_one_hot_i[118];
  assign data_masked[15136] = data_i[15136] & sel_one_hot_i[118];
  assign data_masked[15135] = data_i[15135] & sel_one_hot_i[118];
  assign data_masked[15134] = data_i[15134] & sel_one_hot_i[118];
  assign data_masked[15133] = data_i[15133] & sel_one_hot_i[118];
  assign data_masked[15132] = data_i[15132] & sel_one_hot_i[118];
  assign data_masked[15131] = data_i[15131] & sel_one_hot_i[118];
  assign data_masked[15130] = data_i[15130] & sel_one_hot_i[118];
  assign data_masked[15129] = data_i[15129] & sel_one_hot_i[118];
  assign data_masked[15128] = data_i[15128] & sel_one_hot_i[118];
  assign data_masked[15127] = data_i[15127] & sel_one_hot_i[118];
  assign data_masked[15126] = data_i[15126] & sel_one_hot_i[118];
  assign data_masked[15125] = data_i[15125] & sel_one_hot_i[118];
  assign data_masked[15124] = data_i[15124] & sel_one_hot_i[118];
  assign data_masked[15123] = data_i[15123] & sel_one_hot_i[118];
  assign data_masked[15122] = data_i[15122] & sel_one_hot_i[118];
  assign data_masked[15121] = data_i[15121] & sel_one_hot_i[118];
  assign data_masked[15120] = data_i[15120] & sel_one_hot_i[118];
  assign data_masked[15119] = data_i[15119] & sel_one_hot_i[118];
  assign data_masked[15118] = data_i[15118] & sel_one_hot_i[118];
  assign data_masked[15117] = data_i[15117] & sel_one_hot_i[118];
  assign data_masked[15116] = data_i[15116] & sel_one_hot_i[118];
  assign data_masked[15115] = data_i[15115] & sel_one_hot_i[118];
  assign data_masked[15114] = data_i[15114] & sel_one_hot_i[118];
  assign data_masked[15113] = data_i[15113] & sel_one_hot_i[118];
  assign data_masked[15112] = data_i[15112] & sel_one_hot_i[118];
  assign data_masked[15111] = data_i[15111] & sel_one_hot_i[118];
  assign data_masked[15110] = data_i[15110] & sel_one_hot_i[118];
  assign data_masked[15109] = data_i[15109] & sel_one_hot_i[118];
  assign data_masked[15108] = data_i[15108] & sel_one_hot_i[118];
  assign data_masked[15107] = data_i[15107] & sel_one_hot_i[118];
  assign data_masked[15106] = data_i[15106] & sel_one_hot_i[118];
  assign data_masked[15105] = data_i[15105] & sel_one_hot_i[118];
  assign data_masked[15104] = data_i[15104] & sel_one_hot_i[118];
  assign data_masked[15359] = data_i[15359] & sel_one_hot_i[119];
  assign data_masked[15358] = data_i[15358] & sel_one_hot_i[119];
  assign data_masked[15357] = data_i[15357] & sel_one_hot_i[119];
  assign data_masked[15356] = data_i[15356] & sel_one_hot_i[119];
  assign data_masked[15355] = data_i[15355] & sel_one_hot_i[119];
  assign data_masked[15354] = data_i[15354] & sel_one_hot_i[119];
  assign data_masked[15353] = data_i[15353] & sel_one_hot_i[119];
  assign data_masked[15352] = data_i[15352] & sel_one_hot_i[119];
  assign data_masked[15351] = data_i[15351] & sel_one_hot_i[119];
  assign data_masked[15350] = data_i[15350] & sel_one_hot_i[119];
  assign data_masked[15349] = data_i[15349] & sel_one_hot_i[119];
  assign data_masked[15348] = data_i[15348] & sel_one_hot_i[119];
  assign data_masked[15347] = data_i[15347] & sel_one_hot_i[119];
  assign data_masked[15346] = data_i[15346] & sel_one_hot_i[119];
  assign data_masked[15345] = data_i[15345] & sel_one_hot_i[119];
  assign data_masked[15344] = data_i[15344] & sel_one_hot_i[119];
  assign data_masked[15343] = data_i[15343] & sel_one_hot_i[119];
  assign data_masked[15342] = data_i[15342] & sel_one_hot_i[119];
  assign data_masked[15341] = data_i[15341] & sel_one_hot_i[119];
  assign data_masked[15340] = data_i[15340] & sel_one_hot_i[119];
  assign data_masked[15339] = data_i[15339] & sel_one_hot_i[119];
  assign data_masked[15338] = data_i[15338] & sel_one_hot_i[119];
  assign data_masked[15337] = data_i[15337] & sel_one_hot_i[119];
  assign data_masked[15336] = data_i[15336] & sel_one_hot_i[119];
  assign data_masked[15335] = data_i[15335] & sel_one_hot_i[119];
  assign data_masked[15334] = data_i[15334] & sel_one_hot_i[119];
  assign data_masked[15333] = data_i[15333] & sel_one_hot_i[119];
  assign data_masked[15332] = data_i[15332] & sel_one_hot_i[119];
  assign data_masked[15331] = data_i[15331] & sel_one_hot_i[119];
  assign data_masked[15330] = data_i[15330] & sel_one_hot_i[119];
  assign data_masked[15329] = data_i[15329] & sel_one_hot_i[119];
  assign data_masked[15328] = data_i[15328] & sel_one_hot_i[119];
  assign data_masked[15327] = data_i[15327] & sel_one_hot_i[119];
  assign data_masked[15326] = data_i[15326] & sel_one_hot_i[119];
  assign data_masked[15325] = data_i[15325] & sel_one_hot_i[119];
  assign data_masked[15324] = data_i[15324] & sel_one_hot_i[119];
  assign data_masked[15323] = data_i[15323] & sel_one_hot_i[119];
  assign data_masked[15322] = data_i[15322] & sel_one_hot_i[119];
  assign data_masked[15321] = data_i[15321] & sel_one_hot_i[119];
  assign data_masked[15320] = data_i[15320] & sel_one_hot_i[119];
  assign data_masked[15319] = data_i[15319] & sel_one_hot_i[119];
  assign data_masked[15318] = data_i[15318] & sel_one_hot_i[119];
  assign data_masked[15317] = data_i[15317] & sel_one_hot_i[119];
  assign data_masked[15316] = data_i[15316] & sel_one_hot_i[119];
  assign data_masked[15315] = data_i[15315] & sel_one_hot_i[119];
  assign data_masked[15314] = data_i[15314] & sel_one_hot_i[119];
  assign data_masked[15313] = data_i[15313] & sel_one_hot_i[119];
  assign data_masked[15312] = data_i[15312] & sel_one_hot_i[119];
  assign data_masked[15311] = data_i[15311] & sel_one_hot_i[119];
  assign data_masked[15310] = data_i[15310] & sel_one_hot_i[119];
  assign data_masked[15309] = data_i[15309] & sel_one_hot_i[119];
  assign data_masked[15308] = data_i[15308] & sel_one_hot_i[119];
  assign data_masked[15307] = data_i[15307] & sel_one_hot_i[119];
  assign data_masked[15306] = data_i[15306] & sel_one_hot_i[119];
  assign data_masked[15305] = data_i[15305] & sel_one_hot_i[119];
  assign data_masked[15304] = data_i[15304] & sel_one_hot_i[119];
  assign data_masked[15303] = data_i[15303] & sel_one_hot_i[119];
  assign data_masked[15302] = data_i[15302] & sel_one_hot_i[119];
  assign data_masked[15301] = data_i[15301] & sel_one_hot_i[119];
  assign data_masked[15300] = data_i[15300] & sel_one_hot_i[119];
  assign data_masked[15299] = data_i[15299] & sel_one_hot_i[119];
  assign data_masked[15298] = data_i[15298] & sel_one_hot_i[119];
  assign data_masked[15297] = data_i[15297] & sel_one_hot_i[119];
  assign data_masked[15296] = data_i[15296] & sel_one_hot_i[119];
  assign data_masked[15295] = data_i[15295] & sel_one_hot_i[119];
  assign data_masked[15294] = data_i[15294] & sel_one_hot_i[119];
  assign data_masked[15293] = data_i[15293] & sel_one_hot_i[119];
  assign data_masked[15292] = data_i[15292] & sel_one_hot_i[119];
  assign data_masked[15291] = data_i[15291] & sel_one_hot_i[119];
  assign data_masked[15290] = data_i[15290] & sel_one_hot_i[119];
  assign data_masked[15289] = data_i[15289] & sel_one_hot_i[119];
  assign data_masked[15288] = data_i[15288] & sel_one_hot_i[119];
  assign data_masked[15287] = data_i[15287] & sel_one_hot_i[119];
  assign data_masked[15286] = data_i[15286] & sel_one_hot_i[119];
  assign data_masked[15285] = data_i[15285] & sel_one_hot_i[119];
  assign data_masked[15284] = data_i[15284] & sel_one_hot_i[119];
  assign data_masked[15283] = data_i[15283] & sel_one_hot_i[119];
  assign data_masked[15282] = data_i[15282] & sel_one_hot_i[119];
  assign data_masked[15281] = data_i[15281] & sel_one_hot_i[119];
  assign data_masked[15280] = data_i[15280] & sel_one_hot_i[119];
  assign data_masked[15279] = data_i[15279] & sel_one_hot_i[119];
  assign data_masked[15278] = data_i[15278] & sel_one_hot_i[119];
  assign data_masked[15277] = data_i[15277] & sel_one_hot_i[119];
  assign data_masked[15276] = data_i[15276] & sel_one_hot_i[119];
  assign data_masked[15275] = data_i[15275] & sel_one_hot_i[119];
  assign data_masked[15274] = data_i[15274] & sel_one_hot_i[119];
  assign data_masked[15273] = data_i[15273] & sel_one_hot_i[119];
  assign data_masked[15272] = data_i[15272] & sel_one_hot_i[119];
  assign data_masked[15271] = data_i[15271] & sel_one_hot_i[119];
  assign data_masked[15270] = data_i[15270] & sel_one_hot_i[119];
  assign data_masked[15269] = data_i[15269] & sel_one_hot_i[119];
  assign data_masked[15268] = data_i[15268] & sel_one_hot_i[119];
  assign data_masked[15267] = data_i[15267] & sel_one_hot_i[119];
  assign data_masked[15266] = data_i[15266] & sel_one_hot_i[119];
  assign data_masked[15265] = data_i[15265] & sel_one_hot_i[119];
  assign data_masked[15264] = data_i[15264] & sel_one_hot_i[119];
  assign data_masked[15263] = data_i[15263] & sel_one_hot_i[119];
  assign data_masked[15262] = data_i[15262] & sel_one_hot_i[119];
  assign data_masked[15261] = data_i[15261] & sel_one_hot_i[119];
  assign data_masked[15260] = data_i[15260] & sel_one_hot_i[119];
  assign data_masked[15259] = data_i[15259] & sel_one_hot_i[119];
  assign data_masked[15258] = data_i[15258] & sel_one_hot_i[119];
  assign data_masked[15257] = data_i[15257] & sel_one_hot_i[119];
  assign data_masked[15256] = data_i[15256] & sel_one_hot_i[119];
  assign data_masked[15255] = data_i[15255] & sel_one_hot_i[119];
  assign data_masked[15254] = data_i[15254] & sel_one_hot_i[119];
  assign data_masked[15253] = data_i[15253] & sel_one_hot_i[119];
  assign data_masked[15252] = data_i[15252] & sel_one_hot_i[119];
  assign data_masked[15251] = data_i[15251] & sel_one_hot_i[119];
  assign data_masked[15250] = data_i[15250] & sel_one_hot_i[119];
  assign data_masked[15249] = data_i[15249] & sel_one_hot_i[119];
  assign data_masked[15248] = data_i[15248] & sel_one_hot_i[119];
  assign data_masked[15247] = data_i[15247] & sel_one_hot_i[119];
  assign data_masked[15246] = data_i[15246] & sel_one_hot_i[119];
  assign data_masked[15245] = data_i[15245] & sel_one_hot_i[119];
  assign data_masked[15244] = data_i[15244] & sel_one_hot_i[119];
  assign data_masked[15243] = data_i[15243] & sel_one_hot_i[119];
  assign data_masked[15242] = data_i[15242] & sel_one_hot_i[119];
  assign data_masked[15241] = data_i[15241] & sel_one_hot_i[119];
  assign data_masked[15240] = data_i[15240] & sel_one_hot_i[119];
  assign data_masked[15239] = data_i[15239] & sel_one_hot_i[119];
  assign data_masked[15238] = data_i[15238] & sel_one_hot_i[119];
  assign data_masked[15237] = data_i[15237] & sel_one_hot_i[119];
  assign data_masked[15236] = data_i[15236] & sel_one_hot_i[119];
  assign data_masked[15235] = data_i[15235] & sel_one_hot_i[119];
  assign data_masked[15234] = data_i[15234] & sel_one_hot_i[119];
  assign data_masked[15233] = data_i[15233] & sel_one_hot_i[119];
  assign data_masked[15232] = data_i[15232] & sel_one_hot_i[119];
  assign data_masked[15487] = data_i[15487] & sel_one_hot_i[120];
  assign data_masked[15486] = data_i[15486] & sel_one_hot_i[120];
  assign data_masked[15485] = data_i[15485] & sel_one_hot_i[120];
  assign data_masked[15484] = data_i[15484] & sel_one_hot_i[120];
  assign data_masked[15483] = data_i[15483] & sel_one_hot_i[120];
  assign data_masked[15482] = data_i[15482] & sel_one_hot_i[120];
  assign data_masked[15481] = data_i[15481] & sel_one_hot_i[120];
  assign data_masked[15480] = data_i[15480] & sel_one_hot_i[120];
  assign data_masked[15479] = data_i[15479] & sel_one_hot_i[120];
  assign data_masked[15478] = data_i[15478] & sel_one_hot_i[120];
  assign data_masked[15477] = data_i[15477] & sel_one_hot_i[120];
  assign data_masked[15476] = data_i[15476] & sel_one_hot_i[120];
  assign data_masked[15475] = data_i[15475] & sel_one_hot_i[120];
  assign data_masked[15474] = data_i[15474] & sel_one_hot_i[120];
  assign data_masked[15473] = data_i[15473] & sel_one_hot_i[120];
  assign data_masked[15472] = data_i[15472] & sel_one_hot_i[120];
  assign data_masked[15471] = data_i[15471] & sel_one_hot_i[120];
  assign data_masked[15470] = data_i[15470] & sel_one_hot_i[120];
  assign data_masked[15469] = data_i[15469] & sel_one_hot_i[120];
  assign data_masked[15468] = data_i[15468] & sel_one_hot_i[120];
  assign data_masked[15467] = data_i[15467] & sel_one_hot_i[120];
  assign data_masked[15466] = data_i[15466] & sel_one_hot_i[120];
  assign data_masked[15465] = data_i[15465] & sel_one_hot_i[120];
  assign data_masked[15464] = data_i[15464] & sel_one_hot_i[120];
  assign data_masked[15463] = data_i[15463] & sel_one_hot_i[120];
  assign data_masked[15462] = data_i[15462] & sel_one_hot_i[120];
  assign data_masked[15461] = data_i[15461] & sel_one_hot_i[120];
  assign data_masked[15460] = data_i[15460] & sel_one_hot_i[120];
  assign data_masked[15459] = data_i[15459] & sel_one_hot_i[120];
  assign data_masked[15458] = data_i[15458] & sel_one_hot_i[120];
  assign data_masked[15457] = data_i[15457] & sel_one_hot_i[120];
  assign data_masked[15456] = data_i[15456] & sel_one_hot_i[120];
  assign data_masked[15455] = data_i[15455] & sel_one_hot_i[120];
  assign data_masked[15454] = data_i[15454] & sel_one_hot_i[120];
  assign data_masked[15453] = data_i[15453] & sel_one_hot_i[120];
  assign data_masked[15452] = data_i[15452] & sel_one_hot_i[120];
  assign data_masked[15451] = data_i[15451] & sel_one_hot_i[120];
  assign data_masked[15450] = data_i[15450] & sel_one_hot_i[120];
  assign data_masked[15449] = data_i[15449] & sel_one_hot_i[120];
  assign data_masked[15448] = data_i[15448] & sel_one_hot_i[120];
  assign data_masked[15447] = data_i[15447] & sel_one_hot_i[120];
  assign data_masked[15446] = data_i[15446] & sel_one_hot_i[120];
  assign data_masked[15445] = data_i[15445] & sel_one_hot_i[120];
  assign data_masked[15444] = data_i[15444] & sel_one_hot_i[120];
  assign data_masked[15443] = data_i[15443] & sel_one_hot_i[120];
  assign data_masked[15442] = data_i[15442] & sel_one_hot_i[120];
  assign data_masked[15441] = data_i[15441] & sel_one_hot_i[120];
  assign data_masked[15440] = data_i[15440] & sel_one_hot_i[120];
  assign data_masked[15439] = data_i[15439] & sel_one_hot_i[120];
  assign data_masked[15438] = data_i[15438] & sel_one_hot_i[120];
  assign data_masked[15437] = data_i[15437] & sel_one_hot_i[120];
  assign data_masked[15436] = data_i[15436] & sel_one_hot_i[120];
  assign data_masked[15435] = data_i[15435] & sel_one_hot_i[120];
  assign data_masked[15434] = data_i[15434] & sel_one_hot_i[120];
  assign data_masked[15433] = data_i[15433] & sel_one_hot_i[120];
  assign data_masked[15432] = data_i[15432] & sel_one_hot_i[120];
  assign data_masked[15431] = data_i[15431] & sel_one_hot_i[120];
  assign data_masked[15430] = data_i[15430] & sel_one_hot_i[120];
  assign data_masked[15429] = data_i[15429] & sel_one_hot_i[120];
  assign data_masked[15428] = data_i[15428] & sel_one_hot_i[120];
  assign data_masked[15427] = data_i[15427] & sel_one_hot_i[120];
  assign data_masked[15426] = data_i[15426] & sel_one_hot_i[120];
  assign data_masked[15425] = data_i[15425] & sel_one_hot_i[120];
  assign data_masked[15424] = data_i[15424] & sel_one_hot_i[120];
  assign data_masked[15423] = data_i[15423] & sel_one_hot_i[120];
  assign data_masked[15422] = data_i[15422] & sel_one_hot_i[120];
  assign data_masked[15421] = data_i[15421] & sel_one_hot_i[120];
  assign data_masked[15420] = data_i[15420] & sel_one_hot_i[120];
  assign data_masked[15419] = data_i[15419] & sel_one_hot_i[120];
  assign data_masked[15418] = data_i[15418] & sel_one_hot_i[120];
  assign data_masked[15417] = data_i[15417] & sel_one_hot_i[120];
  assign data_masked[15416] = data_i[15416] & sel_one_hot_i[120];
  assign data_masked[15415] = data_i[15415] & sel_one_hot_i[120];
  assign data_masked[15414] = data_i[15414] & sel_one_hot_i[120];
  assign data_masked[15413] = data_i[15413] & sel_one_hot_i[120];
  assign data_masked[15412] = data_i[15412] & sel_one_hot_i[120];
  assign data_masked[15411] = data_i[15411] & sel_one_hot_i[120];
  assign data_masked[15410] = data_i[15410] & sel_one_hot_i[120];
  assign data_masked[15409] = data_i[15409] & sel_one_hot_i[120];
  assign data_masked[15408] = data_i[15408] & sel_one_hot_i[120];
  assign data_masked[15407] = data_i[15407] & sel_one_hot_i[120];
  assign data_masked[15406] = data_i[15406] & sel_one_hot_i[120];
  assign data_masked[15405] = data_i[15405] & sel_one_hot_i[120];
  assign data_masked[15404] = data_i[15404] & sel_one_hot_i[120];
  assign data_masked[15403] = data_i[15403] & sel_one_hot_i[120];
  assign data_masked[15402] = data_i[15402] & sel_one_hot_i[120];
  assign data_masked[15401] = data_i[15401] & sel_one_hot_i[120];
  assign data_masked[15400] = data_i[15400] & sel_one_hot_i[120];
  assign data_masked[15399] = data_i[15399] & sel_one_hot_i[120];
  assign data_masked[15398] = data_i[15398] & sel_one_hot_i[120];
  assign data_masked[15397] = data_i[15397] & sel_one_hot_i[120];
  assign data_masked[15396] = data_i[15396] & sel_one_hot_i[120];
  assign data_masked[15395] = data_i[15395] & sel_one_hot_i[120];
  assign data_masked[15394] = data_i[15394] & sel_one_hot_i[120];
  assign data_masked[15393] = data_i[15393] & sel_one_hot_i[120];
  assign data_masked[15392] = data_i[15392] & sel_one_hot_i[120];
  assign data_masked[15391] = data_i[15391] & sel_one_hot_i[120];
  assign data_masked[15390] = data_i[15390] & sel_one_hot_i[120];
  assign data_masked[15389] = data_i[15389] & sel_one_hot_i[120];
  assign data_masked[15388] = data_i[15388] & sel_one_hot_i[120];
  assign data_masked[15387] = data_i[15387] & sel_one_hot_i[120];
  assign data_masked[15386] = data_i[15386] & sel_one_hot_i[120];
  assign data_masked[15385] = data_i[15385] & sel_one_hot_i[120];
  assign data_masked[15384] = data_i[15384] & sel_one_hot_i[120];
  assign data_masked[15383] = data_i[15383] & sel_one_hot_i[120];
  assign data_masked[15382] = data_i[15382] & sel_one_hot_i[120];
  assign data_masked[15381] = data_i[15381] & sel_one_hot_i[120];
  assign data_masked[15380] = data_i[15380] & sel_one_hot_i[120];
  assign data_masked[15379] = data_i[15379] & sel_one_hot_i[120];
  assign data_masked[15378] = data_i[15378] & sel_one_hot_i[120];
  assign data_masked[15377] = data_i[15377] & sel_one_hot_i[120];
  assign data_masked[15376] = data_i[15376] & sel_one_hot_i[120];
  assign data_masked[15375] = data_i[15375] & sel_one_hot_i[120];
  assign data_masked[15374] = data_i[15374] & sel_one_hot_i[120];
  assign data_masked[15373] = data_i[15373] & sel_one_hot_i[120];
  assign data_masked[15372] = data_i[15372] & sel_one_hot_i[120];
  assign data_masked[15371] = data_i[15371] & sel_one_hot_i[120];
  assign data_masked[15370] = data_i[15370] & sel_one_hot_i[120];
  assign data_masked[15369] = data_i[15369] & sel_one_hot_i[120];
  assign data_masked[15368] = data_i[15368] & sel_one_hot_i[120];
  assign data_masked[15367] = data_i[15367] & sel_one_hot_i[120];
  assign data_masked[15366] = data_i[15366] & sel_one_hot_i[120];
  assign data_masked[15365] = data_i[15365] & sel_one_hot_i[120];
  assign data_masked[15364] = data_i[15364] & sel_one_hot_i[120];
  assign data_masked[15363] = data_i[15363] & sel_one_hot_i[120];
  assign data_masked[15362] = data_i[15362] & sel_one_hot_i[120];
  assign data_masked[15361] = data_i[15361] & sel_one_hot_i[120];
  assign data_masked[15360] = data_i[15360] & sel_one_hot_i[120];
  assign data_masked[15615] = data_i[15615] & sel_one_hot_i[121];
  assign data_masked[15614] = data_i[15614] & sel_one_hot_i[121];
  assign data_masked[15613] = data_i[15613] & sel_one_hot_i[121];
  assign data_masked[15612] = data_i[15612] & sel_one_hot_i[121];
  assign data_masked[15611] = data_i[15611] & sel_one_hot_i[121];
  assign data_masked[15610] = data_i[15610] & sel_one_hot_i[121];
  assign data_masked[15609] = data_i[15609] & sel_one_hot_i[121];
  assign data_masked[15608] = data_i[15608] & sel_one_hot_i[121];
  assign data_masked[15607] = data_i[15607] & sel_one_hot_i[121];
  assign data_masked[15606] = data_i[15606] & sel_one_hot_i[121];
  assign data_masked[15605] = data_i[15605] & sel_one_hot_i[121];
  assign data_masked[15604] = data_i[15604] & sel_one_hot_i[121];
  assign data_masked[15603] = data_i[15603] & sel_one_hot_i[121];
  assign data_masked[15602] = data_i[15602] & sel_one_hot_i[121];
  assign data_masked[15601] = data_i[15601] & sel_one_hot_i[121];
  assign data_masked[15600] = data_i[15600] & sel_one_hot_i[121];
  assign data_masked[15599] = data_i[15599] & sel_one_hot_i[121];
  assign data_masked[15598] = data_i[15598] & sel_one_hot_i[121];
  assign data_masked[15597] = data_i[15597] & sel_one_hot_i[121];
  assign data_masked[15596] = data_i[15596] & sel_one_hot_i[121];
  assign data_masked[15595] = data_i[15595] & sel_one_hot_i[121];
  assign data_masked[15594] = data_i[15594] & sel_one_hot_i[121];
  assign data_masked[15593] = data_i[15593] & sel_one_hot_i[121];
  assign data_masked[15592] = data_i[15592] & sel_one_hot_i[121];
  assign data_masked[15591] = data_i[15591] & sel_one_hot_i[121];
  assign data_masked[15590] = data_i[15590] & sel_one_hot_i[121];
  assign data_masked[15589] = data_i[15589] & sel_one_hot_i[121];
  assign data_masked[15588] = data_i[15588] & sel_one_hot_i[121];
  assign data_masked[15587] = data_i[15587] & sel_one_hot_i[121];
  assign data_masked[15586] = data_i[15586] & sel_one_hot_i[121];
  assign data_masked[15585] = data_i[15585] & sel_one_hot_i[121];
  assign data_masked[15584] = data_i[15584] & sel_one_hot_i[121];
  assign data_masked[15583] = data_i[15583] & sel_one_hot_i[121];
  assign data_masked[15582] = data_i[15582] & sel_one_hot_i[121];
  assign data_masked[15581] = data_i[15581] & sel_one_hot_i[121];
  assign data_masked[15580] = data_i[15580] & sel_one_hot_i[121];
  assign data_masked[15579] = data_i[15579] & sel_one_hot_i[121];
  assign data_masked[15578] = data_i[15578] & sel_one_hot_i[121];
  assign data_masked[15577] = data_i[15577] & sel_one_hot_i[121];
  assign data_masked[15576] = data_i[15576] & sel_one_hot_i[121];
  assign data_masked[15575] = data_i[15575] & sel_one_hot_i[121];
  assign data_masked[15574] = data_i[15574] & sel_one_hot_i[121];
  assign data_masked[15573] = data_i[15573] & sel_one_hot_i[121];
  assign data_masked[15572] = data_i[15572] & sel_one_hot_i[121];
  assign data_masked[15571] = data_i[15571] & sel_one_hot_i[121];
  assign data_masked[15570] = data_i[15570] & sel_one_hot_i[121];
  assign data_masked[15569] = data_i[15569] & sel_one_hot_i[121];
  assign data_masked[15568] = data_i[15568] & sel_one_hot_i[121];
  assign data_masked[15567] = data_i[15567] & sel_one_hot_i[121];
  assign data_masked[15566] = data_i[15566] & sel_one_hot_i[121];
  assign data_masked[15565] = data_i[15565] & sel_one_hot_i[121];
  assign data_masked[15564] = data_i[15564] & sel_one_hot_i[121];
  assign data_masked[15563] = data_i[15563] & sel_one_hot_i[121];
  assign data_masked[15562] = data_i[15562] & sel_one_hot_i[121];
  assign data_masked[15561] = data_i[15561] & sel_one_hot_i[121];
  assign data_masked[15560] = data_i[15560] & sel_one_hot_i[121];
  assign data_masked[15559] = data_i[15559] & sel_one_hot_i[121];
  assign data_masked[15558] = data_i[15558] & sel_one_hot_i[121];
  assign data_masked[15557] = data_i[15557] & sel_one_hot_i[121];
  assign data_masked[15556] = data_i[15556] & sel_one_hot_i[121];
  assign data_masked[15555] = data_i[15555] & sel_one_hot_i[121];
  assign data_masked[15554] = data_i[15554] & sel_one_hot_i[121];
  assign data_masked[15553] = data_i[15553] & sel_one_hot_i[121];
  assign data_masked[15552] = data_i[15552] & sel_one_hot_i[121];
  assign data_masked[15551] = data_i[15551] & sel_one_hot_i[121];
  assign data_masked[15550] = data_i[15550] & sel_one_hot_i[121];
  assign data_masked[15549] = data_i[15549] & sel_one_hot_i[121];
  assign data_masked[15548] = data_i[15548] & sel_one_hot_i[121];
  assign data_masked[15547] = data_i[15547] & sel_one_hot_i[121];
  assign data_masked[15546] = data_i[15546] & sel_one_hot_i[121];
  assign data_masked[15545] = data_i[15545] & sel_one_hot_i[121];
  assign data_masked[15544] = data_i[15544] & sel_one_hot_i[121];
  assign data_masked[15543] = data_i[15543] & sel_one_hot_i[121];
  assign data_masked[15542] = data_i[15542] & sel_one_hot_i[121];
  assign data_masked[15541] = data_i[15541] & sel_one_hot_i[121];
  assign data_masked[15540] = data_i[15540] & sel_one_hot_i[121];
  assign data_masked[15539] = data_i[15539] & sel_one_hot_i[121];
  assign data_masked[15538] = data_i[15538] & sel_one_hot_i[121];
  assign data_masked[15537] = data_i[15537] & sel_one_hot_i[121];
  assign data_masked[15536] = data_i[15536] & sel_one_hot_i[121];
  assign data_masked[15535] = data_i[15535] & sel_one_hot_i[121];
  assign data_masked[15534] = data_i[15534] & sel_one_hot_i[121];
  assign data_masked[15533] = data_i[15533] & sel_one_hot_i[121];
  assign data_masked[15532] = data_i[15532] & sel_one_hot_i[121];
  assign data_masked[15531] = data_i[15531] & sel_one_hot_i[121];
  assign data_masked[15530] = data_i[15530] & sel_one_hot_i[121];
  assign data_masked[15529] = data_i[15529] & sel_one_hot_i[121];
  assign data_masked[15528] = data_i[15528] & sel_one_hot_i[121];
  assign data_masked[15527] = data_i[15527] & sel_one_hot_i[121];
  assign data_masked[15526] = data_i[15526] & sel_one_hot_i[121];
  assign data_masked[15525] = data_i[15525] & sel_one_hot_i[121];
  assign data_masked[15524] = data_i[15524] & sel_one_hot_i[121];
  assign data_masked[15523] = data_i[15523] & sel_one_hot_i[121];
  assign data_masked[15522] = data_i[15522] & sel_one_hot_i[121];
  assign data_masked[15521] = data_i[15521] & sel_one_hot_i[121];
  assign data_masked[15520] = data_i[15520] & sel_one_hot_i[121];
  assign data_masked[15519] = data_i[15519] & sel_one_hot_i[121];
  assign data_masked[15518] = data_i[15518] & sel_one_hot_i[121];
  assign data_masked[15517] = data_i[15517] & sel_one_hot_i[121];
  assign data_masked[15516] = data_i[15516] & sel_one_hot_i[121];
  assign data_masked[15515] = data_i[15515] & sel_one_hot_i[121];
  assign data_masked[15514] = data_i[15514] & sel_one_hot_i[121];
  assign data_masked[15513] = data_i[15513] & sel_one_hot_i[121];
  assign data_masked[15512] = data_i[15512] & sel_one_hot_i[121];
  assign data_masked[15511] = data_i[15511] & sel_one_hot_i[121];
  assign data_masked[15510] = data_i[15510] & sel_one_hot_i[121];
  assign data_masked[15509] = data_i[15509] & sel_one_hot_i[121];
  assign data_masked[15508] = data_i[15508] & sel_one_hot_i[121];
  assign data_masked[15507] = data_i[15507] & sel_one_hot_i[121];
  assign data_masked[15506] = data_i[15506] & sel_one_hot_i[121];
  assign data_masked[15505] = data_i[15505] & sel_one_hot_i[121];
  assign data_masked[15504] = data_i[15504] & sel_one_hot_i[121];
  assign data_masked[15503] = data_i[15503] & sel_one_hot_i[121];
  assign data_masked[15502] = data_i[15502] & sel_one_hot_i[121];
  assign data_masked[15501] = data_i[15501] & sel_one_hot_i[121];
  assign data_masked[15500] = data_i[15500] & sel_one_hot_i[121];
  assign data_masked[15499] = data_i[15499] & sel_one_hot_i[121];
  assign data_masked[15498] = data_i[15498] & sel_one_hot_i[121];
  assign data_masked[15497] = data_i[15497] & sel_one_hot_i[121];
  assign data_masked[15496] = data_i[15496] & sel_one_hot_i[121];
  assign data_masked[15495] = data_i[15495] & sel_one_hot_i[121];
  assign data_masked[15494] = data_i[15494] & sel_one_hot_i[121];
  assign data_masked[15493] = data_i[15493] & sel_one_hot_i[121];
  assign data_masked[15492] = data_i[15492] & sel_one_hot_i[121];
  assign data_masked[15491] = data_i[15491] & sel_one_hot_i[121];
  assign data_masked[15490] = data_i[15490] & sel_one_hot_i[121];
  assign data_masked[15489] = data_i[15489] & sel_one_hot_i[121];
  assign data_masked[15488] = data_i[15488] & sel_one_hot_i[121];
  assign data_masked[15743] = data_i[15743] & sel_one_hot_i[122];
  assign data_masked[15742] = data_i[15742] & sel_one_hot_i[122];
  assign data_masked[15741] = data_i[15741] & sel_one_hot_i[122];
  assign data_masked[15740] = data_i[15740] & sel_one_hot_i[122];
  assign data_masked[15739] = data_i[15739] & sel_one_hot_i[122];
  assign data_masked[15738] = data_i[15738] & sel_one_hot_i[122];
  assign data_masked[15737] = data_i[15737] & sel_one_hot_i[122];
  assign data_masked[15736] = data_i[15736] & sel_one_hot_i[122];
  assign data_masked[15735] = data_i[15735] & sel_one_hot_i[122];
  assign data_masked[15734] = data_i[15734] & sel_one_hot_i[122];
  assign data_masked[15733] = data_i[15733] & sel_one_hot_i[122];
  assign data_masked[15732] = data_i[15732] & sel_one_hot_i[122];
  assign data_masked[15731] = data_i[15731] & sel_one_hot_i[122];
  assign data_masked[15730] = data_i[15730] & sel_one_hot_i[122];
  assign data_masked[15729] = data_i[15729] & sel_one_hot_i[122];
  assign data_masked[15728] = data_i[15728] & sel_one_hot_i[122];
  assign data_masked[15727] = data_i[15727] & sel_one_hot_i[122];
  assign data_masked[15726] = data_i[15726] & sel_one_hot_i[122];
  assign data_masked[15725] = data_i[15725] & sel_one_hot_i[122];
  assign data_masked[15724] = data_i[15724] & sel_one_hot_i[122];
  assign data_masked[15723] = data_i[15723] & sel_one_hot_i[122];
  assign data_masked[15722] = data_i[15722] & sel_one_hot_i[122];
  assign data_masked[15721] = data_i[15721] & sel_one_hot_i[122];
  assign data_masked[15720] = data_i[15720] & sel_one_hot_i[122];
  assign data_masked[15719] = data_i[15719] & sel_one_hot_i[122];
  assign data_masked[15718] = data_i[15718] & sel_one_hot_i[122];
  assign data_masked[15717] = data_i[15717] & sel_one_hot_i[122];
  assign data_masked[15716] = data_i[15716] & sel_one_hot_i[122];
  assign data_masked[15715] = data_i[15715] & sel_one_hot_i[122];
  assign data_masked[15714] = data_i[15714] & sel_one_hot_i[122];
  assign data_masked[15713] = data_i[15713] & sel_one_hot_i[122];
  assign data_masked[15712] = data_i[15712] & sel_one_hot_i[122];
  assign data_masked[15711] = data_i[15711] & sel_one_hot_i[122];
  assign data_masked[15710] = data_i[15710] & sel_one_hot_i[122];
  assign data_masked[15709] = data_i[15709] & sel_one_hot_i[122];
  assign data_masked[15708] = data_i[15708] & sel_one_hot_i[122];
  assign data_masked[15707] = data_i[15707] & sel_one_hot_i[122];
  assign data_masked[15706] = data_i[15706] & sel_one_hot_i[122];
  assign data_masked[15705] = data_i[15705] & sel_one_hot_i[122];
  assign data_masked[15704] = data_i[15704] & sel_one_hot_i[122];
  assign data_masked[15703] = data_i[15703] & sel_one_hot_i[122];
  assign data_masked[15702] = data_i[15702] & sel_one_hot_i[122];
  assign data_masked[15701] = data_i[15701] & sel_one_hot_i[122];
  assign data_masked[15700] = data_i[15700] & sel_one_hot_i[122];
  assign data_masked[15699] = data_i[15699] & sel_one_hot_i[122];
  assign data_masked[15698] = data_i[15698] & sel_one_hot_i[122];
  assign data_masked[15697] = data_i[15697] & sel_one_hot_i[122];
  assign data_masked[15696] = data_i[15696] & sel_one_hot_i[122];
  assign data_masked[15695] = data_i[15695] & sel_one_hot_i[122];
  assign data_masked[15694] = data_i[15694] & sel_one_hot_i[122];
  assign data_masked[15693] = data_i[15693] & sel_one_hot_i[122];
  assign data_masked[15692] = data_i[15692] & sel_one_hot_i[122];
  assign data_masked[15691] = data_i[15691] & sel_one_hot_i[122];
  assign data_masked[15690] = data_i[15690] & sel_one_hot_i[122];
  assign data_masked[15689] = data_i[15689] & sel_one_hot_i[122];
  assign data_masked[15688] = data_i[15688] & sel_one_hot_i[122];
  assign data_masked[15687] = data_i[15687] & sel_one_hot_i[122];
  assign data_masked[15686] = data_i[15686] & sel_one_hot_i[122];
  assign data_masked[15685] = data_i[15685] & sel_one_hot_i[122];
  assign data_masked[15684] = data_i[15684] & sel_one_hot_i[122];
  assign data_masked[15683] = data_i[15683] & sel_one_hot_i[122];
  assign data_masked[15682] = data_i[15682] & sel_one_hot_i[122];
  assign data_masked[15681] = data_i[15681] & sel_one_hot_i[122];
  assign data_masked[15680] = data_i[15680] & sel_one_hot_i[122];
  assign data_masked[15679] = data_i[15679] & sel_one_hot_i[122];
  assign data_masked[15678] = data_i[15678] & sel_one_hot_i[122];
  assign data_masked[15677] = data_i[15677] & sel_one_hot_i[122];
  assign data_masked[15676] = data_i[15676] & sel_one_hot_i[122];
  assign data_masked[15675] = data_i[15675] & sel_one_hot_i[122];
  assign data_masked[15674] = data_i[15674] & sel_one_hot_i[122];
  assign data_masked[15673] = data_i[15673] & sel_one_hot_i[122];
  assign data_masked[15672] = data_i[15672] & sel_one_hot_i[122];
  assign data_masked[15671] = data_i[15671] & sel_one_hot_i[122];
  assign data_masked[15670] = data_i[15670] & sel_one_hot_i[122];
  assign data_masked[15669] = data_i[15669] & sel_one_hot_i[122];
  assign data_masked[15668] = data_i[15668] & sel_one_hot_i[122];
  assign data_masked[15667] = data_i[15667] & sel_one_hot_i[122];
  assign data_masked[15666] = data_i[15666] & sel_one_hot_i[122];
  assign data_masked[15665] = data_i[15665] & sel_one_hot_i[122];
  assign data_masked[15664] = data_i[15664] & sel_one_hot_i[122];
  assign data_masked[15663] = data_i[15663] & sel_one_hot_i[122];
  assign data_masked[15662] = data_i[15662] & sel_one_hot_i[122];
  assign data_masked[15661] = data_i[15661] & sel_one_hot_i[122];
  assign data_masked[15660] = data_i[15660] & sel_one_hot_i[122];
  assign data_masked[15659] = data_i[15659] & sel_one_hot_i[122];
  assign data_masked[15658] = data_i[15658] & sel_one_hot_i[122];
  assign data_masked[15657] = data_i[15657] & sel_one_hot_i[122];
  assign data_masked[15656] = data_i[15656] & sel_one_hot_i[122];
  assign data_masked[15655] = data_i[15655] & sel_one_hot_i[122];
  assign data_masked[15654] = data_i[15654] & sel_one_hot_i[122];
  assign data_masked[15653] = data_i[15653] & sel_one_hot_i[122];
  assign data_masked[15652] = data_i[15652] & sel_one_hot_i[122];
  assign data_masked[15651] = data_i[15651] & sel_one_hot_i[122];
  assign data_masked[15650] = data_i[15650] & sel_one_hot_i[122];
  assign data_masked[15649] = data_i[15649] & sel_one_hot_i[122];
  assign data_masked[15648] = data_i[15648] & sel_one_hot_i[122];
  assign data_masked[15647] = data_i[15647] & sel_one_hot_i[122];
  assign data_masked[15646] = data_i[15646] & sel_one_hot_i[122];
  assign data_masked[15645] = data_i[15645] & sel_one_hot_i[122];
  assign data_masked[15644] = data_i[15644] & sel_one_hot_i[122];
  assign data_masked[15643] = data_i[15643] & sel_one_hot_i[122];
  assign data_masked[15642] = data_i[15642] & sel_one_hot_i[122];
  assign data_masked[15641] = data_i[15641] & sel_one_hot_i[122];
  assign data_masked[15640] = data_i[15640] & sel_one_hot_i[122];
  assign data_masked[15639] = data_i[15639] & sel_one_hot_i[122];
  assign data_masked[15638] = data_i[15638] & sel_one_hot_i[122];
  assign data_masked[15637] = data_i[15637] & sel_one_hot_i[122];
  assign data_masked[15636] = data_i[15636] & sel_one_hot_i[122];
  assign data_masked[15635] = data_i[15635] & sel_one_hot_i[122];
  assign data_masked[15634] = data_i[15634] & sel_one_hot_i[122];
  assign data_masked[15633] = data_i[15633] & sel_one_hot_i[122];
  assign data_masked[15632] = data_i[15632] & sel_one_hot_i[122];
  assign data_masked[15631] = data_i[15631] & sel_one_hot_i[122];
  assign data_masked[15630] = data_i[15630] & sel_one_hot_i[122];
  assign data_masked[15629] = data_i[15629] & sel_one_hot_i[122];
  assign data_masked[15628] = data_i[15628] & sel_one_hot_i[122];
  assign data_masked[15627] = data_i[15627] & sel_one_hot_i[122];
  assign data_masked[15626] = data_i[15626] & sel_one_hot_i[122];
  assign data_masked[15625] = data_i[15625] & sel_one_hot_i[122];
  assign data_masked[15624] = data_i[15624] & sel_one_hot_i[122];
  assign data_masked[15623] = data_i[15623] & sel_one_hot_i[122];
  assign data_masked[15622] = data_i[15622] & sel_one_hot_i[122];
  assign data_masked[15621] = data_i[15621] & sel_one_hot_i[122];
  assign data_masked[15620] = data_i[15620] & sel_one_hot_i[122];
  assign data_masked[15619] = data_i[15619] & sel_one_hot_i[122];
  assign data_masked[15618] = data_i[15618] & sel_one_hot_i[122];
  assign data_masked[15617] = data_i[15617] & sel_one_hot_i[122];
  assign data_masked[15616] = data_i[15616] & sel_one_hot_i[122];
  assign data_masked[15871] = data_i[15871] & sel_one_hot_i[123];
  assign data_masked[15870] = data_i[15870] & sel_one_hot_i[123];
  assign data_masked[15869] = data_i[15869] & sel_one_hot_i[123];
  assign data_masked[15868] = data_i[15868] & sel_one_hot_i[123];
  assign data_masked[15867] = data_i[15867] & sel_one_hot_i[123];
  assign data_masked[15866] = data_i[15866] & sel_one_hot_i[123];
  assign data_masked[15865] = data_i[15865] & sel_one_hot_i[123];
  assign data_masked[15864] = data_i[15864] & sel_one_hot_i[123];
  assign data_masked[15863] = data_i[15863] & sel_one_hot_i[123];
  assign data_masked[15862] = data_i[15862] & sel_one_hot_i[123];
  assign data_masked[15861] = data_i[15861] & sel_one_hot_i[123];
  assign data_masked[15860] = data_i[15860] & sel_one_hot_i[123];
  assign data_masked[15859] = data_i[15859] & sel_one_hot_i[123];
  assign data_masked[15858] = data_i[15858] & sel_one_hot_i[123];
  assign data_masked[15857] = data_i[15857] & sel_one_hot_i[123];
  assign data_masked[15856] = data_i[15856] & sel_one_hot_i[123];
  assign data_masked[15855] = data_i[15855] & sel_one_hot_i[123];
  assign data_masked[15854] = data_i[15854] & sel_one_hot_i[123];
  assign data_masked[15853] = data_i[15853] & sel_one_hot_i[123];
  assign data_masked[15852] = data_i[15852] & sel_one_hot_i[123];
  assign data_masked[15851] = data_i[15851] & sel_one_hot_i[123];
  assign data_masked[15850] = data_i[15850] & sel_one_hot_i[123];
  assign data_masked[15849] = data_i[15849] & sel_one_hot_i[123];
  assign data_masked[15848] = data_i[15848] & sel_one_hot_i[123];
  assign data_masked[15847] = data_i[15847] & sel_one_hot_i[123];
  assign data_masked[15846] = data_i[15846] & sel_one_hot_i[123];
  assign data_masked[15845] = data_i[15845] & sel_one_hot_i[123];
  assign data_masked[15844] = data_i[15844] & sel_one_hot_i[123];
  assign data_masked[15843] = data_i[15843] & sel_one_hot_i[123];
  assign data_masked[15842] = data_i[15842] & sel_one_hot_i[123];
  assign data_masked[15841] = data_i[15841] & sel_one_hot_i[123];
  assign data_masked[15840] = data_i[15840] & sel_one_hot_i[123];
  assign data_masked[15839] = data_i[15839] & sel_one_hot_i[123];
  assign data_masked[15838] = data_i[15838] & sel_one_hot_i[123];
  assign data_masked[15837] = data_i[15837] & sel_one_hot_i[123];
  assign data_masked[15836] = data_i[15836] & sel_one_hot_i[123];
  assign data_masked[15835] = data_i[15835] & sel_one_hot_i[123];
  assign data_masked[15834] = data_i[15834] & sel_one_hot_i[123];
  assign data_masked[15833] = data_i[15833] & sel_one_hot_i[123];
  assign data_masked[15832] = data_i[15832] & sel_one_hot_i[123];
  assign data_masked[15831] = data_i[15831] & sel_one_hot_i[123];
  assign data_masked[15830] = data_i[15830] & sel_one_hot_i[123];
  assign data_masked[15829] = data_i[15829] & sel_one_hot_i[123];
  assign data_masked[15828] = data_i[15828] & sel_one_hot_i[123];
  assign data_masked[15827] = data_i[15827] & sel_one_hot_i[123];
  assign data_masked[15826] = data_i[15826] & sel_one_hot_i[123];
  assign data_masked[15825] = data_i[15825] & sel_one_hot_i[123];
  assign data_masked[15824] = data_i[15824] & sel_one_hot_i[123];
  assign data_masked[15823] = data_i[15823] & sel_one_hot_i[123];
  assign data_masked[15822] = data_i[15822] & sel_one_hot_i[123];
  assign data_masked[15821] = data_i[15821] & sel_one_hot_i[123];
  assign data_masked[15820] = data_i[15820] & sel_one_hot_i[123];
  assign data_masked[15819] = data_i[15819] & sel_one_hot_i[123];
  assign data_masked[15818] = data_i[15818] & sel_one_hot_i[123];
  assign data_masked[15817] = data_i[15817] & sel_one_hot_i[123];
  assign data_masked[15816] = data_i[15816] & sel_one_hot_i[123];
  assign data_masked[15815] = data_i[15815] & sel_one_hot_i[123];
  assign data_masked[15814] = data_i[15814] & sel_one_hot_i[123];
  assign data_masked[15813] = data_i[15813] & sel_one_hot_i[123];
  assign data_masked[15812] = data_i[15812] & sel_one_hot_i[123];
  assign data_masked[15811] = data_i[15811] & sel_one_hot_i[123];
  assign data_masked[15810] = data_i[15810] & sel_one_hot_i[123];
  assign data_masked[15809] = data_i[15809] & sel_one_hot_i[123];
  assign data_masked[15808] = data_i[15808] & sel_one_hot_i[123];
  assign data_masked[15807] = data_i[15807] & sel_one_hot_i[123];
  assign data_masked[15806] = data_i[15806] & sel_one_hot_i[123];
  assign data_masked[15805] = data_i[15805] & sel_one_hot_i[123];
  assign data_masked[15804] = data_i[15804] & sel_one_hot_i[123];
  assign data_masked[15803] = data_i[15803] & sel_one_hot_i[123];
  assign data_masked[15802] = data_i[15802] & sel_one_hot_i[123];
  assign data_masked[15801] = data_i[15801] & sel_one_hot_i[123];
  assign data_masked[15800] = data_i[15800] & sel_one_hot_i[123];
  assign data_masked[15799] = data_i[15799] & sel_one_hot_i[123];
  assign data_masked[15798] = data_i[15798] & sel_one_hot_i[123];
  assign data_masked[15797] = data_i[15797] & sel_one_hot_i[123];
  assign data_masked[15796] = data_i[15796] & sel_one_hot_i[123];
  assign data_masked[15795] = data_i[15795] & sel_one_hot_i[123];
  assign data_masked[15794] = data_i[15794] & sel_one_hot_i[123];
  assign data_masked[15793] = data_i[15793] & sel_one_hot_i[123];
  assign data_masked[15792] = data_i[15792] & sel_one_hot_i[123];
  assign data_masked[15791] = data_i[15791] & sel_one_hot_i[123];
  assign data_masked[15790] = data_i[15790] & sel_one_hot_i[123];
  assign data_masked[15789] = data_i[15789] & sel_one_hot_i[123];
  assign data_masked[15788] = data_i[15788] & sel_one_hot_i[123];
  assign data_masked[15787] = data_i[15787] & sel_one_hot_i[123];
  assign data_masked[15786] = data_i[15786] & sel_one_hot_i[123];
  assign data_masked[15785] = data_i[15785] & sel_one_hot_i[123];
  assign data_masked[15784] = data_i[15784] & sel_one_hot_i[123];
  assign data_masked[15783] = data_i[15783] & sel_one_hot_i[123];
  assign data_masked[15782] = data_i[15782] & sel_one_hot_i[123];
  assign data_masked[15781] = data_i[15781] & sel_one_hot_i[123];
  assign data_masked[15780] = data_i[15780] & sel_one_hot_i[123];
  assign data_masked[15779] = data_i[15779] & sel_one_hot_i[123];
  assign data_masked[15778] = data_i[15778] & sel_one_hot_i[123];
  assign data_masked[15777] = data_i[15777] & sel_one_hot_i[123];
  assign data_masked[15776] = data_i[15776] & sel_one_hot_i[123];
  assign data_masked[15775] = data_i[15775] & sel_one_hot_i[123];
  assign data_masked[15774] = data_i[15774] & sel_one_hot_i[123];
  assign data_masked[15773] = data_i[15773] & sel_one_hot_i[123];
  assign data_masked[15772] = data_i[15772] & sel_one_hot_i[123];
  assign data_masked[15771] = data_i[15771] & sel_one_hot_i[123];
  assign data_masked[15770] = data_i[15770] & sel_one_hot_i[123];
  assign data_masked[15769] = data_i[15769] & sel_one_hot_i[123];
  assign data_masked[15768] = data_i[15768] & sel_one_hot_i[123];
  assign data_masked[15767] = data_i[15767] & sel_one_hot_i[123];
  assign data_masked[15766] = data_i[15766] & sel_one_hot_i[123];
  assign data_masked[15765] = data_i[15765] & sel_one_hot_i[123];
  assign data_masked[15764] = data_i[15764] & sel_one_hot_i[123];
  assign data_masked[15763] = data_i[15763] & sel_one_hot_i[123];
  assign data_masked[15762] = data_i[15762] & sel_one_hot_i[123];
  assign data_masked[15761] = data_i[15761] & sel_one_hot_i[123];
  assign data_masked[15760] = data_i[15760] & sel_one_hot_i[123];
  assign data_masked[15759] = data_i[15759] & sel_one_hot_i[123];
  assign data_masked[15758] = data_i[15758] & sel_one_hot_i[123];
  assign data_masked[15757] = data_i[15757] & sel_one_hot_i[123];
  assign data_masked[15756] = data_i[15756] & sel_one_hot_i[123];
  assign data_masked[15755] = data_i[15755] & sel_one_hot_i[123];
  assign data_masked[15754] = data_i[15754] & sel_one_hot_i[123];
  assign data_masked[15753] = data_i[15753] & sel_one_hot_i[123];
  assign data_masked[15752] = data_i[15752] & sel_one_hot_i[123];
  assign data_masked[15751] = data_i[15751] & sel_one_hot_i[123];
  assign data_masked[15750] = data_i[15750] & sel_one_hot_i[123];
  assign data_masked[15749] = data_i[15749] & sel_one_hot_i[123];
  assign data_masked[15748] = data_i[15748] & sel_one_hot_i[123];
  assign data_masked[15747] = data_i[15747] & sel_one_hot_i[123];
  assign data_masked[15746] = data_i[15746] & sel_one_hot_i[123];
  assign data_masked[15745] = data_i[15745] & sel_one_hot_i[123];
  assign data_masked[15744] = data_i[15744] & sel_one_hot_i[123];
  assign data_masked[15999] = data_i[15999] & sel_one_hot_i[124];
  assign data_masked[15998] = data_i[15998] & sel_one_hot_i[124];
  assign data_masked[15997] = data_i[15997] & sel_one_hot_i[124];
  assign data_masked[15996] = data_i[15996] & sel_one_hot_i[124];
  assign data_masked[15995] = data_i[15995] & sel_one_hot_i[124];
  assign data_masked[15994] = data_i[15994] & sel_one_hot_i[124];
  assign data_masked[15993] = data_i[15993] & sel_one_hot_i[124];
  assign data_masked[15992] = data_i[15992] & sel_one_hot_i[124];
  assign data_masked[15991] = data_i[15991] & sel_one_hot_i[124];
  assign data_masked[15990] = data_i[15990] & sel_one_hot_i[124];
  assign data_masked[15989] = data_i[15989] & sel_one_hot_i[124];
  assign data_masked[15988] = data_i[15988] & sel_one_hot_i[124];
  assign data_masked[15987] = data_i[15987] & sel_one_hot_i[124];
  assign data_masked[15986] = data_i[15986] & sel_one_hot_i[124];
  assign data_masked[15985] = data_i[15985] & sel_one_hot_i[124];
  assign data_masked[15984] = data_i[15984] & sel_one_hot_i[124];
  assign data_masked[15983] = data_i[15983] & sel_one_hot_i[124];
  assign data_masked[15982] = data_i[15982] & sel_one_hot_i[124];
  assign data_masked[15981] = data_i[15981] & sel_one_hot_i[124];
  assign data_masked[15980] = data_i[15980] & sel_one_hot_i[124];
  assign data_masked[15979] = data_i[15979] & sel_one_hot_i[124];
  assign data_masked[15978] = data_i[15978] & sel_one_hot_i[124];
  assign data_masked[15977] = data_i[15977] & sel_one_hot_i[124];
  assign data_masked[15976] = data_i[15976] & sel_one_hot_i[124];
  assign data_masked[15975] = data_i[15975] & sel_one_hot_i[124];
  assign data_masked[15974] = data_i[15974] & sel_one_hot_i[124];
  assign data_masked[15973] = data_i[15973] & sel_one_hot_i[124];
  assign data_masked[15972] = data_i[15972] & sel_one_hot_i[124];
  assign data_masked[15971] = data_i[15971] & sel_one_hot_i[124];
  assign data_masked[15970] = data_i[15970] & sel_one_hot_i[124];
  assign data_masked[15969] = data_i[15969] & sel_one_hot_i[124];
  assign data_masked[15968] = data_i[15968] & sel_one_hot_i[124];
  assign data_masked[15967] = data_i[15967] & sel_one_hot_i[124];
  assign data_masked[15966] = data_i[15966] & sel_one_hot_i[124];
  assign data_masked[15965] = data_i[15965] & sel_one_hot_i[124];
  assign data_masked[15964] = data_i[15964] & sel_one_hot_i[124];
  assign data_masked[15963] = data_i[15963] & sel_one_hot_i[124];
  assign data_masked[15962] = data_i[15962] & sel_one_hot_i[124];
  assign data_masked[15961] = data_i[15961] & sel_one_hot_i[124];
  assign data_masked[15960] = data_i[15960] & sel_one_hot_i[124];
  assign data_masked[15959] = data_i[15959] & sel_one_hot_i[124];
  assign data_masked[15958] = data_i[15958] & sel_one_hot_i[124];
  assign data_masked[15957] = data_i[15957] & sel_one_hot_i[124];
  assign data_masked[15956] = data_i[15956] & sel_one_hot_i[124];
  assign data_masked[15955] = data_i[15955] & sel_one_hot_i[124];
  assign data_masked[15954] = data_i[15954] & sel_one_hot_i[124];
  assign data_masked[15953] = data_i[15953] & sel_one_hot_i[124];
  assign data_masked[15952] = data_i[15952] & sel_one_hot_i[124];
  assign data_masked[15951] = data_i[15951] & sel_one_hot_i[124];
  assign data_masked[15950] = data_i[15950] & sel_one_hot_i[124];
  assign data_masked[15949] = data_i[15949] & sel_one_hot_i[124];
  assign data_masked[15948] = data_i[15948] & sel_one_hot_i[124];
  assign data_masked[15947] = data_i[15947] & sel_one_hot_i[124];
  assign data_masked[15946] = data_i[15946] & sel_one_hot_i[124];
  assign data_masked[15945] = data_i[15945] & sel_one_hot_i[124];
  assign data_masked[15944] = data_i[15944] & sel_one_hot_i[124];
  assign data_masked[15943] = data_i[15943] & sel_one_hot_i[124];
  assign data_masked[15942] = data_i[15942] & sel_one_hot_i[124];
  assign data_masked[15941] = data_i[15941] & sel_one_hot_i[124];
  assign data_masked[15940] = data_i[15940] & sel_one_hot_i[124];
  assign data_masked[15939] = data_i[15939] & sel_one_hot_i[124];
  assign data_masked[15938] = data_i[15938] & sel_one_hot_i[124];
  assign data_masked[15937] = data_i[15937] & sel_one_hot_i[124];
  assign data_masked[15936] = data_i[15936] & sel_one_hot_i[124];
  assign data_masked[15935] = data_i[15935] & sel_one_hot_i[124];
  assign data_masked[15934] = data_i[15934] & sel_one_hot_i[124];
  assign data_masked[15933] = data_i[15933] & sel_one_hot_i[124];
  assign data_masked[15932] = data_i[15932] & sel_one_hot_i[124];
  assign data_masked[15931] = data_i[15931] & sel_one_hot_i[124];
  assign data_masked[15930] = data_i[15930] & sel_one_hot_i[124];
  assign data_masked[15929] = data_i[15929] & sel_one_hot_i[124];
  assign data_masked[15928] = data_i[15928] & sel_one_hot_i[124];
  assign data_masked[15927] = data_i[15927] & sel_one_hot_i[124];
  assign data_masked[15926] = data_i[15926] & sel_one_hot_i[124];
  assign data_masked[15925] = data_i[15925] & sel_one_hot_i[124];
  assign data_masked[15924] = data_i[15924] & sel_one_hot_i[124];
  assign data_masked[15923] = data_i[15923] & sel_one_hot_i[124];
  assign data_masked[15922] = data_i[15922] & sel_one_hot_i[124];
  assign data_masked[15921] = data_i[15921] & sel_one_hot_i[124];
  assign data_masked[15920] = data_i[15920] & sel_one_hot_i[124];
  assign data_masked[15919] = data_i[15919] & sel_one_hot_i[124];
  assign data_masked[15918] = data_i[15918] & sel_one_hot_i[124];
  assign data_masked[15917] = data_i[15917] & sel_one_hot_i[124];
  assign data_masked[15916] = data_i[15916] & sel_one_hot_i[124];
  assign data_masked[15915] = data_i[15915] & sel_one_hot_i[124];
  assign data_masked[15914] = data_i[15914] & sel_one_hot_i[124];
  assign data_masked[15913] = data_i[15913] & sel_one_hot_i[124];
  assign data_masked[15912] = data_i[15912] & sel_one_hot_i[124];
  assign data_masked[15911] = data_i[15911] & sel_one_hot_i[124];
  assign data_masked[15910] = data_i[15910] & sel_one_hot_i[124];
  assign data_masked[15909] = data_i[15909] & sel_one_hot_i[124];
  assign data_masked[15908] = data_i[15908] & sel_one_hot_i[124];
  assign data_masked[15907] = data_i[15907] & sel_one_hot_i[124];
  assign data_masked[15906] = data_i[15906] & sel_one_hot_i[124];
  assign data_masked[15905] = data_i[15905] & sel_one_hot_i[124];
  assign data_masked[15904] = data_i[15904] & sel_one_hot_i[124];
  assign data_masked[15903] = data_i[15903] & sel_one_hot_i[124];
  assign data_masked[15902] = data_i[15902] & sel_one_hot_i[124];
  assign data_masked[15901] = data_i[15901] & sel_one_hot_i[124];
  assign data_masked[15900] = data_i[15900] & sel_one_hot_i[124];
  assign data_masked[15899] = data_i[15899] & sel_one_hot_i[124];
  assign data_masked[15898] = data_i[15898] & sel_one_hot_i[124];
  assign data_masked[15897] = data_i[15897] & sel_one_hot_i[124];
  assign data_masked[15896] = data_i[15896] & sel_one_hot_i[124];
  assign data_masked[15895] = data_i[15895] & sel_one_hot_i[124];
  assign data_masked[15894] = data_i[15894] & sel_one_hot_i[124];
  assign data_masked[15893] = data_i[15893] & sel_one_hot_i[124];
  assign data_masked[15892] = data_i[15892] & sel_one_hot_i[124];
  assign data_masked[15891] = data_i[15891] & sel_one_hot_i[124];
  assign data_masked[15890] = data_i[15890] & sel_one_hot_i[124];
  assign data_masked[15889] = data_i[15889] & sel_one_hot_i[124];
  assign data_masked[15888] = data_i[15888] & sel_one_hot_i[124];
  assign data_masked[15887] = data_i[15887] & sel_one_hot_i[124];
  assign data_masked[15886] = data_i[15886] & sel_one_hot_i[124];
  assign data_masked[15885] = data_i[15885] & sel_one_hot_i[124];
  assign data_masked[15884] = data_i[15884] & sel_one_hot_i[124];
  assign data_masked[15883] = data_i[15883] & sel_one_hot_i[124];
  assign data_masked[15882] = data_i[15882] & sel_one_hot_i[124];
  assign data_masked[15881] = data_i[15881] & sel_one_hot_i[124];
  assign data_masked[15880] = data_i[15880] & sel_one_hot_i[124];
  assign data_masked[15879] = data_i[15879] & sel_one_hot_i[124];
  assign data_masked[15878] = data_i[15878] & sel_one_hot_i[124];
  assign data_masked[15877] = data_i[15877] & sel_one_hot_i[124];
  assign data_masked[15876] = data_i[15876] & sel_one_hot_i[124];
  assign data_masked[15875] = data_i[15875] & sel_one_hot_i[124];
  assign data_masked[15874] = data_i[15874] & sel_one_hot_i[124];
  assign data_masked[15873] = data_i[15873] & sel_one_hot_i[124];
  assign data_masked[15872] = data_i[15872] & sel_one_hot_i[124];
  assign data_masked[16127] = data_i[16127] & sel_one_hot_i[125];
  assign data_masked[16126] = data_i[16126] & sel_one_hot_i[125];
  assign data_masked[16125] = data_i[16125] & sel_one_hot_i[125];
  assign data_masked[16124] = data_i[16124] & sel_one_hot_i[125];
  assign data_masked[16123] = data_i[16123] & sel_one_hot_i[125];
  assign data_masked[16122] = data_i[16122] & sel_one_hot_i[125];
  assign data_masked[16121] = data_i[16121] & sel_one_hot_i[125];
  assign data_masked[16120] = data_i[16120] & sel_one_hot_i[125];
  assign data_masked[16119] = data_i[16119] & sel_one_hot_i[125];
  assign data_masked[16118] = data_i[16118] & sel_one_hot_i[125];
  assign data_masked[16117] = data_i[16117] & sel_one_hot_i[125];
  assign data_masked[16116] = data_i[16116] & sel_one_hot_i[125];
  assign data_masked[16115] = data_i[16115] & sel_one_hot_i[125];
  assign data_masked[16114] = data_i[16114] & sel_one_hot_i[125];
  assign data_masked[16113] = data_i[16113] & sel_one_hot_i[125];
  assign data_masked[16112] = data_i[16112] & sel_one_hot_i[125];
  assign data_masked[16111] = data_i[16111] & sel_one_hot_i[125];
  assign data_masked[16110] = data_i[16110] & sel_one_hot_i[125];
  assign data_masked[16109] = data_i[16109] & sel_one_hot_i[125];
  assign data_masked[16108] = data_i[16108] & sel_one_hot_i[125];
  assign data_masked[16107] = data_i[16107] & sel_one_hot_i[125];
  assign data_masked[16106] = data_i[16106] & sel_one_hot_i[125];
  assign data_masked[16105] = data_i[16105] & sel_one_hot_i[125];
  assign data_masked[16104] = data_i[16104] & sel_one_hot_i[125];
  assign data_masked[16103] = data_i[16103] & sel_one_hot_i[125];
  assign data_masked[16102] = data_i[16102] & sel_one_hot_i[125];
  assign data_masked[16101] = data_i[16101] & sel_one_hot_i[125];
  assign data_masked[16100] = data_i[16100] & sel_one_hot_i[125];
  assign data_masked[16099] = data_i[16099] & sel_one_hot_i[125];
  assign data_masked[16098] = data_i[16098] & sel_one_hot_i[125];
  assign data_masked[16097] = data_i[16097] & sel_one_hot_i[125];
  assign data_masked[16096] = data_i[16096] & sel_one_hot_i[125];
  assign data_masked[16095] = data_i[16095] & sel_one_hot_i[125];
  assign data_masked[16094] = data_i[16094] & sel_one_hot_i[125];
  assign data_masked[16093] = data_i[16093] & sel_one_hot_i[125];
  assign data_masked[16092] = data_i[16092] & sel_one_hot_i[125];
  assign data_masked[16091] = data_i[16091] & sel_one_hot_i[125];
  assign data_masked[16090] = data_i[16090] & sel_one_hot_i[125];
  assign data_masked[16089] = data_i[16089] & sel_one_hot_i[125];
  assign data_masked[16088] = data_i[16088] & sel_one_hot_i[125];
  assign data_masked[16087] = data_i[16087] & sel_one_hot_i[125];
  assign data_masked[16086] = data_i[16086] & sel_one_hot_i[125];
  assign data_masked[16085] = data_i[16085] & sel_one_hot_i[125];
  assign data_masked[16084] = data_i[16084] & sel_one_hot_i[125];
  assign data_masked[16083] = data_i[16083] & sel_one_hot_i[125];
  assign data_masked[16082] = data_i[16082] & sel_one_hot_i[125];
  assign data_masked[16081] = data_i[16081] & sel_one_hot_i[125];
  assign data_masked[16080] = data_i[16080] & sel_one_hot_i[125];
  assign data_masked[16079] = data_i[16079] & sel_one_hot_i[125];
  assign data_masked[16078] = data_i[16078] & sel_one_hot_i[125];
  assign data_masked[16077] = data_i[16077] & sel_one_hot_i[125];
  assign data_masked[16076] = data_i[16076] & sel_one_hot_i[125];
  assign data_masked[16075] = data_i[16075] & sel_one_hot_i[125];
  assign data_masked[16074] = data_i[16074] & sel_one_hot_i[125];
  assign data_masked[16073] = data_i[16073] & sel_one_hot_i[125];
  assign data_masked[16072] = data_i[16072] & sel_one_hot_i[125];
  assign data_masked[16071] = data_i[16071] & sel_one_hot_i[125];
  assign data_masked[16070] = data_i[16070] & sel_one_hot_i[125];
  assign data_masked[16069] = data_i[16069] & sel_one_hot_i[125];
  assign data_masked[16068] = data_i[16068] & sel_one_hot_i[125];
  assign data_masked[16067] = data_i[16067] & sel_one_hot_i[125];
  assign data_masked[16066] = data_i[16066] & sel_one_hot_i[125];
  assign data_masked[16065] = data_i[16065] & sel_one_hot_i[125];
  assign data_masked[16064] = data_i[16064] & sel_one_hot_i[125];
  assign data_masked[16063] = data_i[16063] & sel_one_hot_i[125];
  assign data_masked[16062] = data_i[16062] & sel_one_hot_i[125];
  assign data_masked[16061] = data_i[16061] & sel_one_hot_i[125];
  assign data_masked[16060] = data_i[16060] & sel_one_hot_i[125];
  assign data_masked[16059] = data_i[16059] & sel_one_hot_i[125];
  assign data_masked[16058] = data_i[16058] & sel_one_hot_i[125];
  assign data_masked[16057] = data_i[16057] & sel_one_hot_i[125];
  assign data_masked[16056] = data_i[16056] & sel_one_hot_i[125];
  assign data_masked[16055] = data_i[16055] & sel_one_hot_i[125];
  assign data_masked[16054] = data_i[16054] & sel_one_hot_i[125];
  assign data_masked[16053] = data_i[16053] & sel_one_hot_i[125];
  assign data_masked[16052] = data_i[16052] & sel_one_hot_i[125];
  assign data_masked[16051] = data_i[16051] & sel_one_hot_i[125];
  assign data_masked[16050] = data_i[16050] & sel_one_hot_i[125];
  assign data_masked[16049] = data_i[16049] & sel_one_hot_i[125];
  assign data_masked[16048] = data_i[16048] & sel_one_hot_i[125];
  assign data_masked[16047] = data_i[16047] & sel_one_hot_i[125];
  assign data_masked[16046] = data_i[16046] & sel_one_hot_i[125];
  assign data_masked[16045] = data_i[16045] & sel_one_hot_i[125];
  assign data_masked[16044] = data_i[16044] & sel_one_hot_i[125];
  assign data_masked[16043] = data_i[16043] & sel_one_hot_i[125];
  assign data_masked[16042] = data_i[16042] & sel_one_hot_i[125];
  assign data_masked[16041] = data_i[16041] & sel_one_hot_i[125];
  assign data_masked[16040] = data_i[16040] & sel_one_hot_i[125];
  assign data_masked[16039] = data_i[16039] & sel_one_hot_i[125];
  assign data_masked[16038] = data_i[16038] & sel_one_hot_i[125];
  assign data_masked[16037] = data_i[16037] & sel_one_hot_i[125];
  assign data_masked[16036] = data_i[16036] & sel_one_hot_i[125];
  assign data_masked[16035] = data_i[16035] & sel_one_hot_i[125];
  assign data_masked[16034] = data_i[16034] & sel_one_hot_i[125];
  assign data_masked[16033] = data_i[16033] & sel_one_hot_i[125];
  assign data_masked[16032] = data_i[16032] & sel_one_hot_i[125];
  assign data_masked[16031] = data_i[16031] & sel_one_hot_i[125];
  assign data_masked[16030] = data_i[16030] & sel_one_hot_i[125];
  assign data_masked[16029] = data_i[16029] & sel_one_hot_i[125];
  assign data_masked[16028] = data_i[16028] & sel_one_hot_i[125];
  assign data_masked[16027] = data_i[16027] & sel_one_hot_i[125];
  assign data_masked[16026] = data_i[16026] & sel_one_hot_i[125];
  assign data_masked[16025] = data_i[16025] & sel_one_hot_i[125];
  assign data_masked[16024] = data_i[16024] & sel_one_hot_i[125];
  assign data_masked[16023] = data_i[16023] & sel_one_hot_i[125];
  assign data_masked[16022] = data_i[16022] & sel_one_hot_i[125];
  assign data_masked[16021] = data_i[16021] & sel_one_hot_i[125];
  assign data_masked[16020] = data_i[16020] & sel_one_hot_i[125];
  assign data_masked[16019] = data_i[16019] & sel_one_hot_i[125];
  assign data_masked[16018] = data_i[16018] & sel_one_hot_i[125];
  assign data_masked[16017] = data_i[16017] & sel_one_hot_i[125];
  assign data_masked[16016] = data_i[16016] & sel_one_hot_i[125];
  assign data_masked[16015] = data_i[16015] & sel_one_hot_i[125];
  assign data_masked[16014] = data_i[16014] & sel_one_hot_i[125];
  assign data_masked[16013] = data_i[16013] & sel_one_hot_i[125];
  assign data_masked[16012] = data_i[16012] & sel_one_hot_i[125];
  assign data_masked[16011] = data_i[16011] & sel_one_hot_i[125];
  assign data_masked[16010] = data_i[16010] & sel_one_hot_i[125];
  assign data_masked[16009] = data_i[16009] & sel_one_hot_i[125];
  assign data_masked[16008] = data_i[16008] & sel_one_hot_i[125];
  assign data_masked[16007] = data_i[16007] & sel_one_hot_i[125];
  assign data_masked[16006] = data_i[16006] & sel_one_hot_i[125];
  assign data_masked[16005] = data_i[16005] & sel_one_hot_i[125];
  assign data_masked[16004] = data_i[16004] & sel_one_hot_i[125];
  assign data_masked[16003] = data_i[16003] & sel_one_hot_i[125];
  assign data_masked[16002] = data_i[16002] & sel_one_hot_i[125];
  assign data_masked[16001] = data_i[16001] & sel_one_hot_i[125];
  assign data_masked[16000] = data_i[16000] & sel_one_hot_i[125];
  assign data_masked[16255] = data_i[16255] & sel_one_hot_i[126];
  assign data_masked[16254] = data_i[16254] & sel_one_hot_i[126];
  assign data_masked[16253] = data_i[16253] & sel_one_hot_i[126];
  assign data_masked[16252] = data_i[16252] & sel_one_hot_i[126];
  assign data_masked[16251] = data_i[16251] & sel_one_hot_i[126];
  assign data_masked[16250] = data_i[16250] & sel_one_hot_i[126];
  assign data_masked[16249] = data_i[16249] & sel_one_hot_i[126];
  assign data_masked[16248] = data_i[16248] & sel_one_hot_i[126];
  assign data_masked[16247] = data_i[16247] & sel_one_hot_i[126];
  assign data_masked[16246] = data_i[16246] & sel_one_hot_i[126];
  assign data_masked[16245] = data_i[16245] & sel_one_hot_i[126];
  assign data_masked[16244] = data_i[16244] & sel_one_hot_i[126];
  assign data_masked[16243] = data_i[16243] & sel_one_hot_i[126];
  assign data_masked[16242] = data_i[16242] & sel_one_hot_i[126];
  assign data_masked[16241] = data_i[16241] & sel_one_hot_i[126];
  assign data_masked[16240] = data_i[16240] & sel_one_hot_i[126];
  assign data_masked[16239] = data_i[16239] & sel_one_hot_i[126];
  assign data_masked[16238] = data_i[16238] & sel_one_hot_i[126];
  assign data_masked[16237] = data_i[16237] & sel_one_hot_i[126];
  assign data_masked[16236] = data_i[16236] & sel_one_hot_i[126];
  assign data_masked[16235] = data_i[16235] & sel_one_hot_i[126];
  assign data_masked[16234] = data_i[16234] & sel_one_hot_i[126];
  assign data_masked[16233] = data_i[16233] & sel_one_hot_i[126];
  assign data_masked[16232] = data_i[16232] & sel_one_hot_i[126];
  assign data_masked[16231] = data_i[16231] & sel_one_hot_i[126];
  assign data_masked[16230] = data_i[16230] & sel_one_hot_i[126];
  assign data_masked[16229] = data_i[16229] & sel_one_hot_i[126];
  assign data_masked[16228] = data_i[16228] & sel_one_hot_i[126];
  assign data_masked[16227] = data_i[16227] & sel_one_hot_i[126];
  assign data_masked[16226] = data_i[16226] & sel_one_hot_i[126];
  assign data_masked[16225] = data_i[16225] & sel_one_hot_i[126];
  assign data_masked[16224] = data_i[16224] & sel_one_hot_i[126];
  assign data_masked[16223] = data_i[16223] & sel_one_hot_i[126];
  assign data_masked[16222] = data_i[16222] & sel_one_hot_i[126];
  assign data_masked[16221] = data_i[16221] & sel_one_hot_i[126];
  assign data_masked[16220] = data_i[16220] & sel_one_hot_i[126];
  assign data_masked[16219] = data_i[16219] & sel_one_hot_i[126];
  assign data_masked[16218] = data_i[16218] & sel_one_hot_i[126];
  assign data_masked[16217] = data_i[16217] & sel_one_hot_i[126];
  assign data_masked[16216] = data_i[16216] & sel_one_hot_i[126];
  assign data_masked[16215] = data_i[16215] & sel_one_hot_i[126];
  assign data_masked[16214] = data_i[16214] & sel_one_hot_i[126];
  assign data_masked[16213] = data_i[16213] & sel_one_hot_i[126];
  assign data_masked[16212] = data_i[16212] & sel_one_hot_i[126];
  assign data_masked[16211] = data_i[16211] & sel_one_hot_i[126];
  assign data_masked[16210] = data_i[16210] & sel_one_hot_i[126];
  assign data_masked[16209] = data_i[16209] & sel_one_hot_i[126];
  assign data_masked[16208] = data_i[16208] & sel_one_hot_i[126];
  assign data_masked[16207] = data_i[16207] & sel_one_hot_i[126];
  assign data_masked[16206] = data_i[16206] & sel_one_hot_i[126];
  assign data_masked[16205] = data_i[16205] & sel_one_hot_i[126];
  assign data_masked[16204] = data_i[16204] & sel_one_hot_i[126];
  assign data_masked[16203] = data_i[16203] & sel_one_hot_i[126];
  assign data_masked[16202] = data_i[16202] & sel_one_hot_i[126];
  assign data_masked[16201] = data_i[16201] & sel_one_hot_i[126];
  assign data_masked[16200] = data_i[16200] & sel_one_hot_i[126];
  assign data_masked[16199] = data_i[16199] & sel_one_hot_i[126];
  assign data_masked[16198] = data_i[16198] & sel_one_hot_i[126];
  assign data_masked[16197] = data_i[16197] & sel_one_hot_i[126];
  assign data_masked[16196] = data_i[16196] & sel_one_hot_i[126];
  assign data_masked[16195] = data_i[16195] & sel_one_hot_i[126];
  assign data_masked[16194] = data_i[16194] & sel_one_hot_i[126];
  assign data_masked[16193] = data_i[16193] & sel_one_hot_i[126];
  assign data_masked[16192] = data_i[16192] & sel_one_hot_i[126];
  assign data_masked[16191] = data_i[16191] & sel_one_hot_i[126];
  assign data_masked[16190] = data_i[16190] & sel_one_hot_i[126];
  assign data_masked[16189] = data_i[16189] & sel_one_hot_i[126];
  assign data_masked[16188] = data_i[16188] & sel_one_hot_i[126];
  assign data_masked[16187] = data_i[16187] & sel_one_hot_i[126];
  assign data_masked[16186] = data_i[16186] & sel_one_hot_i[126];
  assign data_masked[16185] = data_i[16185] & sel_one_hot_i[126];
  assign data_masked[16184] = data_i[16184] & sel_one_hot_i[126];
  assign data_masked[16183] = data_i[16183] & sel_one_hot_i[126];
  assign data_masked[16182] = data_i[16182] & sel_one_hot_i[126];
  assign data_masked[16181] = data_i[16181] & sel_one_hot_i[126];
  assign data_masked[16180] = data_i[16180] & sel_one_hot_i[126];
  assign data_masked[16179] = data_i[16179] & sel_one_hot_i[126];
  assign data_masked[16178] = data_i[16178] & sel_one_hot_i[126];
  assign data_masked[16177] = data_i[16177] & sel_one_hot_i[126];
  assign data_masked[16176] = data_i[16176] & sel_one_hot_i[126];
  assign data_masked[16175] = data_i[16175] & sel_one_hot_i[126];
  assign data_masked[16174] = data_i[16174] & sel_one_hot_i[126];
  assign data_masked[16173] = data_i[16173] & sel_one_hot_i[126];
  assign data_masked[16172] = data_i[16172] & sel_one_hot_i[126];
  assign data_masked[16171] = data_i[16171] & sel_one_hot_i[126];
  assign data_masked[16170] = data_i[16170] & sel_one_hot_i[126];
  assign data_masked[16169] = data_i[16169] & sel_one_hot_i[126];
  assign data_masked[16168] = data_i[16168] & sel_one_hot_i[126];
  assign data_masked[16167] = data_i[16167] & sel_one_hot_i[126];
  assign data_masked[16166] = data_i[16166] & sel_one_hot_i[126];
  assign data_masked[16165] = data_i[16165] & sel_one_hot_i[126];
  assign data_masked[16164] = data_i[16164] & sel_one_hot_i[126];
  assign data_masked[16163] = data_i[16163] & sel_one_hot_i[126];
  assign data_masked[16162] = data_i[16162] & sel_one_hot_i[126];
  assign data_masked[16161] = data_i[16161] & sel_one_hot_i[126];
  assign data_masked[16160] = data_i[16160] & sel_one_hot_i[126];
  assign data_masked[16159] = data_i[16159] & sel_one_hot_i[126];
  assign data_masked[16158] = data_i[16158] & sel_one_hot_i[126];
  assign data_masked[16157] = data_i[16157] & sel_one_hot_i[126];
  assign data_masked[16156] = data_i[16156] & sel_one_hot_i[126];
  assign data_masked[16155] = data_i[16155] & sel_one_hot_i[126];
  assign data_masked[16154] = data_i[16154] & sel_one_hot_i[126];
  assign data_masked[16153] = data_i[16153] & sel_one_hot_i[126];
  assign data_masked[16152] = data_i[16152] & sel_one_hot_i[126];
  assign data_masked[16151] = data_i[16151] & sel_one_hot_i[126];
  assign data_masked[16150] = data_i[16150] & sel_one_hot_i[126];
  assign data_masked[16149] = data_i[16149] & sel_one_hot_i[126];
  assign data_masked[16148] = data_i[16148] & sel_one_hot_i[126];
  assign data_masked[16147] = data_i[16147] & sel_one_hot_i[126];
  assign data_masked[16146] = data_i[16146] & sel_one_hot_i[126];
  assign data_masked[16145] = data_i[16145] & sel_one_hot_i[126];
  assign data_masked[16144] = data_i[16144] & sel_one_hot_i[126];
  assign data_masked[16143] = data_i[16143] & sel_one_hot_i[126];
  assign data_masked[16142] = data_i[16142] & sel_one_hot_i[126];
  assign data_masked[16141] = data_i[16141] & sel_one_hot_i[126];
  assign data_masked[16140] = data_i[16140] & sel_one_hot_i[126];
  assign data_masked[16139] = data_i[16139] & sel_one_hot_i[126];
  assign data_masked[16138] = data_i[16138] & sel_one_hot_i[126];
  assign data_masked[16137] = data_i[16137] & sel_one_hot_i[126];
  assign data_masked[16136] = data_i[16136] & sel_one_hot_i[126];
  assign data_masked[16135] = data_i[16135] & sel_one_hot_i[126];
  assign data_masked[16134] = data_i[16134] & sel_one_hot_i[126];
  assign data_masked[16133] = data_i[16133] & sel_one_hot_i[126];
  assign data_masked[16132] = data_i[16132] & sel_one_hot_i[126];
  assign data_masked[16131] = data_i[16131] & sel_one_hot_i[126];
  assign data_masked[16130] = data_i[16130] & sel_one_hot_i[126];
  assign data_masked[16129] = data_i[16129] & sel_one_hot_i[126];
  assign data_masked[16128] = data_i[16128] & sel_one_hot_i[126];
  assign data_masked[16383] = data_i[16383] & sel_one_hot_i[127];
  assign data_masked[16382] = data_i[16382] & sel_one_hot_i[127];
  assign data_masked[16381] = data_i[16381] & sel_one_hot_i[127];
  assign data_masked[16380] = data_i[16380] & sel_one_hot_i[127];
  assign data_masked[16379] = data_i[16379] & sel_one_hot_i[127];
  assign data_masked[16378] = data_i[16378] & sel_one_hot_i[127];
  assign data_masked[16377] = data_i[16377] & sel_one_hot_i[127];
  assign data_masked[16376] = data_i[16376] & sel_one_hot_i[127];
  assign data_masked[16375] = data_i[16375] & sel_one_hot_i[127];
  assign data_masked[16374] = data_i[16374] & sel_one_hot_i[127];
  assign data_masked[16373] = data_i[16373] & sel_one_hot_i[127];
  assign data_masked[16372] = data_i[16372] & sel_one_hot_i[127];
  assign data_masked[16371] = data_i[16371] & sel_one_hot_i[127];
  assign data_masked[16370] = data_i[16370] & sel_one_hot_i[127];
  assign data_masked[16369] = data_i[16369] & sel_one_hot_i[127];
  assign data_masked[16368] = data_i[16368] & sel_one_hot_i[127];
  assign data_masked[16367] = data_i[16367] & sel_one_hot_i[127];
  assign data_masked[16366] = data_i[16366] & sel_one_hot_i[127];
  assign data_masked[16365] = data_i[16365] & sel_one_hot_i[127];
  assign data_masked[16364] = data_i[16364] & sel_one_hot_i[127];
  assign data_masked[16363] = data_i[16363] & sel_one_hot_i[127];
  assign data_masked[16362] = data_i[16362] & sel_one_hot_i[127];
  assign data_masked[16361] = data_i[16361] & sel_one_hot_i[127];
  assign data_masked[16360] = data_i[16360] & sel_one_hot_i[127];
  assign data_masked[16359] = data_i[16359] & sel_one_hot_i[127];
  assign data_masked[16358] = data_i[16358] & sel_one_hot_i[127];
  assign data_masked[16357] = data_i[16357] & sel_one_hot_i[127];
  assign data_masked[16356] = data_i[16356] & sel_one_hot_i[127];
  assign data_masked[16355] = data_i[16355] & sel_one_hot_i[127];
  assign data_masked[16354] = data_i[16354] & sel_one_hot_i[127];
  assign data_masked[16353] = data_i[16353] & sel_one_hot_i[127];
  assign data_masked[16352] = data_i[16352] & sel_one_hot_i[127];
  assign data_masked[16351] = data_i[16351] & sel_one_hot_i[127];
  assign data_masked[16350] = data_i[16350] & sel_one_hot_i[127];
  assign data_masked[16349] = data_i[16349] & sel_one_hot_i[127];
  assign data_masked[16348] = data_i[16348] & sel_one_hot_i[127];
  assign data_masked[16347] = data_i[16347] & sel_one_hot_i[127];
  assign data_masked[16346] = data_i[16346] & sel_one_hot_i[127];
  assign data_masked[16345] = data_i[16345] & sel_one_hot_i[127];
  assign data_masked[16344] = data_i[16344] & sel_one_hot_i[127];
  assign data_masked[16343] = data_i[16343] & sel_one_hot_i[127];
  assign data_masked[16342] = data_i[16342] & sel_one_hot_i[127];
  assign data_masked[16341] = data_i[16341] & sel_one_hot_i[127];
  assign data_masked[16340] = data_i[16340] & sel_one_hot_i[127];
  assign data_masked[16339] = data_i[16339] & sel_one_hot_i[127];
  assign data_masked[16338] = data_i[16338] & sel_one_hot_i[127];
  assign data_masked[16337] = data_i[16337] & sel_one_hot_i[127];
  assign data_masked[16336] = data_i[16336] & sel_one_hot_i[127];
  assign data_masked[16335] = data_i[16335] & sel_one_hot_i[127];
  assign data_masked[16334] = data_i[16334] & sel_one_hot_i[127];
  assign data_masked[16333] = data_i[16333] & sel_one_hot_i[127];
  assign data_masked[16332] = data_i[16332] & sel_one_hot_i[127];
  assign data_masked[16331] = data_i[16331] & sel_one_hot_i[127];
  assign data_masked[16330] = data_i[16330] & sel_one_hot_i[127];
  assign data_masked[16329] = data_i[16329] & sel_one_hot_i[127];
  assign data_masked[16328] = data_i[16328] & sel_one_hot_i[127];
  assign data_masked[16327] = data_i[16327] & sel_one_hot_i[127];
  assign data_masked[16326] = data_i[16326] & sel_one_hot_i[127];
  assign data_masked[16325] = data_i[16325] & sel_one_hot_i[127];
  assign data_masked[16324] = data_i[16324] & sel_one_hot_i[127];
  assign data_masked[16323] = data_i[16323] & sel_one_hot_i[127];
  assign data_masked[16322] = data_i[16322] & sel_one_hot_i[127];
  assign data_masked[16321] = data_i[16321] & sel_one_hot_i[127];
  assign data_masked[16320] = data_i[16320] & sel_one_hot_i[127];
  assign data_masked[16319] = data_i[16319] & sel_one_hot_i[127];
  assign data_masked[16318] = data_i[16318] & sel_one_hot_i[127];
  assign data_masked[16317] = data_i[16317] & sel_one_hot_i[127];
  assign data_masked[16316] = data_i[16316] & sel_one_hot_i[127];
  assign data_masked[16315] = data_i[16315] & sel_one_hot_i[127];
  assign data_masked[16314] = data_i[16314] & sel_one_hot_i[127];
  assign data_masked[16313] = data_i[16313] & sel_one_hot_i[127];
  assign data_masked[16312] = data_i[16312] & sel_one_hot_i[127];
  assign data_masked[16311] = data_i[16311] & sel_one_hot_i[127];
  assign data_masked[16310] = data_i[16310] & sel_one_hot_i[127];
  assign data_masked[16309] = data_i[16309] & sel_one_hot_i[127];
  assign data_masked[16308] = data_i[16308] & sel_one_hot_i[127];
  assign data_masked[16307] = data_i[16307] & sel_one_hot_i[127];
  assign data_masked[16306] = data_i[16306] & sel_one_hot_i[127];
  assign data_masked[16305] = data_i[16305] & sel_one_hot_i[127];
  assign data_masked[16304] = data_i[16304] & sel_one_hot_i[127];
  assign data_masked[16303] = data_i[16303] & sel_one_hot_i[127];
  assign data_masked[16302] = data_i[16302] & sel_one_hot_i[127];
  assign data_masked[16301] = data_i[16301] & sel_one_hot_i[127];
  assign data_masked[16300] = data_i[16300] & sel_one_hot_i[127];
  assign data_masked[16299] = data_i[16299] & sel_one_hot_i[127];
  assign data_masked[16298] = data_i[16298] & sel_one_hot_i[127];
  assign data_masked[16297] = data_i[16297] & sel_one_hot_i[127];
  assign data_masked[16296] = data_i[16296] & sel_one_hot_i[127];
  assign data_masked[16295] = data_i[16295] & sel_one_hot_i[127];
  assign data_masked[16294] = data_i[16294] & sel_one_hot_i[127];
  assign data_masked[16293] = data_i[16293] & sel_one_hot_i[127];
  assign data_masked[16292] = data_i[16292] & sel_one_hot_i[127];
  assign data_masked[16291] = data_i[16291] & sel_one_hot_i[127];
  assign data_masked[16290] = data_i[16290] & sel_one_hot_i[127];
  assign data_masked[16289] = data_i[16289] & sel_one_hot_i[127];
  assign data_masked[16288] = data_i[16288] & sel_one_hot_i[127];
  assign data_masked[16287] = data_i[16287] & sel_one_hot_i[127];
  assign data_masked[16286] = data_i[16286] & sel_one_hot_i[127];
  assign data_masked[16285] = data_i[16285] & sel_one_hot_i[127];
  assign data_masked[16284] = data_i[16284] & sel_one_hot_i[127];
  assign data_masked[16283] = data_i[16283] & sel_one_hot_i[127];
  assign data_masked[16282] = data_i[16282] & sel_one_hot_i[127];
  assign data_masked[16281] = data_i[16281] & sel_one_hot_i[127];
  assign data_masked[16280] = data_i[16280] & sel_one_hot_i[127];
  assign data_masked[16279] = data_i[16279] & sel_one_hot_i[127];
  assign data_masked[16278] = data_i[16278] & sel_one_hot_i[127];
  assign data_masked[16277] = data_i[16277] & sel_one_hot_i[127];
  assign data_masked[16276] = data_i[16276] & sel_one_hot_i[127];
  assign data_masked[16275] = data_i[16275] & sel_one_hot_i[127];
  assign data_masked[16274] = data_i[16274] & sel_one_hot_i[127];
  assign data_masked[16273] = data_i[16273] & sel_one_hot_i[127];
  assign data_masked[16272] = data_i[16272] & sel_one_hot_i[127];
  assign data_masked[16271] = data_i[16271] & sel_one_hot_i[127];
  assign data_masked[16270] = data_i[16270] & sel_one_hot_i[127];
  assign data_masked[16269] = data_i[16269] & sel_one_hot_i[127];
  assign data_masked[16268] = data_i[16268] & sel_one_hot_i[127];
  assign data_masked[16267] = data_i[16267] & sel_one_hot_i[127];
  assign data_masked[16266] = data_i[16266] & sel_one_hot_i[127];
  assign data_masked[16265] = data_i[16265] & sel_one_hot_i[127];
  assign data_masked[16264] = data_i[16264] & sel_one_hot_i[127];
  assign data_masked[16263] = data_i[16263] & sel_one_hot_i[127];
  assign data_masked[16262] = data_i[16262] & sel_one_hot_i[127];
  assign data_masked[16261] = data_i[16261] & sel_one_hot_i[127];
  assign data_masked[16260] = data_i[16260] & sel_one_hot_i[127];
  assign data_masked[16259] = data_i[16259] & sel_one_hot_i[127];
  assign data_masked[16258] = data_i[16258] & sel_one_hot_i[127];
  assign data_masked[16257] = data_i[16257] & sel_one_hot_i[127];
  assign data_masked[16256] = data_i[16256] & sel_one_hot_i[127];
  assign data_o[0] = N125 | data_masked[0];
  assign N125 = N124 | data_masked[128];
  assign N124 = N123 | data_masked[256];
  assign N123 = N122 | data_masked[384];
  assign N122 = N121 | data_masked[512];
  assign N121 = N120 | data_masked[640];
  assign N120 = N119 | data_masked[768];
  assign N119 = N118 | data_masked[896];
  assign N118 = N117 | data_masked[1024];
  assign N117 = N116 | data_masked[1152];
  assign N116 = N115 | data_masked[1280];
  assign N115 = N114 | data_masked[1408];
  assign N114 = N113 | data_masked[1536];
  assign N113 = N112 | data_masked[1664];
  assign N112 = N111 | data_masked[1792];
  assign N111 = N110 | data_masked[1920];
  assign N110 = N109 | data_masked[2048];
  assign N109 = N108 | data_masked[2176];
  assign N108 = N107 | data_masked[2304];
  assign N107 = N106 | data_masked[2432];
  assign N106 = N105 | data_masked[2560];
  assign N105 = N104 | data_masked[2688];
  assign N104 = N103 | data_masked[2816];
  assign N103 = N102 | data_masked[2944];
  assign N102 = N101 | data_masked[3072];
  assign N101 = N100 | data_masked[3200];
  assign N100 = N99 | data_masked[3328];
  assign N99 = N98 | data_masked[3456];
  assign N98 = N97 | data_masked[3584];
  assign N97 = N96 | data_masked[3712];
  assign N96 = N95 | data_masked[3840];
  assign N95 = N94 | data_masked[3968];
  assign N94 = N93 | data_masked[4096];
  assign N93 = N92 | data_masked[4224];
  assign N92 = N91 | data_masked[4352];
  assign N91 = N90 | data_masked[4480];
  assign N90 = N89 | data_masked[4608];
  assign N89 = N88 | data_masked[4736];
  assign N88 = N87 | data_masked[4864];
  assign N87 = N86 | data_masked[4992];
  assign N86 = N85 | data_masked[5120];
  assign N85 = N84 | data_masked[5248];
  assign N84 = N83 | data_masked[5376];
  assign N83 = N82 | data_masked[5504];
  assign N82 = N81 | data_masked[5632];
  assign N81 = N80 | data_masked[5760];
  assign N80 = N79 | data_masked[5888];
  assign N79 = N78 | data_masked[6016];
  assign N78 = N77 | data_masked[6144];
  assign N77 = N76 | data_masked[6272];
  assign N76 = N75 | data_masked[6400];
  assign N75 = N74 | data_masked[6528];
  assign N74 = N73 | data_masked[6656];
  assign N73 = N72 | data_masked[6784];
  assign N72 = N71 | data_masked[6912];
  assign N71 = N70 | data_masked[7040];
  assign N70 = N69 | data_masked[7168];
  assign N69 = N68 | data_masked[7296];
  assign N68 = N67 | data_masked[7424];
  assign N67 = N66 | data_masked[7552];
  assign N66 = N65 | data_masked[7680];
  assign N65 = N64 | data_masked[7808];
  assign N64 = N63 | data_masked[7936];
  assign N63 = N62 | data_masked[8064];
  assign N62 = N61 | data_masked[8192];
  assign N61 = N60 | data_masked[8320];
  assign N60 = N59 | data_masked[8448];
  assign N59 = N58 | data_masked[8576];
  assign N58 = N57 | data_masked[8704];
  assign N57 = N56 | data_masked[8832];
  assign N56 = N55 | data_masked[8960];
  assign N55 = N54 | data_masked[9088];
  assign N54 = N53 | data_masked[9216];
  assign N53 = N52 | data_masked[9344];
  assign N52 = N51 | data_masked[9472];
  assign N51 = N50 | data_masked[9600];
  assign N50 = N49 | data_masked[9728];
  assign N49 = N48 | data_masked[9856];
  assign N48 = N47 | data_masked[9984];
  assign N47 = N46 | data_masked[10112];
  assign N46 = N45 | data_masked[10240];
  assign N45 = N44 | data_masked[10368];
  assign N44 = N43 | data_masked[10496];
  assign N43 = N42 | data_masked[10624];
  assign N42 = N41 | data_masked[10752];
  assign N41 = N40 | data_masked[10880];
  assign N40 = N39 | data_masked[11008];
  assign N39 = N38 | data_masked[11136];
  assign N38 = N37 | data_masked[11264];
  assign N37 = N36 | data_masked[11392];
  assign N36 = N35 | data_masked[11520];
  assign N35 = N34 | data_masked[11648];
  assign N34 = N33 | data_masked[11776];
  assign N33 = N32 | data_masked[11904];
  assign N32 = N31 | data_masked[12032];
  assign N31 = N30 | data_masked[12160];
  assign N30 = N29 | data_masked[12288];
  assign N29 = N28 | data_masked[12416];
  assign N28 = N27 | data_masked[12544];
  assign N27 = N26 | data_masked[12672];
  assign N26 = N25 | data_masked[12800];
  assign N25 = N24 | data_masked[12928];
  assign N24 = N23 | data_masked[13056];
  assign N23 = N22 | data_masked[13184];
  assign N22 = N21 | data_masked[13312];
  assign N21 = N20 | data_masked[13440];
  assign N20 = N19 | data_masked[13568];
  assign N19 = N18 | data_masked[13696];
  assign N18 = N17 | data_masked[13824];
  assign N17 = N16 | data_masked[13952];
  assign N16 = N15 | data_masked[14080];
  assign N15 = N14 | data_masked[14208];
  assign N14 = N13 | data_masked[14336];
  assign N13 = N12 | data_masked[14464];
  assign N12 = N11 | data_masked[14592];
  assign N11 = N10 | data_masked[14720];
  assign N10 = N9 | data_masked[14848];
  assign N9 = N8 | data_masked[14976];
  assign N8 = N7 | data_masked[15104];
  assign N7 = N6 | data_masked[15232];
  assign N6 = N5 | data_masked[15360];
  assign N5 = N4 | data_masked[15488];
  assign N4 = N3 | data_masked[15616];
  assign N3 = N2 | data_masked[15744];
  assign N2 = N1 | data_masked[15872];
  assign N1 = N0 | data_masked[16000];
  assign N0 = data_masked[16256] | data_masked[16128];
  assign data_o[1] = N251 | data_masked[1];
  assign N251 = N250 | data_masked[129];
  assign N250 = N249 | data_masked[257];
  assign N249 = N248 | data_masked[385];
  assign N248 = N247 | data_masked[513];
  assign N247 = N246 | data_masked[641];
  assign N246 = N245 | data_masked[769];
  assign N245 = N244 | data_masked[897];
  assign N244 = N243 | data_masked[1025];
  assign N243 = N242 | data_masked[1153];
  assign N242 = N241 | data_masked[1281];
  assign N241 = N240 | data_masked[1409];
  assign N240 = N239 | data_masked[1537];
  assign N239 = N238 | data_masked[1665];
  assign N238 = N237 | data_masked[1793];
  assign N237 = N236 | data_masked[1921];
  assign N236 = N235 | data_masked[2049];
  assign N235 = N234 | data_masked[2177];
  assign N234 = N233 | data_masked[2305];
  assign N233 = N232 | data_masked[2433];
  assign N232 = N231 | data_masked[2561];
  assign N231 = N230 | data_masked[2689];
  assign N230 = N229 | data_masked[2817];
  assign N229 = N228 | data_masked[2945];
  assign N228 = N227 | data_masked[3073];
  assign N227 = N226 | data_masked[3201];
  assign N226 = N225 | data_masked[3329];
  assign N225 = N224 | data_masked[3457];
  assign N224 = N223 | data_masked[3585];
  assign N223 = N222 | data_masked[3713];
  assign N222 = N221 | data_masked[3841];
  assign N221 = N220 | data_masked[3969];
  assign N220 = N219 | data_masked[4097];
  assign N219 = N218 | data_masked[4225];
  assign N218 = N217 | data_masked[4353];
  assign N217 = N216 | data_masked[4481];
  assign N216 = N215 | data_masked[4609];
  assign N215 = N214 | data_masked[4737];
  assign N214 = N213 | data_masked[4865];
  assign N213 = N212 | data_masked[4993];
  assign N212 = N211 | data_masked[5121];
  assign N211 = N210 | data_masked[5249];
  assign N210 = N209 | data_masked[5377];
  assign N209 = N208 | data_masked[5505];
  assign N208 = N207 | data_masked[5633];
  assign N207 = N206 | data_masked[5761];
  assign N206 = N205 | data_masked[5889];
  assign N205 = N204 | data_masked[6017];
  assign N204 = N203 | data_masked[6145];
  assign N203 = N202 | data_masked[6273];
  assign N202 = N201 | data_masked[6401];
  assign N201 = N200 | data_masked[6529];
  assign N200 = N199 | data_masked[6657];
  assign N199 = N198 | data_masked[6785];
  assign N198 = N197 | data_masked[6913];
  assign N197 = N196 | data_masked[7041];
  assign N196 = N195 | data_masked[7169];
  assign N195 = N194 | data_masked[7297];
  assign N194 = N193 | data_masked[7425];
  assign N193 = N192 | data_masked[7553];
  assign N192 = N191 | data_masked[7681];
  assign N191 = N190 | data_masked[7809];
  assign N190 = N189 | data_masked[7937];
  assign N189 = N188 | data_masked[8065];
  assign N188 = N187 | data_masked[8193];
  assign N187 = N186 | data_masked[8321];
  assign N186 = N185 | data_masked[8449];
  assign N185 = N184 | data_masked[8577];
  assign N184 = N183 | data_masked[8705];
  assign N183 = N182 | data_masked[8833];
  assign N182 = N181 | data_masked[8961];
  assign N181 = N180 | data_masked[9089];
  assign N180 = N179 | data_masked[9217];
  assign N179 = N178 | data_masked[9345];
  assign N178 = N177 | data_masked[9473];
  assign N177 = N176 | data_masked[9601];
  assign N176 = N175 | data_masked[9729];
  assign N175 = N174 | data_masked[9857];
  assign N174 = N173 | data_masked[9985];
  assign N173 = N172 | data_masked[10113];
  assign N172 = N171 | data_masked[10241];
  assign N171 = N170 | data_masked[10369];
  assign N170 = N169 | data_masked[10497];
  assign N169 = N168 | data_masked[10625];
  assign N168 = N167 | data_masked[10753];
  assign N167 = N166 | data_masked[10881];
  assign N166 = N165 | data_masked[11009];
  assign N165 = N164 | data_masked[11137];
  assign N164 = N163 | data_masked[11265];
  assign N163 = N162 | data_masked[11393];
  assign N162 = N161 | data_masked[11521];
  assign N161 = N160 | data_masked[11649];
  assign N160 = N159 | data_masked[11777];
  assign N159 = N158 | data_masked[11905];
  assign N158 = N157 | data_masked[12033];
  assign N157 = N156 | data_masked[12161];
  assign N156 = N155 | data_masked[12289];
  assign N155 = N154 | data_masked[12417];
  assign N154 = N153 | data_masked[12545];
  assign N153 = N152 | data_masked[12673];
  assign N152 = N151 | data_masked[12801];
  assign N151 = N150 | data_masked[12929];
  assign N150 = N149 | data_masked[13057];
  assign N149 = N148 | data_masked[13185];
  assign N148 = N147 | data_masked[13313];
  assign N147 = N146 | data_masked[13441];
  assign N146 = N145 | data_masked[13569];
  assign N145 = N144 | data_masked[13697];
  assign N144 = N143 | data_masked[13825];
  assign N143 = N142 | data_masked[13953];
  assign N142 = N141 | data_masked[14081];
  assign N141 = N140 | data_masked[14209];
  assign N140 = N139 | data_masked[14337];
  assign N139 = N138 | data_masked[14465];
  assign N138 = N137 | data_masked[14593];
  assign N137 = N136 | data_masked[14721];
  assign N136 = N135 | data_masked[14849];
  assign N135 = N134 | data_masked[14977];
  assign N134 = N133 | data_masked[15105];
  assign N133 = N132 | data_masked[15233];
  assign N132 = N131 | data_masked[15361];
  assign N131 = N130 | data_masked[15489];
  assign N130 = N129 | data_masked[15617];
  assign N129 = N128 | data_masked[15745];
  assign N128 = N127 | data_masked[15873];
  assign N127 = N126 | data_masked[16001];
  assign N126 = data_masked[16257] | data_masked[16129];
  assign data_o[2] = N377 | data_masked[2];
  assign N377 = N376 | data_masked[130];
  assign N376 = N375 | data_masked[258];
  assign N375 = N374 | data_masked[386];
  assign N374 = N373 | data_masked[514];
  assign N373 = N372 | data_masked[642];
  assign N372 = N371 | data_masked[770];
  assign N371 = N370 | data_masked[898];
  assign N370 = N369 | data_masked[1026];
  assign N369 = N368 | data_masked[1154];
  assign N368 = N367 | data_masked[1282];
  assign N367 = N366 | data_masked[1410];
  assign N366 = N365 | data_masked[1538];
  assign N365 = N364 | data_masked[1666];
  assign N364 = N363 | data_masked[1794];
  assign N363 = N362 | data_masked[1922];
  assign N362 = N361 | data_masked[2050];
  assign N361 = N360 | data_masked[2178];
  assign N360 = N359 | data_masked[2306];
  assign N359 = N358 | data_masked[2434];
  assign N358 = N357 | data_masked[2562];
  assign N357 = N356 | data_masked[2690];
  assign N356 = N355 | data_masked[2818];
  assign N355 = N354 | data_masked[2946];
  assign N354 = N353 | data_masked[3074];
  assign N353 = N352 | data_masked[3202];
  assign N352 = N351 | data_masked[3330];
  assign N351 = N350 | data_masked[3458];
  assign N350 = N349 | data_masked[3586];
  assign N349 = N348 | data_masked[3714];
  assign N348 = N347 | data_masked[3842];
  assign N347 = N346 | data_masked[3970];
  assign N346 = N345 | data_masked[4098];
  assign N345 = N344 | data_masked[4226];
  assign N344 = N343 | data_masked[4354];
  assign N343 = N342 | data_masked[4482];
  assign N342 = N341 | data_masked[4610];
  assign N341 = N340 | data_masked[4738];
  assign N340 = N339 | data_masked[4866];
  assign N339 = N338 | data_masked[4994];
  assign N338 = N337 | data_masked[5122];
  assign N337 = N336 | data_masked[5250];
  assign N336 = N335 | data_masked[5378];
  assign N335 = N334 | data_masked[5506];
  assign N334 = N333 | data_masked[5634];
  assign N333 = N332 | data_masked[5762];
  assign N332 = N331 | data_masked[5890];
  assign N331 = N330 | data_masked[6018];
  assign N330 = N329 | data_masked[6146];
  assign N329 = N328 | data_masked[6274];
  assign N328 = N327 | data_masked[6402];
  assign N327 = N326 | data_masked[6530];
  assign N326 = N325 | data_masked[6658];
  assign N325 = N324 | data_masked[6786];
  assign N324 = N323 | data_masked[6914];
  assign N323 = N322 | data_masked[7042];
  assign N322 = N321 | data_masked[7170];
  assign N321 = N320 | data_masked[7298];
  assign N320 = N319 | data_masked[7426];
  assign N319 = N318 | data_masked[7554];
  assign N318 = N317 | data_masked[7682];
  assign N317 = N316 | data_masked[7810];
  assign N316 = N315 | data_masked[7938];
  assign N315 = N314 | data_masked[8066];
  assign N314 = N313 | data_masked[8194];
  assign N313 = N312 | data_masked[8322];
  assign N312 = N311 | data_masked[8450];
  assign N311 = N310 | data_masked[8578];
  assign N310 = N309 | data_masked[8706];
  assign N309 = N308 | data_masked[8834];
  assign N308 = N307 | data_masked[8962];
  assign N307 = N306 | data_masked[9090];
  assign N306 = N305 | data_masked[9218];
  assign N305 = N304 | data_masked[9346];
  assign N304 = N303 | data_masked[9474];
  assign N303 = N302 | data_masked[9602];
  assign N302 = N301 | data_masked[9730];
  assign N301 = N300 | data_masked[9858];
  assign N300 = N299 | data_masked[9986];
  assign N299 = N298 | data_masked[10114];
  assign N298 = N297 | data_masked[10242];
  assign N297 = N296 | data_masked[10370];
  assign N296 = N295 | data_masked[10498];
  assign N295 = N294 | data_masked[10626];
  assign N294 = N293 | data_masked[10754];
  assign N293 = N292 | data_masked[10882];
  assign N292 = N291 | data_masked[11010];
  assign N291 = N290 | data_masked[11138];
  assign N290 = N289 | data_masked[11266];
  assign N289 = N288 | data_masked[11394];
  assign N288 = N287 | data_masked[11522];
  assign N287 = N286 | data_masked[11650];
  assign N286 = N285 | data_masked[11778];
  assign N285 = N284 | data_masked[11906];
  assign N284 = N283 | data_masked[12034];
  assign N283 = N282 | data_masked[12162];
  assign N282 = N281 | data_masked[12290];
  assign N281 = N280 | data_masked[12418];
  assign N280 = N279 | data_masked[12546];
  assign N279 = N278 | data_masked[12674];
  assign N278 = N277 | data_masked[12802];
  assign N277 = N276 | data_masked[12930];
  assign N276 = N275 | data_masked[13058];
  assign N275 = N274 | data_masked[13186];
  assign N274 = N273 | data_masked[13314];
  assign N273 = N272 | data_masked[13442];
  assign N272 = N271 | data_masked[13570];
  assign N271 = N270 | data_masked[13698];
  assign N270 = N269 | data_masked[13826];
  assign N269 = N268 | data_masked[13954];
  assign N268 = N267 | data_masked[14082];
  assign N267 = N266 | data_masked[14210];
  assign N266 = N265 | data_masked[14338];
  assign N265 = N264 | data_masked[14466];
  assign N264 = N263 | data_masked[14594];
  assign N263 = N262 | data_masked[14722];
  assign N262 = N261 | data_masked[14850];
  assign N261 = N260 | data_masked[14978];
  assign N260 = N259 | data_masked[15106];
  assign N259 = N258 | data_masked[15234];
  assign N258 = N257 | data_masked[15362];
  assign N257 = N256 | data_masked[15490];
  assign N256 = N255 | data_masked[15618];
  assign N255 = N254 | data_masked[15746];
  assign N254 = N253 | data_masked[15874];
  assign N253 = N252 | data_masked[16002];
  assign N252 = data_masked[16258] | data_masked[16130];
  assign data_o[3] = N503 | data_masked[3];
  assign N503 = N502 | data_masked[131];
  assign N502 = N501 | data_masked[259];
  assign N501 = N500 | data_masked[387];
  assign N500 = N499 | data_masked[515];
  assign N499 = N498 | data_masked[643];
  assign N498 = N497 | data_masked[771];
  assign N497 = N496 | data_masked[899];
  assign N496 = N495 | data_masked[1027];
  assign N495 = N494 | data_masked[1155];
  assign N494 = N493 | data_masked[1283];
  assign N493 = N492 | data_masked[1411];
  assign N492 = N491 | data_masked[1539];
  assign N491 = N490 | data_masked[1667];
  assign N490 = N489 | data_masked[1795];
  assign N489 = N488 | data_masked[1923];
  assign N488 = N487 | data_masked[2051];
  assign N487 = N486 | data_masked[2179];
  assign N486 = N485 | data_masked[2307];
  assign N485 = N484 | data_masked[2435];
  assign N484 = N483 | data_masked[2563];
  assign N483 = N482 | data_masked[2691];
  assign N482 = N481 | data_masked[2819];
  assign N481 = N480 | data_masked[2947];
  assign N480 = N479 | data_masked[3075];
  assign N479 = N478 | data_masked[3203];
  assign N478 = N477 | data_masked[3331];
  assign N477 = N476 | data_masked[3459];
  assign N476 = N475 | data_masked[3587];
  assign N475 = N474 | data_masked[3715];
  assign N474 = N473 | data_masked[3843];
  assign N473 = N472 | data_masked[3971];
  assign N472 = N471 | data_masked[4099];
  assign N471 = N470 | data_masked[4227];
  assign N470 = N469 | data_masked[4355];
  assign N469 = N468 | data_masked[4483];
  assign N468 = N467 | data_masked[4611];
  assign N467 = N466 | data_masked[4739];
  assign N466 = N465 | data_masked[4867];
  assign N465 = N464 | data_masked[4995];
  assign N464 = N463 | data_masked[5123];
  assign N463 = N462 | data_masked[5251];
  assign N462 = N461 | data_masked[5379];
  assign N461 = N460 | data_masked[5507];
  assign N460 = N459 | data_masked[5635];
  assign N459 = N458 | data_masked[5763];
  assign N458 = N457 | data_masked[5891];
  assign N457 = N456 | data_masked[6019];
  assign N456 = N455 | data_masked[6147];
  assign N455 = N454 | data_masked[6275];
  assign N454 = N453 | data_masked[6403];
  assign N453 = N452 | data_masked[6531];
  assign N452 = N451 | data_masked[6659];
  assign N451 = N450 | data_masked[6787];
  assign N450 = N449 | data_masked[6915];
  assign N449 = N448 | data_masked[7043];
  assign N448 = N447 | data_masked[7171];
  assign N447 = N446 | data_masked[7299];
  assign N446 = N445 | data_masked[7427];
  assign N445 = N444 | data_masked[7555];
  assign N444 = N443 | data_masked[7683];
  assign N443 = N442 | data_masked[7811];
  assign N442 = N441 | data_masked[7939];
  assign N441 = N440 | data_masked[8067];
  assign N440 = N439 | data_masked[8195];
  assign N439 = N438 | data_masked[8323];
  assign N438 = N437 | data_masked[8451];
  assign N437 = N436 | data_masked[8579];
  assign N436 = N435 | data_masked[8707];
  assign N435 = N434 | data_masked[8835];
  assign N434 = N433 | data_masked[8963];
  assign N433 = N432 | data_masked[9091];
  assign N432 = N431 | data_masked[9219];
  assign N431 = N430 | data_masked[9347];
  assign N430 = N429 | data_masked[9475];
  assign N429 = N428 | data_masked[9603];
  assign N428 = N427 | data_masked[9731];
  assign N427 = N426 | data_masked[9859];
  assign N426 = N425 | data_masked[9987];
  assign N425 = N424 | data_masked[10115];
  assign N424 = N423 | data_masked[10243];
  assign N423 = N422 | data_masked[10371];
  assign N422 = N421 | data_masked[10499];
  assign N421 = N420 | data_masked[10627];
  assign N420 = N419 | data_masked[10755];
  assign N419 = N418 | data_masked[10883];
  assign N418 = N417 | data_masked[11011];
  assign N417 = N416 | data_masked[11139];
  assign N416 = N415 | data_masked[11267];
  assign N415 = N414 | data_masked[11395];
  assign N414 = N413 | data_masked[11523];
  assign N413 = N412 | data_masked[11651];
  assign N412 = N411 | data_masked[11779];
  assign N411 = N410 | data_masked[11907];
  assign N410 = N409 | data_masked[12035];
  assign N409 = N408 | data_masked[12163];
  assign N408 = N407 | data_masked[12291];
  assign N407 = N406 | data_masked[12419];
  assign N406 = N405 | data_masked[12547];
  assign N405 = N404 | data_masked[12675];
  assign N404 = N403 | data_masked[12803];
  assign N403 = N402 | data_masked[12931];
  assign N402 = N401 | data_masked[13059];
  assign N401 = N400 | data_masked[13187];
  assign N400 = N399 | data_masked[13315];
  assign N399 = N398 | data_masked[13443];
  assign N398 = N397 | data_masked[13571];
  assign N397 = N396 | data_masked[13699];
  assign N396 = N395 | data_masked[13827];
  assign N395 = N394 | data_masked[13955];
  assign N394 = N393 | data_masked[14083];
  assign N393 = N392 | data_masked[14211];
  assign N392 = N391 | data_masked[14339];
  assign N391 = N390 | data_masked[14467];
  assign N390 = N389 | data_masked[14595];
  assign N389 = N388 | data_masked[14723];
  assign N388 = N387 | data_masked[14851];
  assign N387 = N386 | data_masked[14979];
  assign N386 = N385 | data_masked[15107];
  assign N385 = N384 | data_masked[15235];
  assign N384 = N383 | data_masked[15363];
  assign N383 = N382 | data_masked[15491];
  assign N382 = N381 | data_masked[15619];
  assign N381 = N380 | data_masked[15747];
  assign N380 = N379 | data_masked[15875];
  assign N379 = N378 | data_masked[16003];
  assign N378 = data_masked[16259] | data_masked[16131];
  assign data_o[4] = N629 | data_masked[4];
  assign N629 = N628 | data_masked[132];
  assign N628 = N627 | data_masked[260];
  assign N627 = N626 | data_masked[388];
  assign N626 = N625 | data_masked[516];
  assign N625 = N624 | data_masked[644];
  assign N624 = N623 | data_masked[772];
  assign N623 = N622 | data_masked[900];
  assign N622 = N621 | data_masked[1028];
  assign N621 = N620 | data_masked[1156];
  assign N620 = N619 | data_masked[1284];
  assign N619 = N618 | data_masked[1412];
  assign N618 = N617 | data_masked[1540];
  assign N617 = N616 | data_masked[1668];
  assign N616 = N615 | data_masked[1796];
  assign N615 = N614 | data_masked[1924];
  assign N614 = N613 | data_masked[2052];
  assign N613 = N612 | data_masked[2180];
  assign N612 = N611 | data_masked[2308];
  assign N611 = N610 | data_masked[2436];
  assign N610 = N609 | data_masked[2564];
  assign N609 = N608 | data_masked[2692];
  assign N608 = N607 | data_masked[2820];
  assign N607 = N606 | data_masked[2948];
  assign N606 = N605 | data_masked[3076];
  assign N605 = N604 | data_masked[3204];
  assign N604 = N603 | data_masked[3332];
  assign N603 = N602 | data_masked[3460];
  assign N602 = N601 | data_masked[3588];
  assign N601 = N600 | data_masked[3716];
  assign N600 = N599 | data_masked[3844];
  assign N599 = N598 | data_masked[3972];
  assign N598 = N597 | data_masked[4100];
  assign N597 = N596 | data_masked[4228];
  assign N596 = N595 | data_masked[4356];
  assign N595 = N594 | data_masked[4484];
  assign N594 = N593 | data_masked[4612];
  assign N593 = N592 | data_masked[4740];
  assign N592 = N591 | data_masked[4868];
  assign N591 = N590 | data_masked[4996];
  assign N590 = N589 | data_masked[5124];
  assign N589 = N588 | data_masked[5252];
  assign N588 = N587 | data_masked[5380];
  assign N587 = N586 | data_masked[5508];
  assign N586 = N585 | data_masked[5636];
  assign N585 = N584 | data_masked[5764];
  assign N584 = N583 | data_masked[5892];
  assign N583 = N582 | data_masked[6020];
  assign N582 = N581 | data_masked[6148];
  assign N581 = N580 | data_masked[6276];
  assign N580 = N579 | data_masked[6404];
  assign N579 = N578 | data_masked[6532];
  assign N578 = N577 | data_masked[6660];
  assign N577 = N576 | data_masked[6788];
  assign N576 = N575 | data_masked[6916];
  assign N575 = N574 | data_masked[7044];
  assign N574 = N573 | data_masked[7172];
  assign N573 = N572 | data_masked[7300];
  assign N572 = N571 | data_masked[7428];
  assign N571 = N570 | data_masked[7556];
  assign N570 = N569 | data_masked[7684];
  assign N569 = N568 | data_masked[7812];
  assign N568 = N567 | data_masked[7940];
  assign N567 = N566 | data_masked[8068];
  assign N566 = N565 | data_masked[8196];
  assign N565 = N564 | data_masked[8324];
  assign N564 = N563 | data_masked[8452];
  assign N563 = N562 | data_masked[8580];
  assign N562 = N561 | data_masked[8708];
  assign N561 = N560 | data_masked[8836];
  assign N560 = N559 | data_masked[8964];
  assign N559 = N558 | data_masked[9092];
  assign N558 = N557 | data_masked[9220];
  assign N557 = N556 | data_masked[9348];
  assign N556 = N555 | data_masked[9476];
  assign N555 = N554 | data_masked[9604];
  assign N554 = N553 | data_masked[9732];
  assign N553 = N552 | data_masked[9860];
  assign N552 = N551 | data_masked[9988];
  assign N551 = N550 | data_masked[10116];
  assign N550 = N549 | data_masked[10244];
  assign N549 = N548 | data_masked[10372];
  assign N548 = N547 | data_masked[10500];
  assign N547 = N546 | data_masked[10628];
  assign N546 = N545 | data_masked[10756];
  assign N545 = N544 | data_masked[10884];
  assign N544 = N543 | data_masked[11012];
  assign N543 = N542 | data_masked[11140];
  assign N542 = N541 | data_masked[11268];
  assign N541 = N540 | data_masked[11396];
  assign N540 = N539 | data_masked[11524];
  assign N539 = N538 | data_masked[11652];
  assign N538 = N537 | data_masked[11780];
  assign N537 = N536 | data_masked[11908];
  assign N536 = N535 | data_masked[12036];
  assign N535 = N534 | data_masked[12164];
  assign N534 = N533 | data_masked[12292];
  assign N533 = N532 | data_masked[12420];
  assign N532 = N531 | data_masked[12548];
  assign N531 = N530 | data_masked[12676];
  assign N530 = N529 | data_masked[12804];
  assign N529 = N528 | data_masked[12932];
  assign N528 = N527 | data_masked[13060];
  assign N527 = N526 | data_masked[13188];
  assign N526 = N525 | data_masked[13316];
  assign N525 = N524 | data_masked[13444];
  assign N524 = N523 | data_masked[13572];
  assign N523 = N522 | data_masked[13700];
  assign N522 = N521 | data_masked[13828];
  assign N521 = N520 | data_masked[13956];
  assign N520 = N519 | data_masked[14084];
  assign N519 = N518 | data_masked[14212];
  assign N518 = N517 | data_masked[14340];
  assign N517 = N516 | data_masked[14468];
  assign N516 = N515 | data_masked[14596];
  assign N515 = N514 | data_masked[14724];
  assign N514 = N513 | data_masked[14852];
  assign N513 = N512 | data_masked[14980];
  assign N512 = N511 | data_masked[15108];
  assign N511 = N510 | data_masked[15236];
  assign N510 = N509 | data_masked[15364];
  assign N509 = N508 | data_masked[15492];
  assign N508 = N507 | data_masked[15620];
  assign N507 = N506 | data_masked[15748];
  assign N506 = N505 | data_masked[15876];
  assign N505 = N504 | data_masked[16004];
  assign N504 = data_masked[16260] | data_masked[16132];
  assign data_o[5] = N755 | data_masked[5];
  assign N755 = N754 | data_masked[133];
  assign N754 = N753 | data_masked[261];
  assign N753 = N752 | data_masked[389];
  assign N752 = N751 | data_masked[517];
  assign N751 = N750 | data_masked[645];
  assign N750 = N749 | data_masked[773];
  assign N749 = N748 | data_masked[901];
  assign N748 = N747 | data_masked[1029];
  assign N747 = N746 | data_masked[1157];
  assign N746 = N745 | data_masked[1285];
  assign N745 = N744 | data_masked[1413];
  assign N744 = N743 | data_masked[1541];
  assign N743 = N742 | data_masked[1669];
  assign N742 = N741 | data_masked[1797];
  assign N741 = N740 | data_masked[1925];
  assign N740 = N739 | data_masked[2053];
  assign N739 = N738 | data_masked[2181];
  assign N738 = N737 | data_masked[2309];
  assign N737 = N736 | data_masked[2437];
  assign N736 = N735 | data_masked[2565];
  assign N735 = N734 | data_masked[2693];
  assign N734 = N733 | data_masked[2821];
  assign N733 = N732 | data_masked[2949];
  assign N732 = N731 | data_masked[3077];
  assign N731 = N730 | data_masked[3205];
  assign N730 = N729 | data_masked[3333];
  assign N729 = N728 | data_masked[3461];
  assign N728 = N727 | data_masked[3589];
  assign N727 = N726 | data_masked[3717];
  assign N726 = N725 | data_masked[3845];
  assign N725 = N724 | data_masked[3973];
  assign N724 = N723 | data_masked[4101];
  assign N723 = N722 | data_masked[4229];
  assign N722 = N721 | data_masked[4357];
  assign N721 = N720 | data_masked[4485];
  assign N720 = N719 | data_masked[4613];
  assign N719 = N718 | data_masked[4741];
  assign N718 = N717 | data_masked[4869];
  assign N717 = N716 | data_masked[4997];
  assign N716 = N715 | data_masked[5125];
  assign N715 = N714 | data_masked[5253];
  assign N714 = N713 | data_masked[5381];
  assign N713 = N712 | data_masked[5509];
  assign N712 = N711 | data_masked[5637];
  assign N711 = N710 | data_masked[5765];
  assign N710 = N709 | data_masked[5893];
  assign N709 = N708 | data_masked[6021];
  assign N708 = N707 | data_masked[6149];
  assign N707 = N706 | data_masked[6277];
  assign N706 = N705 | data_masked[6405];
  assign N705 = N704 | data_masked[6533];
  assign N704 = N703 | data_masked[6661];
  assign N703 = N702 | data_masked[6789];
  assign N702 = N701 | data_masked[6917];
  assign N701 = N700 | data_masked[7045];
  assign N700 = N699 | data_masked[7173];
  assign N699 = N698 | data_masked[7301];
  assign N698 = N697 | data_masked[7429];
  assign N697 = N696 | data_masked[7557];
  assign N696 = N695 | data_masked[7685];
  assign N695 = N694 | data_masked[7813];
  assign N694 = N693 | data_masked[7941];
  assign N693 = N692 | data_masked[8069];
  assign N692 = N691 | data_masked[8197];
  assign N691 = N690 | data_masked[8325];
  assign N690 = N689 | data_masked[8453];
  assign N689 = N688 | data_masked[8581];
  assign N688 = N687 | data_masked[8709];
  assign N687 = N686 | data_masked[8837];
  assign N686 = N685 | data_masked[8965];
  assign N685 = N684 | data_masked[9093];
  assign N684 = N683 | data_masked[9221];
  assign N683 = N682 | data_masked[9349];
  assign N682 = N681 | data_masked[9477];
  assign N681 = N680 | data_masked[9605];
  assign N680 = N679 | data_masked[9733];
  assign N679 = N678 | data_masked[9861];
  assign N678 = N677 | data_masked[9989];
  assign N677 = N676 | data_masked[10117];
  assign N676 = N675 | data_masked[10245];
  assign N675 = N674 | data_masked[10373];
  assign N674 = N673 | data_masked[10501];
  assign N673 = N672 | data_masked[10629];
  assign N672 = N671 | data_masked[10757];
  assign N671 = N670 | data_masked[10885];
  assign N670 = N669 | data_masked[11013];
  assign N669 = N668 | data_masked[11141];
  assign N668 = N667 | data_masked[11269];
  assign N667 = N666 | data_masked[11397];
  assign N666 = N665 | data_masked[11525];
  assign N665 = N664 | data_masked[11653];
  assign N664 = N663 | data_masked[11781];
  assign N663 = N662 | data_masked[11909];
  assign N662 = N661 | data_masked[12037];
  assign N661 = N660 | data_masked[12165];
  assign N660 = N659 | data_masked[12293];
  assign N659 = N658 | data_masked[12421];
  assign N658 = N657 | data_masked[12549];
  assign N657 = N656 | data_masked[12677];
  assign N656 = N655 | data_masked[12805];
  assign N655 = N654 | data_masked[12933];
  assign N654 = N653 | data_masked[13061];
  assign N653 = N652 | data_masked[13189];
  assign N652 = N651 | data_masked[13317];
  assign N651 = N650 | data_masked[13445];
  assign N650 = N649 | data_masked[13573];
  assign N649 = N648 | data_masked[13701];
  assign N648 = N647 | data_masked[13829];
  assign N647 = N646 | data_masked[13957];
  assign N646 = N645 | data_masked[14085];
  assign N645 = N644 | data_masked[14213];
  assign N644 = N643 | data_masked[14341];
  assign N643 = N642 | data_masked[14469];
  assign N642 = N641 | data_masked[14597];
  assign N641 = N640 | data_masked[14725];
  assign N640 = N639 | data_masked[14853];
  assign N639 = N638 | data_masked[14981];
  assign N638 = N637 | data_masked[15109];
  assign N637 = N636 | data_masked[15237];
  assign N636 = N635 | data_masked[15365];
  assign N635 = N634 | data_masked[15493];
  assign N634 = N633 | data_masked[15621];
  assign N633 = N632 | data_masked[15749];
  assign N632 = N631 | data_masked[15877];
  assign N631 = N630 | data_masked[16005];
  assign N630 = data_masked[16261] | data_masked[16133];
  assign data_o[6] = N881 | data_masked[6];
  assign N881 = N880 | data_masked[134];
  assign N880 = N879 | data_masked[262];
  assign N879 = N878 | data_masked[390];
  assign N878 = N877 | data_masked[518];
  assign N877 = N876 | data_masked[646];
  assign N876 = N875 | data_masked[774];
  assign N875 = N874 | data_masked[902];
  assign N874 = N873 | data_masked[1030];
  assign N873 = N872 | data_masked[1158];
  assign N872 = N871 | data_masked[1286];
  assign N871 = N870 | data_masked[1414];
  assign N870 = N869 | data_masked[1542];
  assign N869 = N868 | data_masked[1670];
  assign N868 = N867 | data_masked[1798];
  assign N867 = N866 | data_masked[1926];
  assign N866 = N865 | data_masked[2054];
  assign N865 = N864 | data_masked[2182];
  assign N864 = N863 | data_masked[2310];
  assign N863 = N862 | data_masked[2438];
  assign N862 = N861 | data_masked[2566];
  assign N861 = N860 | data_masked[2694];
  assign N860 = N859 | data_masked[2822];
  assign N859 = N858 | data_masked[2950];
  assign N858 = N857 | data_masked[3078];
  assign N857 = N856 | data_masked[3206];
  assign N856 = N855 | data_masked[3334];
  assign N855 = N854 | data_masked[3462];
  assign N854 = N853 | data_masked[3590];
  assign N853 = N852 | data_masked[3718];
  assign N852 = N851 | data_masked[3846];
  assign N851 = N850 | data_masked[3974];
  assign N850 = N849 | data_masked[4102];
  assign N849 = N848 | data_masked[4230];
  assign N848 = N847 | data_masked[4358];
  assign N847 = N846 | data_masked[4486];
  assign N846 = N845 | data_masked[4614];
  assign N845 = N844 | data_masked[4742];
  assign N844 = N843 | data_masked[4870];
  assign N843 = N842 | data_masked[4998];
  assign N842 = N841 | data_masked[5126];
  assign N841 = N840 | data_masked[5254];
  assign N840 = N839 | data_masked[5382];
  assign N839 = N838 | data_masked[5510];
  assign N838 = N837 | data_masked[5638];
  assign N837 = N836 | data_masked[5766];
  assign N836 = N835 | data_masked[5894];
  assign N835 = N834 | data_masked[6022];
  assign N834 = N833 | data_masked[6150];
  assign N833 = N832 | data_masked[6278];
  assign N832 = N831 | data_masked[6406];
  assign N831 = N830 | data_masked[6534];
  assign N830 = N829 | data_masked[6662];
  assign N829 = N828 | data_masked[6790];
  assign N828 = N827 | data_masked[6918];
  assign N827 = N826 | data_masked[7046];
  assign N826 = N825 | data_masked[7174];
  assign N825 = N824 | data_masked[7302];
  assign N824 = N823 | data_masked[7430];
  assign N823 = N822 | data_masked[7558];
  assign N822 = N821 | data_masked[7686];
  assign N821 = N820 | data_masked[7814];
  assign N820 = N819 | data_masked[7942];
  assign N819 = N818 | data_masked[8070];
  assign N818 = N817 | data_masked[8198];
  assign N817 = N816 | data_masked[8326];
  assign N816 = N815 | data_masked[8454];
  assign N815 = N814 | data_masked[8582];
  assign N814 = N813 | data_masked[8710];
  assign N813 = N812 | data_masked[8838];
  assign N812 = N811 | data_masked[8966];
  assign N811 = N810 | data_masked[9094];
  assign N810 = N809 | data_masked[9222];
  assign N809 = N808 | data_masked[9350];
  assign N808 = N807 | data_masked[9478];
  assign N807 = N806 | data_masked[9606];
  assign N806 = N805 | data_masked[9734];
  assign N805 = N804 | data_masked[9862];
  assign N804 = N803 | data_masked[9990];
  assign N803 = N802 | data_masked[10118];
  assign N802 = N801 | data_masked[10246];
  assign N801 = N800 | data_masked[10374];
  assign N800 = N799 | data_masked[10502];
  assign N799 = N798 | data_masked[10630];
  assign N798 = N797 | data_masked[10758];
  assign N797 = N796 | data_masked[10886];
  assign N796 = N795 | data_masked[11014];
  assign N795 = N794 | data_masked[11142];
  assign N794 = N793 | data_masked[11270];
  assign N793 = N792 | data_masked[11398];
  assign N792 = N791 | data_masked[11526];
  assign N791 = N790 | data_masked[11654];
  assign N790 = N789 | data_masked[11782];
  assign N789 = N788 | data_masked[11910];
  assign N788 = N787 | data_masked[12038];
  assign N787 = N786 | data_masked[12166];
  assign N786 = N785 | data_masked[12294];
  assign N785 = N784 | data_masked[12422];
  assign N784 = N783 | data_masked[12550];
  assign N783 = N782 | data_masked[12678];
  assign N782 = N781 | data_masked[12806];
  assign N781 = N780 | data_masked[12934];
  assign N780 = N779 | data_masked[13062];
  assign N779 = N778 | data_masked[13190];
  assign N778 = N777 | data_masked[13318];
  assign N777 = N776 | data_masked[13446];
  assign N776 = N775 | data_masked[13574];
  assign N775 = N774 | data_masked[13702];
  assign N774 = N773 | data_masked[13830];
  assign N773 = N772 | data_masked[13958];
  assign N772 = N771 | data_masked[14086];
  assign N771 = N770 | data_masked[14214];
  assign N770 = N769 | data_masked[14342];
  assign N769 = N768 | data_masked[14470];
  assign N768 = N767 | data_masked[14598];
  assign N767 = N766 | data_masked[14726];
  assign N766 = N765 | data_masked[14854];
  assign N765 = N764 | data_masked[14982];
  assign N764 = N763 | data_masked[15110];
  assign N763 = N762 | data_masked[15238];
  assign N762 = N761 | data_masked[15366];
  assign N761 = N760 | data_masked[15494];
  assign N760 = N759 | data_masked[15622];
  assign N759 = N758 | data_masked[15750];
  assign N758 = N757 | data_masked[15878];
  assign N757 = N756 | data_masked[16006];
  assign N756 = data_masked[16262] | data_masked[16134];
  assign data_o[7] = N1007 | data_masked[7];
  assign N1007 = N1006 | data_masked[135];
  assign N1006 = N1005 | data_masked[263];
  assign N1005 = N1004 | data_masked[391];
  assign N1004 = N1003 | data_masked[519];
  assign N1003 = N1002 | data_masked[647];
  assign N1002 = N1001 | data_masked[775];
  assign N1001 = N1000 | data_masked[903];
  assign N1000 = N999 | data_masked[1031];
  assign N999 = N998 | data_masked[1159];
  assign N998 = N997 | data_masked[1287];
  assign N997 = N996 | data_masked[1415];
  assign N996 = N995 | data_masked[1543];
  assign N995 = N994 | data_masked[1671];
  assign N994 = N993 | data_masked[1799];
  assign N993 = N992 | data_masked[1927];
  assign N992 = N991 | data_masked[2055];
  assign N991 = N990 | data_masked[2183];
  assign N990 = N989 | data_masked[2311];
  assign N989 = N988 | data_masked[2439];
  assign N988 = N987 | data_masked[2567];
  assign N987 = N986 | data_masked[2695];
  assign N986 = N985 | data_masked[2823];
  assign N985 = N984 | data_masked[2951];
  assign N984 = N983 | data_masked[3079];
  assign N983 = N982 | data_masked[3207];
  assign N982 = N981 | data_masked[3335];
  assign N981 = N980 | data_masked[3463];
  assign N980 = N979 | data_masked[3591];
  assign N979 = N978 | data_masked[3719];
  assign N978 = N977 | data_masked[3847];
  assign N977 = N976 | data_masked[3975];
  assign N976 = N975 | data_masked[4103];
  assign N975 = N974 | data_masked[4231];
  assign N974 = N973 | data_masked[4359];
  assign N973 = N972 | data_masked[4487];
  assign N972 = N971 | data_masked[4615];
  assign N971 = N970 | data_masked[4743];
  assign N970 = N969 | data_masked[4871];
  assign N969 = N968 | data_masked[4999];
  assign N968 = N967 | data_masked[5127];
  assign N967 = N966 | data_masked[5255];
  assign N966 = N965 | data_masked[5383];
  assign N965 = N964 | data_masked[5511];
  assign N964 = N963 | data_masked[5639];
  assign N963 = N962 | data_masked[5767];
  assign N962 = N961 | data_masked[5895];
  assign N961 = N960 | data_masked[6023];
  assign N960 = N959 | data_masked[6151];
  assign N959 = N958 | data_masked[6279];
  assign N958 = N957 | data_masked[6407];
  assign N957 = N956 | data_masked[6535];
  assign N956 = N955 | data_masked[6663];
  assign N955 = N954 | data_masked[6791];
  assign N954 = N953 | data_masked[6919];
  assign N953 = N952 | data_masked[7047];
  assign N952 = N951 | data_masked[7175];
  assign N951 = N950 | data_masked[7303];
  assign N950 = N949 | data_masked[7431];
  assign N949 = N948 | data_masked[7559];
  assign N948 = N947 | data_masked[7687];
  assign N947 = N946 | data_masked[7815];
  assign N946 = N945 | data_masked[7943];
  assign N945 = N944 | data_masked[8071];
  assign N944 = N943 | data_masked[8199];
  assign N943 = N942 | data_masked[8327];
  assign N942 = N941 | data_masked[8455];
  assign N941 = N940 | data_masked[8583];
  assign N940 = N939 | data_masked[8711];
  assign N939 = N938 | data_masked[8839];
  assign N938 = N937 | data_masked[8967];
  assign N937 = N936 | data_masked[9095];
  assign N936 = N935 | data_masked[9223];
  assign N935 = N934 | data_masked[9351];
  assign N934 = N933 | data_masked[9479];
  assign N933 = N932 | data_masked[9607];
  assign N932 = N931 | data_masked[9735];
  assign N931 = N930 | data_masked[9863];
  assign N930 = N929 | data_masked[9991];
  assign N929 = N928 | data_masked[10119];
  assign N928 = N927 | data_masked[10247];
  assign N927 = N926 | data_masked[10375];
  assign N926 = N925 | data_masked[10503];
  assign N925 = N924 | data_masked[10631];
  assign N924 = N923 | data_masked[10759];
  assign N923 = N922 | data_masked[10887];
  assign N922 = N921 | data_masked[11015];
  assign N921 = N920 | data_masked[11143];
  assign N920 = N919 | data_masked[11271];
  assign N919 = N918 | data_masked[11399];
  assign N918 = N917 | data_masked[11527];
  assign N917 = N916 | data_masked[11655];
  assign N916 = N915 | data_masked[11783];
  assign N915 = N914 | data_masked[11911];
  assign N914 = N913 | data_masked[12039];
  assign N913 = N912 | data_masked[12167];
  assign N912 = N911 | data_masked[12295];
  assign N911 = N910 | data_masked[12423];
  assign N910 = N909 | data_masked[12551];
  assign N909 = N908 | data_masked[12679];
  assign N908 = N907 | data_masked[12807];
  assign N907 = N906 | data_masked[12935];
  assign N906 = N905 | data_masked[13063];
  assign N905 = N904 | data_masked[13191];
  assign N904 = N903 | data_masked[13319];
  assign N903 = N902 | data_masked[13447];
  assign N902 = N901 | data_masked[13575];
  assign N901 = N900 | data_masked[13703];
  assign N900 = N899 | data_masked[13831];
  assign N899 = N898 | data_masked[13959];
  assign N898 = N897 | data_masked[14087];
  assign N897 = N896 | data_masked[14215];
  assign N896 = N895 | data_masked[14343];
  assign N895 = N894 | data_masked[14471];
  assign N894 = N893 | data_masked[14599];
  assign N893 = N892 | data_masked[14727];
  assign N892 = N891 | data_masked[14855];
  assign N891 = N890 | data_masked[14983];
  assign N890 = N889 | data_masked[15111];
  assign N889 = N888 | data_masked[15239];
  assign N888 = N887 | data_masked[15367];
  assign N887 = N886 | data_masked[15495];
  assign N886 = N885 | data_masked[15623];
  assign N885 = N884 | data_masked[15751];
  assign N884 = N883 | data_masked[15879];
  assign N883 = N882 | data_masked[16007];
  assign N882 = data_masked[16263] | data_masked[16135];
  assign data_o[8] = N1133 | data_masked[8];
  assign N1133 = N1132 | data_masked[136];
  assign N1132 = N1131 | data_masked[264];
  assign N1131 = N1130 | data_masked[392];
  assign N1130 = N1129 | data_masked[520];
  assign N1129 = N1128 | data_masked[648];
  assign N1128 = N1127 | data_masked[776];
  assign N1127 = N1126 | data_masked[904];
  assign N1126 = N1125 | data_masked[1032];
  assign N1125 = N1124 | data_masked[1160];
  assign N1124 = N1123 | data_masked[1288];
  assign N1123 = N1122 | data_masked[1416];
  assign N1122 = N1121 | data_masked[1544];
  assign N1121 = N1120 | data_masked[1672];
  assign N1120 = N1119 | data_masked[1800];
  assign N1119 = N1118 | data_masked[1928];
  assign N1118 = N1117 | data_masked[2056];
  assign N1117 = N1116 | data_masked[2184];
  assign N1116 = N1115 | data_masked[2312];
  assign N1115 = N1114 | data_masked[2440];
  assign N1114 = N1113 | data_masked[2568];
  assign N1113 = N1112 | data_masked[2696];
  assign N1112 = N1111 | data_masked[2824];
  assign N1111 = N1110 | data_masked[2952];
  assign N1110 = N1109 | data_masked[3080];
  assign N1109 = N1108 | data_masked[3208];
  assign N1108 = N1107 | data_masked[3336];
  assign N1107 = N1106 | data_masked[3464];
  assign N1106 = N1105 | data_masked[3592];
  assign N1105 = N1104 | data_masked[3720];
  assign N1104 = N1103 | data_masked[3848];
  assign N1103 = N1102 | data_masked[3976];
  assign N1102 = N1101 | data_masked[4104];
  assign N1101 = N1100 | data_masked[4232];
  assign N1100 = N1099 | data_masked[4360];
  assign N1099 = N1098 | data_masked[4488];
  assign N1098 = N1097 | data_masked[4616];
  assign N1097 = N1096 | data_masked[4744];
  assign N1096 = N1095 | data_masked[4872];
  assign N1095 = N1094 | data_masked[5000];
  assign N1094 = N1093 | data_masked[5128];
  assign N1093 = N1092 | data_masked[5256];
  assign N1092 = N1091 | data_masked[5384];
  assign N1091 = N1090 | data_masked[5512];
  assign N1090 = N1089 | data_masked[5640];
  assign N1089 = N1088 | data_masked[5768];
  assign N1088 = N1087 | data_masked[5896];
  assign N1087 = N1086 | data_masked[6024];
  assign N1086 = N1085 | data_masked[6152];
  assign N1085 = N1084 | data_masked[6280];
  assign N1084 = N1083 | data_masked[6408];
  assign N1083 = N1082 | data_masked[6536];
  assign N1082 = N1081 | data_masked[6664];
  assign N1081 = N1080 | data_masked[6792];
  assign N1080 = N1079 | data_masked[6920];
  assign N1079 = N1078 | data_masked[7048];
  assign N1078 = N1077 | data_masked[7176];
  assign N1077 = N1076 | data_masked[7304];
  assign N1076 = N1075 | data_masked[7432];
  assign N1075 = N1074 | data_masked[7560];
  assign N1074 = N1073 | data_masked[7688];
  assign N1073 = N1072 | data_masked[7816];
  assign N1072 = N1071 | data_masked[7944];
  assign N1071 = N1070 | data_masked[8072];
  assign N1070 = N1069 | data_masked[8200];
  assign N1069 = N1068 | data_masked[8328];
  assign N1068 = N1067 | data_masked[8456];
  assign N1067 = N1066 | data_masked[8584];
  assign N1066 = N1065 | data_masked[8712];
  assign N1065 = N1064 | data_masked[8840];
  assign N1064 = N1063 | data_masked[8968];
  assign N1063 = N1062 | data_masked[9096];
  assign N1062 = N1061 | data_masked[9224];
  assign N1061 = N1060 | data_masked[9352];
  assign N1060 = N1059 | data_masked[9480];
  assign N1059 = N1058 | data_masked[9608];
  assign N1058 = N1057 | data_masked[9736];
  assign N1057 = N1056 | data_masked[9864];
  assign N1056 = N1055 | data_masked[9992];
  assign N1055 = N1054 | data_masked[10120];
  assign N1054 = N1053 | data_masked[10248];
  assign N1053 = N1052 | data_masked[10376];
  assign N1052 = N1051 | data_masked[10504];
  assign N1051 = N1050 | data_masked[10632];
  assign N1050 = N1049 | data_masked[10760];
  assign N1049 = N1048 | data_masked[10888];
  assign N1048 = N1047 | data_masked[11016];
  assign N1047 = N1046 | data_masked[11144];
  assign N1046 = N1045 | data_masked[11272];
  assign N1045 = N1044 | data_masked[11400];
  assign N1044 = N1043 | data_masked[11528];
  assign N1043 = N1042 | data_masked[11656];
  assign N1042 = N1041 | data_masked[11784];
  assign N1041 = N1040 | data_masked[11912];
  assign N1040 = N1039 | data_masked[12040];
  assign N1039 = N1038 | data_masked[12168];
  assign N1038 = N1037 | data_masked[12296];
  assign N1037 = N1036 | data_masked[12424];
  assign N1036 = N1035 | data_masked[12552];
  assign N1035 = N1034 | data_masked[12680];
  assign N1034 = N1033 | data_masked[12808];
  assign N1033 = N1032 | data_masked[12936];
  assign N1032 = N1031 | data_masked[13064];
  assign N1031 = N1030 | data_masked[13192];
  assign N1030 = N1029 | data_masked[13320];
  assign N1029 = N1028 | data_masked[13448];
  assign N1028 = N1027 | data_masked[13576];
  assign N1027 = N1026 | data_masked[13704];
  assign N1026 = N1025 | data_masked[13832];
  assign N1025 = N1024 | data_masked[13960];
  assign N1024 = N1023 | data_masked[14088];
  assign N1023 = N1022 | data_masked[14216];
  assign N1022 = N1021 | data_masked[14344];
  assign N1021 = N1020 | data_masked[14472];
  assign N1020 = N1019 | data_masked[14600];
  assign N1019 = N1018 | data_masked[14728];
  assign N1018 = N1017 | data_masked[14856];
  assign N1017 = N1016 | data_masked[14984];
  assign N1016 = N1015 | data_masked[15112];
  assign N1015 = N1014 | data_masked[15240];
  assign N1014 = N1013 | data_masked[15368];
  assign N1013 = N1012 | data_masked[15496];
  assign N1012 = N1011 | data_masked[15624];
  assign N1011 = N1010 | data_masked[15752];
  assign N1010 = N1009 | data_masked[15880];
  assign N1009 = N1008 | data_masked[16008];
  assign N1008 = data_masked[16264] | data_masked[16136];
  assign data_o[9] = N1259 | data_masked[9];
  assign N1259 = N1258 | data_masked[137];
  assign N1258 = N1257 | data_masked[265];
  assign N1257 = N1256 | data_masked[393];
  assign N1256 = N1255 | data_masked[521];
  assign N1255 = N1254 | data_masked[649];
  assign N1254 = N1253 | data_masked[777];
  assign N1253 = N1252 | data_masked[905];
  assign N1252 = N1251 | data_masked[1033];
  assign N1251 = N1250 | data_masked[1161];
  assign N1250 = N1249 | data_masked[1289];
  assign N1249 = N1248 | data_masked[1417];
  assign N1248 = N1247 | data_masked[1545];
  assign N1247 = N1246 | data_masked[1673];
  assign N1246 = N1245 | data_masked[1801];
  assign N1245 = N1244 | data_masked[1929];
  assign N1244 = N1243 | data_masked[2057];
  assign N1243 = N1242 | data_masked[2185];
  assign N1242 = N1241 | data_masked[2313];
  assign N1241 = N1240 | data_masked[2441];
  assign N1240 = N1239 | data_masked[2569];
  assign N1239 = N1238 | data_masked[2697];
  assign N1238 = N1237 | data_masked[2825];
  assign N1237 = N1236 | data_masked[2953];
  assign N1236 = N1235 | data_masked[3081];
  assign N1235 = N1234 | data_masked[3209];
  assign N1234 = N1233 | data_masked[3337];
  assign N1233 = N1232 | data_masked[3465];
  assign N1232 = N1231 | data_masked[3593];
  assign N1231 = N1230 | data_masked[3721];
  assign N1230 = N1229 | data_masked[3849];
  assign N1229 = N1228 | data_masked[3977];
  assign N1228 = N1227 | data_masked[4105];
  assign N1227 = N1226 | data_masked[4233];
  assign N1226 = N1225 | data_masked[4361];
  assign N1225 = N1224 | data_masked[4489];
  assign N1224 = N1223 | data_masked[4617];
  assign N1223 = N1222 | data_masked[4745];
  assign N1222 = N1221 | data_masked[4873];
  assign N1221 = N1220 | data_masked[5001];
  assign N1220 = N1219 | data_masked[5129];
  assign N1219 = N1218 | data_masked[5257];
  assign N1218 = N1217 | data_masked[5385];
  assign N1217 = N1216 | data_masked[5513];
  assign N1216 = N1215 | data_masked[5641];
  assign N1215 = N1214 | data_masked[5769];
  assign N1214 = N1213 | data_masked[5897];
  assign N1213 = N1212 | data_masked[6025];
  assign N1212 = N1211 | data_masked[6153];
  assign N1211 = N1210 | data_masked[6281];
  assign N1210 = N1209 | data_masked[6409];
  assign N1209 = N1208 | data_masked[6537];
  assign N1208 = N1207 | data_masked[6665];
  assign N1207 = N1206 | data_masked[6793];
  assign N1206 = N1205 | data_masked[6921];
  assign N1205 = N1204 | data_masked[7049];
  assign N1204 = N1203 | data_masked[7177];
  assign N1203 = N1202 | data_masked[7305];
  assign N1202 = N1201 | data_masked[7433];
  assign N1201 = N1200 | data_masked[7561];
  assign N1200 = N1199 | data_masked[7689];
  assign N1199 = N1198 | data_masked[7817];
  assign N1198 = N1197 | data_masked[7945];
  assign N1197 = N1196 | data_masked[8073];
  assign N1196 = N1195 | data_masked[8201];
  assign N1195 = N1194 | data_masked[8329];
  assign N1194 = N1193 | data_masked[8457];
  assign N1193 = N1192 | data_masked[8585];
  assign N1192 = N1191 | data_masked[8713];
  assign N1191 = N1190 | data_masked[8841];
  assign N1190 = N1189 | data_masked[8969];
  assign N1189 = N1188 | data_masked[9097];
  assign N1188 = N1187 | data_masked[9225];
  assign N1187 = N1186 | data_masked[9353];
  assign N1186 = N1185 | data_masked[9481];
  assign N1185 = N1184 | data_masked[9609];
  assign N1184 = N1183 | data_masked[9737];
  assign N1183 = N1182 | data_masked[9865];
  assign N1182 = N1181 | data_masked[9993];
  assign N1181 = N1180 | data_masked[10121];
  assign N1180 = N1179 | data_masked[10249];
  assign N1179 = N1178 | data_masked[10377];
  assign N1178 = N1177 | data_masked[10505];
  assign N1177 = N1176 | data_masked[10633];
  assign N1176 = N1175 | data_masked[10761];
  assign N1175 = N1174 | data_masked[10889];
  assign N1174 = N1173 | data_masked[11017];
  assign N1173 = N1172 | data_masked[11145];
  assign N1172 = N1171 | data_masked[11273];
  assign N1171 = N1170 | data_masked[11401];
  assign N1170 = N1169 | data_masked[11529];
  assign N1169 = N1168 | data_masked[11657];
  assign N1168 = N1167 | data_masked[11785];
  assign N1167 = N1166 | data_masked[11913];
  assign N1166 = N1165 | data_masked[12041];
  assign N1165 = N1164 | data_masked[12169];
  assign N1164 = N1163 | data_masked[12297];
  assign N1163 = N1162 | data_masked[12425];
  assign N1162 = N1161 | data_masked[12553];
  assign N1161 = N1160 | data_masked[12681];
  assign N1160 = N1159 | data_masked[12809];
  assign N1159 = N1158 | data_masked[12937];
  assign N1158 = N1157 | data_masked[13065];
  assign N1157 = N1156 | data_masked[13193];
  assign N1156 = N1155 | data_masked[13321];
  assign N1155 = N1154 | data_masked[13449];
  assign N1154 = N1153 | data_masked[13577];
  assign N1153 = N1152 | data_masked[13705];
  assign N1152 = N1151 | data_masked[13833];
  assign N1151 = N1150 | data_masked[13961];
  assign N1150 = N1149 | data_masked[14089];
  assign N1149 = N1148 | data_masked[14217];
  assign N1148 = N1147 | data_masked[14345];
  assign N1147 = N1146 | data_masked[14473];
  assign N1146 = N1145 | data_masked[14601];
  assign N1145 = N1144 | data_masked[14729];
  assign N1144 = N1143 | data_masked[14857];
  assign N1143 = N1142 | data_masked[14985];
  assign N1142 = N1141 | data_masked[15113];
  assign N1141 = N1140 | data_masked[15241];
  assign N1140 = N1139 | data_masked[15369];
  assign N1139 = N1138 | data_masked[15497];
  assign N1138 = N1137 | data_masked[15625];
  assign N1137 = N1136 | data_masked[15753];
  assign N1136 = N1135 | data_masked[15881];
  assign N1135 = N1134 | data_masked[16009];
  assign N1134 = data_masked[16265] | data_masked[16137];
  assign data_o[10] = N1385 | data_masked[10];
  assign N1385 = N1384 | data_masked[138];
  assign N1384 = N1383 | data_masked[266];
  assign N1383 = N1382 | data_masked[394];
  assign N1382 = N1381 | data_masked[522];
  assign N1381 = N1380 | data_masked[650];
  assign N1380 = N1379 | data_masked[778];
  assign N1379 = N1378 | data_masked[906];
  assign N1378 = N1377 | data_masked[1034];
  assign N1377 = N1376 | data_masked[1162];
  assign N1376 = N1375 | data_masked[1290];
  assign N1375 = N1374 | data_masked[1418];
  assign N1374 = N1373 | data_masked[1546];
  assign N1373 = N1372 | data_masked[1674];
  assign N1372 = N1371 | data_masked[1802];
  assign N1371 = N1370 | data_masked[1930];
  assign N1370 = N1369 | data_masked[2058];
  assign N1369 = N1368 | data_masked[2186];
  assign N1368 = N1367 | data_masked[2314];
  assign N1367 = N1366 | data_masked[2442];
  assign N1366 = N1365 | data_masked[2570];
  assign N1365 = N1364 | data_masked[2698];
  assign N1364 = N1363 | data_masked[2826];
  assign N1363 = N1362 | data_masked[2954];
  assign N1362 = N1361 | data_masked[3082];
  assign N1361 = N1360 | data_masked[3210];
  assign N1360 = N1359 | data_masked[3338];
  assign N1359 = N1358 | data_masked[3466];
  assign N1358 = N1357 | data_masked[3594];
  assign N1357 = N1356 | data_masked[3722];
  assign N1356 = N1355 | data_masked[3850];
  assign N1355 = N1354 | data_masked[3978];
  assign N1354 = N1353 | data_masked[4106];
  assign N1353 = N1352 | data_masked[4234];
  assign N1352 = N1351 | data_masked[4362];
  assign N1351 = N1350 | data_masked[4490];
  assign N1350 = N1349 | data_masked[4618];
  assign N1349 = N1348 | data_masked[4746];
  assign N1348 = N1347 | data_masked[4874];
  assign N1347 = N1346 | data_masked[5002];
  assign N1346 = N1345 | data_masked[5130];
  assign N1345 = N1344 | data_masked[5258];
  assign N1344 = N1343 | data_masked[5386];
  assign N1343 = N1342 | data_masked[5514];
  assign N1342 = N1341 | data_masked[5642];
  assign N1341 = N1340 | data_masked[5770];
  assign N1340 = N1339 | data_masked[5898];
  assign N1339 = N1338 | data_masked[6026];
  assign N1338 = N1337 | data_masked[6154];
  assign N1337 = N1336 | data_masked[6282];
  assign N1336 = N1335 | data_masked[6410];
  assign N1335 = N1334 | data_masked[6538];
  assign N1334 = N1333 | data_masked[6666];
  assign N1333 = N1332 | data_masked[6794];
  assign N1332 = N1331 | data_masked[6922];
  assign N1331 = N1330 | data_masked[7050];
  assign N1330 = N1329 | data_masked[7178];
  assign N1329 = N1328 | data_masked[7306];
  assign N1328 = N1327 | data_masked[7434];
  assign N1327 = N1326 | data_masked[7562];
  assign N1326 = N1325 | data_masked[7690];
  assign N1325 = N1324 | data_masked[7818];
  assign N1324 = N1323 | data_masked[7946];
  assign N1323 = N1322 | data_masked[8074];
  assign N1322 = N1321 | data_masked[8202];
  assign N1321 = N1320 | data_masked[8330];
  assign N1320 = N1319 | data_masked[8458];
  assign N1319 = N1318 | data_masked[8586];
  assign N1318 = N1317 | data_masked[8714];
  assign N1317 = N1316 | data_masked[8842];
  assign N1316 = N1315 | data_masked[8970];
  assign N1315 = N1314 | data_masked[9098];
  assign N1314 = N1313 | data_masked[9226];
  assign N1313 = N1312 | data_masked[9354];
  assign N1312 = N1311 | data_masked[9482];
  assign N1311 = N1310 | data_masked[9610];
  assign N1310 = N1309 | data_masked[9738];
  assign N1309 = N1308 | data_masked[9866];
  assign N1308 = N1307 | data_masked[9994];
  assign N1307 = N1306 | data_masked[10122];
  assign N1306 = N1305 | data_masked[10250];
  assign N1305 = N1304 | data_masked[10378];
  assign N1304 = N1303 | data_masked[10506];
  assign N1303 = N1302 | data_masked[10634];
  assign N1302 = N1301 | data_masked[10762];
  assign N1301 = N1300 | data_masked[10890];
  assign N1300 = N1299 | data_masked[11018];
  assign N1299 = N1298 | data_masked[11146];
  assign N1298 = N1297 | data_masked[11274];
  assign N1297 = N1296 | data_masked[11402];
  assign N1296 = N1295 | data_masked[11530];
  assign N1295 = N1294 | data_masked[11658];
  assign N1294 = N1293 | data_masked[11786];
  assign N1293 = N1292 | data_masked[11914];
  assign N1292 = N1291 | data_masked[12042];
  assign N1291 = N1290 | data_masked[12170];
  assign N1290 = N1289 | data_masked[12298];
  assign N1289 = N1288 | data_masked[12426];
  assign N1288 = N1287 | data_masked[12554];
  assign N1287 = N1286 | data_masked[12682];
  assign N1286 = N1285 | data_masked[12810];
  assign N1285 = N1284 | data_masked[12938];
  assign N1284 = N1283 | data_masked[13066];
  assign N1283 = N1282 | data_masked[13194];
  assign N1282 = N1281 | data_masked[13322];
  assign N1281 = N1280 | data_masked[13450];
  assign N1280 = N1279 | data_masked[13578];
  assign N1279 = N1278 | data_masked[13706];
  assign N1278 = N1277 | data_masked[13834];
  assign N1277 = N1276 | data_masked[13962];
  assign N1276 = N1275 | data_masked[14090];
  assign N1275 = N1274 | data_masked[14218];
  assign N1274 = N1273 | data_masked[14346];
  assign N1273 = N1272 | data_masked[14474];
  assign N1272 = N1271 | data_masked[14602];
  assign N1271 = N1270 | data_masked[14730];
  assign N1270 = N1269 | data_masked[14858];
  assign N1269 = N1268 | data_masked[14986];
  assign N1268 = N1267 | data_masked[15114];
  assign N1267 = N1266 | data_masked[15242];
  assign N1266 = N1265 | data_masked[15370];
  assign N1265 = N1264 | data_masked[15498];
  assign N1264 = N1263 | data_masked[15626];
  assign N1263 = N1262 | data_masked[15754];
  assign N1262 = N1261 | data_masked[15882];
  assign N1261 = N1260 | data_masked[16010];
  assign N1260 = data_masked[16266] | data_masked[16138];
  assign data_o[11] = N1511 | data_masked[11];
  assign N1511 = N1510 | data_masked[139];
  assign N1510 = N1509 | data_masked[267];
  assign N1509 = N1508 | data_masked[395];
  assign N1508 = N1507 | data_masked[523];
  assign N1507 = N1506 | data_masked[651];
  assign N1506 = N1505 | data_masked[779];
  assign N1505 = N1504 | data_masked[907];
  assign N1504 = N1503 | data_masked[1035];
  assign N1503 = N1502 | data_masked[1163];
  assign N1502 = N1501 | data_masked[1291];
  assign N1501 = N1500 | data_masked[1419];
  assign N1500 = N1499 | data_masked[1547];
  assign N1499 = N1498 | data_masked[1675];
  assign N1498 = N1497 | data_masked[1803];
  assign N1497 = N1496 | data_masked[1931];
  assign N1496 = N1495 | data_masked[2059];
  assign N1495 = N1494 | data_masked[2187];
  assign N1494 = N1493 | data_masked[2315];
  assign N1493 = N1492 | data_masked[2443];
  assign N1492 = N1491 | data_masked[2571];
  assign N1491 = N1490 | data_masked[2699];
  assign N1490 = N1489 | data_masked[2827];
  assign N1489 = N1488 | data_masked[2955];
  assign N1488 = N1487 | data_masked[3083];
  assign N1487 = N1486 | data_masked[3211];
  assign N1486 = N1485 | data_masked[3339];
  assign N1485 = N1484 | data_masked[3467];
  assign N1484 = N1483 | data_masked[3595];
  assign N1483 = N1482 | data_masked[3723];
  assign N1482 = N1481 | data_masked[3851];
  assign N1481 = N1480 | data_masked[3979];
  assign N1480 = N1479 | data_masked[4107];
  assign N1479 = N1478 | data_masked[4235];
  assign N1478 = N1477 | data_masked[4363];
  assign N1477 = N1476 | data_masked[4491];
  assign N1476 = N1475 | data_masked[4619];
  assign N1475 = N1474 | data_masked[4747];
  assign N1474 = N1473 | data_masked[4875];
  assign N1473 = N1472 | data_masked[5003];
  assign N1472 = N1471 | data_masked[5131];
  assign N1471 = N1470 | data_masked[5259];
  assign N1470 = N1469 | data_masked[5387];
  assign N1469 = N1468 | data_masked[5515];
  assign N1468 = N1467 | data_masked[5643];
  assign N1467 = N1466 | data_masked[5771];
  assign N1466 = N1465 | data_masked[5899];
  assign N1465 = N1464 | data_masked[6027];
  assign N1464 = N1463 | data_masked[6155];
  assign N1463 = N1462 | data_masked[6283];
  assign N1462 = N1461 | data_masked[6411];
  assign N1461 = N1460 | data_masked[6539];
  assign N1460 = N1459 | data_masked[6667];
  assign N1459 = N1458 | data_masked[6795];
  assign N1458 = N1457 | data_masked[6923];
  assign N1457 = N1456 | data_masked[7051];
  assign N1456 = N1455 | data_masked[7179];
  assign N1455 = N1454 | data_masked[7307];
  assign N1454 = N1453 | data_masked[7435];
  assign N1453 = N1452 | data_masked[7563];
  assign N1452 = N1451 | data_masked[7691];
  assign N1451 = N1450 | data_masked[7819];
  assign N1450 = N1449 | data_masked[7947];
  assign N1449 = N1448 | data_masked[8075];
  assign N1448 = N1447 | data_masked[8203];
  assign N1447 = N1446 | data_masked[8331];
  assign N1446 = N1445 | data_masked[8459];
  assign N1445 = N1444 | data_masked[8587];
  assign N1444 = N1443 | data_masked[8715];
  assign N1443 = N1442 | data_masked[8843];
  assign N1442 = N1441 | data_masked[8971];
  assign N1441 = N1440 | data_masked[9099];
  assign N1440 = N1439 | data_masked[9227];
  assign N1439 = N1438 | data_masked[9355];
  assign N1438 = N1437 | data_masked[9483];
  assign N1437 = N1436 | data_masked[9611];
  assign N1436 = N1435 | data_masked[9739];
  assign N1435 = N1434 | data_masked[9867];
  assign N1434 = N1433 | data_masked[9995];
  assign N1433 = N1432 | data_masked[10123];
  assign N1432 = N1431 | data_masked[10251];
  assign N1431 = N1430 | data_masked[10379];
  assign N1430 = N1429 | data_masked[10507];
  assign N1429 = N1428 | data_masked[10635];
  assign N1428 = N1427 | data_masked[10763];
  assign N1427 = N1426 | data_masked[10891];
  assign N1426 = N1425 | data_masked[11019];
  assign N1425 = N1424 | data_masked[11147];
  assign N1424 = N1423 | data_masked[11275];
  assign N1423 = N1422 | data_masked[11403];
  assign N1422 = N1421 | data_masked[11531];
  assign N1421 = N1420 | data_masked[11659];
  assign N1420 = N1419 | data_masked[11787];
  assign N1419 = N1418 | data_masked[11915];
  assign N1418 = N1417 | data_masked[12043];
  assign N1417 = N1416 | data_masked[12171];
  assign N1416 = N1415 | data_masked[12299];
  assign N1415 = N1414 | data_masked[12427];
  assign N1414 = N1413 | data_masked[12555];
  assign N1413 = N1412 | data_masked[12683];
  assign N1412 = N1411 | data_masked[12811];
  assign N1411 = N1410 | data_masked[12939];
  assign N1410 = N1409 | data_masked[13067];
  assign N1409 = N1408 | data_masked[13195];
  assign N1408 = N1407 | data_masked[13323];
  assign N1407 = N1406 | data_masked[13451];
  assign N1406 = N1405 | data_masked[13579];
  assign N1405 = N1404 | data_masked[13707];
  assign N1404 = N1403 | data_masked[13835];
  assign N1403 = N1402 | data_masked[13963];
  assign N1402 = N1401 | data_masked[14091];
  assign N1401 = N1400 | data_masked[14219];
  assign N1400 = N1399 | data_masked[14347];
  assign N1399 = N1398 | data_masked[14475];
  assign N1398 = N1397 | data_masked[14603];
  assign N1397 = N1396 | data_masked[14731];
  assign N1396 = N1395 | data_masked[14859];
  assign N1395 = N1394 | data_masked[14987];
  assign N1394 = N1393 | data_masked[15115];
  assign N1393 = N1392 | data_masked[15243];
  assign N1392 = N1391 | data_masked[15371];
  assign N1391 = N1390 | data_masked[15499];
  assign N1390 = N1389 | data_masked[15627];
  assign N1389 = N1388 | data_masked[15755];
  assign N1388 = N1387 | data_masked[15883];
  assign N1387 = N1386 | data_masked[16011];
  assign N1386 = data_masked[16267] | data_masked[16139];
  assign data_o[12] = N1637 | data_masked[12];
  assign N1637 = N1636 | data_masked[140];
  assign N1636 = N1635 | data_masked[268];
  assign N1635 = N1634 | data_masked[396];
  assign N1634 = N1633 | data_masked[524];
  assign N1633 = N1632 | data_masked[652];
  assign N1632 = N1631 | data_masked[780];
  assign N1631 = N1630 | data_masked[908];
  assign N1630 = N1629 | data_masked[1036];
  assign N1629 = N1628 | data_masked[1164];
  assign N1628 = N1627 | data_masked[1292];
  assign N1627 = N1626 | data_masked[1420];
  assign N1626 = N1625 | data_masked[1548];
  assign N1625 = N1624 | data_masked[1676];
  assign N1624 = N1623 | data_masked[1804];
  assign N1623 = N1622 | data_masked[1932];
  assign N1622 = N1621 | data_masked[2060];
  assign N1621 = N1620 | data_masked[2188];
  assign N1620 = N1619 | data_masked[2316];
  assign N1619 = N1618 | data_masked[2444];
  assign N1618 = N1617 | data_masked[2572];
  assign N1617 = N1616 | data_masked[2700];
  assign N1616 = N1615 | data_masked[2828];
  assign N1615 = N1614 | data_masked[2956];
  assign N1614 = N1613 | data_masked[3084];
  assign N1613 = N1612 | data_masked[3212];
  assign N1612 = N1611 | data_masked[3340];
  assign N1611 = N1610 | data_masked[3468];
  assign N1610 = N1609 | data_masked[3596];
  assign N1609 = N1608 | data_masked[3724];
  assign N1608 = N1607 | data_masked[3852];
  assign N1607 = N1606 | data_masked[3980];
  assign N1606 = N1605 | data_masked[4108];
  assign N1605 = N1604 | data_masked[4236];
  assign N1604 = N1603 | data_masked[4364];
  assign N1603 = N1602 | data_masked[4492];
  assign N1602 = N1601 | data_masked[4620];
  assign N1601 = N1600 | data_masked[4748];
  assign N1600 = N1599 | data_masked[4876];
  assign N1599 = N1598 | data_masked[5004];
  assign N1598 = N1597 | data_masked[5132];
  assign N1597 = N1596 | data_masked[5260];
  assign N1596 = N1595 | data_masked[5388];
  assign N1595 = N1594 | data_masked[5516];
  assign N1594 = N1593 | data_masked[5644];
  assign N1593 = N1592 | data_masked[5772];
  assign N1592 = N1591 | data_masked[5900];
  assign N1591 = N1590 | data_masked[6028];
  assign N1590 = N1589 | data_masked[6156];
  assign N1589 = N1588 | data_masked[6284];
  assign N1588 = N1587 | data_masked[6412];
  assign N1587 = N1586 | data_masked[6540];
  assign N1586 = N1585 | data_masked[6668];
  assign N1585 = N1584 | data_masked[6796];
  assign N1584 = N1583 | data_masked[6924];
  assign N1583 = N1582 | data_masked[7052];
  assign N1582 = N1581 | data_masked[7180];
  assign N1581 = N1580 | data_masked[7308];
  assign N1580 = N1579 | data_masked[7436];
  assign N1579 = N1578 | data_masked[7564];
  assign N1578 = N1577 | data_masked[7692];
  assign N1577 = N1576 | data_masked[7820];
  assign N1576 = N1575 | data_masked[7948];
  assign N1575 = N1574 | data_masked[8076];
  assign N1574 = N1573 | data_masked[8204];
  assign N1573 = N1572 | data_masked[8332];
  assign N1572 = N1571 | data_masked[8460];
  assign N1571 = N1570 | data_masked[8588];
  assign N1570 = N1569 | data_masked[8716];
  assign N1569 = N1568 | data_masked[8844];
  assign N1568 = N1567 | data_masked[8972];
  assign N1567 = N1566 | data_masked[9100];
  assign N1566 = N1565 | data_masked[9228];
  assign N1565 = N1564 | data_masked[9356];
  assign N1564 = N1563 | data_masked[9484];
  assign N1563 = N1562 | data_masked[9612];
  assign N1562 = N1561 | data_masked[9740];
  assign N1561 = N1560 | data_masked[9868];
  assign N1560 = N1559 | data_masked[9996];
  assign N1559 = N1558 | data_masked[10124];
  assign N1558 = N1557 | data_masked[10252];
  assign N1557 = N1556 | data_masked[10380];
  assign N1556 = N1555 | data_masked[10508];
  assign N1555 = N1554 | data_masked[10636];
  assign N1554 = N1553 | data_masked[10764];
  assign N1553 = N1552 | data_masked[10892];
  assign N1552 = N1551 | data_masked[11020];
  assign N1551 = N1550 | data_masked[11148];
  assign N1550 = N1549 | data_masked[11276];
  assign N1549 = N1548 | data_masked[11404];
  assign N1548 = N1547 | data_masked[11532];
  assign N1547 = N1546 | data_masked[11660];
  assign N1546 = N1545 | data_masked[11788];
  assign N1545 = N1544 | data_masked[11916];
  assign N1544 = N1543 | data_masked[12044];
  assign N1543 = N1542 | data_masked[12172];
  assign N1542 = N1541 | data_masked[12300];
  assign N1541 = N1540 | data_masked[12428];
  assign N1540 = N1539 | data_masked[12556];
  assign N1539 = N1538 | data_masked[12684];
  assign N1538 = N1537 | data_masked[12812];
  assign N1537 = N1536 | data_masked[12940];
  assign N1536 = N1535 | data_masked[13068];
  assign N1535 = N1534 | data_masked[13196];
  assign N1534 = N1533 | data_masked[13324];
  assign N1533 = N1532 | data_masked[13452];
  assign N1532 = N1531 | data_masked[13580];
  assign N1531 = N1530 | data_masked[13708];
  assign N1530 = N1529 | data_masked[13836];
  assign N1529 = N1528 | data_masked[13964];
  assign N1528 = N1527 | data_masked[14092];
  assign N1527 = N1526 | data_masked[14220];
  assign N1526 = N1525 | data_masked[14348];
  assign N1525 = N1524 | data_masked[14476];
  assign N1524 = N1523 | data_masked[14604];
  assign N1523 = N1522 | data_masked[14732];
  assign N1522 = N1521 | data_masked[14860];
  assign N1521 = N1520 | data_masked[14988];
  assign N1520 = N1519 | data_masked[15116];
  assign N1519 = N1518 | data_masked[15244];
  assign N1518 = N1517 | data_masked[15372];
  assign N1517 = N1516 | data_masked[15500];
  assign N1516 = N1515 | data_masked[15628];
  assign N1515 = N1514 | data_masked[15756];
  assign N1514 = N1513 | data_masked[15884];
  assign N1513 = N1512 | data_masked[16012];
  assign N1512 = data_masked[16268] | data_masked[16140];
  assign data_o[13] = N1763 | data_masked[13];
  assign N1763 = N1762 | data_masked[141];
  assign N1762 = N1761 | data_masked[269];
  assign N1761 = N1760 | data_masked[397];
  assign N1760 = N1759 | data_masked[525];
  assign N1759 = N1758 | data_masked[653];
  assign N1758 = N1757 | data_masked[781];
  assign N1757 = N1756 | data_masked[909];
  assign N1756 = N1755 | data_masked[1037];
  assign N1755 = N1754 | data_masked[1165];
  assign N1754 = N1753 | data_masked[1293];
  assign N1753 = N1752 | data_masked[1421];
  assign N1752 = N1751 | data_masked[1549];
  assign N1751 = N1750 | data_masked[1677];
  assign N1750 = N1749 | data_masked[1805];
  assign N1749 = N1748 | data_masked[1933];
  assign N1748 = N1747 | data_masked[2061];
  assign N1747 = N1746 | data_masked[2189];
  assign N1746 = N1745 | data_masked[2317];
  assign N1745 = N1744 | data_masked[2445];
  assign N1744 = N1743 | data_masked[2573];
  assign N1743 = N1742 | data_masked[2701];
  assign N1742 = N1741 | data_masked[2829];
  assign N1741 = N1740 | data_masked[2957];
  assign N1740 = N1739 | data_masked[3085];
  assign N1739 = N1738 | data_masked[3213];
  assign N1738 = N1737 | data_masked[3341];
  assign N1737 = N1736 | data_masked[3469];
  assign N1736 = N1735 | data_masked[3597];
  assign N1735 = N1734 | data_masked[3725];
  assign N1734 = N1733 | data_masked[3853];
  assign N1733 = N1732 | data_masked[3981];
  assign N1732 = N1731 | data_masked[4109];
  assign N1731 = N1730 | data_masked[4237];
  assign N1730 = N1729 | data_masked[4365];
  assign N1729 = N1728 | data_masked[4493];
  assign N1728 = N1727 | data_masked[4621];
  assign N1727 = N1726 | data_masked[4749];
  assign N1726 = N1725 | data_masked[4877];
  assign N1725 = N1724 | data_masked[5005];
  assign N1724 = N1723 | data_masked[5133];
  assign N1723 = N1722 | data_masked[5261];
  assign N1722 = N1721 | data_masked[5389];
  assign N1721 = N1720 | data_masked[5517];
  assign N1720 = N1719 | data_masked[5645];
  assign N1719 = N1718 | data_masked[5773];
  assign N1718 = N1717 | data_masked[5901];
  assign N1717 = N1716 | data_masked[6029];
  assign N1716 = N1715 | data_masked[6157];
  assign N1715 = N1714 | data_masked[6285];
  assign N1714 = N1713 | data_masked[6413];
  assign N1713 = N1712 | data_masked[6541];
  assign N1712 = N1711 | data_masked[6669];
  assign N1711 = N1710 | data_masked[6797];
  assign N1710 = N1709 | data_masked[6925];
  assign N1709 = N1708 | data_masked[7053];
  assign N1708 = N1707 | data_masked[7181];
  assign N1707 = N1706 | data_masked[7309];
  assign N1706 = N1705 | data_masked[7437];
  assign N1705 = N1704 | data_masked[7565];
  assign N1704 = N1703 | data_masked[7693];
  assign N1703 = N1702 | data_masked[7821];
  assign N1702 = N1701 | data_masked[7949];
  assign N1701 = N1700 | data_masked[8077];
  assign N1700 = N1699 | data_masked[8205];
  assign N1699 = N1698 | data_masked[8333];
  assign N1698 = N1697 | data_masked[8461];
  assign N1697 = N1696 | data_masked[8589];
  assign N1696 = N1695 | data_masked[8717];
  assign N1695 = N1694 | data_masked[8845];
  assign N1694 = N1693 | data_masked[8973];
  assign N1693 = N1692 | data_masked[9101];
  assign N1692 = N1691 | data_masked[9229];
  assign N1691 = N1690 | data_masked[9357];
  assign N1690 = N1689 | data_masked[9485];
  assign N1689 = N1688 | data_masked[9613];
  assign N1688 = N1687 | data_masked[9741];
  assign N1687 = N1686 | data_masked[9869];
  assign N1686 = N1685 | data_masked[9997];
  assign N1685 = N1684 | data_masked[10125];
  assign N1684 = N1683 | data_masked[10253];
  assign N1683 = N1682 | data_masked[10381];
  assign N1682 = N1681 | data_masked[10509];
  assign N1681 = N1680 | data_masked[10637];
  assign N1680 = N1679 | data_masked[10765];
  assign N1679 = N1678 | data_masked[10893];
  assign N1678 = N1677 | data_masked[11021];
  assign N1677 = N1676 | data_masked[11149];
  assign N1676 = N1675 | data_masked[11277];
  assign N1675 = N1674 | data_masked[11405];
  assign N1674 = N1673 | data_masked[11533];
  assign N1673 = N1672 | data_masked[11661];
  assign N1672 = N1671 | data_masked[11789];
  assign N1671 = N1670 | data_masked[11917];
  assign N1670 = N1669 | data_masked[12045];
  assign N1669 = N1668 | data_masked[12173];
  assign N1668 = N1667 | data_masked[12301];
  assign N1667 = N1666 | data_masked[12429];
  assign N1666 = N1665 | data_masked[12557];
  assign N1665 = N1664 | data_masked[12685];
  assign N1664 = N1663 | data_masked[12813];
  assign N1663 = N1662 | data_masked[12941];
  assign N1662 = N1661 | data_masked[13069];
  assign N1661 = N1660 | data_masked[13197];
  assign N1660 = N1659 | data_masked[13325];
  assign N1659 = N1658 | data_masked[13453];
  assign N1658 = N1657 | data_masked[13581];
  assign N1657 = N1656 | data_masked[13709];
  assign N1656 = N1655 | data_masked[13837];
  assign N1655 = N1654 | data_masked[13965];
  assign N1654 = N1653 | data_masked[14093];
  assign N1653 = N1652 | data_masked[14221];
  assign N1652 = N1651 | data_masked[14349];
  assign N1651 = N1650 | data_masked[14477];
  assign N1650 = N1649 | data_masked[14605];
  assign N1649 = N1648 | data_masked[14733];
  assign N1648 = N1647 | data_masked[14861];
  assign N1647 = N1646 | data_masked[14989];
  assign N1646 = N1645 | data_masked[15117];
  assign N1645 = N1644 | data_masked[15245];
  assign N1644 = N1643 | data_masked[15373];
  assign N1643 = N1642 | data_masked[15501];
  assign N1642 = N1641 | data_masked[15629];
  assign N1641 = N1640 | data_masked[15757];
  assign N1640 = N1639 | data_masked[15885];
  assign N1639 = N1638 | data_masked[16013];
  assign N1638 = data_masked[16269] | data_masked[16141];
  assign data_o[14] = N1889 | data_masked[14];
  assign N1889 = N1888 | data_masked[142];
  assign N1888 = N1887 | data_masked[270];
  assign N1887 = N1886 | data_masked[398];
  assign N1886 = N1885 | data_masked[526];
  assign N1885 = N1884 | data_masked[654];
  assign N1884 = N1883 | data_masked[782];
  assign N1883 = N1882 | data_masked[910];
  assign N1882 = N1881 | data_masked[1038];
  assign N1881 = N1880 | data_masked[1166];
  assign N1880 = N1879 | data_masked[1294];
  assign N1879 = N1878 | data_masked[1422];
  assign N1878 = N1877 | data_masked[1550];
  assign N1877 = N1876 | data_masked[1678];
  assign N1876 = N1875 | data_masked[1806];
  assign N1875 = N1874 | data_masked[1934];
  assign N1874 = N1873 | data_masked[2062];
  assign N1873 = N1872 | data_masked[2190];
  assign N1872 = N1871 | data_masked[2318];
  assign N1871 = N1870 | data_masked[2446];
  assign N1870 = N1869 | data_masked[2574];
  assign N1869 = N1868 | data_masked[2702];
  assign N1868 = N1867 | data_masked[2830];
  assign N1867 = N1866 | data_masked[2958];
  assign N1866 = N1865 | data_masked[3086];
  assign N1865 = N1864 | data_masked[3214];
  assign N1864 = N1863 | data_masked[3342];
  assign N1863 = N1862 | data_masked[3470];
  assign N1862 = N1861 | data_masked[3598];
  assign N1861 = N1860 | data_masked[3726];
  assign N1860 = N1859 | data_masked[3854];
  assign N1859 = N1858 | data_masked[3982];
  assign N1858 = N1857 | data_masked[4110];
  assign N1857 = N1856 | data_masked[4238];
  assign N1856 = N1855 | data_masked[4366];
  assign N1855 = N1854 | data_masked[4494];
  assign N1854 = N1853 | data_masked[4622];
  assign N1853 = N1852 | data_masked[4750];
  assign N1852 = N1851 | data_masked[4878];
  assign N1851 = N1850 | data_masked[5006];
  assign N1850 = N1849 | data_masked[5134];
  assign N1849 = N1848 | data_masked[5262];
  assign N1848 = N1847 | data_masked[5390];
  assign N1847 = N1846 | data_masked[5518];
  assign N1846 = N1845 | data_masked[5646];
  assign N1845 = N1844 | data_masked[5774];
  assign N1844 = N1843 | data_masked[5902];
  assign N1843 = N1842 | data_masked[6030];
  assign N1842 = N1841 | data_masked[6158];
  assign N1841 = N1840 | data_masked[6286];
  assign N1840 = N1839 | data_masked[6414];
  assign N1839 = N1838 | data_masked[6542];
  assign N1838 = N1837 | data_masked[6670];
  assign N1837 = N1836 | data_masked[6798];
  assign N1836 = N1835 | data_masked[6926];
  assign N1835 = N1834 | data_masked[7054];
  assign N1834 = N1833 | data_masked[7182];
  assign N1833 = N1832 | data_masked[7310];
  assign N1832 = N1831 | data_masked[7438];
  assign N1831 = N1830 | data_masked[7566];
  assign N1830 = N1829 | data_masked[7694];
  assign N1829 = N1828 | data_masked[7822];
  assign N1828 = N1827 | data_masked[7950];
  assign N1827 = N1826 | data_masked[8078];
  assign N1826 = N1825 | data_masked[8206];
  assign N1825 = N1824 | data_masked[8334];
  assign N1824 = N1823 | data_masked[8462];
  assign N1823 = N1822 | data_masked[8590];
  assign N1822 = N1821 | data_masked[8718];
  assign N1821 = N1820 | data_masked[8846];
  assign N1820 = N1819 | data_masked[8974];
  assign N1819 = N1818 | data_masked[9102];
  assign N1818 = N1817 | data_masked[9230];
  assign N1817 = N1816 | data_masked[9358];
  assign N1816 = N1815 | data_masked[9486];
  assign N1815 = N1814 | data_masked[9614];
  assign N1814 = N1813 | data_masked[9742];
  assign N1813 = N1812 | data_masked[9870];
  assign N1812 = N1811 | data_masked[9998];
  assign N1811 = N1810 | data_masked[10126];
  assign N1810 = N1809 | data_masked[10254];
  assign N1809 = N1808 | data_masked[10382];
  assign N1808 = N1807 | data_masked[10510];
  assign N1807 = N1806 | data_masked[10638];
  assign N1806 = N1805 | data_masked[10766];
  assign N1805 = N1804 | data_masked[10894];
  assign N1804 = N1803 | data_masked[11022];
  assign N1803 = N1802 | data_masked[11150];
  assign N1802 = N1801 | data_masked[11278];
  assign N1801 = N1800 | data_masked[11406];
  assign N1800 = N1799 | data_masked[11534];
  assign N1799 = N1798 | data_masked[11662];
  assign N1798 = N1797 | data_masked[11790];
  assign N1797 = N1796 | data_masked[11918];
  assign N1796 = N1795 | data_masked[12046];
  assign N1795 = N1794 | data_masked[12174];
  assign N1794 = N1793 | data_masked[12302];
  assign N1793 = N1792 | data_masked[12430];
  assign N1792 = N1791 | data_masked[12558];
  assign N1791 = N1790 | data_masked[12686];
  assign N1790 = N1789 | data_masked[12814];
  assign N1789 = N1788 | data_masked[12942];
  assign N1788 = N1787 | data_masked[13070];
  assign N1787 = N1786 | data_masked[13198];
  assign N1786 = N1785 | data_masked[13326];
  assign N1785 = N1784 | data_masked[13454];
  assign N1784 = N1783 | data_masked[13582];
  assign N1783 = N1782 | data_masked[13710];
  assign N1782 = N1781 | data_masked[13838];
  assign N1781 = N1780 | data_masked[13966];
  assign N1780 = N1779 | data_masked[14094];
  assign N1779 = N1778 | data_masked[14222];
  assign N1778 = N1777 | data_masked[14350];
  assign N1777 = N1776 | data_masked[14478];
  assign N1776 = N1775 | data_masked[14606];
  assign N1775 = N1774 | data_masked[14734];
  assign N1774 = N1773 | data_masked[14862];
  assign N1773 = N1772 | data_masked[14990];
  assign N1772 = N1771 | data_masked[15118];
  assign N1771 = N1770 | data_masked[15246];
  assign N1770 = N1769 | data_masked[15374];
  assign N1769 = N1768 | data_masked[15502];
  assign N1768 = N1767 | data_masked[15630];
  assign N1767 = N1766 | data_masked[15758];
  assign N1766 = N1765 | data_masked[15886];
  assign N1765 = N1764 | data_masked[16014];
  assign N1764 = data_masked[16270] | data_masked[16142];
  assign data_o[15] = N2015 | data_masked[15];
  assign N2015 = N2014 | data_masked[143];
  assign N2014 = N2013 | data_masked[271];
  assign N2013 = N2012 | data_masked[399];
  assign N2012 = N2011 | data_masked[527];
  assign N2011 = N2010 | data_masked[655];
  assign N2010 = N2009 | data_masked[783];
  assign N2009 = N2008 | data_masked[911];
  assign N2008 = N2007 | data_masked[1039];
  assign N2007 = N2006 | data_masked[1167];
  assign N2006 = N2005 | data_masked[1295];
  assign N2005 = N2004 | data_masked[1423];
  assign N2004 = N2003 | data_masked[1551];
  assign N2003 = N2002 | data_masked[1679];
  assign N2002 = N2001 | data_masked[1807];
  assign N2001 = N2000 | data_masked[1935];
  assign N2000 = N1999 | data_masked[2063];
  assign N1999 = N1998 | data_masked[2191];
  assign N1998 = N1997 | data_masked[2319];
  assign N1997 = N1996 | data_masked[2447];
  assign N1996 = N1995 | data_masked[2575];
  assign N1995 = N1994 | data_masked[2703];
  assign N1994 = N1993 | data_masked[2831];
  assign N1993 = N1992 | data_masked[2959];
  assign N1992 = N1991 | data_masked[3087];
  assign N1991 = N1990 | data_masked[3215];
  assign N1990 = N1989 | data_masked[3343];
  assign N1989 = N1988 | data_masked[3471];
  assign N1988 = N1987 | data_masked[3599];
  assign N1987 = N1986 | data_masked[3727];
  assign N1986 = N1985 | data_masked[3855];
  assign N1985 = N1984 | data_masked[3983];
  assign N1984 = N1983 | data_masked[4111];
  assign N1983 = N1982 | data_masked[4239];
  assign N1982 = N1981 | data_masked[4367];
  assign N1981 = N1980 | data_masked[4495];
  assign N1980 = N1979 | data_masked[4623];
  assign N1979 = N1978 | data_masked[4751];
  assign N1978 = N1977 | data_masked[4879];
  assign N1977 = N1976 | data_masked[5007];
  assign N1976 = N1975 | data_masked[5135];
  assign N1975 = N1974 | data_masked[5263];
  assign N1974 = N1973 | data_masked[5391];
  assign N1973 = N1972 | data_masked[5519];
  assign N1972 = N1971 | data_masked[5647];
  assign N1971 = N1970 | data_masked[5775];
  assign N1970 = N1969 | data_masked[5903];
  assign N1969 = N1968 | data_masked[6031];
  assign N1968 = N1967 | data_masked[6159];
  assign N1967 = N1966 | data_masked[6287];
  assign N1966 = N1965 | data_masked[6415];
  assign N1965 = N1964 | data_masked[6543];
  assign N1964 = N1963 | data_masked[6671];
  assign N1963 = N1962 | data_masked[6799];
  assign N1962 = N1961 | data_masked[6927];
  assign N1961 = N1960 | data_masked[7055];
  assign N1960 = N1959 | data_masked[7183];
  assign N1959 = N1958 | data_masked[7311];
  assign N1958 = N1957 | data_masked[7439];
  assign N1957 = N1956 | data_masked[7567];
  assign N1956 = N1955 | data_masked[7695];
  assign N1955 = N1954 | data_masked[7823];
  assign N1954 = N1953 | data_masked[7951];
  assign N1953 = N1952 | data_masked[8079];
  assign N1952 = N1951 | data_masked[8207];
  assign N1951 = N1950 | data_masked[8335];
  assign N1950 = N1949 | data_masked[8463];
  assign N1949 = N1948 | data_masked[8591];
  assign N1948 = N1947 | data_masked[8719];
  assign N1947 = N1946 | data_masked[8847];
  assign N1946 = N1945 | data_masked[8975];
  assign N1945 = N1944 | data_masked[9103];
  assign N1944 = N1943 | data_masked[9231];
  assign N1943 = N1942 | data_masked[9359];
  assign N1942 = N1941 | data_masked[9487];
  assign N1941 = N1940 | data_masked[9615];
  assign N1940 = N1939 | data_masked[9743];
  assign N1939 = N1938 | data_masked[9871];
  assign N1938 = N1937 | data_masked[9999];
  assign N1937 = N1936 | data_masked[10127];
  assign N1936 = N1935 | data_masked[10255];
  assign N1935 = N1934 | data_masked[10383];
  assign N1934 = N1933 | data_masked[10511];
  assign N1933 = N1932 | data_masked[10639];
  assign N1932 = N1931 | data_masked[10767];
  assign N1931 = N1930 | data_masked[10895];
  assign N1930 = N1929 | data_masked[11023];
  assign N1929 = N1928 | data_masked[11151];
  assign N1928 = N1927 | data_masked[11279];
  assign N1927 = N1926 | data_masked[11407];
  assign N1926 = N1925 | data_masked[11535];
  assign N1925 = N1924 | data_masked[11663];
  assign N1924 = N1923 | data_masked[11791];
  assign N1923 = N1922 | data_masked[11919];
  assign N1922 = N1921 | data_masked[12047];
  assign N1921 = N1920 | data_masked[12175];
  assign N1920 = N1919 | data_masked[12303];
  assign N1919 = N1918 | data_masked[12431];
  assign N1918 = N1917 | data_masked[12559];
  assign N1917 = N1916 | data_masked[12687];
  assign N1916 = N1915 | data_masked[12815];
  assign N1915 = N1914 | data_masked[12943];
  assign N1914 = N1913 | data_masked[13071];
  assign N1913 = N1912 | data_masked[13199];
  assign N1912 = N1911 | data_masked[13327];
  assign N1911 = N1910 | data_masked[13455];
  assign N1910 = N1909 | data_masked[13583];
  assign N1909 = N1908 | data_masked[13711];
  assign N1908 = N1907 | data_masked[13839];
  assign N1907 = N1906 | data_masked[13967];
  assign N1906 = N1905 | data_masked[14095];
  assign N1905 = N1904 | data_masked[14223];
  assign N1904 = N1903 | data_masked[14351];
  assign N1903 = N1902 | data_masked[14479];
  assign N1902 = N1901 | data_masked[14607];
  assign N1901 = N1900 | data_masked[14735];
  assign N1900 = N1899 | data_masked[14863];
  assign N1899 = N1898 | data_masked[14991];
  assign N1898 = N1897 | data_masked[15119];
  assign N1897 = N1896 | data_masked[15247];
  assign N1896 = N1895 | data_masked[15375];
  assign N1895 = N1894 | data_masked[15503];
  assign N1894 = N1893 | data_masked[15631];
  assign N1893 = N1892 | data_masked[15759];
  assign N1892 = N1891 | data_masked[15887];
  assign N1891 = N1890 | data_masked[16015];
  assign N1890 = data_masked[16271] | data_masked[16143];
  assign data_o[16] = N2141 | data_masked[16];
  assign N2141 = N2140 | data_masked[144];
  assign N2140 = N2139 | data_masked[272];
  assign N2139 = N2138 | data_masked[400];
  assign N2138 = N2137 | data_masked[528];
  assign N2137 = N2136 | data_masked[656];
  assign N2136 = N2135 | data_masked[784];
  assign N2135 = N2134 | data_masked[912];
  assign N2134 = N2133 | data_masked[1040];
  assign N2133 = N2132 | data_masked[1168];
  assign N2132 = N2131 | data_masked[1296];
  assign N2131 = N2130 | data_masked[1424];
  assign N2130 = N2129 | data_masked[1552];
  assign N2129 = N2128 | data_masked[1680];
  assign N2128 = N2127 | data_masked[1808];
  assign N2127 = N2126 | data_masked[1936];
  assign N2126 = N2125 | data_masked[2064];
  assign N2125 = N2124 | data_masked[2192];
  assign N2124 = N2123 | data_masked[2320];
  assign N2123 = N2122 | data_masked[2448];
  assign N2122 = N2121 | data_masked[2576];
  assign N2121 = N2120 | data_masked[2704];
  assign N2120 = N2119 | data_masked[2832];
  assign N2119 = N2118 | data_masked[2960];
  assign N2118 = N2117 | data_masked[3088];
  assign N2117 = N2116 | data_masked[3216];
  assign N2116 = N2115 | data_masked[3344];
  assign N2115 = N2114 | data_masked[3472];
  assign N2114 = N2113 | data_masked[3600];
  assign N2113 = N2112 | data_masked[3728];
  assign N2112 = N2111 | data_masked[3856];
  assign N2111 = N2110 | data_masked[3984];
  assign N2110 = N2109 | data_masked[4112];
  assign N2109 = N2108 | data_masked[4240];
  assign N2108 = N2107 | data_masked[4368];
  assign N2107 = N2106 | data_masked[4496];
  assign N2106 = N2105 | data_masked[4624];
  assign N2105 = N2104 | data_masked[4752];
  assign N2104 = N2103 | data_masked[4880];
  assign N2103 = N2102 | data_masked[5008];
  assign N2102 = N2101 | data_masked[5136];
  assign N2101 = N2100 | data_masked[5264];
  assign N2100 = N2099 | data_masked[5392];
  assign N2099 = N2098 | data_masked[5520];
  assign N2098 = N2097 | data_masked[5648];
  assign N2097 = N2096 | data_masked[5776];
  assign N2096 = N2095 | data_masked[5904];
  assign N2095 = N2094 | data_masked[6032];
  assign N2094 = N2093 | data_masked[6160];
  assign N2093 = N2092 | data_masked[6288];
  assign N2092 = N2091 | data_masked[6416];
  assign N2091 = N2090 | data_masked[6544];
  assign N2090 = N2089 | data_masked[6672];
  assign N2089 = N2088 | data_masked[6800];
  assign N2088 = N2087 | data_masked[6928];
  assign N2087 = N2086 | data_masked[7056];
  assign N2086 = N2085 | data_masked[7184];
  assign N2085 = N2084 | data_masked[7312];
  assign N2084 = N2083 | data_masked[7440];
  assign N2083 = N2082 | data_masked[7568];
  assign N2082 = N2081 | data_masked[7696];
  assign N2081 = N2080 | data_masked[7824];
  assign N2080 = N2079 | data_masked[7952];
  assign N2079 = N2078 | data_masked[8080];
  assign N2078 = N2077 | data_masked[8208];
  assign N2077 = N2076 | data_masked[8336];
  assign N2076 = N2075 | data_masked[8464];
  assign N2075 = N2074 | data_masked[8592];
  assign N2074 = N2073 | data_masked[8720];
  assign N2073 = N2072 | data_masked[8848];
  assign N2072 = N2071 | data_masked[8976];
  assign N2071 = N2070 | data_masked[9104];
  assign N2070 = N2069 | data_masked[9232];
  assign N2069 = N2068 | data_masked[9360];
  assign N2068 = N2067 | data_masked[9488];
  assign N2067 = N2066 | data_masked[9616];
  assign N2066 = N2065 | data_masked[9744];
  assign N2065 = N2064 | data_masked[9872];
  assign N2064 = N2063 | data_masked[10000];
  assign N2063 = N2062 | data_masked[10128];
  assign N2062 = N2061 | data_masked[10256];
  assign N2061 = N2060 | data_masked[10384];
  assign N2060 = N2059 | data_masked[10512];
  assign N2059 = N2058 | data_masked[10640];
  assign N2058 = N2057 | data_masked[10768];
  assign N2057 = N2056 | data_masked[10896];
  assign N2056 = N2055 | data_masked[11024];
  assign N2055 = N2054 | data_masked[11152];
  assign N2054 = N2053 | data_masked[11280];
  assign N2053 = N2052 | data_masked[11408];
  assign N2052 = N2051 | data_masked[11536];
  assign N2051 = N2050 | data_masked[11664];
  assign N2050 = N2049 | data_masked[11792];
  assign N2049 = N2048 | data_masked[11920];
  assign N2048 = N2047 | data_masked[12048];
  assign N2047 = N2046 | data_masked[12176];
  assign N2046 = N2045 | data_masked[12304];
  assign N2045 = N2044 | data_masked[12432];
  assign N2044 = N2043 | data_masked[12560];
  assign N2043 = N2042 | data_masked[12688];
  assign N2042 = N2041 | data_masked[12816];
  assign N2041 = N2040 | data_masked[12944];
  assign N2040 = N2039 | data_masked[13072];
  assign N2039 = N2038 | data_masked[13200];
  assign N2038 = N2037 | data_masked[13328];
  assign N2037 = N2036 | data_masked[13456];
  assign N2036 = N2035 | data_masked[13584];
  assign N2035 = N2034 | data_masked[13712];
  assign N2034 = N2033 | data_masked[13840];
  assign N2033 = N2032 | data_masked[13968];
  assign N2032 = N2031 | data_masked[14096];
  assign N2031 = N2030 | data_masked[14224];
  assign N2030 = N2029 | data_masked[14352];
  assign N2029 = N2028 | data_masked[14480];
  assign N2028 = N2027 | data_masked[14608];
  assign N2027 = N2026 | data_masked[14736];
  assign N2026 = N2025 | data_masked[14864];
  assign N2025 = N2024 | data_masked[14992];
  assign N2024 = N2023 | data_masked[15120];
  assign N2023 = N2022 | data_masked[15248];
  assign N2022 = N2021 | data_masked[15376];
  assign N2021 = N2020 | data_masked[15504];
  assign N2020 = N2019 | data_masked[15632];
  assign N2019 = N2018 | data_masked[15760];
  assign N2018 = N2017 | data_masked[15888];
  assign N2017 = N2016 | data_masked[16016];
  assign N2016 = data_masked[16272] | data_masked[16144];
  assign data_o[17] = N2267 | data_masked[17];
  assign N2267 = N2266 | data_masked[145];
  assign N2266 = N2265 | data_masked[273];
  assign N2265 = N2264 | data_masked[401];
  assign N2264 = N2263 | data_masked[529];
  assign N2263 = N2262 | data_masked[657];
  assign N2262 = N2261 | data_masked[785];
  assign N2261 = N2260 | data_masked[913];
  assign N2260 = N2259 | data_masked[1041];
  assign N2259 = N2258 | data_masked[1169];
  assign N2258 = N2257 | data_masked[1297];
  assign N2257 = N2256 | data_masked[1425];
  assign N2256 = N2255 | data_masked[1553];
  assign N2255 = N2254 | data_masked[1681];
  assign N2254 = N2253 | data_masked[1809];
  assign N2253 = N2252 | data_masked[1937];
  assign N2252 = N2251 | data_masked[2065];
  assign N2251 = N2250 | data_masked[2193];
  assign N2250 = N2249 | data_masked[2321];
  assign N2249 = N2248 | data_masked[2449];
  assign N2248 = N2247 | data_masked[2577];
  assign N2247 = N2246 | data_masked[2705];
  assign N2246 = N2245 | data_masked[2833];
  assign N2245 = N2244 | data_masked[2961];
  assign N2244 = N2243 | data_masked[3089];
  assign N2243 = N2242 | data_masked[3217];
  assign N2242 = N2241 | data_masked[3345];
  assign N2241 = N2240 | data_masked[3473];
  assign N2240 = N2239 | data_masked[3601];
  assign N2239 = N2238 | data_masked[3729];
  assign N2238 = N2237 | data_masked[3857];
  assign N2237 = N2236 | data_masked[3985];
  assign N2236 = N2235 | data_masked[4113];
  assign N2235 = N2234 | data_masked[4241];
  assign N2234 = N2233 | data_masked[4369];
  assign N2233 = N2232 | data_masked[4497];
  assign N2232 = N2231 | data_masked[4625];
  assign N2231 = N2230 | data_masked[4753];
  assign N2230 = N2229 | data_masked[4881];
  assign N2229 = N2228 | data_masked[5009];
  assign N2228 = N2227 | data_masked[5137];
  assign N2227 = N2226 | data_masked[5265];
  assign N2226 = N2225 | data_masked[5393];
  assign N2225 = N2224 | data_masked[5521];
  assign N2224 = N2223 | data_masked[5649];
  assign N2223 = N2222 | data_masked[5777];
  assign N2222 = N2221 | data_masked[5905];
  assign N2221 = N2220 | data_masked[6033];
  assign N2220 = N2219 | data_masked[6161];
  assign N2219 = N2218 | data_masked[6289];
  assign N2218 = N2217 | data_masked[6417];
  assign N2217 = N2216 | data_masked[6545];
  assign N2216 = N2215 | data_masked[6673];
  assign N2215 = N2214 | data_masked[6801];
  assign N2214 = N2213 | data_masked[6929];
  assign N2213 = N2212 | data_masked[7057];
  assign N2212 = N2211 | data_masked[7185];
  assign N2211 = N2210 | data_masked[7313];
  assign N2210 = N2209 | data_masked[7441];
  assign N2209 = N2208 | data_masked[7569];
  assign N2208 = N2207 | data_masked[7697];
  assign N2207 = N2206 | data_masked[7825];
  assign N2206 = N2205 | data_masked[7953];
  assign N2205 = N2204 | data_masked[8081];
  assign N2204 = N2203 | data_masked[8209];
  assign N2203 = N2202 | data_masked[8337];
  assign N2202 = N2201 | data_masked[8465];
  assign N2201 = N2200 | data_masked[8593];
  assign N2200 = N2199 | data_masked[8721];
  assign N2199 = N2198 | data_masked[8849];
  assign N2198 = N2197 | data_masked[8977];
  assign N2197 = N2196 | data_masked[9105];
  assign N2196 = N2195 | data_masked[9233];
  assign N2195 = N2194 | data_masked[9361];
  assign N2194 = N2193 | data_masked[9489];
  assign N2193 = N2192 | data_masked[9617];
  assign N2192 = N2191 | data_masked[9745];
  assign N2191 = N2190 | data_masked[9873];
  assign N2190 = N2189 | data_masked[10001];
  assign N2189 = N2188 | data_masked[10129];
  assign N2188 = N2187 | data_masked[10257];
  assign N2187 = N2186 | data_masked[10385];
  assign N2186 = N2185 | data_masked[10513];
  assign N2185 = N2184 | data_masked[10641];
  assign N2184 = N2183 | data_masked[10769];
  assign N2183 = N2182 | data_masked[10897];
  assign N2182 = N2181 | data_masked[11025];
  assign N2181 = N2180 | data_masked[11153];
  assign N2180 = N2179 | data_masked[11281];
  assign N2179 = N2178 | data_masked[11409];
  assign N2178 = N2177 | data_masked[11537];
  assign N2177 = N2176 | data_masked[11665];
  assign N2176 = N2175 | data_masked[11793];
  assign N2175 = N2174 | data_masked[11921];
  assign N2174 = N2173 | data_masked[12049];
  assign N2173 = N2172 | data_masked[12177];
  assign N2172 = N2171 | data_masked[12305];
  assign N2171 = N2170 | data_masked[12433];
  assign N2170 = N2169 | data_masked[12561];
  assign N2169 = N2168 | data_masked[12689];
  assign N2168 = N2167 | data_masked[12817];
  assign N2167 = N2166 | data_masked[12945];
  assign N2166 = N2165 | data_masked[13073];
  assign N2165 = N2164 | data_masked[13201];
  assign N2164 = N2163 | data_masked[13329];
  assign N2163 = N2162 | data_masked[13457];
  assign N2162 = N2161 | data_masked[13585];
  assign N2161 = N2160 | data_masked[13713];
  assign N2160 = N2159 | data_masked[13841];
  assign N2159 = N2158 | data_masked[13969];
  assign N2158 = N2157 | data_masked[14097];
  assign N2157 = N2156 | data_masked[14225];
  assign N2156 = N2155 | data_masked[14353];
  assign N2155 = N2154 | data_masked[14481];
  assign N2154 = N2153 | data_masked[14609];
  assign N2153 = N2152 | data_masked[14737];
  assign N2152 = N2151 | data_masked[14865];
  assign N2151 = N2150 | data_masked[14993];
  assign N2150 = N2149 | data_masked[15121];
  assign N2149 = N2148 | data_masked[15249];
  assign N2148 = N2147 | data_masked[15377];
  assign N2147 = N2146 | data_masked[15505];
  assign N2146 = N2145 | data_masked[15633];
  assign N2145 = N2144 | data_masked[15761];
  assign N2144 = N2143 | data_masked[15889];
  assign N2143 = N2142 | data_masked[16017];
  assign N2142 = data_masked[16273] | data_masked[16145];
  assign data_o[18] = N2393 | data_masked[18];
  assign N2393 = N2392 | data_masked[146];
  assign N2392 = N2391 | data_masked[274];
  assign N2391 = N2390 | data_masked[402];
  assign N2390 = N2389 | data_masked[530];
  assign N2389 = N2388 | data_masked[658];
  assign N2388 = N2387 | data_masked[786];
  assign N2387 = N2386 | data_masked[914];
  assign N2386 = N2385 | data_masked[1042];
  assign N2385 = N2384 | data_masked[1170];
  assign N2384 = N2383 | data_masked[1298];
  assign N2383 = N2382 | data_masked[1426];
  assign N2382 = N2381 | data_masked[1554];
  assign N2381 = N2380 | data_masked[1682];
  assign N2380 = N2379 | data_masked[1810];
  assign N2379 = N2378 | data_masked[1938];
  assign N2378 = N2377 | data_masked[2066];
  assign N2377 = N2376 | data_masked[2194];
  assign N2376 = N2375 | data_masked[2322];
  assign N2375 = N2374 | data_masked[2450];
  assign N2374 = N2373 | data_masked[2578];
  assign N2373 = N2372 | data_masked[2706];
  assign N2372 = N2371 | data_masked[2834];
  assign N2371 = N2370 | data_masked[2962];
  assign N2370 = N2369 | data_masked[3090];
  assign N2369 = N2368 | data_masked[3218];
  assign N2368 = N2367 | data_masked[3346];
  assign N2367 = N2366 | data_masked[3474];
  assign N2366 = N2365 | data_masked[3602];
  assign N2365 = N2364 | data_masked[3730];
  assign N2364 = N2363 | data_masked[3858];
  assign N2363 = N2362 | data_masked[3986];
  assign N2362 = N2361 | data_masked[4114];
  assign N2361 = N2360 | data_masked[4242];
  assign N2360 = N2359 | data_masked[4370];
  assign N2359 = N2358 | data_masked[4498];
  assign N2358 = N2357 | data_masked[4626];
  assign N2357 = N2356 | data_masked[4754];
  assign N2356 = N2355 | data_masked[4882];
  assign N2355 = N2354 | data_masked[5010];
  assign N2354 = N2353 | data_masked[5138];
  assign N2353 = N2352 | data_masked[5266];
  assign N2352 = N2351 | data_masked[5394];
  assign N2351 = N2350 | data_masked[5522];
  assign N2350 = N2349 | data_masked[5650];
  assign N2349 = N2348 | data_masked[5778];
  assign N2348 = N2347 | data_masked[5906];
  assign N2347 = N2346 | data_masked[6034];
  assign N2346 = N2345 | data_masked[6162];
  assign N2345 = N2344 | data_masked[6290];
  assign N2344 = N2343 | data_masked[6418];
  assign N2343 = N2342 | data_masked[6546];
  assign N2342 = N2341 | data_masked[6674];
  assign N2341 = N2340 | data_masked[6802];
  assign N2340 = N2339 | data_masked[6930];
  assign N2339 = N2338 | data_masked[7058];
  assign N2338 = N2337 | data_masked[7186];
  assign N2337 = N2336 | data_masked[7314];
  assign N2336 = N2335 | data_masked[7442];
  assign N2335 = N2334 | data_masked[7570];
  assign N2334 = N2333 | data_masked[7698];
  assign N2333 = N2332 | data_masked[7826];
  assign N2332 = N2331 | data_masked[7954];
  assign N2331 = N2330 | data_masked[8082];
  assign N2330 = N2329 | data_masked[8210];
  assign N2329 = N2328 | data_masked[8338];
  assign N2328 = N2327 | data_masked[8466];
  assign N2327 = N2326 | data_masked[8594];
  assign N2326 = N2325 | data_masked[8722];
  assign N2325 = N2324 | data_masked[8850];
  assign N2324 = N2323 | data_masked[8978];
  assign N2323 = N2322 | data_masked[9106];
  assign N2322 = N2321 | data_masked[9234];
  assign N2321 = N2320 | data_masked[9362];
  assign N2320 = N2319 | data_masked[9490];
  assign N2319 = N2318 | data_masked[9618];
  assign N2318 = N2317 | data_masked[9746];
  assign N2317 = N2316 | data_masked[9874];
  assign N2316 = N2315 | data_masked[10002];
  assign N2315 = N2314 | data_masked[10130];
  assign N2314 = N2313 | data_masked[10258];
  assign N2313 = N2312 | data_masked[10386];
  assign N2312 = N2311 | data_masked[10514];
  assign N2311 = N2310 | data_masked[10642];
  assign N2310 = N2309 | data_masked[10770];
  assign N2309 = N2308 | data_masked[10898];
  assign N2308 = N2307 | data_masked[11026];
  assign N2307 = N2306 | data_masked[11154];
  assign N2306 = N2305 | data_masked[11282];
  assign N2305 = N2304 | data_masked[11410];
  assign N2304 = N2303 | data_masked[11538];
  assign N2303 = N2302 | data_masked[11666];
  assign N2302 = N2301 | data_masked[11794];
  assign N2301 = N2300 | data_masked[11922];
  assign N2300 = N2299 | data_masked[12050];
  assign N2299 = N2298 | data_masked[12178];
  assign N2298 = N2297 | data_masked[12306];
  assign N2297 = N2296 | data_masked[12434];
  assign N2296 = N2295 | data_masked[12562];
  assign N2295 = N2294 | data_masked[12690];
  assign N2294 = N2293 | data_masked[12818];
  assign N2293 = N2292 | data_masked[12946];
  assign N2292 = N2291 | data_masked[13074];
  assign N2291 = N2290 | data_masked[13202];
  assign N2290 = N2289 | data_masked[13330];
  assign N2289 = N2288 | data_masked[13458];
  assign N2288 = N2287 | data_masked[13586];
  assign N2287 = N2286 | data_masked[13714];
  assign N2286 = N2285 | data_masked[13842];
  assign N2285 = N2284 | data_masked[13970];
  assign N2284 = N2283 | data_masked[14098];
  assign N2283 = N2282 | data_masked[14226];
  assign N2282 = N2281 | data_masked[14354];
  assign N2281 = N2280 | data_masked[14482];
  assign N2280 = N2279 | data_masked[14610];
  assign N2279 = N2278 | data_masked[14738];
  assign N2278 = N2277 | data_masked[14866];
  assign N2277 = N2276 | data_masked[14994];
  assign N2276 = N2275 | data_masked[15122];
  assign N2275 = N2274 | data_masked[15250];
  assign N2274 = N2273 | data_masked[15378];
  assign N2273 = N2272 | data_masked[15506];
  assign N2272 = N2271 | data_masked[15634];
  assign N2271 = N2270 | data_masked[15762];
  assign N2270 = N2269 | data_masked[15890];
  assign N2269 = N2268 | data_masked[16018];
  assign N2268 = data_masked[16274] | data_masked[16146];
  assign data_o[19] = N2519 | data_masked[19];
  assign N2519 = N2518 | data_masked[147];
  assign N2518 = N2517 | data_masked[275];
  assign N2517 = N2516 | data_masked[403];
  assign N2516 = N2515 | data_masked[531];
  assign N2515 = N2514 | data_masked[659];
  assign N2514 = N2513 | data_masked[787];
  assign N2513 = N2512 | data_masked[915];
  assign N2512 = N2511 | data_masked[1043];
  assign N2511 = N2510 | data_masked[1171];
  assign N2510 = N2509 | data_masked[1299];
  assign N2509 = N2508 | data_masked[1427];
  assign N2508 = N2507 | data_masked[1555];
  assign N2507 = N2506 | data_masked[1683];
  assign N2506 = N2505 | data_masked[1811];
  assign N2505 = N2504 | data_masked[1939];
  assign N2504 = N2503 | data_masked[2067];
  assign N2503 = N2502 | data_masked[2195];
  assign N2502 = N2501 | data_masked[2323];
  assign N2501 = N2500 | data_masked[2451];
  assign N2500 = N2499 | data_masked[2579];
  assign N2499 = N2498 | data_masked[2707];
  assign N2498 = N2497 | data_masked[2835];
  assign N2497 = N2496 | data_masked[2963];
  assign N2496 = N2495 | data_masked[3091];
  assign N2495 = N2494 | data_masked[3219];
  assign N2494 = N2493 | data_masked[3347];
  assign N2493 = N2492 | data_masked[3475];
  assign N2492 = N2491 | data_masked[3603];
  assign N2491 = N2490 | data_masked[3731];
  assign N2490 = N2489 | data_masked[3859];
  assign N2489 = N2488 | data_masked[3987];
  assign N2488 = N2487 | data_masked[4115];
  assign N2487 = N2486 | data_masked[4243];
  assign N2486 = N2485 | data_masked[4371];
  assign N2485 = N2484 | data_masked[4499];
  assign N2484 = N2483 | data_masked[4627];
  assign N2483 = N2482 | data_masked[4755];
  assign N2482 = N2481 | data_masked[4883];
  assign N2481 = N2480 | data_masked[5011];
  assign N2480 = N2479 | data_masked[5139];
  assign N2479 = N2478 | data_masked[5267];
  assign N2478 = N2477 | data_masked[5395];
  assign N2477 = N2476 | data_masked[5523];
  assign N2476 = N2475 | data_masked[5651];
  assign N2475 = N2474 | data_masked[5779];
  assign N2474 = N2473 | data_masked[5907];
  assign N2473 = N2472 | data_masked[6035];
  assign N2472 = N2471 | data_masked[6163];
  assign N2471 = N2470 | data_masked[6291];
  assign N2470 = N2469 | data_masked[6419];
  assign N2469 = N2468 | data_masked[6547];
  assign N2468 = N2467 | data_masked[6675];
  assign N2467 = N2466 | data_masked[6803];
  assign N2466 = N2465 | data_masked[6931];
  assign N2465 = N2464 | data_masked[7059];
  assign N2464 = N2463 | data_masked[7187];
  assign N2463 = N2462 | data_masked[7315];
  assign N2462 = N2461 | data_masked[7443];
  assign N2461 = N2460 | data_masked[7571];
  assign N2460 = N2459 | data_masked[7699];
  assign N2459 = N2458 | data_masked[7827];
  assign N2458 = N2457 | data_masked[7955];
  assign N2457 = N2456 | data_masked[8083];
  assign N2456 = N2455 | data_masked[8211];
  assign N2455 = N2454 | data_masked[8339];
  assign N2454 = N2453 | data_masked[8467];
  assign N2453 = N2452 | data_masked[8595];
  assign N2452 = N2451 | data_masked[8723];
  assign N2451 = N2450 | data_masked[8851];
  assign N2450 = N2449 | data_masked[8979];
  assign N2449 = N2448 | data_masked[9107];
  assign N2448 = N2447 | data_masked[9235];
  assign N2447 = N2446 | data_masked[9363];
  assign N2446 = N2445 | data_masked[9491];
  assign N2445 = N2444 | data_masked[9619];
  assign N2444 = N2443 | data_masked[9747];
  assign N2443 = N2442 | data_masked[9875];
  assign N2442 = N2441 | data_masked[10003];
  assign N2441 = N2440 | data_masked[10131];
  assign N2440 = N2439 | data_masked[10259];
  assign N2439 = N2438 | data_masked[10387];
  assign N2438 = N2437 | data_masked[10515];
  assign N2437 = N2436 | data_masked[10643];
  assign N2436 = N2435 | data_masked[10771];
  assign N2435 = N2434 | data_masked[10899];
  assign N2434 = N2433 | data_masked[11027];
  assign N2433 = N2432 | data_masked[11155];
  assign N2432 = N2431 | data_masked[11283];
  assign N2431 = N2430 | data_masked[11411];
  assign N2430 = N2429 | data_masked[11539];
  assign N2429 = N2428 | data_masked[11667];
  assign N2428 = N2427 | data_masked[11795];
  assign N2427 = N2426 | data_masked[11923];
  assign N2426 = N2425 | data_masked[12051];
  assign N2425 = N2424 | data_masked[12179];
  assign N2424 = N2423 | data_masked[12307];
  assign N2423 = N2422 | data_masked[12435];
  assign N2422 = N2421 | data_masked[12563];
  assign N2421 = N2420 | data_masked[12691];
  assign N2420 = N2419 | data_masked[12819];
  assign N2419 = N2418 | data_masked[12947];
  assign N2418 = N2417 | data_masked[13075];
  assign N2417 = N2416 | data_masked[13203];
  assign N2416 = N2415 | data_masked[13331];
  assign N2415 = N2414 | data_masked[13459];
  assign N2414 = N2413 | data_masked[13587];
  assign N2413 = N2412 | data_masked[13715];
  assign N2412 = N2411 | data_masked[13843];
  assign N2411 = N2410 | data_masked[13971];
  assign N2410 = N2409 | data_masked[14099];
  assign N2409 = N2408 | data_masked[14227];
  assign N2408 = N2407 | data_masked[14355];
  assign N2407 = N2406 | data_masked[14483];
  assign N2406 = N2405 | data_masked[14611];
  assign N2405 = N2404 | data_masked[14739];
  assign N2404 = N2403 | data_masked[14867];
  assign N2403 = N2402 | data_masked[14995];
  assign N2402 = N2401 | data_masked[15123];
  assign N2401 = N2400 | data_masked[15251];
  assign N2400 = N2399 | data_masked[15379];
  assign N2399 = N2398 | data_masked[15507];
  assign N2398 = N2397 | data_masked[15635];
  assign N2397 = N2396 | data_masked[15763];
  assign N2396 = N2395 | data_masked[15891];
  assign N2395 = N2394 | data_masked[16019];
  assign N2394 = data_masked[16275] | data_masked[16147];
  assign data_o[20] = N2645 | data_masked[20];
  assign N2645 = N2644 | data_masked[148];
  assign N2644 = N2643 | data_masked[276];
  assign N2643 = N2642 | data_masked[404];
  assign N2642 = N2641 | data_masked[532];
  assign N2641 = N2640 | data_masked[660];
  assign N2640 = N2639 | data_masked[788];
  assign N2639 = N2638 | data_masked[916];
  assign N2638 = N2637 | data_masked[1044];
  assign N2637 = N2636 | data_masked[1172];
  assign N2636 = N2635 | data_masked[1300];
  assign N2635 = N2634 | data_masked[1428];
  assign N2634 = N2633 | data_masked[1556];
  assign N2633 = N2632 | data_masked[1684];
  assign N2632 = N2631 | data_masked[1812];
  assign N2631 = N2630 | data_masked[1940];
  assign N2630 = N2629 | data_masked[2068];
  assign N2629 = N2628 | data_masked[2196];
  assign N2628 = N2627 | data_masked[2324];
  assign N2627 = N2626 | data_masked[2452];
  assign N2626 = N2625 | data_masked[2580];
  assign N2625 = N2624 | data_masked[2708];
  assign N2624 = N2623 | data_masked[2836];
  assign N2623 = N2622 | data_masked[2964];
  assign N2622 = N2621 | data_masked[3092];
  assign N2621 = N2620 | data_masked[3220];
  assign N2620 = N2619 | data_masked[3348];
  assign N2619 = N2618 | data_masked[3476];
  assign N2618 = N2617 | data_masked[3604];
  assign N2617 = N2616 | data_masked[3732];
  assign N2616 = N2615 | data_masked[3860];
  assign N2615 = N2614 | data_masked[3988];
  assign N2614 = N2613 | data_masked[4116];
  assign N2613 = N2612 | data_masked[4244];
  assign N2612 = N2611 | data_masked[4372];
  assign N2611 = N2610 | data_masked[4500];
  assign N2610 = N2609 | data_masked[4628];
  assign N2609 = N2608 | data_masked[4756];
  assign N2608 = N2607 | data_masked[4884];
  assign N2607 = N2606 | data_masked[5012];
  assign N2606 = N2605 | data_masked[5140];
  assign N2605 = N2604 | data_masked[5268];
  assign N2604 = N2603 | data_masked[5396];
  assign N2603 = N2602 | data_masked[5524];
  assign N2602 = N2601 | data_masked[5652];
  assign N2601 = N2600 | data_masked[5780];
  assign N2600 = N2599 | data_masked[5908];
  assign N2599 = N2598 | data_masked[6036];
  assign N2598 = N2597 | data_masked[6164];
  assign N2597 = N2596 | data_masked[6292];
  assign N2596 = N2595 | data_masked[6420];
  assign N2595 = N2594 | data_masked[6548];
  assign N2594 = N2593 | data_masked[6676];
  assign N2593 = N2592 | data_masked[6804];
  assign N2592 = N2591 | data_masked[6932];
  assign N2591 = N2590 | data_masked[7060];
  assign N2590 = N2589 | data_masked[7188];
  assign N2589 = N2588 | data_masked[7316];
  assign N2588 = N2587 | data_masked[7444];
  assign N2587 = N2586 | data_masked[7572];
  assign N2586 = N2585 | data_masked[7700];
  assign N2585 = N2584 | data_masked[7828];
  assign N2584 = N2583 | data_masked[7956];
  assign N2583 = N2582 | data_masked[8084];
  assign N2582 = N2581 | data_masked[8212];
  assign N2581 = N2580 | data_masked[8340];
  assign N2580 = N2579 | data_masked[8468];
  assign N2579 = N2578 | data_masked[8596];
  assign N2578 = N2577 | data_masked[8724];
  assign N2577 = N2576 | data_masked[8852];
  assign N2576 = N2575 | data_masked[8980];
  assign N2575 = N2574 | data_masked[9108];
  assign N2574 = N2573 | data_masked[9236];
  assign N2573 = N2572 | data_masked[9364];
  assign N2572 = N2571 | data_masked[9492];
  assign N2571 = N2570 | data_masked[9620];
  assign N2570 = N2569 | data_masked[9748];
  assign N2569 = N2568 | data_masked[9876];
  assign N2568 = N2567 | data_masked[10004];
  assign N2567 = N2566 | data_masked[10132];
  assign N2566 = N2565 | data_masked[10260];
  assign N2565 = N2564 | data_masked[10388];
  assign N2564 = N2563 | data_masked[10516];
  assign N2563 = N2562 | data_masked[10644];
  assign N2562 = N2561 | data_masked[10772];
  assign N2561 = N2560 | data_masked[10900];
  assign N2560 = N2559 | data_masked[11028];
  assign N2559 = N2558 | data_masked[11156];
  assign N2558 = N2557 | data_masked[11284];
  assign N2557 = N2556 | data_masked[11412];
  assign N2556 = N2555 | data_masked[11540];
  assign N2555 = N2554 | data_masked[11668];
  assign N2554 = N2553 | data_masked[11796];
  assign N2553 = N2552 | data_masked[11924];
  assign N2552 = N2551 | data_masked[12052];
  assign N2551 = N2550 | data_masked[12180];
  assign N2550 = N2549 | data_masked[12308];
  assign N2549 = N2548 | data_masked[12436];
  assign N2548 = N2547 | data_masked[12564];
  assign N2547 = N2546 | data_masked[12692];
  assign N2546 = N2545 | data_masked[12820];
  assign N2545 = N2544 | data_masked[12948];
  assign N2544 = N2543 | data_masked[13076];
  assign N2543 = N2542 | data_masked[13204];
  assign N2542 = N2541 | data_masked[13332];
  assign N2541 = N2540 | data_masked[13460];
  assign N2540 = N2539 | data_masked[13588];
  assign N2539 = N2538 | data_masked[13716];
  assign N2538 = N2537 | data_masked[13844];
  assign N2537 = N2536 | data_masked[13972];
  assign N2536 = N2535 | data_masked[14100];
  assign N2535 = N2534 | data_masked[14228];
  assign N2534 = N2533 | data_masked[14356];
  assign N2533 = N2532 | data_masked[14484];
  assign N2532 = N2531 | data_masked[14612];
  assign N2531 = N2530 | data_masked[14740];
  assign N2530 = N2529 | data_masked[14868];
  assign N2529 = N2528 | data_masked[14996];
  assign N2528 = N2527 | data_masked[15124];
  assign N2527 = N2526 | data_masked[15252];
  assign N2526 = N2525 | data_masked[15380];
  assign N2525 = N2524 | data_masked[15508];
  assign N2524 = N2523 | data_masked[15636];
  assign N2523 = N2522 | data_masked[15764];
  assign N2522 = N2521 | data_masked[15892];
  assign N2521 = N2520 | data_masked[16020];
  assign N2520 = data_masked[16276] | data_masked[16148];
  assign data_o[21] = N2771 | data_masked[21];
  assign N2771 = N2770 | data_masked[149];
  assign N2770 = N2769 | data_masked[277];
  assign N2769 = N2768 | data_masked[405];
  assign N2768 = N2767 | data_masked[533];
  assign N2767 = N2766 | data_masked[661];
  assign N2766 = N2765 | data_masked[789];
  assign N2765 = N2764 | data_masked[917];
  assign N2764 = N2763 | data_masked[1045];
  assign N2763 = N2762 | data_masked[1173];
  assign N2762 = N2761 | data_masked[1301];
  assign N2761 = N2760 | data_masked[1429];
  assign N2760 = N2759 | data_masked[1557];
  assign N2759 = N2758 | data_masked[1685];
  assign N2758 = N2757 | data_masked[1813];
  assign N2757 = N2756 | data_masked[1941];
  assign N2756 = N2755 | data_masked[2069];
  assign N2755 = N2754 | data_masked[2197];
  assign N2754 = N2753 | data_masked[2325];
  assign N2753 = N2752 | data_masked[2453];
  assign N2752 = N2751 | data_masked[2581];
  assign N2751 = N2750 | data_masked[2709];
  assign N2750 = N2749 | data_masked[2837];
  assign N2749 = N2748 | data_masked[2965];
  assign N2748 = N2747 | data_masked[3093];
  assign N2747 = N2746 | data_masked[3221];
  assign N2746 = N2745 | data_masked[3349];
  assign N2745 = N2744 | data_masked[3477];
  assign N2744 = N2743 | data_masked[3605];
  assign N2743 = N2742 | data_masked[3733];
  assign N2742 = N2741 | data_masked[3861];
  assign N2741 = N2740 | data_masked[3989];
  assign N2740 = N2739 | data_masked[4117];
  assign N2739 = N2738 | data_masked[4245];
  assign N2738 = N2737 | data_masked[4373];
  assign N2737 = N2736 | data_masked[4501];
  assign N2736 = N2735 | data_masked[4629];
  assign N2735 = N2734 | data_masked[4757];
  assign N2734 = N2733 | data_masked[4885];
  assign N2733 = N2732 | data_masked[5013];
  assign N2732 = N2731 | data_masked[5141];
  assign N2731 = N2730 | data_masked[5269];
  assign N2730 = N2729 | data_masked[5397];
  assign N2729 = N2728 | data_masked[5525];
  assign N2728 = N2727 | data_masked[5653];
  assign N2727 = N2726 | data_masked[5781];
  assign N2726 = N2725 | data_masked[5909];
  assign N2725 = N2724 | data_masked[6037];
  assign N2724 = N2723 | data_masked[6165];
  assign N2723 = N2722 | data_masked[6293];
  assign N2722 = N2721 | data_masked[6421];
  assign N2721 = N2720 | data_masked[6549];
  assign N2720 = N2719 | data_masked[6677];
  assign N2719 = N2718 | data_masked[6805];
  assign N2718 = N2717 | data_masked[6933];
  assign N2717 = N2716 | data_masked[7061];
  assign N2716 = N2715 | data_masked[7189];
  assign N2715 = N2714 | data_masked[7317];
  assign N2714 = N2713 | data_masked[7445];
  assign N2713 = N2712 | data_masked[7573];
  assign N2712 = N2711 | data_masked[7701];
  assign N2711 = N2710 | data_masked[7829];
  assign N2710 = N2709 | data_masked[7957];
  assign N2709 = N2708 | data_masked[8085];
  assign N2708 = N2707 | data_masked[8213];
  assign N2707 = N2706 | data_masked[8341];
  assign N2706 = N2705 | data_masked[8469];
  assign N2705 = N2704 | data_masked[8597];
  assign N2704 = N2703 | data_masked[8725];
  assign N2703 = N2702 | data_masked[8853];
  assign N2702 = N2701 | data_masked[8981];
  assign N2701 = N2700 | data_masked[9109];
  assign N2700 = N2699 | data_masked[9237];
  assign N2699 = N2698 | data_masked[9365];
  assign N2698 = N2697 | data_masked[9493];
  assign N2697 = N2696 | data_masked[9621];
  assign N2696 = N2695 | data_masked[9749];
  assign N2695 = N2694 | data_masked[9877];
  assign N2694 = N2693 | data_masked[10005];
  assign N2693 = N2692 | data_masked[10133];
  assign N2692 = N2691 | data_masked[10261];
  assign N2691 = N2690 | data_masked[10389];
  assign N2690 = N2689 | data_masked[10517];
  assign N2689 = N2688 | data_masked[10645];
  assign N2688 = N2687 | data_masked[10773];
  assign N2687 = N2686 | data_masked[10901];
  assign N2686 = N2685 | data_masked[11029];
  assign N2685 = N2684 | data_masked[11157];
  assign N2684 = N2683 | data_masked[11285];
  assign N2683 = N2682 | data_masked[11413];
  assign N2682 = N2681 | data_masked[11541];
  assign N2681 = N2680 | data_masked[11669];
  assign N2680 = N2679 | data_masked[11797];
  assign N2679 = N2678 | data_masked[11925];
  assign N2678 = N2677 | data_masked[12053];
  assign N2677 = N2676 | data_masked[12181];
  assign N2676 = N2675 | data_masked[12309];
  assign N2675 = N2674 | data_masked[12437];
  assign N2674 = N2673 | data_masked[12565];
  assign N2673 = N2672 | data_masked[12693];
  assign N2672 = N2671 | data_masked[12821];
  assign N2671 = N2670 | data_masked[12949];
  assign N2670 = N2669 | data_masked[13077];
  assign N2669 = N2668 | data_masked[13205];
  assign N2668 = N2667 | data_masked[13333];
  assign N2667 = N2666 | data_masked[13461];
  assign N2666 = N2665 | data_masked[13589];
  assign N2665 = N2664 | data_masked[13717];
  assign N2664 = N2663 | data_masked[13845];
  assign N2663 = N2662 | data_masked[13973];
  assign N2662 = N2661 | data_masked[14101];
  assign N2661 = N2660 | data_masked[14229];
  assign N2660 = N2659 | data_masked[14357];
  assign N2659 = N2658 | data_masked[14485];
  assign N2658 = N2657 | data_masked[14613];
  assign N2657 = N2656 | data_masked[14741];
  assign N2656 = N2655 | data_masked[14869];
  assign N2655 = N2654 | data_masked[14997];
  assign N2654 = N2653 | data_masked[15125];
  assign N2653 = N2652 | data_masked[15253];
  assign N2652 = N2651 | data_masked[15381];
  assign N2651 = N2650 | data_masked[15509];
  assign N2650 = N2649 | data_masked[15637];
  assign N2649 = N2648 | data_masked[15765];
  assign N2648 = N2647 | data_masked[15893];
  assign N2647 = N2646 | data_masked[16021];
  assign N2646 = data_masked[16277] | data_masked[16149];
  assign data_o[22] = N2897 | data_masked[22];
  assign N2897 = N2896 | data_masked[150];
  assign N2896 = N2895 | data_masked[278];
  assign N2895 = N2894 | data_masked[406];
  assign N2894 = N2893 | data_masked[534];
  assign N2893 = N2892 | data_masked[662];
  assign N2892 = N2891 | data_masked[790];
  assign N2891 = N2890 | data_masked[918];
  assign N2890 = N2889 | data_masked[1046];
  assign N2889 = N2888 | data_masked[1174];
  assign N2888 = N2887 | data_masked[1302];
  assign N2887 = N2886 | data_masked[1430];
  assign N2886 = N2885 | data_masked[1558];
  assign N2885 = N2884 | data_masked[1686];
  assign N2884 = N2883 | data_masked[1814];
  assign N2883 = N2882 | data_masked[1942];
  assign N2882 = N2881 | data_masked[2070];
  assign N2881 = N2880 | data_masked[2198];
  assign N2880 = N2879 | data_masked[2326];
  assign N2879 = N2878 | data_masked[2454];
  assign N2878 = N2877 | data_masked[2582];
  assign N2877 = N2876 | data_masked[2710];
  assign N2876 = N2875 | data_masked[2838];
  assign N2875 = N2874 | data_masked[2966];
  assign N2874 = N2873 | data_masked[3094];
  assign N2873 = N2872 | data_masked[3222];
  assign N2872 = N2871 | data_masked[3350];
  assign N2871 = N2870 | data_masked[3478];
  assign N2870 = N2869 | data_masked[3606];
  assign N2869 = N2868 | data_masked[3734];
  assign N2868 = N2867 | data_masked[3862];
  assign N2867 = N2866 | data_masked[3990];
  assign N2866 = N2865 | data_masked[4118];
  assign N2865 = N2864 | data_masked[4246];
  assign N2864 = N2863 | data_masked[4374];
  assign N2863 = N2862 | data_masked[4502];
  assign N2862 = N2861 | data_masked[4630];
  assign N2861 = N2860 | data_masked[4758];
  assign N2860 = N2859 | data_masked[4886];
  assign N2859 = N2858 | data_masked[5014];
  assign N2858 = N2857 | data_masked[5142];
  assign N2857 = N2856 | data_masked[5270];
  assign N2856 = N2855 | data_masked[5398];
  assign N2855 = N2854 | data_masked[5526];
  assign N2854 = N2853 | data_masked[5654];
  assign N2853 = N2852 | data_masked[5782];
  assign N2852 = N2851 | data_masked[5910];
  assign N2851 = N2850 | data_masked[6038];
  assign N2850 = N2849 | data_masked[6166];
  assign N2849 = N2848 | data_masked[6294];
  assign N2848 = N2847 | data_masked[6422];
  assign N2847 = N2846 | data_masked[6550];
  assign N2846 = N2845 | data_masked[6678];
  assign N2845 = N2844 | data_masked[6806];
  assign N2844 = N2843 | data_masked[6934];
  assign N2843 = N2842 | data_masked[7062];
  assign N2842 = N2841 | data_masked[7190];
  assign N2841 = N2840 | data_masked[7318];
  assign N2840 = N2839 | data_masked[7446];
  assign N2839 = N2838 | data_masked[7574];
  assign N2838 = N2837 | data_masked[7702];
  assign N2837 = N2836 | data_masked[7830];
  assign N2836 = N2835 | data_masked[7958];
  assign N2835 = N2834 | data_masked[8086];
  assign N2834 = N2833 | data_masked[8214];
  assign N2833 = N2832 | data_masked[8342];
  assign N2832 = N2831 | data_masked[8470];
  assign N2831 = N2830 | data_masked[8598];
  assign N2830 = N2829 | data_masked[8726];
  assign N2829 = N2828 | data_masked[8854];
  assign N2828 = N2827 | data_masked[8982];
  assign N2827 = N2826 | data_masked[9110];
  assign N2826 = N2825 | data_masked[9238];
  assign N2825 = N2824 | data_masked[9366];
  assign N2824 = N2823 | data_masked[9494];
  assign N2823 = N2822 | data_masked[9622];
  assign N2822 = N2821 | data_masked[9750];
  assign N2821 = N2820 | data_masked[9878];
  assign N2820 = N2819 | data_masked[10006];
  assign N2819 = N2818 | data_masked[10134];
  assign N2818 = N2817 | data_masked[10262];
  assign N2817 = N2816 | data_masked[10390];
  assign N2816 = N2815 | data_masked[10518];
  assign N2815 = N2814 | data_masked[10646];
  assign N2814 = N2813 | data_masked[10774];
  assign N2813 = N2812 | data_masked[10902];
  assign N2812 = N2811 | data_masked[11030];
  assign N2811 = N2810 | data_masked[11158];
  assign N2810 = N2809 | data_masked[11286];
  assign N2809 = N2808 | data_masked[11414];
  assign N2808 = N2807 | data_masked[11542];
  assign N2807 = N2806 | data_masked[11670];
  assign N2806 = N2805 | data_masked[11798];
  assign N2805 = N2804 | data_masked[11926];
  assign N2804 = N2803 | data_masked[12054];
  assign N2803 = N2802 | data_masked[12182];
  assign N2802 = N2801 | data_masked[12310];
  assign N2801 = N2800 | data_masked[12438];
  assign N2800 = N2799 | data_masked[12566];
  assign N2799 = N2798 | data_masked[12694];
  assign N2798 = N2797 | data_masked[12822];
  assign N2797 = N2796 | data_masked[12950];
  assign N2796 = N2795 | data_masked[13078];
  assign N2795 = N2794 | data_masked[13206];
  assign N2794 = N2793 | data_masked[13334];
  assign N2793 = N2792 | data_masked[13462];
  assign N2792 = N2791 | data_masked[13590];
  assign N2791 = N2790 | data_masked[13718];
  assign N2790 = N2789 | data_masked[13846];
  assign N2789 = N2788 | data_masked[13974];
  assign N2788 = N2787 | data_masked[14102];
  assign N2787 = N2786 | data_masked[14230];
  assign N2786 = N2785 | data_masked[14358];
  assign N2785 = N2784 | data_masked[14486];
  assign N2784 = N2783 | data_masked[14614];
  assign N2783 = N2782 | data_masked[14742];
  assign N2782 = N2781 | data_masked[14870];
  assign N2781 = N2780 | data_masked[14998];
  assign N2780 = N2779 | data_masked[15126];
  assign N2779 = N2778 | data_masked[15254];
  assign N2778 = N2777 | data_masked[15382];
  assign N2777 = N2776 | data_masked[15510];
  assign N2776 = N2775 | data_masked[15638];
  assign N2775 = N2774 | data_masked[15766];
  assign N2774 = N2773 | data_masked[15894];
  assign N2773 = N2772 | data_masked[16022];
  assign N2772 = data_masked[16278] | data_masked[16150];
  assign data_o[23] = N3023 | data_masked[23];
  assign N3023 = N3022 | data_masked[151];
  assign N3022 = N3021 | data_masked[279];
  assign N3021 = N3020 | data_masked[407];
  assign N3020 = N3019 | data_masked[535];
  assign N3019 = N3018 | data_masked[663];
  assign N3018 = N3017 | data_masked[791];
  assign N3017 = N3016 | data_masked[919];
  assign N3016 = N3015 | data_masked[1047];
  assign N3015 = N3014 | data_masked[1175];
  assign N3014 = N3013 | data_masked[1303];
  assign N3013 = N3012 | data_masked[1431];
  assign N3012 = N3011 | data_masked[1559];
  assign N3011 = N3010 | data_masked[1687];
  assign N3010 = N3009 | data_masked[1815];
  assign N3009 = N3008 | data_masked[1943];
  assign N3008 = N3007 | data_masked[2071];
  assign N3007 = N3006 | data_masked[2199];
  assign N3006 = N3005 | data_masked[2327];
  assign N3005 = N3004 | data_masked[2455];
  assign N3004 = N3003 | data_masked[2583];
  assign N3003 = N3002 | data_masked[2711];
  assign N3002 = N3001 | data_masked[2839];
  assign N3001 = N3000 | data_masked[2967];
  assign N3000 = N2999 | data_masked[3095];
  assign N2999 = N2998 | data_masked[3223];
  assign N2998 = N2997 | data_masked[3351];
  assign N2997 = N2996 | data_masked[3479];
  assign N2996 = N2995 | data_masked[3607];
  assign N2995 = N2994 | data_masked[3735];
  assign N2994 = N2993 | data_masked[3863];
  assign N2993 = N2992 | data_masked[3991];
  assign N2992 = N2991 | data_masked[4119];
  assign N2991 = N2990 | data_masked[4247];
  assign N2990 = N2989 | data_masked[4375];
  assign N2989 = N2988 | data_masked[4503];
  assign N2988 = N2987 | data_masked[4631];
  assign N2987 = N2986 | data_masked[4759];
  assign N2986 = N2985 | data_masked[4887];
  assign N2985 = N2984 | data_masked[5015];
  assign N2984 = N2983 | data_masked[5143];
  assign N2983 = N2982 | data_masked[5271];
  assign N2982 = N2981 | data_masked[5399];
  assign N2981 = N2980 | data_masked[5527];
  assign N2980 = N2979 | data_masked[5655];
  assign N2979 = N2978 | data_masked[5783];
  assign N2978 = N2977 | data_masked[5911];
  assign N2977 = N2976 | data_masked[6039];
  assign N2976 = N2975 | data_masked[6167];
  assign N2975 = N2974 | data_masked[6295];
  assign N2974 = N2973 | data_masked[6423];
  assign N2973 = N2972 | data_masked[6551];
  assign N2972 = N2971 | data_masked[6679];
  assign N2971 = N2970 | data_masked[6807];
  assign N2970 = N2969 | data_masked[6935];
  assign N2969 = N2968 | data_masked[7063];
  assign N2968 = N2967 | data_masked[7191];
  assign N2967 = N2966 | data_masked[7319];
  assign N2966 = N2965 | data_masked[7447];
  assign N2965 = N2964 | data_masked[7575];
  assign N2964 = N2963 | data_masked[7703];
  assign N2963 = N2962 | data_masked[7831];
  assign N2962 = N2961 | data_masked[7959];
  assign N2961 = N2960 | data_masked[8087];
  assign N2960 = N2959 | data_masked[8215];
  assign N2959 = N2958 | data_masked[8343];
  assign N2958 = N2957 | data_masked[8471];
  assign N2957 = N2956 | data_masked[8599];
  assign N2956 = N2955 | data_masked[8727];
  assign N2955 = N2954 | data_masked[8855];
  assign N2954 = N2953 | data_masked[8983];
  assign N2953 = N2952 | data_masked[9111];
  assign N2952 = N2951 | data_masked[9239];
  assign N2951 = N2950 | data_masked[9367];
  assign N2950 = N2949 | data_masked[9495];
  assign N2949 = N2948 | data_masked[9623];
  assign N2948 = N2947 | data_masked[9751];
  assign N2947 = N2946 | data_masked[9879];
  assign N2946 = N2945 | data_masked[10007];
  assign N2945 = N2944 | data_masked[10135];
  assign N2944 = N2943 | data_masked[10263];
  assign N2943 = N2942 | data_masked[10391];
  assign N2942 = N2941 | data_masked[10519];
  assign N2941 = N2940 | data_masked[10647];
  assign N2940 = N2939 | data_masked[10775];
  assign N2939 = N2938 | data_masked[10903];
  assign N2938 = N2937 | data_masked[11031];
  assign N2937 = N2936 | data_masked[11159];
  assign N2936 = N2935 | data_masked[11287];
  assign N2935 = N2934 | data_masked[11415];
  assign N2934 = N2933 | data_masked[11543];
  assign N2933 = N2932 | data_masked[11671];
  assign N2932 = N2931 | data_masked[11799];
  assign N2931 = N2930 | data_masked[11927];
  assign N2930 = N2929 | data_masked[12055];
  assign N2929 = N2928 | data_masked[12183];
  assign N2928 = N2927 | data_masked[12311];
  assign N2927 = N2926 | data_masked[12439];
  assign N2926 = N2925 | data_masked[12567];
  assign N2925 = N2924 | data_masked[12695];
  assign N2924 = N2923 | data_masked[12823];
  assign N2923 = N2922 | data_masked[12951];
  assign N2922 = N2921 | data_masked[13079];
  assign N2921 = N2920 | data_masked[13207];
  assign N2920 = N2919 | data_masked[13335];
  assign N2919 = N2918 | data_masked[13463];
  assign N2918 = N2917 | data_masked[13591];
  assign N2917 = N2916 | data_masked[13719];
  assign N2916 = N2915 | data_masked[13847];
  assign N2915 = N2914 | data_masked[13975];
  assign N2914 = N2913 | data_masked[14103];
  assign N2913 = N2912 | data_masked[14231];
  assign N2912 = N2911 | data_masked[14359];
  assign N2911 = N2910 | data_masked[14487];
  assign N2910 = N2909 | data_masked[14615];
  assign N2909 = N2908 | data_masked[14743];
  assign N2908 = N2907 | data_masked[14871];
  assign N2907 = N2906 | data_masked[14999];
  assign N2906 = N2905 | data_masked[15127];
  assign N2905 = N2904 | data_masked[15255];
  assign N2904 = N2903 | data_masked[15383];
  assign N2903 = N2902 | data_masked[15511];
  assign N2902 = N2901 | data_masked[15639];
  assign N2901 = N2900 | data_masked[15767];
  assign N2900 = N2899 | data_masked[15895];
  assign N2899 = N2898 | data_masked[16023];
  assign N2898 = data_masked[16279] | data_masked[16151];
  assign data_o[24] = N3149 | data_masked[24];
  assign N3149 = N3148 | data_masked[152];
  assign N3148 = N3147 | data_masked[280];
  assign N3147 = N3146 | data_masked[408];
  assign N3146 = N3145 | data_masked[536];
  assign N3145 = N3144 | data_masked[664];
  assign N3144 = N3143 | data_masked[792];
  assign N3143 = N3142 | data_masked[920];
  assign N3142 = N3141 | data_masked[1048];
  assign N3141 = N3140 | data_masked[1176];
  assign N3140 = N3139 | data_masked[1304];
  assign N3139 = N3138 | data_masked[1432];
  assign N3138 = N3137 | data_masked[1560];
  assign N3137 = N3136 | data_masked[1688];
  assign N3136 = N3135 | data_masked[1816];
  assign N3135 = N3134 | data_masked[1944];
  assign N3134 = N3133 | data_masked[2072];
  assign N3133 = N3132 | data_masked[2200];
  assign N3132 = N3131 | data_masked[2328];
  assign N3131 = N3130 | data_masked[2456];
  assign N3130 = N3129 | data_masked[2584];
  assign N3129 = N3128 | data_masked[2712];
  assign N3128 = N3127 | data_masked[2840];
  assign N3127 = N3126 | data_masked[2968];
  assign N3126 = N3125 | data_masked[3096];
  assign N3125 = N3124 | data_masked[3224];
  assign N3124 = N3123 | data_masked[3352];
  assign N3123 = N3122 | data_masked[3480];
  assign N3122 = N3121 | data_masked[3608];
  assign N3121 = N3120 | data_masked[3736];
  assign N3120 = N3119 | data_masked[3864];
  assign N3119 = N3118 | data_masked[3992];
  assign N3118 = N3117 | data_masked[4120];
  assign N3117 = N3116 | data_masked[4248];
  assign N3116 = N3115 | data_masked[4376];
  assign N3115 = N3114 | data_masked[4504];
  assign N3114 = N3113 | data_masked[4632];
  assign N3113 = N3112 | data_masked[4760];
  assign N3112 = N3111 | data_masked[4888];
  assign N3111 = N3110 | data_masked[5016];
  assign N3110 = N3109 | data_masked[5144];
  assign N3109 = N3108 | data_masked[5272];
  assign N3108 = N3107 | data_masked[5400];
  assign N3107 = N3106 | data_masked[5528];
  assign N3106 = N3105 | data_masked[5656];
  assign N3105 = N3104 | data_masked[5784];
  assign N3104 = N3103 | data_masked[5912];
  assign N3103 = N3102 | data_masked[6040];
  assign N3102 = N3101 | data_masked[6168];
  assign N3101 = N3100 | data_masked[6296];
  assign N3100 = N3099 | data_masked[6424];
  assign N3099 = N3098 | data_masked[6552];
  assign N3098 = N3097 | data_masked[6680];
  assign N3097 = N3096 | data_masked[6808];
  assign N3096 = N3095 | data_masked[6936];
  assign N3095 = N3094 | data_masked[7064];
  assign N3094 = N3093 | data_masked[7192];
  assign N3093 = N3092 | data_masked[7320];
  assign N3092 = N3091 | data_masked[7448];
  assign N3091 = N3090 | data_masked[7576];
  assign N3090 = N3089 | data_masked[7704];
  assign N3089 = N3088 | data_masked[7832];
  assign N3088 = N3087 | data_masked[7960];
  assign N3087 = N3086 | data_masked[8088];
  assign N3086 = N3085 | data_masked[8216];
  assign N3085 = N3084 | data_masked[8344];
  assign N3084 = N3083 | data_masked[8472];
  assign N3083 = N3082 | data_masked[8600];
  assign N3082 = N3081 | data_masked[8728];
  assign N3081 = N3080 | data_masked[8856];
  assign N3080 = N3079 | data_masked[8984];
  assign N3079 = N3078 | data_masked[9112];
  assign N3078 = N3077 | data_masked[9240];
  assign N3077 = N3076 | data_masked[9368];
  assign N3076 = N3075 | data_masked[9496];
  assign N3075 = N3074 | data_masked[9624];
  assign N3074 = N3073 | data_masked[9752];
  assign N3073 = N3072 | data_masked[9880];
  assign N3072 = N3071 | data_masked[10008];
  assign N3071 = N3070 | data_masked[10136];
  assign N3070 = N3069 | data_masked[10264];
  assign N3069 = N3068 | data_masked[10392];
  assign N3068 = N3067 | data_masked[10520];
  assign N3067 = N3066 | data_masked[10648];
  assign N3066 = N3065 | data_masked[10776];
  assign N3065 = N3064 | data_masked[10904];
  assign N3064 = N3063 | data_masked[11032];
  assign N3063 = N3062 | data_masked[11160];
  assign N3062 = N3061 | data_masked[11288];
  assign N3061 = N3060 | data_masked[11416];
  assign N3060 = N3059 | data_masked[11544];
  assign N3059 = N3058 | data_masked[11672];
  assign N3058 = N3057 | data_masked[11800];
  assign N3057 = N3056 | data_masked[11928];
  assign N3056 = N3055 | data_masked[12056];
  assign N3055 = N3054 | data_masked[12184];
  assign N3054 = N3053 | data_masked[12312];
  assign N3053 = N3052 | data_masked[12440];
  assign N3052 = N3051 | data_masked[12568];
  assign N3051 = N3050 | data_masked[12696];
  assign N3050 = N3049 | data_masked[12824];
  assign N3049 = N3048 | data_masked[12952];
  assign N3048 = N3047 | data_masked[13080];
  assign N3047 = N3046 | data_masked[13208];
  assign N3046 = N3045 | data_masked[13336];
  assign N3045 = N3044 | data_masked[13464];
  assign N3044 = N3043 | data_masked[13592];
  assign N3043 = N3042 | data_masked[13720];
  assign N3042 = N3041 | data_masked[13848];
  assign N3041 = N3040 | data_masked[13976];
  assign N3040 = N3039 | data_masked[14104];
  assign N3039 = N3038 | data_masked[14232];
  assign N3038 = N3037 | data_masked[14360];
  assign N3037 = N3036 | data_masked[14488];
  assign N3036 = N3035 | data_masked[14616];
  assign N3035 = N3034 | data_masked[14744];
  assign N3034 = N3033 | data_masked[14872];
  assign N3033 = N3032 | data_masked[15000];
  assign N3032 = N3031 | data_masked[15128];
  assign N3031 = N3030 | data_masked[15256];
  assign N3030 = N3029 | data_masked[15384];
  assign N3029 = N3028 | data_masked[15512];
  assign N3028 = N3027 | data_masked[15640];
  assign N3027 = N3026 | data_masked[15768];
  assign N3026 = N3025 | data_masked[15896];
  assign N3025 = N3024 | data_masked[16024];
  assign N3024 = data_masked[16280] | data_masked[16152];
  assign data_o[25] = N3275 | data_masked[25];
  assign N3275 = N3274 | data_masked[153];
  assign N3274 = N3273 | data_masked[281];
  assign N3273 = N3272 | data_masked[409];
  assign N3272 = N3271 | data_masked[537];
  assign N3271 = N3270 | data_masked[665];
  assign N3270 = N3269 | data_masked[793];
  assign N3269 = N3268 | data_masked[921];
  assign N3268 = N3267 | data_masked[1049];
  assign N3267 = N3266 | data_masked[1177];
  assign N3266 = N3265 | data_masked[1305];
  assign N3265 = N3264 | data_masked[1433];
  assign N3264 = N3263 | data_masked[1561];
  assign N3263 = N3262 | data_masked[1689];
  assign N3262 = N3261 | data_masked[1817];
  assign N3261 = N3260 | data_masked[1945];
  assign N3260 = N3259 | data_masked[2073];
  assign N3259 = N3258 | data_masked[2201];
  assign N3258 = N3257 | data_masked[2329];
  assign N3257 = N3256 | data_masked[2457];
  assign N3256 = N3255 | data_masked[2585];
  assign N3255 = N3254 | data_masked[2713];
  assign N3254 = N3253 | data_masked[2841];
  assign N3253 = N3252 | data_masked[2969];
  assign N3252 = N3251 | data_masked[3097];
  assign N3251 = N3250 | data_masked[3225];
  assign N3250 = N3249 | data_masked[3353];
  assign N3249 = N3248 | data_masked[3481];
  assign N3248 = N3247 | data_masked[3609];
  assign N3247 = N3246 | data_masked[3737];
  assign N3246 = N3245 | data_masked[3865];
  assign N3245 = N3244 | data_masked[3993];
  assign N3244 = N3243 | data_masked[4121];
  assign N3243 = N3242 | data_masked[4249];
  assign N3242 = N3241 | data_masked[4377];
  assign N3241 = N3240 | data_masked[4505];
  assign N3240 = N3239 | data_masked[4633];
  assign N3239 = N3238 | data_masked[4761];
  assign N3238 = N3237 | data_masked[4889];
  assign N3237 = N3236 | data_masked[5017];
  assign N3236 = N3235 | data_masked[5145];
  assign N3235 = N3234 | data_masked[5273];
  assign N3234 = N3233 | data_masked[5401];
  assign N3233 = N3232 | data_masked[5529];
  assign N3232 = N3231 | data_masked[5657];
  assign N3231 = N3230 | data_masked[5785];
  assign N3230 = N3229 | data_masked[5913];
  assign N3229 = N3228 | data_masked[6041];
  assign N3228 = N3227 | data_masked[6169];
  assign N3227 = N3226 | data_masked[6297];
  assign N3226 = N3225 | data_masked[6425];
  assign N3225 = N3224 | data_masked[6553];
  assign N3224 = N3223 | data_masked[6681];
  assign N3223 = N3222 | data_masked[6809];
  assign N3222 = N3221 | data_masked[6937];
  assign N3221 = N3220 | data_masked[7065];
  assign N3220 = N3219 | data_masked[7193];
  assign N3219 = N3218 | data_masked[7321];
  assign N3218 = N3217 | data_masked[7449];
  assign N3217 = N3216 | data_masked[7577];
  assign N3216 = N3215 | data_masked[7705];
  assign N3215 = N3214 | data_masked[7833];
  assign N3214 = N3213 | data_masked[7961];
  assign N3213 = N3212 | data_masked[8089];
  assign N3212 = N3211 | data_masked[8217];
  assign N3211 = N3210 | data_masked[8345];
  assign N3210 = N3209 | data_masked[8473];
  assign N3209 = N3208 | data_masked[8601];
  assign N3208 = N3207 | data_masked[8729];
  assign N3207 = N3206 | data_masked[8857];
  assign N3206 = N3205 | data_masked[8985];
  assign N3205 = N3204 | data_masked[9113];
  assign N3204 = N3203 | data_masked[9241];
  assign N3203 = N3202 | data_masked[9369];
  assign N3202 = N3201 | data_masked[9497];
  assign N3201 = N3200 | data_masked[9625];
  assign N3200 = N3199 | data_masked[9753];
  assign N3199 = N3198 | data_masked[9881];
  assign N3198 = N3197 | data_masked[10009];
  assign N3197 = N3196 | data_masked[10137];
  assign N3196 = N3195 | data_masked[10265];
  assign N3195 = N3194 | data_masked[10393];
  assign N3194 = N3193 | data_masked[10521];
  assign N3193 = N3192 | data_masked[10649];
  assign N3192 = N3191 | data_masked[10777];
  assign N3191 = N3190 | data_masked[10905];
  assign N3190 = N3189 | data_masked[11033];
  assign N3189 = N3188 | data_masked[11161];
  assign N3188 = N3187 | data_masked[11289];
  assign N3187 = N3186 | data_masked[11417];
  assign N3186 = N3185 | data_masked[11545];
  assign N3185 = N3184 | data_masked[11673];
  assign N3184 = N3183 | data_masked[11801];
  assign N3183 = N3182 | data_masked[11929];
  assign N3182 = N3181 | data_masked[12057];
  assign N3181 = N3180 | data_masked[12185];
  assign N3180 = N3179 | data_masked[12313];
  assign N3179 = N3178 | data_masked[12441];
  assign N3178 = N3177 | data_masked[12569];
  assign N3177 = N3176 | data_masked[12697];
  assign N3176 = N3175 | data_masked[12825];
  assign N3175 = N3174 | data_masked[12953];
  assign N3174 = N3173 | data_masked[13081];
  assign N3173 = N3172 | data_masked[13209];
  assign N3172 = N3171 | data_masked[13337];
  assign N3171 = N3170 | data_masked[13465];
  assign N3170 = N3169 | data_masked[13593];
  assign N3169 = N3168 | data_masked[13721];
  assign N3168 = N3167 | data_masked[13849];
  assign N3167 = N3166 | data_masked[13977];
  assign N3166 = N3165 | data_masked[14105];
  assign N3165 = N3164 | data_masked[14233];
  assign N3164 = N3163 | data_masked[14361];
  assign N3163 = N3162 | data_masked[14489];
  assign N3162 = N3161 | data_masked[14617];
  assign N3161 = N3160 | data_masked[14745];
  assign N3160 = N3159 | data_masked[14873];
  assign N3159 = N3158 | data_masked[15001];
  assign N3158 = N3157 | data_masked[15129];
  assign N3157 = N3156 | data_masked[15257];
  assign N3156 = N3155 | data_masked[15385];
  assign N3155 = N3154 | data_masked[15513];
  assign N3154 = N3153 | data_masked[15641];
  assign N3153 = N3152 | data_masked[15769];
  assign N3152 = N3151 | data_masked[15897];
  assign N3151 = N3150 | data_masked[16025];
  assign N3150 = data_masked[16281] | data_masked[16153];
  assign data_o[26] = N3401 | data_masked[26];
  assign N3401 = N3400 | data_masked[154];
  assign N3400 = N3399 | data_masked[282];
  assign N3399 = N3398 | data_masked[410];
  assign N3398 = N3397 | data_masked[538];
  assign N3397 = N3396 | data_masked[666];
  assign N3396 = N3395 | data_masked[794];
  assign N3395 = N3394 | data_masked[922];
  assign N3394 = N3393 | data_masked[1050];
  assign N3393 = N3392 | data_masked[1178];
  assign N3392 = N3391 | data_masked[1306];
  assign N3391 = N3390 | data_masked[1434];
  assign N3390 = N3389 | data_masked[1562];
  assign N3389 = N3388 | data_masked[1690];
  assign N3388 = N3387 | data_masked[1818];
  assign N3387 = N3386 | data_masked[1946];
  assign N3386 = N3385 | data_masked[2074];
  assign N3385 = N3384 | data_masked[2202];
  assign N3384 = N3383 | data_masked[2330];
  assign N3383 = N3382 | data_masked[2458];
  assign N3382 = N3381 | data_masked[2586];
  assign N3381 = N3380 | data_masked[2714];
  assign N3380 = N3379 | data_masked[2842];
  assign N3379 = N3378 | data_masked[2970];
  assign N3378 = N3377 | data_masked[3098];
  assign N3377 = N3376 | data_masked[3226];
  assign N3376 = N3375 | data_masked[3354];
  assign N3375 = N3374 | data_masked[3482];
  assign N3374 = N3373 | data_masked[3610];
  assign N3373 = N3372 | data_masked[3738];
  assign N3372 = N3371 | data_masked[3866];
  assign N3371 = N3370 | data_masked[3994];
  assign N3370 = N3369 | data_masked[4122];
  assign N3369 = N3368 | data_masked[4250];
  assign N3368 = N3367 | data_masked[4378];
  assign N3367 = N3366 | data_masked[4506];
  assign N3366 = N3365 | data_masked[4634];
  assign N3365 = N3364 | data_masked[4762];
  assign N3364 = N3363 | data_masked[4890];
  assign N3363 = N3362 | data_masked[5018];
  assign N3362 = N3361 | data_masked[5146];
  assign N3361 = N3360 | data_masked[5274];
  assign N3360 = N3359 | data_masked[5402];
  assign N3359 = N3358 | data_masked[5530];
  assign N3358 = N3357 | data_masked[5658];
  assign N3357 = N3356 | data_masked[5786];
  assign N3356 = N3355 | data_masked[5914];
  assign N3355 = N3354 | data_masked[6042];
  assign N3354 = N3353 | data_masked[6170];
  assign N3353 = N3352 | data_masked[6298];
  assign N3352 = N3351 | data_masked[6426];
  assign N3351 = N3350 | data_masked[6554];
  assign N3350 = N3349 | data_masked[6682];
  assign N3349 = N3348 | data_masked[6810];
  assign N3348 = N3347 | data_masked[6938];
  assign N3347 = N3346 | data_masked[7066];
  assign N3346 = N3345 | data_masked[7194];
  assign N3345 = N3344 | data_masked[7322];
  assign N3344 = N3343 | data_masked[7450];
  assign N3343 = N3342 | data_masked[7578];
  assign N3342 = N3341 | data_masked[7706];
  assign N3341 = N3340 | data_masked[7834];
  assign N3340 = N3339 | data_masked[7962];
  assign N3339 = N3338 | data_masked[8090];
  assign N3338 = N3337 | data_masked[8218];
  assign N3337 = N3336 | data_masked[8346];
  assign N3336 = N3335 | data_masked[8474];
  assign N3335 = N3334 | data_masked[8602];
  assign N3334 = N3333 | data_masked[8730];
  assign N3333 = N3332 | data_masked[8858];
  assign N3332 = N3331 | data_masked[8986];
  assign N3331 = N3330 | data_masked[9114];
  assign N3330 = N3329 | data_masked[9242];
  assign N3329 = N3328 | data_masked[9370];
  assign N3328 = N3327 | data_masked[9498];
  assign N3327 = N3326 | data_masked[9626];
  assign N3326 = N3325 | data_masked[9754];
  assign N3325 = N3324 | data_masked[9882];
  assign N3324 = N3323 | data_masked[10010];
  assign N3323 = N3322 | data_masked[10138];
  assign N3322 = N3321 | data_masked[10266];
  assign N3321 = N3320 | data_masked[10394];
  assign N3320 = N3319 | data_masked[10522];
  assign N3319 = N3318 | data_masked[10650];
  assign N3318 = N3317 | data_masked[10778];
  assign N3317 = N3316 | data_masked[10906];
  assign N3316 = N3315 | data_masked[11034];
  assign N3315 = N3314 | data_masked[11162];
  assign N3314 = N3313 | data_masked[11290];
  assign N3313 = N3312 | data_masked[11418];
  assign N3312 = N3311 | data_masked[11546];
  assign N3311 = N3310 | data_masked[11674];
  assign N3310 = N3309 | data_masked[11802];
  assign N3309 = N3308 | data_masked[11930];
  assign N3308 = N3307 | data_masked[12058];
  assign N3307 = N3306 | data_masked[12186];
  assign N3306 = N3305 | data_masked[12314];
  assign N3305 = N3304 | data_masked[12442];
  assign N3304 = N3303 | data_masked[12570];
  assign N3303 = N3302 | data_masked[12698];
  assign N3302 = N3301 | data_masked[12826];
  assign N3301 = N3300 | data_masked[12954];
  assign N3300 = N3299 | data_masked[13082];
  assign N3299 = N3298 | data_masked[13210];
  assign N3298 = N3297 | data_masked[13338];
  assign N3297 = N3296 | data_masked[13466];
  assign N3296 = N3295 | data_masked[13594];
  assign N3295 = N3294 | data_masked[13722];
  assign N3294 = N3293 | data_masked[13850];
  assign N3293 = N3292 | data_masked[13978];
  assign N3292 = N3291 | data_masked[14106];
  assign N3291 = N3290 | data_masked[14234];
  assign N3290 = N3289 | data_masked[14362];
  assign N3289 = N3288 | data_masked[14490];
  assign N3288 = N3287 | data_masked[14618];
  assign N3287 = N3286 | data_masked[14746];
  assign N3286 = N3285 | data_masked[14874];
  assign N3285 = N3284 | data_masked[15002];
  assign N3284 = N3283 | data_masked[15130];
  assign N3283 = N3282 | data_masked[15258];
  assign N3282 = N3281 | data_masked[15386];
  assign N3281 = N3280 | data_masked[15514];
  assign N3280 = N3279 | data_masked[15642];
  assign N3279 = N3278 | data_masked[15770];
  assign N3278 = N3277 | data_masked[15898];
  assign N3277 = N3276 | data_masked[16026];
  assign N3276 = data_masked[16282] | data_masked[16154];
  assign data_o[27] = N3527 | data_masked[27];
  assign N3527 = N3526 | data_masked[155];
  assign N3526 = N3525 | data_masked[283];
  assign N3525 = N3524 | data_masked[411];
  assign N3524 = N3523 | data_masked[539];
  assign N3523 = N3522 | data_masked[667];
  assign N3522 = N3521 | data_masked[795];
  assign N3521 = N3520 | data_masked[923];
  assign N3520 = N3519 | data_masked[1051];
  assign N3519 = N3518 | data_masked[1179];
  assign N3518 = N3517 | data_masked[1307];
  assign N3517 = N3516 | data_masked[1435];
  assign N3516 = N3515 | data_masked[1563];
  assign N3515 = N3514 | data_masked[1691];
  assign N3514 = N3513 | data_masked[1819];
  assign N3513 = N3512 | data_masked[1947];
  assign N3512 = N3511 | data_masked[2075];
  assign N3511 = N3510 | data_masked[2203];
  assign N3510 = N3509 | data_masked[2331];
  assign N3509 = N3508 | data_masked[2459];
  assign N3508 = N3507 | data_masked[2587];
  assign N3507 = N3506 | data_masked[2715];
  assign N3506 = N3505 | data_masked[2843];
  assign N3505 = N3504 | data_masked[2971];
  assign N3504 = N3503 | data_masked[3099];
  assign N3503 = N3502 | data_masked[3227];
  assign N3502 = N3501 | data_masked[3355];
  assign N3501 = N3500 | data_masked[3483];
  assign N3500 = N3499 | data_masked[3611];
  assign N3499 = N3498 | data_masked[3739];
  assign N3498 = N3497 | data_masked[3867];
  assign N3497 = N3496 | data_masked[3995];
  assign N3496 = N3495 | data_masked[4123];
  assign N3495 = N3494 | data_masked[4251];
  assign N3494 = N3493 | data_masked[4379];
  assign N3493 = N3492 | data_masked[4507];
  assign N3492 = N3491 | data_masked[4635];
  assign N3491 = N3490 | data_masked[4763];
  assign N3490 = N3489 | data_masked[4891];
  assign N3489 = N3488 | data_masked[5019];
  assign N3488 = N3487 | data_masked[5147];
  assign N3487 = N3486 | data_masked[5275];
  assign N3486 = N3485 | data_masked[5403];
  assign N3485 = N3484 | data_masked[5531];
  assign N3484 = N3483 | data_masked[5659];
  assign N3483 = N3482 | data_masked[5787];
  assign N3482 = N3481 | data_masked[5915];
  assign N3481 = N3480 | data_masked[6043];
  assign N3480 = N3479 | data_masked[6171];
  assign N3479 = N3478 | data_masked[6299];
  assign N3478 = N3477 | data_masked[6427];
  assign N3477 = N3476 | data_masked[6555];
  assign N3476 = N3475 | data_masked[6683];
  assign N3475 = N3474 | data_masked[6811];
  assign N3474 = N3473 | data_masked[6939];
  assign N3473 = N3472 | data_masked[7067];
  assign N3472 = N3471 | data_masked[7195];
  assign N3471 = N3470 | data_masked[7323];
  assign N3470 = N3469 | data_masked[7451];
  assign N3469 = N3468 | data_masked[7579];
  assign N3468 = N3467 | data_masked[7707];
  assign N3467 = N3466 | data_masked[7835];
  assign N3466 = N3465 | data_masked[7963];
  assign N3465 = N3464 | data_masked[8091];
  assign N3464 = N3463 | data_masked[8219];
  assign N3463 = N3462 | data_masked[8347];
  assign N3462 = N3461 | data_masked[8475];
  assign N3461 = N3460 | data_masked[8603];
  assign N3460 = N3459 | data_masked[8731];
  assign N3459 = N3458 | data_masked[8859];
  assign N3458 = N3457 | data_masked[8987];
  assign N3457 = N3456 | data_masked[9115];
  assign N3456 = N3455 | data_masked[9243];
  assign N3455 = N3454 | data_masked[9371];
  assign N3454 = N3453 | data_masked[9499];
  assign N3453 = N3452 | data_masked[9627];
  assign N3452 = N3451 | data_masked[9755];
  assign N3451 = N3450 | data_masked[9883];
  assign N3450 = N3449 | data_masked[10011];
  assign N3449 = N3448 | data_masked[10139];
  assign N3448 = N3447 | data_masked[10267];
  assign N3447 = N3446 | data_masked[10395];
  assign N3446 = N3445 | data_masked[10523];
  assign N3445 = N3444 | data_masked[10651];
  assign N3444 = N3443 | data_masked[10779];
  assign N3443 = N3442 | data_masked[10907];
  assign N3442 = N3441 | data_masked[11035];
  assign N3441 = N3440 | data_masked[11163];
  assign N3440 = N3439 | data_masked[11291];
  assign N3439 = N3438 | data_masked[11419];
  assign N3438 = N3437 | data_masked[11547];
  assign N3437 = N3436 | data_masked[11675];
  assign N3436 = N3435 | data_masked[11803];
  assign N3435 = N3434 | data_masked[11931];
  assign N3434 = N3433 | data_masked[12059];
  assign N3433 = N3432 | data_masked[12187];
  assign N3432 = N3431 | data_masked[12315];
  assign N3431 = N3430 | data_masked[12443];
  assign N3430 = N3429 | data_masked[12571];
  assign N3429 = N3428 | data_masked[12699];
  assign N3428 = N3427 | data_masked[12827];
  assign N3427 = N3426 | data_masked[12955];
  assign N3426 = N3425 | data_masked[13083];
  assign N3425 = N3424 | data_masked[13211];
  assign N3424 = N3423 | data_masked[13339];
  assign N3423 = N3422 | data_masked[13467];
  assign N3422 = N3421 | data_masked[13595];
  assign N3421 = N3420 | data_masked[13723];
  assign N3420 = N3419 | data_masked[13851];
  assign N3419 = N3418 | data_masked[13979];
  assign N3418 = N3417 | data_masked[14107];
  assign N3417 = N3416 | data_masked[14235];
  assign N3416 = N3415 | data_masked[14363];
  assign N3415 = N3414 | data_masked[14491];
  assign N3414 = N3413 | data_masked[14619];
  assign N3413 = N3412 | data_masked[14747];
  assign N3412 = N3411 | data_masked[14875];
  assign N3411 = N3410 | data_masked[15003];
  assign N3410 = N3409 | data_masked[15131];
  assign N3409 = N3408 | data_masked[15259];
  assign N3408 = N3407 | data_masked[15387];
  assign N3407 = N3406 | data_masked[15515];
  assign N3406 = N3405 | data_masked[15643];
  assign N3405 = N3404 | data_masked[15771];
  assign N3404 = N3403 | data_masked[15899];
  assign N3403 = N3402 | data_masked[16027];
  assign N3402 = data_masked[16283] | data_masked[16155];
  assign data_o[28] = N3653 | data_masked[28];
  assign N3653 = N3652 | data_masked[156];
  assign N3652 = N3651 | data_masked[284];
  assign N3651 = N3650 | data_masked[412];
  assign N3650 = N3649 | data_masked[540];
  assign N3649 = N3648 | data_masked[668];
  assign N3648 = N3647 | data_masked[796];
  assign N3647 = N3646 | data_masked[924];
  assign N3646 = N3645 | data_masked[1052];
  assign N3645 = N3644 | data_masked[1180];
  assign N3644 = N3643 | data_masked[1308];
  assign N3643 = N3642 | data_masked[1436];
  assign N3642 = N3641 | data_masked[1564];
  assign N3641 = N3640 | data_masked[1692];
  assign N3640 = N3639 | data_masked[1820];
  assign N3639 = N3638 | data_masked[1948];
  assign N3638 = N3637 | data_masked[2076];
  assign N3637 = N3636 | data_masked[2204];
  assign N3636 = N3635 | data_masked[2332];
  assign N3635 = N3634 | data_masked[2460];
  assign N3634 = N3633 | data_masked[2588];
  assign N3633 = N3632 | data_masked[2716];
  assign N3632 = N3631 | data_masked[2844];
  assign N3631 = N3630 | data_masked[2972];
  assign N3630 = N3629 | data_masked[3100];
  assign N3629 = N3628 | data_masked[3228];
  assign N3628 = N3627 | data_masked[3356];
  assign N3627 = N3626 | data_masked[3484];
  assign N3626 = N3625 | data_masked[3612];
  assign N3625 = N3624 | data_masked[3740];
  assign N3624 = N3623 | data_masked[3868];
  assign N3623 = N3622 | data_masked[3996];
  assign N3622 = N3621 | data_masked[4124];
  assign N3621 = N3620 | data_masked[4252];
  assign N3620 = N3619 | data_masked[4380];
  assign N3619 = N3618 | data_masked[4508];
  assign N3618 = N3617 | data_masked[4636];
  assign N3617 = N3616 | data_masked[4764];
  assign N3616 = N3615 | data_masked[4892];
  assign N3615 = N3614 | data_masked[5020];
  assign N3614 = N3613 | data_masked[5148];
  assign N3613 = N3612 | data_masked[5276];
  assign N3612 = N3611 | data_masked[5404];
  assign N3611 = N3610 | data_masked[5532];
  assign N3610 = N3609 | data_masked[5660];
  assign N3609 = N3608 | data_masked[5788];
  assign N3608 = N3607 | data_masked[5916];
  assign N3607 = N3606 | data_masked[6044];
  assign N3606 = N3605 | data_masked[6172];
  assign N3605 = N3604 | data_masked[6300];
  assign N3604 = N3603 | data_masked[6428];
  assign N3603 = N3602 | data_masked[6556];
  assign N3602 = N3601 | data_masked[6684];
  assign N3601 = N3600 | data_masked[6812];
  assign N3600 = N3599 | data_masked[6940];
  assign N3599 = N3598 | data_masked[7068];
  assign N3598 = N3597 | data_masked[7196];
  assign N3597 = N3596 | data_masked[7324];
  assign N3596 = N3595 | data_masked[7452];
  assign N3595 = N3594 | data_masked[7580];
  assign N3594 = N3593 | data_masked[7708];
  assign N3593 = N3592 | data_masked[7836];
  assign N3592 = N3591 | data_masked[7964];
  assign N3591 = N3590 | data_masked[8092];
  assign N3590 = N3589 | data_masked[8220];
  assign N3589 = N3588 | data_masked[8348];
  assign N3588 = N3587 | data_masked[8476];
  assign N3587 = N3586 | data_masked[8604];
  assign N3586 = N3585 | data_masked[8732];
  assign N3585 = N3584 | data_masked[8860];
  assign N3584 = N3583 | data_masked[8988];
  assign N3583 = N3582 | data_masked[9116];
  assign N3582 = N3581 | data_masked[9244];
  assign N3581 = N3580 | data_masked[9372];
  assign N3580 = N3579 | data_masked[9500];
  assign N3579 = N3578 | data_masked[9628];
  assign N3578 = N3577 | data_masked[9756];
  assign N3577 = N3576 | data_masked[9884];
  assign N3576 = N3575 | data_masked[10012];
  assign N3575 = N3574 | data_masked[10140];
  assign N3574 = N3573 | data_masked[10268];
  assign N3573 = N3572 | data_masked[10396];
  assign N3572 = N3571 | data_masked[10524];
  assign N3571 = N3570 | data_masked[10652];
  assign N3570 = N3569 | data_masked[10780];
  assign N3569 = N3568 | data_masked[10908];
  assign N3568 = N3567 | data_masked[11036];
  assign N3567 = N3566 | data_masked[11164];
  assign N3566 = N3565 | data_masked[11292];
  assign N3565 = N3564 | data_masked[11420];
  assign N3564 = N3563 | data_masked[11548];
  assign N3563 = N3562 | data_masked[11676];
  assign N3562 = N3561 | data_masked[11804];
  assign N3561 = N3560 | data_masked[11932];
  assign N3560 = N3559 | data_masked[12060];
  assign N3559 = N3558 | data_masked[12188];
  assign N3558 = N3557 | data_masked[12316];
  assign N3557 = N3556 | data_masked[12444];
  assign N3556 = N3555 | data_masked[12572];
  assign N3555 = N3554 | data_masked[12700];
  assign N3554 = N3553 | data_masked[12828];
  assign N3553 = N3552 | data_masked[12956];
  assign N3552 = N3551 | data_masked[13084];
  assign N3551 = N3550 | data_masked[13212];
  assign N3550 = N3549 | data_masked[13340];
  assign N3549 = N3548 | data_masked[13468];
  assign N3548 = N3547 | data_masked[13596];
  assign N3547 = N3546 | data_masked[13724];
  assign N3546 = N3545 | data_masked[13852];
  assign N3545 = N3544 | data_masked[13980];
  assign N3544 = N3543 | data_masked[14108];
  assign N3543 = N3542 | data_masked[14236];
  assign N3542 = N3541 | data_masked[14364];
  assign N3541 = N3540 | data_masked[14492];
  assign N3540 = N3539 | data_masked[14620];
  assign N3539 = N3538 | data_masked[14748];
  assign N3538 = N3537 | data_masked[14876];
  assign N3537 = N3536 | data_masked[15004];
  assign N3536 = N3535 | data_masked[15132];
  assign N3535 = N3534 | data_masked[15260];
  assign N3534 = N3533 | data_masked[15388];
  assign N3533 = N3532 | data_masked[15516];
  assign N3532 = N3531 | data_masked[15644];
  assign N3531 = N3530 | data_masked[15772];
  assign N3530 = N3529 | data_masked[15900];
  assign N3529 = N3528 | data_masked[16028];
  assign N3528 = data_masked[16284] | data_masked[16156];
  assign data_o[29] = N3779 | data_masked[29];
  assign N3779 = N3778 | data_masked[157];
  assign N3778 = N3777 | data_masked[285];
  assign N3777 = N3776 | data_masked[413];
  assign N3776 = N3775 | data_masked[541];
  assign N3775 = N3774 | data_masked[669];
  assign N3774 = N3773 | data_masked[797];
  assign N3773 = N3772 | data_masked[925];
  assign N3772 = N3771 | data_masked[1053];
  assign N3771 = N3770 | data_masked[1181];
  assign N3770 = N3769 | data_masked[1309];
  assign N3769 = N3768 | data_masked[1437];
  assign N3768 = N3767 | data_masked[1565];
  assign N3767 = N3766 | data_masked[1693];
  assign N3766 = N3765 | data_masked[1821];
  assign N3765 = N3764 | data_masked[1949];
  assign N3764 = N3763 | data_masked[2077];
  assign N3763 = N3762 | data_masked[2205];
  assign N3762 = N3761 | data_masked[2333];
  assign N3761 = N3760 | data_masked[2461];
  assign N3760 = N3759 | data_masked[2589];
  assign N3759 = N3758 | data_masked[2717];
  assign N3758 = N3757 | data_masked[2845];
  assign N3757 = N3756 | data_masked[2973];
  assign N3756 = N3755 | data_masked[3101];
  assign N3755 = N3754 | data_masked[3229];
  assign N3754 = N3753 | data_masked[3357];
  assign N3753 = N3752 | data_masked[3485];
  assign N3752 = N3751 | data_masked[3613];
  assign N3751 = N3750 | data_masked[3741];
  assign N3750 = N3749 | data_masked[3869];
  assign N3749 = N3748 | data_masked[3997];
  assign N3748 = N3747 | data_masked[4125];
  assign N3747 = N3746 | data_masked[4253];
  assign N3746 = N3745 | data_masked[4381];
  assign N3745 = N3744 | data_masked[4509];
  assign N3744 = N3743 | data_masked[4637];
  assign N3743 = N3742 | data_masked[4765];
  assign N3742 = N3741 | data_masked[4893];
  assign N3741 = N3740 | data_masked[5021];
  assign N3740 = N3739 | data_masked[5149];
  assign N3739 = N3738 | data_masked[5277];
  assign N3738 = N3737 | data_masked[5405];
  assign N3737 = N3736 | data_masked[5533];
  assign N3736 = N3735 | data_masked[5661];
  assign N3735 = N3734 | data_masked[5789];
  assign N3734 = N3733 | data_masked[5917];
  assign N3733 = N3732 | data_masked[6045];
  assign N3732 = N3731 | data_masked[6173];
  assign N3731 = N3730 | data_masked[6301];
  assign N3730 = N3729 | data_masked[6429];
  assign N3729 = N3728 | data_masked[6557];
  assign N3728 = N3727 | data_masked[6685];
  assign N3727 = N3726 | data_masked[6813];
  assign N3726 = N3725 | data_masked[6941];
  assign N3725 = N3724 | data_masked[7069];
  assign N3724 = N3723 | data_masked[7197];
  assign N3723 = N3722 | data_masked[7325];
  assign N3722 = N3721 | data_masked[7453];
  assign N3721 = N3720 | data_masked[7581];
  assign N3720 = N3719 | data_masked[7709];
  assign N3719 = N3718 | data_masked[7837];
  assign N3718 = N3717 | data_masked[7965];
  assign N3717 = N3716 | data_masked[8093];
  assign N3716 = N3715 | data_masked[8221];
  assign N3715 = N3714 | data_masked[8349];
  assign N3714 = N3713 | data_masked[8477];
  assign N3713 = N3712 | data_masked[8605];
  assign N3712 = N3711 | data_masked[8733];
  assign N3711 = N3710 | data_masked[8861];
  assign N3710 = N3709 | data_masked[8989];
  assign N3709 = N3708 | data_masked[9117];
  assign N3708 = N3707 | data_masked[9245];
  assign N3707 = N3706 | data_masked[9373];
  assign N3706 = N3705 | data_masked[9501];
  assign N3705 = N3704 | data_masked[9629];
  assign N3704 = N3703 | data_masked[9757];
  assign N3703 = N3702 | data_masked[9885];
  assign N3702 = N3701 | data_masked[10013];
  assign N3701 = N3700 | data_masked[10141];
  assign N3700 = N3699 | data_masked[10269];
  assign N3699 = N3698 | data_masked[10397];
  assign N3698 = N3697 | data_masked[10525];
  assign N3697 = N3696 | data_masked[10653];
  assign N3696 = N3695 | data_masked[10781];
  assign N3695 = N3694 | data_masked[10909];
  assign N3694 = N3693 | data_masked[11037];
  assign N3693 = N3692 | data_masked[11165];
  assign N3692 = N3691 | data_masked[11293];
  assign N3691 = N3690 | data_masked[11421];
  assign N3690 = N3689 | data_masked[11549];
  assign N3689 = N3688 | data_masked[11677];
  assign N3688 = N3687 | data_masked[11805];
  assign N3687 = N3686 | data_masked[11933];
  assign N3686 = N3685 | data_masked[12061];
  assign N3685 = N3684 | data_masked[12189];
  assign N3684 = N3683 | data_masked[12317];
  assign N3683 = N3682 | data_masked[12445];
  assign N3682 = N3681 | data_masked[12573];
  assign N3681 = N3680 | data_masked[12701];
  assign N3680 = N3679 | data_masked[12829];
  assign N3679 = N3678 | data_masked[12957];
  assign N3678 = N3677 | data_masked[13085];
  assign N3677 = N3676 | data_masked[13213];
  assign N3676 = N3675 | data_masked[13341];
  assign N3675 = N3674 | data_masked[13469];
  assign N3674 = N3673 | data_masked[13597];
  assign N3673 = N3672 | data_masked[13725];
  assign N3672 = N3671 | data_masked[13853];
  assign N3671 = N3670 | data_masked[13981];
  assign N3670 = N3669 | data_masked[14109];
  assign N3669 = N3668 | data_masked[14237];
  assign N3668 = N3667 | data_masked[14365];
  assign N3667 = N3666 | data_masked[14493];
  assign N3666 = N3665 | data_masked[14621];
  assign N3665 = N3664 | data_masked[14749];
  assign N3664 = N3663 | data_masked[14877];
  assign N3663 = N3662 | data_masked[15005];
  assign N3662 = N3661 | data_masked[15133];
  assign N3661 = N3660 | data_masked[15261];
  assign N3660 = N3659 | data_masked[15389];
  assign N3659 = N3658 | data_masked[15517];
  assign N3658 = N3657 | data_masked[15645];
  assign N3657 = N3656 | data_masked[15773];
  assign N3656 = N3655 | data_masked[15901];
  assign N3655 = N3654 | data_masked[16029];
  assign N3654 = data_masked[16285] | data_masked[16157];
  assign data_o[30] = N3905 | data_masked[30];
  assign N3905 = N3904 | data_masked[158];
  assign N3904 = N3903 | data_masked[286];
  assign N3903 = N3902 | data_masked[414];
  assign N3902 = N3901 | data_masked[542];
  assign N3901 = N3900 | data_masked[670];
  assign N3900 = N3899 | data_masked[798];
  assign N3899 = N3898 | data_masked[926];
  assign N3898 = N3897 | data_masked[1054];
  assign N3897 = N3896 | data_masked[1182];
  assign N3896 = N3895 | data_masked[1310];
  assign N3895 = N3894 | data_masked[1438];
  assign N3894 = N3893 | data_masked[1566];
  assign N3893 = N3892 | data_masked[1694];
  assign N3892 = N3891 | data_masked[1822];
  assign N3891 = N3890 | data_masked[1950];
  assign N3890 = N3889 | data_masked[2078];
  assign N3889 = N3888 | data_masked[2206];
  assign N3888 = N3887 | data_masked[2334];
  assign N3887 = N3886 | data_masked[2462];
  assign N3886 = N3885 | data_masked[2590];
  assign N3885 = N3884 | data_masked[2718];
  assign N3884 = N3883 | data_masked[2846];
  assign N3883 = N3882 | data_masked[2974];
  assign N3882 = N3881 | data_masked[3102];
  assign N3881 = N3880 | data_masked[3230];
  assign N3880 = N3879 | data_masked[3358];
  assign N3879 = N3878 | data_masked[3486];
  assign N3878 = N3877 | data_masked[3614];
  assign N3877 = N3876 | data_masked[3742];
  assign N3876 = N3875 | data_masked[3870];
  assign N3875 = N3874 | data_masked[3998];
  assign N3874 = N3873 | data_masked[4126];
  assign N3873 = N3872 | data_masked[4254];
  assign N3872 = N3871 | data_masked[4382];
  assign N3871 = N3870 | data_masked[4510];
  assign N3870 = N3869 | data_masked[4638];
  assign N3869 = N3868 | data_masked[4766];
  assign N3868 = N3867 | data_masked[4894];
  assign N3867 = N3866 | data_masked[5022];
  assign N3866 = N3865 | data_masked[5150];
  assign N3865 = N3864 | data_masked[5278];
  assign N3864 = N3863 | data_masked[5406];
  assign N3863 = N3862 | data_masked[5534];
  assign N3862 = N3861 | data_masked[5662];
  assign N3861 = N3860 | data_masked[5790];
  assign N3860 = N3859 | data_masked[5918];
  assign N3859 = N3858 | data_masked[6046];
  assign N3858 = N3857 | data_masked[6174];
  assign N3857 = N3856 | data_masked[6302];
  assign N3856 = N3855 | data_masked[6430];
  assign N3855 = N3854 | data_masked[6558];
  assign N3854 = N3853 | data_masked[6686];
  assign N3853 = N3852 | data_masked[6814];
  assign N3852 = N3851 | data_masked[6942];
  assign N3851 = N3850 | data_masked[7070];
  assign N3850 = N3849 | data_masked[7198];
  assign N3849 = N3848 | data_masked[7326];
  assign N3848 = N3847 | data_masked[7454];
  assign N3847 = N3846 | data_masked[7582];
  assign N3846 = N3845 | data_masked[7710];
  assign N3845 = N3844 | data_masked[7838];
  assign N3844 = N3843 | data_masked[7966];
  assign N3843 = N3842 | data_masked[8094];
  assign N3842 = N3841 | data_masked[8222];
  assign N3841 = N3840 | data_masked[8350];
  assign N3840 = N3839 | data_masked[8478];
  assign N3839 = N3838 | data_masked[8606];
  assign N3838 = N3837 | data_masked[8734];
  assign N3837 = N3836 | data_masked[8862];
  assign N3836 = N3835 | data_masked[8990];
  assign N3835 = N3834 | data_masked[9118];
  assign N3834 = N3833 | data_masked[9246];
  assign N3833 = N3832 | data_masked[9374];
  assign N3832 = N3831 | data_masked[9502];
  assign N3831 = N3830 | data_masked[9630];
  assign N3830 = N3829 | data_masked[9758];
  assign N3829 = N3828 | data_masked[9886];
  assign N3828 = N3827 | data_masked[10014];
  assign N3827 = N3826 | data_masked[10142];
  assign N3826 = N3825 | data_masked[10270];
  assign N3825 = N3824 | data_masked[10398];
  assign N3824 = N3823 | data_masked[10526];
  assign N3823 = N3822 | data_masked[10654];
  assign N3822 = N3821 | data_masked[10782];
  assign N3821 = N3820 | data_masked[10910];
  assign N3820 = N3819 | data_masked[11038];
  assign N3819 = N3818 | data_masked[11166];
  assign N3818 = N3817 | data_masked[11294];
  assign N3817 = N3816 | data_masked[11422];
  assign N3816 = N3815 | data_masked[11550];
  assign N3815 = N3814 | data_masked[11678];
  assign N3814 = N3813 | data_masked[11806];
  assign N3813 = N3812 | data_masked[11934];
  assign N3812 = N3811 | data_masked[12062];
  assign N3811 = N3810 | data_masked[12190];
  assign N3810 = N3809 | data_masked[12318];
  assign N3809 = N3808 | data_masked[12446];
  assign N3808 = N3807 | data_masked[12574];
  assign N3807 = N3806 | data_masked[12702];
  assign N3806 = N3805 | data_masked[12830];
  assign N3805 = N3804 | data_masked[12958];
  assign N3804 = N3803 | data_masked[13086];
  assign N3803 = N3802 | data_masked[13214];
  assign N3802 = N3801 | data_masked[13342];
  assign N3801 = N3800 | data_masked[13470];
  assign N3800 = N3799 | data_masked[13598];
  assign N3799 = N3798 | data_masked[13726];
  assign N3798 = N3797 | data_masked[13854];
  assign N3797 = N3796 | data_masked[13982];
  assign N3796 = N3795 | data_masked[14110];
  assign N3795 = N3794 | data_masked[14238];
  assign N3794 = N3793 | data_masked[14366];
  assign N3793 = N3792 | data_masked[14494];
  assign N3792 = N3791 | data_masked[14622];
  assign N3791 = N3790 | data_masked[14750];
  assign N3790 = N3789 | data_masked[14878];
  assign N3789 = N3788 | data_masked[15006];
  assign N3788 = N3787 | data_masked[15134];
  assign N3787 = N3786 | data_masked[15262];
  assign N3786 = N3785 | data_masked[15390];
  assign N3785 = N3784 | data_masked[15518];
  assign N3784 = N3783 | data_masked[15646];
  assign N3783 = N3782 | data_masked[15774];
  assign N3782 = N3781 | data_masked[15902];
  assign N3781 = N3780 | data_masked[16030];
  assign N3780 = data_masked[16286] | data_masked[16158];
  assign data_o[31] = N4031 | data_masked[31];
  assign N4031 = N4030 | data_masked[159];
  assign N4030 = N4029 | data_masked[287];
  assign N4029 = N4028 | data_masked[415];
  assign N4028 = N4027 | data_masked[543];
  assign N4027 = N4026 | data_masked[671];
  assign N4026 = N4025 | data_masked[799];
  assign N4025 = N4024 | data_masked[927];
  assign N4024 = N4023 | data_masked[1055];
  assign N4023 = N4022 | data_masked[1183];
  assign N4022 = N4021 | data_masked[1311];
  assign N4021 = N4020 | data_masked[1439];
  assign N4020 = N4019 | data_masked[1567];
  assign N4019 = N4018 | data_masked[1695];
  assign N4018 = N4017 | data_masked[1823];
  assign N4017 = N4016 | data_masked[1951];
  assign N4016 = N4015 | data_masked[2079];
  assign N4015 = N4014 | data_masked[2207];
  assign N4014 = N4013 | data_masked[2335];
  assign N4013 = N4012 | data_masked[2463];
  assign N4012 = N4011 | data_masked[2591];
  assign N4011 = N4010 | data_masked[2719];
  assign N4010 = N4009 | data_masked[2847];
  assign N4009 = N4008 | data_masked[2975];
  assign N4008 = N4007 | data_masked[3103];
  assign N4007 = N4006 | data_masked[3231];
  assign N4006 = N4005 | data_masked[3359];
  assign N4005 = N4004 | data_masked[3487];
  assign N4004 = N4003 | data_masked[3615];
  assign N4003 = N4002 | data_masked[3743];
  assign N4002 = N4001 | data_masked[3871];
  assign N4001 = N4000 | data_masked[3999];
  assign N4000 = N3999 | data_masked[4127];
  assign N3999 = N3998 | data_masked[4255];
  assign N3998 = N3997 | data_masked[4383];
  assign N3997 = N3996 | data_masked[4511];
  assign N3996 = N3995 | data_masked[4639];
  assign N3995 = N3994 | data_masked[4767];
  assign N3994 = N3993 | data_masked[4895];
  assign N3993 = N3992 | data_masked[5023];
  assign N3992 = N3991 | data_masked[5151];
  assign N3991 = N3990 | data_masked[5279];
  assign N3990 = N3989 | data_masked[5407];
  assign N3989 = N3988 | data_masked[5535];
  assign N3988 = N3987 | data_masked[5663];
  assign N3987 = N3986 | data_masked[5791];
  assign N3986 = N3985 | data_masked[5919];
  assign N3985 = N3984 | data_masked[6047];
  assign N3984 = N3983 | data_masked[6175];
  assign N3983 = N3982 | data_masked[6303];
  assign N3982 = N3981 | data_masked[6431];
  assign N3981 = N3980 | data_masked[6559];
  assign N3980 = N3979 | data_masked[6687];
  assign N3979 = N3978 | data_masked[6815];
  assign N3978 = N3977 | data_masked[6943];
  assign N3977 = N3976 | data_masked[7071];
  assign N3976 = N3975 | data_masked[7199];
  assign N3975 = N3974 | data_masked[7327];
  assign N3974 = N3973 | data_masked[7455];
  assign N3973 = N3972 | data_masked[7583];
  assign N3972 = N3971 | data_masked[7711];
  assign N3971 = N3970 | data_masked[7839];
  assign N3970 = N3969 | data_masked[7967];
  assign N3969 = N3968 | data_masked[8095];
  assign N3968 = N3967 | data_masked[8223];
  assign N3967 = N3966 | data_masked[8351];
  assign N3966 = N3965 | data_masked[8479];
  assign N3965 = N3964 | data_masked[8607];
  assign N3964 = N3963 | data_masked[8735];
  assign N3963 = N3962 | data_masked[8863];
  assign N3962 = N3961 | data_masked[8991];
  assign N3961 = N3960 | data_masked[9119];
  assign N3960 = N3959 | data_masked[9247];
  assign N3959 = N3958 | data_masked[9375];
  assign N3958 = N3957 | data_masked[9503];
  assign N3957 = N3956 | data_masked[9631];
  assign N3956 = N3955 | data_masked[9759];
  assign N3955 = N3954 | data_masked[9887];
  assign N3954 = N3953 | data_masked[10015];
  assign N3953 = N3952 | data_masked[10143];
  assign N3952 = N3951 | data_masked[10271];
  assign N3951 = N3950 | data_masked[10399];
  assign N3950 = N3949 | data_masked[10527];
  assign N3949 = N3948 | data_masked[10655];
  assign N3948 = N3947 | data_masked[10783];
  assign N3947 = N3946 | data_masked[10911];
  assign N3946 = N3945 | data_masked[11039];
  assign N3945 = N3944 | data_masked[11167];
  assign N3944 = N3943 | data_masked[11295];
  assign N3943 = N3942 | data_masked[11423];
  assign N3942 = N3941 | data_masked[11551];
  assign N3941 = N3940 | data_masked[11679];
  assign N3940 = N3939 | data_masked[11807];
  assign N3939 = N3938 | data_masked[11935];
  assign N3938 = N3937 | data_masked[12063];
  assign N3937 = N3936 | data_masked[12191];
  assign N3936 = N3935 | data_masked[12319];
  assign N3935 = N3934 | data_masked[12447];
  assign N3934 = N3933 | data_masked[12575];
  assign N3933 = N3932 | data_masked[12703];
  assign N3932 = N3931 | data_masked[12831];
  assign N3931 = N3930 | data_masked[12959];
  assign N3930 = N3929 | data_masked[13087];
  assign N3929 = N3928 | data_masked[13215];
  assign N3928 = N3927 | data_masked[13343];
  assign N3927 = N3926 | data_masked[13471];
  assign N3926 = N3925 | data_masked[13599];
  assign N3925 = N3924 | data_masked[13727];
  assign N3924 = N3923 | data_masked[13855];
  assign N3923 = N3922 | data_masked[13983];
  assign N3922 = N3921 | data_masked[14111];
  assign N3921 = N3920 | data_masked[14239];
  assign N3920 = N3919 | data_masked[14367];
  assign N3919 = N3918 | data_masked[14495];
  assign N3918 = N3917 | data_masked[14623];
  assign N3917 = N3916 | data_masked[14751];
  assign N3916 = N3915 | data_masked[14879];
  assign N3915 = N3914 | data_masked[15007];
  assign N3914 = N3913 | data_masked[15135];
  assign N3913 = N3912 | data_masked[15263];
  assign N3912 = N3911 | data_masked[15391];
  assign N3911 = N3910 | data_masked[15519];
  assign N3910 = N3909 | data_masked[15647];
  assign N3909 = N3908 | data_masked[15775];
  assign N3908 = N3907 | data_masked[15903];
  assign N3907 = N3906 | data_masked[16031];
  assign N3906 = data_masked[16287] | data_masked[16159];
  assign data_o[32] = N4157 | data_masked[32];
  assign N4157 = N4156 | data_masked[160];
  assign N4156 = N4155 | data_masked[288];
  assign N4155 = N4154 | data_masked[416];
  assign N4154 = N4153 | data_masked[544];
  assign N4153 = N4152 | data_masked[672];
  assign N4152 = N4151 | data_masked[800];
  assign N4151 = N4150 | data_masked[928];
  assign N4150 = N4149 | data_masked[1056];
  assign N4149 = N4148 | data_masked[1184];
  assign N4148 = N4147 | data_masked[1312];
  assign N4147 = N4146 | data_masked[1440];
  assign N4146 = N4145 | data_masked[1568];
  assign N4145 = N4144 | data_masked[1696];
  assign N4144 = N4143 | data_masked[1824];
  assign N4143 = N4142 | data_masked[1952];
  assign N4142 = N4141 | data_masked[2080];
  assign N4141 = N4140 | data_masked[2208];
  assign N4140 = N4139 | data_masked[2336];
  assign N4139 = N4138 | data_masked[2464];
  assign N4138 = N4137 | data_masked[2592];
  assign N4137 = N4136 | data_masked[2720];
  assign N4136 = N4135 | data_masked[2848];
  assign N4135 = N4134 | data_masked[2976];
  assign N4134 = N4133 | data_masked[3104];
  assign N4133 = N4132 | data_masked[3232];
  assign N4132 = N4131 | data_masked[3360];
  assign N4131 = N4130 | data_masked[3488];
  assign N4130 = N4129 | data_masked[3616];
  assign N4129 = N4128 | data_masked[3744];
  assign N4128 = N4127 | data_masked[3872];
  assign N4127 = N4126 | data_masked[4000];
  assign N4126 = N4125 | data_masked[4128];
  assign N4125 = N4124 | data_masked[4256];
  assign N4124 = N4123 | data_masked[4384];
  assign N4123 = N4122 | data_masked[4512];
  assign N4122 = N4121 | data_masked[4640];
  assign N4121 = N4120 | data_masked[4768];
  assign N4120 = N4119 | data_masked[4896];
  assign N4119 = N4118 | data_masked[5024];
  assign N4118 = N4117 | data_masked[5152];
  assign N4117 = N4116 | data_masked[5280];
  assign N4116 = N4115 | data_masked[5408];
  assign N4115 = N4114 | data_masked[5536];
  assign N4114 = N4113 | data_masked[5664];
  assign N4113 = N4112 | data_masked[5792];
  assign N4112 = N4111 | data_masked[5920];
  assign N4111 = N4110 | data_masked[6048];
  assign N4110 = N4109 | data_masked[6176];
  assign N4109 = N4108 | data_masked[6304];
  assign N4108 = N4107 | data_masked[6432];
  assign N4107 = N4106 | data_masked[6560];
  assign N4106 = N4105 | data_masked[6688];
  assign N4105 = N4104 | data_masked[6816];
  assign N4104 = N4103 | data_masked[6944];
  assign N4103 = N4102 | data_masked[7072];
  assign N4102 = N4101 | data_masked[7200];
  assign N4101 = N4100 | data_masked[7328];
  assign N4100 = N4099 | data_masked[7456];
  assign N4099 = N4098 | data_masked[7584];
  assign N4098 = N4097 | data_masked[7712];
  assign N4097 = N4096 | data_masked[7840];
  assign N4096 = N4095 | data_masked[7968];
  assign N4095 = N4094 | data_masked[8096];
  assign N4094 = N4093 | data_masked[8224];
  assign N4093 = N4092 | data_masked[8352];
  assign N4092 = N4091 | data_masked[8480];
  assign N4091 = N4090 | data_masked[8608];
  assign N4090 = N4089 | data_masked[8736];
  assign N4089 = N4088 | data_masked[8864];
  assign N4088 = N4087 | data_masked[8992];
  assign N4087 = N4086 | data_masked[9120];
  assign N4086 = N4085 | data_masked[9248];
  assign N4085 = N4084 | data_masked[9376];
  assign N4084 = N4083 | data_masked[9504];
  assign N4083 = N4082 | data_masked[9632];
  assign N4082 = N4081 | data_masked[9760];
  assign N4081 = N4080 | data_masked[9888];
  assign N4080 = N4079 | data_masked[10016];
  assign N4079 = N4078 | data_masked[10144];
  assign N4078 = N4077 | data_masked[10272];
  assign N4077 = N4076 | data_masked[10400];
  assign N4076 = N4075 | data_masked[10528];
  assign N4075 = N4074 | data_masked[10656];
  assign N4074 = N4073 | data_masked[10784];
  assign N4073 = N4072 | data_masked[10912];
  assign N4072 = N4071 | data_masked[11040];
  assign N4071 = N4070 | data_masked[11168];
  assign N4070 = N4069 | data_masked[11296];
  assign N4069 = N4068 | data_masked[11424];
  assign N4068 = N4067 | data_masked[11552];
  assign N4067 = N4066 | data_masked[11680];
  assign N4066 = N4065 | data_masked[11808];
  assign N4065 = N4064 | data_masked[11936];
  assign N4064 = N4063 | data_masked[12064];
  assign N4063 = N4062 | data_masked[12192];
  assign N4062 = N4061 | data_masked[12320];
  assign N4061 = N4060 | data_masked[12448];
  assign N4060 = N4059 | data_masked[12576];
  assign N4059 = N4058 | data_masked[12704];
  assign N4058 = N4057 | data_masked[12832];
  assign N4057 = N4056 | data_masked[12960];
  assign N4056 = N4055 | data_masked[13088];
  assign N4055 = N4054 | data_masked[13216];
  assign N4054 = N4053 | data_masked[13344];
  assign N4053 = N4052 | data_masked[13472];
  assign N4052 = N4051 | data_masked[13600];
  assign N4051 = N4050 | data_masked[13728];
  assign N4050 = N4049 | data_masked[13856];
  assign N4049 = N4048 | data_masked[13984];
  assign N4048 = N4047 | data_masked[14112];
  assign N4047 = N4046 | data_masked[14240];
  assign N4046 = N4045 | data_masked[14368];
  assign N4045 = N4044 | data_masked[14496];
  assign N4044 = N4043 | data_masked[14624];
  assign N4043 = N4042 | data_masked[14752];
  assign N4042 = N4041 | data_masked[14880];
  assign N4041 = N4040 | data_masked[15008];
  assign N4040 = N4039 | data_masked[15136];
  assign N4039 = N4038 | data_masked[15264];
  assign N4038 = N4037 | data_masked[15392];
  assign N4037 = N4036 | data_masked[15520];
  assign N4036 = N4035 | data_masked[15648];
  assign N4035 = N4034 | data_masked[15776];
  assign N4034 = N4033 | data_masked[15904];
  assign N4033 = N4032 | data_masked[16032];
  assign N4032 = data_masked[16288] | data_masked[16160];
  assign data_o[33] = N4283 | data_masked[33];
  assign N4283 = N4282 | data_masked[161];
  assign N4282 = N4281 | data_masked[289];
  assign N4281 = N4280 | data_masked[417];
  assign N4280 = N4279 | data_masked[545];
  assign N4279 = N4278 | data_masked[673];
  assign N4278 = N4277 | data_masked[801];
  assign N4277 = N4276 | data_masked[929];
  assign N4276 = N4275 | data_masked[1057];
  assign N4275 = N4274 | data_masked[1185];
  assign N4274 = N4273 | data_masked[1313];
  assign N4273 = N4272 | data_masked[1441];
  assign N4272 = N4271 | data_masked[1569];
  assign N4271 = N4270 | data_masked[1697];
  assign N4270 = N4269 | data_masked[1825];
  assign N4269 = N4268 | data_masked[1953];
  assign N4268 = N4267 | data_masked[2081];
  assign N4267 = N4266 | data_masked[2209];
  assign N4266 = N4265 | data_masked[2337];
  assign N4265 = N4264 | data_masked[2465];
  assign N4264 = N4263 | data_masked[2593];
  assign N4263 = N4262 | data_masked[2721];
  assign N4262 = N4261 | data_masked[2849];
  assign N4261 = N4260 | data_masked[2977];
  assign N4260 = N4259 | data_masked[3105];
  assign N4259 = N4258 | data_masked[3233];
  assign N4258 = N4257 | data_masked[3361];
  assign N4257 = N4256 | data_masked[3489];
  assign N4256 = N4255 | data_masked[3617];
  assign N4255 = N4254 | data_masked[3745];
  assign N4254 = N4253 | data_masked[3873];
  assign N4253 = N4252 | data_masked[4001];
  assign N4252 = N4251 | data_masked[4129];
  assign N4251 = N4250 | data_masked[4257];
  assign N4250 = N4249 | data_masked[4385];
  assign N4249 = N4248 | data_masked[4513];
  assign N4248 = N4247 | data_masked[4641];
  assign N4247 = N4246 | data_masked[4769];
  assign N4246 = N4245 | data_masked[4897];
  assign N4245 = N4244 | data_masked[5025];
  assign N4244 = N4243 | data_masked[5153];
  assign N4243 = N4242 | data_masked[5281];
  assign N4242 = N4241 | data_masked[5409];
  assign N4241 = N4240 | data_masked[5537];
  assign N4240 = N4239 | data_masked[5665];
  assign N4239 = N4238 | data_masked[5793];
  assign N4238 = N4237 | data_masked[5921];
  assign N4237 = N4236 | data_masked[6049];
  assign N4236 = N4235 | data_masked[6177];
  assign N4235 = N4234 | data_masked[6305];
  assign N4234 = N4233 | data_masked[6433];
  assign N4233 = N4232 | data_masked[6561];
  assign N4232 = N4231 | data_masked[6689];
  assign N4231 = N4230 | data_masked[6817];
  assign N4230 = N4229 | data_masked[6945];
  assign N4229 = N4228 | data_masked[7073];
  assign N4228 = N4227 | data_masked[7201];
  assign N4227 = N4226 | data_masked[7329];
  assign N4226 = N4225 | data_masked[7457];
  assign N4225 = N4224 | data_masked[7585];
  assign N4224 = N4223 | data_masked[7713];
  assign N4223 = N4222 | data_masked[7841];
  assign N4222 = N4221 | data_masked[7969];
  assign N4221 = N4220 | data_masked[8097];
  assign N4220 = N4219 | data_masked[8225];
  assign N4219 = N4218 | data_masked[8353];
  assign N4218 = N4217 | data_masked[8481];
  assign N4217 = N4216 | data_masked[8609];
  assign N4216 = N4215 | data_masked[8737];
  assign N4215 = N4214 | data_masked[8865];
  assign N4214 = N4213 | data_masked[8993];
  assign N4213 = N4212 | data_masked[9121];
  assign N4212 = N4211 | data_masked[9249];
  assign N4211 = N4210 | data_masked[9377];
  assign N4210 = N4209 | data_masked[9505];
  assign N4209 = N4208 | data_masked[9633];
  assign N4208 = N4207 | data_masked[9761];
  assign N4207 = N4206 | data_masked[9889];
  assign N4206 = N4205 | data_masked[10017];
  assign N4205 = N4204 | data_masked[10145];
  assign N4204 = N4203 | data_masked[10273];
  assign N4203 = N4202 | data_masked[10401];
  assign N4202 = N4201 | data_masked[10529];
  assign N4201 = N4200 | data_masked[10657];
  assign N4200 = N4199 | data_masked[10785];
  assign N4199 = N4198 | data_masked[10913];
  assign N4198 = N4197 | data_masked[11041];
  assign N4197 = N4196 | data_masked[11169];
  assign N4196 = N4195 | data_masked[11297];
  assign N4195 = N4194 | data_masked[11425];
  assign N4194 = N4193 | data_masked[11553];
  assign N4193 = N4192 | data_masked[11681];
  assign N4192 = N4191 | data_masked[11809];
  assign N4191 = N4190 | data_masked[11937];
  assign N4190 = N4189 | data_masked[12065];
  assign N4189 = N4188 | data_masked[12193];
  assign N4188 = N4187 | data_masked[12321];
  assign N4187 = N4186 | data_masked[12449];
  assign N4186 = N4185 | data_masked[12577];
  assign N4185 = N4184 | data_masked[12705];
  assign N4184 = N4183 | data_masked[12833];
  assign N4183 = N4182 | data_masked[12961];
  assign N4182 = N4181 | data_masked[13089];
  assign N4181 = N4180 | data_masked[13217];
  assign N4180 = N4179 | data_masked[13345];
  assign N4179 = N4178 | data_masked[13473];
  assign N4178 = N4177 | data_masked[13601];
  assign N4177 = N4176 | data_masked[13729];
  assign N4176 = N4175 | data_masked[13857];
  assign N4175 = N4174 | data_masked[13985];
  assign N4174 = N4173 | data_masked[14113];
  assign N4173 = N4172 | data_masked[14241];
  assign N4172 = N4171 | data_masked[14369];
  assign N4171 = N4170 | data_masked[14497];
  assign N4170 = N4169 | data_masked[14625];
  assign N4169 = N4168 | data_masked[14753];
  assign N4168 = N4167 | data_masked[14881];
  assign N4167 = N4166 | data_masked[15009];
  assign N4166 = N4165 | data_masked[15137];
  assign N4165 = N4164 | data_masked[15265];
  assign N4164 = N4163 | data_masked[15393];
  assign N4163 = N4162 | data_masked[15521];
  assign N4162 = N4161 | data_masked[15649];
  assign N4161 = N4160 | data_masked[15777];
  assign N4160 = N4159 | data_masked[15905];
  assign N4159 = N4158 | data_masked[16033];
  assign N4158 = data_masked[16289] | data_masked[16161];
  assign data_o[34] = N4409 | data_masked[34];
  assign N4409 = N4408 | data_masked[162];
  assign N4408 = N4407 | data_masked[290];
  assign N4407 = N4406 | data_masked[418];
  assign N4406 = N4405 | data_masked[546];
  assign N4405 = N4404 | data_masked[674];
  assign N4404 = N4403 | data_masked[802];
  assign N4403 = N4402 | data_masked[930];
  assign N4402 = N4401 | data_masked[1058];
  assign N4401 = N4400 | data_masked[1186];
  assign N4400 = N4399 | data_masked[1314];
  assign N4399 = N4398 | data_masked[1442];
  assign N4398 = N4397 | data_masked[1570];
  assign N4397 = N4396 | data_masked[1698];
  assign N4396 = N4395 | data_masked[1826];
  assign N4395 = N4394 | data_masked[1954];
  assign N4394 = N4393 | data_masked[2082];
  assign N4393 = N4392 | data_masked[2210];
  assign N4392 = N4391 | data_masked[2338];
  assign N4391 = N4390 | data_masked[2466];
  assign N4390 = N4389 | data_masked[2594];
  assign N4389 = N4388 | data_masked[2722];
  assign N4388 = N4387 | data_masked[2850];
  assign N4387 = N4386 | data_masked[2978];
  assign N4386 = N4385 | data_masked[3106];
  assign N4385 = N4384 | data_masked[3234];
  assign N4384 = N4383 | data_masked[3362];
  assign N4383 = N4382 | data_masked[3490];
  assign N4382 = N4381 | data_masked[3618];
  assign N4381 = N4380 | data_masked[3746];
  assign N4380 = N4379 | data_masked[3874];
  assign N4379 = N4378 | data_masked[4002];
  assign N4378 = N4377 | data_masked[4130];
  assign N4377 = N4376 | data_masked[4258];
  assign N4376 = N4375 | data_masked[4386];
  assign N4375 = N4374 | data_masked[4514];
  assign N4374 = N4373 | data_masked[4642];
  assign N4373 = N4372 | data_masked[4770];
  assign N4372 = N4371 | data_masked[4898];
  assign N4371 = N4370 | data_masked[5026];
  assign N4370 = N4369 | data_masked[5154];
  assign N4369 = N4368 | data_masked[5282];
  assign N4368 = N4367 | data_masked[5410];
  assign N4367 = N4366 | data_masked[5538];
  assign N4366 = N4365 | data_masked[5666];
  assign N4365 = N4364 | data_masked[5794];
  assign N4364 = N4363 | data_masked[5922];
  assign N4363 = N4362 | data_masked[6050];
  assign N4362 = N4361 | data_masked[6178];
  assign N4361 = N4360 | data_masked[6306];
  assign N4360 = N4359 | data_masked[6434];
  assign N4359 = N4358 | data_masked[6562];
  assign N4358 = N4357 | data_masked[6690];
  assign N4357 = N4356 | data_masked[6818];
  assign N4356 = N4355 | data_masked[6946];
  assign N4355 = N4354 | data_masked[7074];
  assign N4354 = N4353 | data_masked[7202];
  assign N4353 = N4352 | data_masked[7330];
  assign N4352 = N4351 | data_masked[7458];
  assign N4351 = N4350 | data_masked[7586];
  assign N4350 = N4349 | data_masked[7714];
  assign N4349 = N4348 | data_masked[7842];
  assign N4348 = N4347 | data_masked[7970];
  assign N4347 = N4346 | data_masked[8098];
  assign N4346 = N4345 | data_masked[8226];
  assign N4345 = N4344 | data_masked[8354];
  assign N4344 = N4343 | data_masked[8482];
  assign N4343 = N4342 | data_masked[8610];
  assign N4342 = N4341 | data_masked[8738];
  assign N4341 = N4340 | data_masked[8866];
  assign N4340 = N4339 | data_masked[8994];
  assign N4339 = N4338 | data_masked[9122];
  assign N4338 = N4337 | data_masked[9250];
  assign N4337 = N4336 | data_masked[9378];
  assign N4336 = N4335 | data_masked[9506];
  assign N4335 = N4334 | data_masked[9634];
  assign N4334 = N4333 | data_masked[9762];
  assign N4333 = N4332 | data_masked[9890];
  assign N4332 = N4331 | data_masked[10018];
  assign N4331 = N4330 | data_masked[10146];
  assign N4330 = N4329 | data_masked[10274];
  assign N4329 = N4328 | data_masked[10402];
  assign N4328 = N4327 | data_masked[10530];
  assign N4327 = N4326 | data_masked[10658];
  assign N4326 = N4325 | data_masked[10786];
  assign N4325 = N4324 | data_masked[10914];
  assign N4324 = N4323 | data_masked[11042];
  assign N4323 = N4322 | data_masked[11170];
  assign N4322 = N4321 | data_masked[11298];
  assign N4321 = N4320 | data_masked[11426];
  assign N4320 = N4319 | data_masked[11554];
  assign N4319 = N4318 | data_masked[11682];
  assign N4318 = N4317 | data_masked[11810];
  assign N4317 = N4316 | data_masked[11938];
  assign N4316 = N4315 | data_masked[12066];
  assign N4315 = N4314 | data_masked[12194];
  assign N4314 = N4313 | data_masked[12322];
  assign N4313 = N4312 | data_masked[12450];
  assign N4312 = N4311 | data_masked[12578];
  assign N4311 = N4310 | data_masked[12706];
  assign N4310 = N4309 | data_masked[12834];
  assign N4309 = N4308 | data_masked[12962];
  assign N4308 = N4307 | data_masked[13090];
  assign N4307 = N4306 | data_masked[13218];
  assign N4306 = N4305 | data_masked[13346];
  assign N4305 = N4304 | data_masked[13474];
  assign N4304 = N4303 | data_masked[13602];
  assign N4303 = N4302 | data_masked[13730];
  assign N4302 = N4301 | data_masked[13858];
  assign N4301 = N4300 | data_masked[13986];
  assign N4300 = N4299 | data_masked[14114];
  assign N4299 = N4298 | data_masked[14242];
  assign N4298 = N4297 | data_masked[14370];
  assign N4297 = N4296 | data_masked[14498];
  assign N4296 = N4295 | data_masked[14626];
  assign N4295 = N4294 | data_masked[14754];
  assign N4294 = N4293 | data_masked[14882];
  assign N4293 = N4292 | data_masked[15010];
  assign N4292 = N4291 | data_masked[15138];
  assign N4291 = N4290 | data_masked[15266];
  assign N4290 = N4289 | data_masked[15394];
  assign N4289 = N4288 | data_masked[15522];
  assign N4288 = N4287 | data_masked[15650];
  assign N4287 = N4286 | data_masked[15778];
  assign N4286 = N4285 | data_masked[15906];
  assign N4285 = N4284 | data_masked[16034];
  assign N4284 = data_masked[16290] | data_masked[16162];
  assign data_o[35] = N4535 | data_masked[35];
  assign N4535 = N4534 | data_masked[163];
  assign N4534 = N4533 | data_masked[291];
  assign N4533 = N4532 | data_masked[419];
  assign N4532 = N4531 | data_masked[547];
  assign N4531 = N4530 | data_masked[675];
  assign N4530 = N4529 | data_masked[803];
  assign N4529 = N4528 | data_masked[931];
  assign N4528 = N4527 | data_masked[1059];
  assign N4527 = N4526 | data_masked[1187];
  assign N4526 = N4525 | data_masked[1315];
  assign N4525 = N4524 | data_masked[1443];
  assign N4524 = N4523 | data_masked[1571];
  assign N4523 = N4522 | data_masked[1699];
  assign N4522 = N4521 | data_masked[1827];
  assign N4521 = N4520 | data_masked[1955];
  assign N4520 = N4519 | data_masked[2083];
  assign N4519 = N4518 | data_masked[2211];
  assign N4518 = N4517 | data_masked[2339];
  assign N4517 = N4516 | data_masked[2467];
  assign N4516 = N4515 | data_masked[2595];
  assign N4515 = N4514 | data_masked[2723];
  assign N4514 = N4513 | data_masked[2851];
  assign N4513 = N4512 | data_masked[2979];
  assign N4512 = N4511 | data_masked[3107];
  assign N4511 = N4510 | data_masked[3235];
  assign N4510 = N4509 | data_masked[3363];
  assign N4509 = N4508 | data_masked[3491];
  assign N4508 = N4507 | data_masked[3619];
  assign N4507 = N4506 | data_masked[3747];
  assign N4506 = N4505 | data_masked[3875];
  assign N4505 = N4504 | data_masked[4003];
  assign N4504 = N4503 | data_masked[4131];
  assign N4503 = N4502 | data_masked[4259];
  assign N4502 = N4501 | data_masked[4387];
  assign N4501 = N4500 | data_masked[4515];
  assign N4500 = N4499 | data_masked[4643];
  assign N4499 = N4498 | data_masked[4771];
  assign N4498 = N4497 | data_masked[4899];
  assign N4497 = N4496 | data_masked[5027];
  assign N4496 = N4495 | data_masked[5155];
  assign N4495 = N4494 | data_masked[5283];
  assign N4494 = N4493 | data_masked[5411];
  assign N4493 = N4492 | data_masked[5539];
  assign N4492 = N4491 | data_masked[5667];
  assign N4491 = N4490 | data_masked[5795];
  assign N4490 = N4489 | data_masked[5923];
  assign N4489 = N4488 | data_masked[6051];
  assign N4488 = N4487 | data_masked[6179];
  assign N4487 = N4486 | data_masked[6307];
  assign N4486 = N4485 | data_masked[6435];
  assign N4485 = N4484 | data_masked[6563];
  assign N4484 = N4483 | data_masked[6691];
  assign N4483 = N4482 | data_masked[6819];
  assign N4482 = N4481 | data_masked[6947];
  assign N4481 = N4480 | data_masked[7075];
  assign N4480 = N4479 | data_masked[7203];
  assign N4479 = N4478 | data_masked[7331];
  assign N4478 = N4477 | data_masked[7459];
  assign N4477 = N4476 | data_masked[7587];
  assign N4476 = N4475 | data_masked[7715];
  assign N4475 = N4474 | data_masked[7843];
  assign N4474 = N4473 | data_masked[7971];
  assign N4473 = N4472 | data_masked[8099];
  assign N4472 = N4471 | data_masked[8227];
  assign N4471 = N4470 | data_masked[8355];
  assign N4470 = N4469 | data_masked[8483];
  assign N4469 = N4468 | data_masked[8611];
  assign N4468 = N4467 | data_masked[8739];
  assign N4467 = N4466 | data_masked[8867];
  assign N4466 = N4465 | data_masked[8995];
  assign N4465 = N4464 | data_masked[9123];
  assign N4464 = N4463 | data_masked[9251];
  assign N4463 = N4462 | data_masked[9379];
  assign N4462 = N4461 | data_masked[9507];
  assign N4461 = N4460 | data_masked[9635];
  assign N4460 = N4459 | data_masked[9763];
  assign N4459 = N4458 | data_masked[9891];
  assign N4458 = N4457 | data_masked[10019];
  assign N4457 = N4456 | data_masked[10147];
  assign N4456 = N4455 | data_masked[10275];
  assign N4455 = N4454 | data_masked[10403];
  assign N4454 = N4453 | data_masked[10531];
  assign N4453 = N4452 | data_masked[10659];
  assign N4452 = N4451 | data_masked[10787];
  assign N4451 = N4450 | data_masked[10915];
  assign N4450 = N4449 | data_masked[11043];
  assign N4449 = N4448 | data_masked[11171];
  assign N4448 = N4447 | data_masked[11299];
  assign N4447 = N4446 | data_masked[11427];
  assign N4446 = N4445 | data_masked[11555];
  assign N4445 = N4444 | data_masked[11683];
  assign N4444 = N4443 | data_masked[11811];
  assign N4443 = N4442 | data_masked[11939];
  assign N4442 = N4441 | data_masked[12067];
  assign N4441 = N4440 | data_masked[12195];
  assign N4440 = N4439 | data_masked[12323];
  assign N4439 = N4438 | data_masked[12451];
  assign N4438 = N4437 | data_masked[12579];
  assign N4437 = N4436 | data_masked[12707];
  assign N4436 = N4435 | data_masked[12835];
  assign N4435 = N4434 | data_masked[12963];
  assign N4434 = N4433 | data_masked[13091];
  assign N4433 = N4432 | data_masked[13219];
  assign N4432 = N4431 | data_masked[13347];
  assign N4431 = N4430 | data_masked[13475];
  assign N4430 = N4429 | data_masked[13603];
  assign N4429 = N4428 | data_masked[13731];
  assign N4428 = N4427 | data_masked[13859];
  assign N4427 = N4426 | data_masked[13987];
  assign N4426 = N4425 | data_masked[14115];
  assign N4425 = N4424 | data_masked[14243];
  assign N4424 = N4423 | data_masked[14371];
  assign N4423 = N4422 | data_masked[14499];
  assign N4422 = N4421 | data_masked[14627];
  assign N4421 = N4420 | data_masked[14755];
  assign N4420 = N4419 | data_masked[14883];
  assign N4419 = N4418 | data_masked[15011];
  assign N4418 = N4417 | data_masked[15139];
  assign N4417 = N4416 | data_masked[15267];
  assign N4416 = N4415 | data_masked[15395];
  assign N4415 = N4414 | data_masked[15523];
  assign N4414 = N4413 | data_masked[15651];
  assign N4413 = N4412 | data_masked[15779];
  assign N4412 = N4411 | data_masked[15907];
  assign N4411 = N4410 | data_masked[16035];
  assign N4410 = data_masked[16291] | data_masked[16163];
  assign data_o[36] = N4661 | data_masked[36];
  assign N4661 = N4660 | data_masked[164];
  assign N4660 = N4659 | data_masked[292];
  assign N4659 = N4658 | data_masked[420];
  assign N4658 = N4657 | data_masked[548];
  assign N4657 = N4656 | data_masked[676];
  assign N4656 = N4655 | data_masked[804];
  assign N4655 = N4654 | data_masked[932];
  assign N4654 = N4653 | data_masked[1060];
  assign N4653 = N4652 | data_masked[1188];
  assign N4652 = N4651 | data_masked[1316];
  assign N4651 = N4650 | data_masked[1444];
  assign N4650 = N4649 | data_masked[1572];
  assign N4649 = N4648 | data_masked[1700];
  assign N4648 = N4647 | data_masked[1828];
  assign N4647 = N4646 | data_masked[1956];
  assign N4646 = N4645 | data_masked[2084];
  assign N4645 = N4644 | data_masked[2212];
  assign N4644 = N4643 | data_masked[2340];
  assign N4643 = N4642 | data_masked[2468];
  assign N4642 = N4641 | data_masked[2596];
  assign N4641 = N4640 | data_masked[2724];
  assign N4640 = N4639 | data_masked[2852];
  assign N4639 = N4638 | data_masked[2980];
  assign N4638 = N4637 | data_masked[3108];
  assign N4637 = N4636 | data_masked[3236];
  assign N4636 = N4635 | data_masked[3364];
  assign N4635 = N4634 | data_masked[3492];
  assign N4634 = N4633 | data_masked[3620];
  assign N4633 = N4632 | data_masked[3748];
  assign N4632 = N4631 | data_masked[3876];
  assign N4631 = N4630 | data_masked[4004];
  assign N4630 = N4629 | data_masked[4132];
  assign N4629 = N4628 | data_masked[4260];
  assign N4628 = N4627 | data_masked[4388];
  assign N4627 = N4626 | data_masked[4516];
  assign N4626 = N4625 | data_masked[4644];
  assign N4625 = N4624 | data_masked[4772];
  assign N4624 = N4623 | data_masked[4900];
  assign N4623 = N4622 | data_masked[5028];
  assign N4622 = N4621 | data_masked[5156];
  assign N4621 = N4620 | data_masked[5284];
  assign N4620 = N4619 | data_masked[5412];
  assign N4619 = N4618 | data_masked[5540];
  assign N4618 = N4617 | data_masked[5668];
  assign N4617 = N4616 | data_masked[5796];
  assign N4616 = N4615 | data_masked[5924];
  assign N4615 = N4614 | data_masked[6052];
  assign N4614 = N4613 | data_masked[6180];
  assign N4613 = N4612 | data_masked[6308];
  assign N4612 = N4611 | data_masked[6436];
  assign N4611 = N4610 | data_masked[6564];
  assign N4610 = N4609 | data_masked[6692];
  assign N4609 = N4608 | data_masked[6820];
  assign N4608 = N4607 | data_masked[6948];
  assign N4607 = N4606 | data_masked[7076];
  assign N4606 = N4605 | data_masked[7204];
  assign N4605 = N4604 | data_masked[7332];
  assign N4604 = N4603 | data_masked[7460];
  assign N4603 = N4602 | data_masked[7588];
  assign N4602 = N4601 | data_masked[7716];
  assign N4601 = N4600 | data_masked[7844];
  assign N4600 = N4599 | data_masked[7972];
  assign N4599 = N4598 | data_masked[8100];
  assign N4598 = N4597 | data_masked[8228];
  assign N4597 = N4596 | data_masked[8356];
  assign N4596 = N4595 | data_masked[8484];
  assign N4595 = N4594 | data_masked[8612];
  assign N4594 = N4593 | data_masked[8740];
  assign N4593 = N4592 | data_masked[8868];
  assign N4592 = N4591 | data_masked[8996];
  assign N4591 = N4590 | data_masked[9124];
  assign N4590 = N4589 | data_masked[9252];
  assign N4589 = N4588 | data_masked[9380];
  assign N4588 = N4587 | data_masked[9508];
  assign N4587 = N4586 | data_masked[9636];
  assign N4586 = N4585 | data_masked[9764];
  assign N4585 = N4584 | data_masked[9892];
  assign N4584 = N4583 | data_masked[10020];
  assign N4583 = N4582 | data_masked[10148];
  assign N4582 = N4581 | data_masked[10276];
  assign N4581 = N4580 | data_masked[10404];
  assign N4580 = N4579 | data_masked[10532];
  assign N4579 = N4578 | data_masked[10660];
  assign N4578 = N4577 | data_masked[10788];
  assign N4577 = N4576 | data_masked[10916];
  assign N4576 = N4575 | data_masked[11044];
  assign N4575 = N4574 | data_masked[11172];
  assign N4574 = N4573 | data_masked[11300];
  assign N4573 = N4572 | data_masked[11428];
  assign N4572 = N4571 | data_masked[11556];
  assign N4571 = N4570 | data_masked[11684];
  assign N4570 = N4569 | data_masked[11812];
  assign N4569 = N4568 | data_masked[11940];
  assign N4568 = N4567 | data_masked[12068];
  assign N4567 = N4566 | data_masked[12196];
  assign N4566 = N4565 | data_masked[12324];
  assign N4565 = N4564 | data_masked[12452];
  assign N4564 = N4563 | data_masked[12580];
  assign N4563 = N4562 | data_masked[12708];
  assign N4562 = N4561 | data_masked[12836];
  assign N4561 = N4560 | data_masked[12964];
  assign N4560 = N4559 | data_masked[13092];
  assign N4559 = N4558 | data_masked[13220];
  assign N4558 = N4557 | data_masked[13348];
  assign N4557 = N4556 | data_masked[13476];
  assign N4556 = N4555 | data_masked[13604];
  assign N4555 = N4554 | data_masked[13732];
  assign N4554 = N4553 | data_masked[13860];
  assign N4553 = N4552 | data_masked[13988];
  assign N4552 = N4551 | data_masked[14116];
  assign N4551 = N4550 | data_masked[14244];
  assign N4550 = N4549 | data_masked[14372];
  assign N4549 = N4548 | data_masked[14500];
  assign N4548 = N4547 | data_masked[14628];
  assign N4547 = N4546 | data_masked[14756];
  assign N4546 = N4545 | data_masked[14884];
  assign N4545 = N4544 | data_masked[15012];
  assign N4544 = N4543 | data_masked[15140];
  assign N4543 = N4542 | data_masked[15268];
  assign N4542 = N4541 | data_masked[15396];
  assign N4541 = N4540 | data_masked[15524];
  assign N4540 = N4539 | data_masked[15652];
  assign N4539 = N4538 | data_masked[15780];
  assign N4538 = N4537 | data_masked[15908];
  assign N4537 = N4536 | data_masked[16036];
  assign N4536 = data_masked[16292] | data_masked[16164];
  assign data_o[37] = N4787 | data_masked[37];
  assign N4787 = N4786 | data_masked[165];
  assign N4786 = N4785 | data_masked[293];
  assign N4785 = N4784 | data_masked[421];
  assign N4784 = N4783 | data_masked[549];
  assign N4783 = N4782 | data_masked[677];
  assign N4782 = N4781 | data_masked[805];
  assign N4781 = N4780 | data_masked[933];
  assign N4780 = N4779 | data_masked[1061];
  assign N4779 = N4778 | data_masked[1189];
  assign N4778 = N4777 | data_masked[1317];
  assign N4777 = N4776 | data_masked[1445];
  assign N4776 = N4775 | data_masked[1573];
  assign N4775 = N4774 | data_masked[1701];
  assign N4774 = N4773 | data_masked[1829];
  assign N4773 = N4772 | data_masked[1957];
  assign N4772 = N4771 | data_masked[2085];
  assign N4771 = N4770 | data_masked[2213];
  assign N4770 = N4769 | data_masked[2341];
  assign N4769 = N4768 | data_masked[2469];
  assign N4768 = N4767 | data_masked[2597];
  assign N4767 = N4766 | data_masked[2725];
  assign N4766 = N4765 | data_masked[2853];
  assign N4765 = N4764 | data_masked[2981];
  assign N4764 = N4763 | data_masked[3109];
  assign N4763 = N4762 | data_masked[3237];
  assign N4762 = N4761 | data_masked[3365];
  assign N4761 = N4760 | data_masked[3493];
  assign N4760 = N4759 | data_masked[3621];
  assign N4759 = N4758 | data_masked[3749];
  assign N4758 = N4757 | data_masked[3877];
  assign N4757 = N4756 | data_masked[4005];
  assign N4756 = N4755 | data_masked[4133];
  assign N4755 = N4754 | data_masked[4261];
  assign N4754 = N4753 | data_masked[4389];
  assign N4753 = N4752 | data_masked[4517];
  assign N4752 = N4751 | data_masked[4645];
  assign N4751 = N4750 | data_masked[4773];
  assign N4750 = N4749 | data_masked[4901];
  assign N4749 = N4748 | data_masked[5029];
  assign N4748 = N4747 | data_masked[5157];
  assign N4747 = N4746 | data_masked[5285];
  assign N4746 = N4745 | data_masked[5413];
  assign N4745 = N4744 | data_masked[5541];
  assign N4744 = N4743 | data_masked[5669];
  assign N4743 = N4742 | data_masked[5797];
  assign N4742 = N4741 | data_masked[5925];
  assign N4741 = N4740 | data_masked[6053];
  assign N4740 = N4739 | data_masked[6181];
  assign N4739 = N4738 | data_masked[6309];
  assign N4738 = N4737 | data_masked[6437];
  assign N4737 = N4736 | data_masked[6565];
  assign N4736 = N4735 | data_masked[6693];
  assign N4735 = N4734 | data_masked[6821];
  assign N4734 = N4733 | data_masked[6949];
  assign N4733 = N4732 | data_masked[7077];
  assign N4732 = N4731 | data_masked[7205];
  assign N4731 = N4730 | data_masked[7333];
  assign N4730 = N4729 | data_masked[7461];
  assign N4729 = N4728 | data_masked[7589];
  assign N4728 = N4727 | data_masked[7717];
  assign N4727 = N4726 | data_masked[7845];
  assign N4726 = N4725 | data_masked[7973];
  assign N4725 = N4724 | data_masked[8101];
  assign N4724 = N4723 | data_masked[8229];
  assign N4723 = N4722 | data_masked[8357];
  assign N4722 = N4721 | data_masked[8485];
  assign N4721 = N4720 | data_masked[8613];
  assign N4720 = N4719 | data_masked[8741];
  assign N4719 = N4718 | data_masked[8869];
  assign N4718 = N4717 | data_masked[8997];
  assign N4717 = N4716 | data_masked[9125];
  assign N4716 = N4715 | data_masked[9253];
  assign N4715 = N4714 | data_masked[9381];
  assign N4714 = N4713 | data_masked[9509];
  assign N4713 = N4712 | data_masked[9637];
  assign N4712 = N4711 | data_masked[9765];
  assign N4711 = N4710 | data_masked[9893];
  assign N4710 = N4709 | data_masked[10021];
  assign N4709 = N4708 | data_masked[10149];
  assign N4708 = N4707 | data_masked[10277];
  assign N4707 = N4706 | data_masked[10405];
  assign N4706 = N4705 | data_masked[10533];
  assign N4705 = N4704 | data_masked[10661];
  assign N4704 = N4703 | data_masked[10789];
  assign N4703 = N4702 | data_masked[10917];
  assign N4702 = N4701 | data_masked[11045];
  assign N4701 = N4700 | data_masked[11173];
  assign N4700 = N4699 | data_masked[11301];
  assign N4699 = N4698 | data_masked[11429];
  assign N4698 = N4697 | data_masked[11557];
  assign N4697 = N4696 | data_masked[11685];
  assign N4696 = N4695 | data_masked[11813];
  assign N4695 = N4694 | data_masked[11941];
  assign N4694 = N4693 | data_masked[12069];
  assign N4693 = N4692 | data_masked[12197];
  assign N4692 = N4691 | data_masked[12325];
  assign N4691 = N4690 | data_masked[12453];
  assign N4690 = N4689 | data_masked[12581];
  assign N4689 = N4688 | data_masked[12709];
  assign N4688 = N4687 | data_masked[12837];
  assign N4687 = N4686 | data_masked[12965];
  assign N4686 = N4685 | data_masked[13093];
  assign N4685 = N4684 | data_masked[13221];
  assign N4684 = N4683 | data_masked[13349];
  assign N4683 = N4682 | data_masked[13477];
  assign N4682 = N4681 | data_masked[13605];
  assign N4681 = N4680 | data_masked[13733];
  assign N4680 = N4679 | data_masked[13861];
  assign N4679 = N4678 | data_masked[13989];
  assign N4678 = N4677 | data_masked[14117];
  assign N4677 = N4676 | data_masked[14245];
  assign N4676 = N4675 | data_masked[14373];
  assign N4675 = N4674 | data_masked[14501];
  assign N4674 = N4673 | data_masked[14629];
  assign N4673 = N4672 | data_masked[14757];
  assign N4672 = N4671 | data_masked[14885];
  assign N4671 = N4670 | data_masked[15013];
  assign N4670 = N4669 | data_masked[15141];
  assign N4669 = N4668 | data_masked[15269];
  assign N4668 = N4667 | data_masked[15397];
  assign N4667 = N4666 | data_masked[15525];
  assign N4666 = N4665 | data_masked[15653];
  assign N4665 = N4664 | data_masked[15781];
  assign N4664 = N4663 | data_masked[15909];
  assign N4663 = N4662 | data_masked[16037];
  assign N4662 = data_masked[16293] | data_masked[16165];
  assign data_o[38] = N4913 | data_masked[38];
  assign N4913 = N4912 | data_masked[166];
  assign N4912 = N4911 | data_masked[294];
  assign N4911 = N4910 | data_masked[422];
  assign N4910 = N4909 | data_masked[550];
  assign N4909 = N4908 | data_masked[678];
  assign N4908 = N4907 | data_masked[806];
  assign N4907 = N4906 | data_masked[934];
  assign N4906 = N4905 | data_masked[1062];
  assign N4905 = N4904 | data_masked[1190];
  assign N4904 = N4903 | data_masked[1318];
  assign N4903 = N4902 | data_masked[1446];
  assign N4902 = N4901 | data_masked[1574];
  assign N4901 = N4900 | data_masked[1702];
  assign N4900 = N4899 | data_masked[1830];
  assign N4899 = N4898 | data_masked[1958];
  assign N4898 = N4897 | data_masked[2086];
  assign N4897 = N4896 | data_masked[2214];
  assign N4896 = N4895 | data_masked[2342];
  assign N4895 = N4894 | data_masked[2470];
  assign N4894 = N4893 | data_masked[2598];
  assign N4893 = N4892 | data_masked[2726];
  assign N4892 = N4891 | data_masked[2854];
  assign N4891 = N4890 | data_masked[2982];
  assign N4890 = N4889 | data_masked[3110];
  assign N4889 = N4888 | data_masked[3238];
  assign N4888 = N4887 | data_masked[3366];
  assign N4887 = N4886 | data_masked[3494];
  assign N4886 = N4885 | data_masked[3622];
  assign N4885 = N4884 | data_masked[3750];
  assign N4884 = N4883 | data_masked[3878];
  assign N4883 = N4882 | data_masked[4006];
  assign N4882 = N4881 | data_masked[4134];
  assign N4881 = N4880 | data_masked[4262];
  assign N4880 = N4879 | data_masked[4390];
  assign N4879 = N4878 | data_masked[4518];
  assign N4878 = N4877 | data_masked[4646];
  assign N4877 = N4876 | data_masked[4774];
  assign N4876 = N4875 | data_masked[4902];
  assign N4875 = N4874 | data_masked[5030];
  assign N4874 = N4873 | data_masked[5158];
  assign N4873 = N4872 | data_masked[5286];
  assign N4872 = N4871 | data_masked[5414];
  assign N4871 = N4870 | data_masked[5542];
  assign N4870 = N4869 | data_masked[5670];
  assign N4869 = N4868 | data_masked[5798];
  assign N4868 = N4867 | data_masked[5926];
  assign N4867 = N4866 | data_masked[6054];
  assign N4866 = N4865 | data_masked[6182];
  assign N4865 = N4864 | data_masked[6310];
  assign N4864 = N4863 | data_masked[6438];
  assign N4863 = N4862 | data_masked[6566];
  assign N4862 = N4861 | data_masked[6694];
  assign N4861 = N4860 | data_masked[6822];
  assign N4860 = N4859 | data_masked[6950];
  assign N4859 = N4858 | data_masked[7078];
  assign N4858 = N4857 | data_masked[7206];
  assign N4857 = N4856 | data_masked[7334];
  assign N4856 = N4855 | data_masked[7462];
  assign N4855 = N4854 | data_masked[7590];
  assign N4854 = N4853 | data_masked[7718];
  assign N4853 = N4852 | data_masked[7846];
  assign N4852 = N4851 | data_masked[7974];
  assign N4851 = N4850 | data_masked[8102];
  assign N4850 = N4849 | data_masked[8230];
  assign N4849 = N4848 | data_masked[8358];
  assign N4848 = N4847 | data_masked[8486];
  assign N4847 = N4846 | data_masked[8614];
  assign N4846 = N4845 | data_masked[8742];
  assign N4845 = N4844 | data_masked[8870];
  assign N4844 = N4843 | data_masked[8998];
  assign N4843 = N4842 | data_masked[9126];
  assign N4842 = N4841 | data_masked[9254];
  assign N4841 = N4840 | data_masked[9382];
  assign N4840 = N4839 | data_masked[9510];
  assign N4839 = N4838 | data_masked[9638];
  assign N4838 = N4837 | data_masked[9766];
  assign N4837 = N4836 | data_masked[9894];
  assign N4836 = N4835 | data_masked[10022];
  assign N4835 = N4834 | data_masked[10150];
  assign N4834 = N4833 | data_masked[10278];
  assign N4833 = N4832 | data_masked[10406];
  assign N4832 = N4831 | data_masked[10534];
  assign N4831 = N4830 | data_masked[10662];
  assign N4830 = N4829 | data_masked[10790];
  assign N4829 = N4828 | data_masked[10918];
  assign N4828 = N4827 | data_masked[11046];
  assign N4827 = N4826 | data_masked[11174];
  assign N4826 = N4825 | data_masked[11302];
  assign N4825 = N4824 | data_masked[11430];
  assign N4824 = N4823 | data_masked[11558];
  assign N4823 = N4822 | data_masked[11686];
  assign N4822 = N4821 | data_masked[11814];
  assign N4821 = N4820 | data_masked[11942];
  assign N4820 = N4819 | data_masked[12070];
  assign N4819 = N4818 | data_masked[12198];
  assign N4818 = N4817 | data_masked[12326];
  assign N4817 = N4816 | data_masked[12454];
  assign N4816 = N4815 | data_masked[12582];
  assign N4815 = N4814 | data_masked[12710];
  assign N4814 = N4813 | data_masked[12838];
  assign N4813 = N4812 | data_masked[12966];
  assign N4812 = N4811 | data_masked[13094];
  assign N4811 = N4810 | data_masked[13222];
  assign N4810 = N4809 | data_masked[13350];
  assign N4809 = N4808 | data_masked[13478];
  assign N4808 = N4807 | data_masked[13606];
  assign N4807 = N4806 | data_masked[13734];
  assign N4806 = N4805 | data_masked[13862];
  assign N4805 = N4804 | data_masked[13990];
  assign N4804 = N4803 | data_masked[14118];
  assign N4803 = N4802 | data_masked[14246];
  assign N4802 = N4801 | data_masked[14374];
  assign N4801 = N4800 | data_masked[14502];
  assign N4800 = N4799 | data_masked[14630];
  assign N4799 = N4798 | data_masked[14758];
  assign N4798 = N4797 | data_masked[14886];
  assign N4797 = N4796 | data_masked[15014];
  assign N4796 = N4795 | data_masked[15142];
  assign N4795 = N4794 | data_masked[15270];
  assign N4794 = N4793 | data_masked[15398];
  assign N4793 = N4792 | data_masked[15526];
  assign N4792 = N4791 | data_masked[15654];
  assign N4791 = N4790 | data_masked[15782];
  assign N4790 = N4789 | data_masked[15910];
  assign N4789 = N4788 | data_masked[16038];
  assign N4788 = data_masked[16294] | data_masked[16166];
  assign data_o[39] = N5039 | data_masked[39];
  assign N5039 = N5038 | data_masked[167];
  assign N5038 = N5037 | data_masked[295];
  assign N5037 = N5036 | data_masked[423];
  assign N5036 = N5035 | data_masked[551];
  assign N5035 = N5034 | data_masked[679];
  assign N5034 = N5033 | data_masked[807];
  assign N5033 = N5032 | data_masked[935];
  assign N5032 = N5031 | data_masked[1063];
  assign N5031 = N5030 | data_masked[1191];
  assign N5030 = N5029 | data_masked[1319];
  assign N5029 = N5028 | data_masked[1447];
  assign N5028 = N5027 | data_masked[1575];
  assign N5027 = N5026 | data_masked[1703];
  assign N5026 = N5025 | data_masked[1831];
  assign N5025 = N5024 | data_masked[1959];
  assign N5024 = N5023 | data_masked[2087];
  assign N5023 = N5022 | data_masked[2215];
  assign N5022 = N5021 | data_masked[2343];
  assign N5021 = N5020 | data_masked[2471];
  assign N5020 = N5019 | data_masked[2599];
  assign N5019 = N5018 | data_masked[2727];
  assign N5018 = N5017 | data_masked[2855];
  assign N5017 = N5016 | data_masked[2983];
  assign N5016 = N5015 | data_masked[3111];
  assign N5015 = N5014 | data_masked[3239];
  assign N5014 = N5013 | data_masked[3367];
  assign N5013 = N5012 | data_masked[3495];
  assign N5012 = N5011 | data_masked[3623];
  assign N5011 = N5010 | data_masked[3751];
  assign N5010 = N5009 | data_masked[3879];
  assign N5009 = N5008 | data_masked[4007];
  assign N5008 = N5007 | data_masked[4135];
  assign N5007 = N5006 | data_masked[4263];
  assign N5006 = N5005 | data_masked[4391];
  assign N5005 = N5004 | data_masked[4519];
  assign N5004 = N5003 | data_masked[4647];
  assign N5003 = N5002 | data_masked[4775];
  assign N5002 = N5001 | data_masked[4903];
  assign N5001 = N5000 | data_masked[5031];
  assign N5000 = N4999 | data_masked[5159];
  assign N4999 = N4998 | data_masked[5287];
  assign N4998 = N4997 | data_masked[5415];
  assign N4997 = N4996 | data_masked[5543];
  assign N4996 = N4995 | data_masked[5671];
  assign N4995 = N4994 | data_masked[5799];
  assign N4994 = N4993 | data_masked[5927];
  assign N4993 = N4992 | data_masked[6055];
  assign N4992 = N4991 | data_masked[6183];
  assign N4991 = N4990 | data_masked[6311];
  assign N4990 = N4989 | data_masked[6439];
  assign N4989 = N4988 | data_masked[6567];
  assign N4988 = N4987 | data_masked[6695];
  assign N4987 = N4986 | data_masked[6823];
  assign N4986 = N4985 | data_masked[6951];
  assign N4985 = N4984 | data_masked[7079];
  assign N4984 = N4983 | data_masked[7207];
  assign N4983 = N4982 | data_masked[7335];
  assign N4982 = N4981 | data_masked[7463];
  assign N4981 = N4980 | data_masked[7591];
  assign N4980 = N4979 | data_masked[7719];
  assign N4979 = N4978 | data_masked[7847];
  assign N4978 = N4977 | data_masked[7975];
  assign N4977 = N4976 | data_masked[8103];
  assign N4976 = N4975 | data_masked[8231];
  assign N4975 = N4974 | data_masked[8359];
  assign N4974 = N4973 | data_masked[8487];
  assign N4973 = N4972 | data_masked[8615];
  assign N4972 = N4971 | data_masked[8743];
  assign N4971 = N4970 | data_masked[8871];
  assign N4970 = N4969 | data_masked[8999];
  assign N4969 = N4968 | data_masked[9127];
  assign N4968 = N4967 | data_masked[9255];
  assign N4967 = N4966 | data_masked[9383];
  assign N4966 = N4965 | data_masked[9511];
  assign N4965 = N4964 | data_masked[9639];
  assign N4964 = N4963 | data_masked[9767];
  assign N4963 = N4962 | data_masked[9895];
  assign N4962 = N4961 | data_masked[10023];
  assign N4961 = N4960 | data_masked[10151];
  assign N4960 = N4959 | data_masked[10279];
  assign N4959 = N4958 | data_masked[10407];
  assign N4958 = N4957 | data_masked[10535];
  assign N4957 = N4956 | data_masked[10663];
  assign N4956 = N4955 | data_masked[10791];
  assign N4955 = N4954 | data_masked[10919];
  assign N4954 = N4953 | data_masked[11047];
  assign N4953 = N4952 | data_masked[11175];
  assign N4952 = N4951 | data_masked[11303];
  assign N4951 = N4950 | data_masked[11431];
  assign N4950 = N4949 | data_masked[11559];
  assign N4949 = N4948 | data_masked[11687];
  assign N4948 = N4947 | data_masked[11815];
  assign N4947 = N4946 | data_masked[11943];
  assign N4946 = N4945 | data_masked[12071];
  assign N4945 = N4944 | data_masked[12199];
  assign N4944 = N4943 | data_masked[12327];
  assign N4943 = N4942 | data_masked[12455];
  assign N4942 = N4941 | data_masked[12583];
  assign N4941 = N4940 | data_masked[12711];
  assign N4940 = N4939 | data_masked[12839];
  assign N4939 = N4938 | data_masked[12967];
  assign N4938 = N4937 | data_masked[13095];
  assign N4937 = N4936 | data_masked[13223];
  assign N4936 = N4935 | data_masked[13351];
  assign N4935 = N4934 | data_masked[13479];
  assign N4934 = N4933 | data_masked[13607];
  assign N4933 = N4932 | data_masked[13735];
  assign N4932 = N4931 | data_masked[13863];
  assign N4931 = N4930 | data_masked[13991];
  assign N4930 = N4929 | data_masked[14119];
  assign N4929 = N4928 | data_masked[14247];
  assign N4928 = N4927 | data_masked[14375];
  assign N4927 = N4926 | data_masked[14503];
  assign N4926 = N4925 | data_masked[14631];
  assign N4925 = N4924 | data_masked[14759];
  assign N4924 = N4923 | data_masked[14887];
  assign N4923 = N4922 | data_masked[15015];
  assign N4922 = N4921 | data_masked[15143];
  assign N4921 = N4920 | data_masked[15271];
  assign N4920 = N4919 | data_masked[15399];
  assign N4919 = N4918 | data_masked[15527];
  assign N4918 = N4917 | data_masked[15655];
  assign N4917 = N4916 | data_masked[15783];
  assign N4916 = N4915 | data_masked[15911];
  assign N4915 = N4914 | data_masked[16039];
  assign N4914 = data_masked[16295] | data_masked[16167];
  assign data_o[40] = N5165 | data_masked[40];
  assign N5165 = N5164 | data_masked[168];
  assign N5164 = N5163 | data_masked[296];
  assign N5163 = N5162 | data_masked[424];
  assign N5162 = N5161 | data_masked[552];
  assign N5161 = N5160 | data_masked[680];
  assign N5160 = N5159 | data_masked[808];
  assign N5159 = N5158 | data_masked[936];
  assign N5158 = N5157 | data_masked[1064];
  assign N5157 = N5156 | data_masked[1192];
  assign N5156 = N5155 | data_masked[1320];
  assign N5155 = N5154 | data_masked[1448];
  assign N5154 = N5153 | data_masked[1576];
  assign N5153 = N5152 | data_masked[1704];
  assign N5152 = N5151 | data_masked[1832];
  assign N5151 = N5150 | data_masked[1960];
  assign N5150 = N5149 | data_masked[2088];
  assign N5149 = N5148 | data_masked[2216];
  assign N5148 = N5147 | data_masked[2344];
  assign N5147 = N5146 | data_masked[2472];
  assign N5146 = N5145 | data_masked[2600];
  assign N5145 = N5144 | data_masked[2728];
  assign N5144 = N5143 | data_masked[2856];
  assign N5143 = N5142 | data_masked[2984];
  assign N5142 = N5141 | data_masked[3112];
  assign N5141 = N5140 | data_masked[3240];
  assign N5140 = N5139 | data_masked[3368];
  assign N5139 = N5138 | data_masked[3496];
  assign N5138 = N5137 | data_masked[3624];
  assign N5137 = N5136 | data_masked[3752];
  assign N5136 = N5135 | data_masked[3880];
  assign N5135 = N5134 | data_masked[4008];
  assign N5134 = N5133 | data_masked[4136];
  assign N5133 = N5132 | data_masked[4264];
  assign N5132 = N5131 | data_masked[4392];
  assign N5131 = N5130 | data_masked[4520];
  assign N5130 = N5129 | data_masked[4648];
  assign N5129 = N5128 | data_masked[4776];
  assign N5128 = N5127 | data_masked[4904];
  assign N5127 = N5126 | data_masked[5032];
  assign N5126 = N5125 | data_masked[5160];
  assign N5125 = N5124 | data_masked[5288];
  assign N5124 = N5123 | data_masked[5416];
  assign N5123 = N5122 | data_masked[5544];
  assign N5122 = N5121 | data_masked[5672];
  assign N5121 = N5120 | data_masked[5800];
  assign N5120 = N5119 | data_masked[5928];
  assign N5119 = N5118 | data_masked[6056];
  assign N5118 = N5117 | data_masked[6184];
  assign N5117 = N5116 | data_masked[6312];
  assign N5116 = N5115 | data_masked[6440];
  assign N5115 = N5114 | data_masked[6568];
  assign N5114 = N5113 | data_masked[6696];
  assign N5113 = N5112 | data_masked[6824];
  assign N5112 = N5111 | data_masked[6952];
  assign N5111 = N5110 | data_masked[7080];
  assign N5110 = N5109 | data_masked[7208];
  assign N5109 = N5108 | data_masked[7336];
  assign N5108 = N5107 | data_masked[7464];
  assign N5107 = N5106 | data_masked[7592];
  assign N5106 = N5105 | data_masked[7720];
  assign N5105 = N5104 | data_masked[7848];
  assign N5104 = N5103 | data_masked[7976];
  assign N5103 = N5102 | data_masked[8104];
  assign N5102 = N5101 | data_masked[8232];
  assign N5101 = N5100 | data_masked[8360];
  assign N5100 = N5099 | data_masked[8488];
  assign N5099 = N5098 | data_masked[8616];
  assign N5098 = N5097 | data_masked[8744];
  assign N5097 = N5096 | data_masked[8872];
  assign N5096 = N5095 | data_masked[9000];
  assign N5095 = N5094 | data_masked[9128];
  assign N5094 = N5093 | data_masked[9256];
  assign N5093 = N5092 | data_masked[9384];
  assign N5092 = N5091 | data_masked[9512];
  assign N5091 = N5090 | data_masked[9640];
  assign N5090 = N5089 | data_masked[9768];
  assign N5089 = N5088 | data_masked[9896];
  assign N5088 = N5087 | data_masked[10024];
  assign N5087 = N5086 | data_masked[10152];
  assign N5086 = N5085 | data_masked[10280];
  assign N5085 = N5084 | data_masked[10408];
  assign N5084 = N5083 | data_masked[10536];
  assign N5083 = N5082 | data_masked[10664];
  assign N5082 = N5081 | data_masked[10792];
  assign N5081 = N5080 | data_masked[10920];
  assign N5080 = N5079 | data_masked[11048];
  assign N5079 = N5078 | data_masked[11176];
  assign N5078 = N5077 | data_masked[11304];
  assign N5077 = N5076 | data_masked[11432];
  assign N5076 = N5075 | data_masked[11560];
  assign N5075 = N5074 | data_masked[11688];
  assign N5074 = N5073 | data_masked[11816];
  assign N5073 = N5072 | data_masked[11944];
  assign N5072 = N5071 | data_masked[12072];
  assign N5071 = N5070 | data_masked[12200];
  assign N5070 = N5069 | data_masked[12328];
  assign N5069 = N5068 | data_masked[12456];
  assign N5068 = N5067 | data_masked[12584];
  assign N5067 = N5066 | data_masked[12712];
  assign N5066 = N5065 | data_masked[12840];
  assign N5065 = N5064 | data_masked[12968];
  assign N5064 = N5063 | data_masked[13096];
  assign N5063 = N5062 | data_masked[13224];
  assign N5062 = N5061 | data_masked[13352];
  assign N5061 = N5060 | data_masked[13480];
  assign N5060 = N5059 | data_masked[13608];
  assign N5059 = N5058 | data_masked[13736];
  assign N5058 = N5057 | data_masked[13864];
  assign N5057 = N5056 | data_masked[13992];
  assign N5056 = N5055 | data_masked[14120];
  assign N5055 = N5054 | data_masked[14248];
  assign N5054 = N5053 | data_masked[14376];
  assign N5053 = N5052 | data_masked[14504];
  assign N5052 = N5051 | data_masked[14632];
  assign N5051 = N5050 | data_masked[14760];
  assign N5050 = N5049 | data_masked[14888];
  assign N5049 = N5048 | data_masked[15016];
  assign N5048 = N5047 | data_masked[15144];
  assign N5047 = N5046 | data_masked[15272];
  assign N5046 = N5045 | data_masked[15400];
  assign N5045 = N5044 | data_masked[15528];
  assign N5044 = N5043 | data_masked[15656];
  assign N5043 = N5042 | data_masked[15784];
  assign N5042 = N5041 | data_masked[15912];
  assign N5041 = N5040 | data_masked[16040];
  assign N5040 = data_masked[16296] | data_masked[16168];
  assign data_o[41] = N5291 | data_masked[41];
  assign N5291 = N5290 | data_masked[169];
  assign N5290 = N5289 | data_masked[297];
  assign N5289 = N5288 | data_masked[425];
  assign N5288 = N5287 | data_masked[553];
  assign N5287 = N5286 | data_masked[681];
  assign N5286 = N5285 | data_masked[809];
  assign N5285 = N5284 | data_masked[937];
  assign N5284 = N5283 | data_masked[1065];
  assign N5283 = N5282 | data_masked[1193];
  assign N5282 = N5281 | data_masked[1321];
  assign N5281 = N5280 | data_masked[1449];
  assign N5280 = N5279 | data_masked[1577];
  assign N5279 = N5278 | data_masked[1705];
  assign N5278 = N5277 | data_masked[1833];
  assign N5277 = N5276 | data_masked[1961];
  assign N5276 = N5275 | data_masked[2089];
  assign N5275 = N5274 | data_masked[2217];
  assign N5274 = N5273 | data_masked[2345];
  assign N5273 = N5272 | data_masked[2473];
  assign N5272 = N5271 | data_masked[2601];
  assign N5271 = N5270 | data_masked[2729];
  assign N5270 = N5269 | data_masked[2857];
  assign N5269 = N5268 | data_masked[2985];
  assign N5268 = N5267 | data_masked[3113];
  assign N5267 = N5266 | data_masked[3241];
  assign N5266 = N5265 | data_masked[3369];
  assign N5265 = N5264 | data_masked[3497];
  assign N5264 = N5263 | data_masked[3625];
  assign N5263 = N5262 | data_masked[3753];
  assign N5262 = N5261 | data_masked[3881];
  assign N5261 = N5260 | data_masked[4009];
  assign N5260 = N5259 | data_masked[4137];
  assign N5259 = N5258 | data_masked[4265];
  assign N5258 = N5257 | data_masked[4393];
  assign N5257 = N5256 | data_masked[4521];
  assign N5256 = N5255 | data_masked[4649];
  assign N5255 = N5254 | data_masked[4777];
  assign N5254 = N5253 | data_masked[4905];
  assign N5253 = N5252 | data_masked[5033];
  assign N5252 = N5251 | data_masked[5161];
  assign N5251 = N5250 | data_masked[5289];
  assign N5250 = N5249 | data_masked[5417];
  assign N5249 = N5248 | data_masked[5545];
  assign N5248 = N5247 | data_masked[5673];
  assign N5247 = N5246 | data_masked[5801];
  assign N5246 = N5245 | data_masked[5929];
  assign N5245 = N5244 | data_masked[6057];
  assign N5244 = N5243 | data_masked[6185];
  assign N5243 = N5242 | data_masked[6313];
  assign N5242 = N5241 | data_masked[6441];
  assign N5241 = N5240 | data_masked[6569];
  assign N5240 = N5239 | data_masked[6697];
  assign N5239 = N5238 | data_masked[6825];
  assign N5238 = N5237 | data_masked[6953];
  assign N5237 = N5236 | data_masked[7081];
  assign N5236 = N5235 | data_masked[7209];
  assign N5235 = N5234 | data_masked[7337];
  assign N5234 = N5233 | data_masked[7465];
  assign N5233 = N5232 | data_masked[7593];
  assign N5232 = N5231 | data_masked[7721];
  assign N5231 = N5230 | data_masked[7849];
  assign N5230 = N5229 | data_masked[7977];
  assign N5229 = N5228 | data_masked[8105];
  assign N5228 = N5227 | data_masked[8233];
  assign N5227 = N5226 | data_masked[8361];
  assign N5226 = N5225 | data_masked[8489];
  assign N5225 = N5224 | data_masked[8617];
  assign N5224 = N5223 | data_masked[8745];
  assign N5223 = N5222 | data_masked[8873];
  assign N5222 = N5221 | data_masked[9001];
  assign N5221 = N5220 | data_masked[9129];
  assign N5220 = N5219 | data_masked[9257];
  assign N5219 = N5218 | data_masked[9385];
  assign N5218 = N5217 | data_masked[9513];
  assign N5217 = N5216 | data_masked[9641];
  assign N5216 = N5215 | data_masked[9769];
  assign N5215 = N5214 | data_masked[9897];
  assign N5214 = N5213 | data_masked[10025];
  assign N5213 = N5212 | data_masked[10153];
  assign N5212 = N5211 | data_masked[10281];
  assign N5211 = N5210 | data_masked[10409];
  assign N5210 = N5209 | data_masked[10537];
  assign N5209 = N5208 | data_masked[10665];
  assign N5208 = N5207 | data_masked[10793];
  assign N5207 = N5206 | data_masked[10921];
  assign N5206 = N5205 | data_masked[11049];
  assign N5205 = N5204 | data_masked[11177];
  assign N5204 = N5203 | data_masked[11305];
  assign N5203 = N5202 | data_masked[11433];
  assign N5202 = N5201 | data_masked[11561];
  assign N5201 = N5200 | data_masked[11689];
  assign N5200 = N5199 | data_masked[11817];
  assign N5199 = N5198 | data_masked[11945];
  assign N5198 = N5197 | data_masked[12073];
  assign N5197 = N5196 | data_masked[12201];
  assign N5196 = N5195 | data_masked[12329];
  assign N5195 = N5194 | data_masked[12457];
  assign N5194 = N5193 | data_masked[12585];
  assign N5193 = N5192 | data_masked[12713];
  assign N5192 = N5191 | data_masked[12841];
  assign N5191 = N5190 | data_masked[12969];
  assign N5190 = N5189 | data_masked[13097];
  assign N5189 = N5188 | data_masked[13225];
  assign N5188 = N5187 | data_masked[13353];
  assign N5187 = N5186 | data_masked[13481];
  assign N5186 = N5185 | data_masked[13609];
  assign N5185 = N5184 | data_masked[13737];
  assign N5184 = N5183 | data_masked[13865];
  assign N5183 = N5182 | data_masked[13993];
  assign N5182 = N5181 | data_masked[14121];
  assign N5181 = N5180 | data_masked[14249];
  assign N5180 = N5179 | data_masked[14377];
  assign N5179 = N5178 | data_masked[14505];
  assign N5178 = N5177 | data_masked[14633];
  assign N5177 = N5176 | data_masked[14761];
  assign N5176 = N5175 | data_masked[14889];
  assign N5175 = N5174 | data_masked[15017];
  assign N5174 = N5173 | data_masked[15145];
  assign N5173 = N5172 | data_masked[15273];
  assign N5172 = N5171 | data_masked[15401];
  assign N5171 = N5170 | data_masked[15529];
  assign N5170 = N5169 | data_masked[15657];
  assign N5169 = N5168 | data_masked[15785];
  assign N5168 = N5167 | data_masked[15913];
  assign N5167 = N5166 | data_masked[16041];
  assign N5166 = data_masked[16297] | data_masked[16169];
  assign data_o[42] = N5417 | data_masked[42];
  assign N5417 = N5416 | data_masked[170];
  assign N5416 = N5415 | data_masked[298];
  assign N5415 = N5414 | data_masked[426];
  assign N5414 = N5413 | data_masked[554];
  assign N5413 = N5412 | data_masked[682];
  assign N5412 = N5411 | data_masked[810];
  assign N5411 = N5410 | data_masked[938];
  assign N5410 = N5409 | data_masked[1066];
  assign N5409 = N5408 | data_masked[1194];
  assign N5408 = N5407 | data_masked[1322];
  assign N5407 = N5406 | data_masked[1450];
  assign N5406 = N5405 | data_masked[1578];
  assign N5405 = N5404 | data_masked[1706];
  assign N5404 = N5403 | data_masked[1834];
  assign N5403 = N5402 | data_masked[1962];
  assign N5402 = N5401 | data_masked[2090];
  assign N5401 = N5400 | data_masked[2218];
  assign N5400 = N5399 | data_masked[2346];
  assign N5399 = N5398 | data_masked[2474];
  assign N5398 = N5397 | data_masked[2602];
  assign N5397 = N5396 | data_masked[2730];
  assign N5396 = N5395 | data_masked[2858];
  assign N5395 = N5394 | data_masked[2986];
  assign N5394 = N5393 | data_masked[3114];
  assign N5393 = N5392 | data_masked[3242];
  assign N5392 = N5391 | data_masked[3370];
  assign N5391 = N5390 | data_masked[3498];
  assign N5390 = N5389 | data_masked[3626];
  assign N5389 = N5388 | data_masked[3754];
  assign N5388 = N5387 | data_masked[3882];
  assign N5387 = N5386 | data_masked[4010];
  assign N5386 = N5385 | data_masked[4138];
  assign N5385 = N5384 | data_masked[4266];
  assign N5384 = N5383 | data_masked[4394];
  assign N5383 = N5382 | data_masked[4522];
  assign N5382 = N5381 | data_masked[4650];
  assign N5381 = N5380 | data_masked[4778];
  assign N5380 = N5379 | data_masked[4906];
  assign N5379 = N5378 | data_masked[5034];
  assign N5378 = N5377 | data_masked[5162];
  assign N5377 = N5376 | data_masked[5290];
  assign N5376 = N5375 | data_masked[5418];
  assign N5375 = N5374 | data_masked[5546];
  assign N5374 = N5373 | data_masked[5674];
  assign N5373 = N5372 | data_masked[5802];
  assign N5372 = N5371 | data_masked[5930];
  assign N5371 = N5370 | data_masked[6058];
  assign N5370 = N5369 | data_masked[6186];
  assign N5369 = N5368 | data_masked[6314];
  assign N5368 = N5367 | data_masked[6442];
  assign N5367 = N5366 | data_masked[6570];
  assign N5366 = N5365 | data_masked[6698];
  assign N5365 = N5364 | data_masked[6826];
  assign N5364 = N5363 | data_masked[6954];
  assign N5363 = N5362 | data_masked[7082];
  assign N5362 = N5361 | data_masked[7210];
  assign N5361 = N5360 | data_masked[7338];
  assign N5360 = N5359 | data_masked[7466];
  assign N5359 = N5358 | data_masked[7594];
  assign N5358 = N5357 | data_masked[7722];
  assign N5357 = N5356 | data_masked[7850];
  assign N5356 = N5355 | data_masked[7978];
  assign N5355 = N5354 | data_masked[8106];
  assign N5354 = N5353 | data_masked[8234];
  assign N5353 = N5352 | data_masked[8362];
  assign N5352 = N5351 | data_masked[8490];
  assign N5351 = N5350 | data_masked[8618];
  assign N5350 = N5349 | data_masked[8746];
  assign N5349 = N5348 | data_masked[8874];
  assign N5348 = N5347 | data_masked[9002];
  assign N5347 = N5346 | data_masked[9130];
  assign N5346 = N5345 | data_masked[9258];
  assign N5345 = N5344 | data_masked[9386];
  assign N5344 = N5343 | data_masked[9514];
  assign N5343 = N5342 | data_masked[9642];
  assign N5342 = N5341 | data_masked[9770];
  assign N5341 = N5340 | data_masked[9898];
  assign N5340 = N5339 | data_masked[10026];
  assign N5339 = N5338 | data_masked[10154];
  assign N5338 = N5337 | data_masked[10282];
  assign N5337 = N5336 | data_masked[10410];
  assign N5336 = N5335 | data_masked[10538];
  assign N5335 = N5334 | data_masked[10666];
  assign N5334 = N5333 | data_masked[10794];
  assign N5333 = N5332 | data_masked[10922];
  assign N5332 = N5331 | data_masked[11050];
  assign N5331 = N5330 | data_masked[11178];
  assign N5330 = N5329 | data_masked[11306];
  assign N5329 = N5328 | data_masked[11434];
  assign N5328 = N5327 | data_masked[11562];
  assign N5327 = N5326 | data_masked[11690];
  assign N5326 = N5325 | data_masked[11818];
  assign N5325 = N5324 | data_masked[11946];
  assign N5324 = N5323 | data_masked[12074];
  assign N5323 = N5322 | data_masked[12202];
  assign N5322 = N5321 | data_masked[12330];
  assign N5321 = N5320 | data_masked[12458];
  assign N5320 = N5319 | data_masked[12586];
  assign N5319 = N5318 | data_masked[12714];
  assign N5318 = N5317 | data_masked[12842];
  assign N5317 = N5316 | data_masked[12970];
  assign N5316 = N5315 | data_masked[13098];
  assign N5315 = N5314 | data_masked[13226];
  assign N5314 = N5313 | data_masked[13354];
  assign N5313 = N5312 | data_masked[13482];
  assign N5312 = N5311 | data_masked[13610];
  assign N5311 = N5310 | data_masked[13738];
  assign N5310 = N5309 | data_masked[13866];
  assign N5309 = N5308 | data_masked[13994];
  assign N5308 = N5307 | data_masked[14122];
  assign N5307 = N5306 | data_masked[14250];
  assign N5306 = N5305 | data_masked[14378];
  assign N5305 = N5304 | data_masked[14506];
  assign N5304 = N5303 | data_masked[14634];
  assign N5303 = N5302 | data_masked[14762];
  assign N5302 = N5301 | data_masked[14890];
  assign N5301 = N5300 | data_masked[15018];
  assign N5300 = N5299 | data_masked[15146];
  assign N5299 = N5298 | data_masked[15274];
  assign N5298 = N5297 | data_masked[15402];
  assign N5297 = N5296 | data_masked[15530];
  assign N5296 = N5295 | data_masked[15658];
  assign N5295 = N5294 | data_masked[15786];
  assign N5294 = N5293 | data_masked[15914];
  assign N5293 = N5292 | data_masked[16042];
  assign N5292 = data_masked[16298] | data_masked[16170];
  assign data_o[43] = N5543 | data_masked[43];
  assign N5543 = N5542 | data_masked[171];
  assign N5542 = N5541 | data_masked[299];
  assign N5541 = N5540 | data_masked[427];
  assign N5540 = N5539 | data_masked[555];
  assign N5539 = N5538 | data_masked[683];
  assign N5538 = N5537 | data_masked[811];
  assign N5537 = N5536 | data_masked[939];
  assign N5536 = N5535 | data_masked[1067];
  assign N5535 = N5534 | data_masked[1195];
  assign N5534 = N5533 | data_masked[1323];
  assign N5533 = N5532 | data_masked[1451];
  assign N5532 = N5531 | data_masked[1579];
  assign N5531 = N5530 | data_masked[1707];
  assign N5530 = N5529 | data_masked[1835];
  assign N5529 = N5528 | data_masked[1963];
  assign N5528 = N5527 | data_masked[2091];
  assign N5527 = N5526 | data_masked[2219];
  assign N5526 = N5525 | data_masked[2347];
  assign N5525 = N5524 | data_masked[2475];
  assign N5524 = N5523 | data_masked[2603];
  assign N5523 = N5522 | data_masked[2731];
  assign N5522 = N5521 | data_masked[2859];
  assign N5521 = N5520 | data_masked[2987];
  assign N5520 = N5519 | data_masked[3115];
  assign N5519 = N5518 | data_masked[3243];
  assign N5518 = N5517 | data_masked[3371];
  assign N5517 = N5516 | data_masked[3499];
  assign N5516 = N5515 | data_masked[3627];
  assign N5515 = N5514 | data_masked[3755];
  assign N5514 = N5513 | data_masked[3883];
  assign N5513 = N5512 | data_masked[4011];
  assign N5512 = N5511 | data_masked[4139];
  assign N5511 = N5510 | data_masked[4267];
  assign N5510 = N5509 | data_masked[4395];
  assign N5509 = N5508 | data_masked[4523];
  assign N5508 = N5507 | data_masked[4651];
  assign N5507 = N5506 | data_masked[4779];
  assign N5506 = N5505 | data_masked[4907];
  assign N5505 = N5504 | data_masked[5035];
  assign N5504 = N5503 | data_masked[5163];
  assign N5503 = N5502 | data_masked[5291];
  assign N5502 = N5501 | data_masked[5419];
  assign N5501 = N5500 | data_masked[5547];
  assign N5500 = N5499 | data_masked[5675];
  assign N5499 = N5498 | data_masked[5803];
  assign N5498 = N5497 | data_masked[5931];
  assign N5497 = N5496 | data_masked[6059];
  assign N5496 = N5495 | data_masked[6187];
  assign N5495 = N5494 | data_masked[6315];
  assign N5494 = N5493 | data_masked[6443];
  assign N5493 = N5492 | data_masked[6571];
  assign N5492 = N5491 | data_masked[6699];
  assign N5491 = N5490 | data_masked[6827];
  assign N5490 = N5489 | data_masked[6955];
  assign N5489 = N5488 | data_masked[7083];
  assign N5488 = N5487 | data_masked[7211];
  assign N5487 = N5486 | data_masked[7339];
  assign N5486 = N5485 | data_masked[7467];
  assign N5485 = N5484 | data_masked[7595];
  assign N5484 = N5483 | data_masked[7723];
  assign N5483 = N5482 | data_masked[7851];
  assign N5482 = N5481 | data_masked[7979];
  assign N5481 = N5480 | data_masked[8107];
  assign N5480 = N5479 | data_masked[8235];
  assign N5479 = N5478 | data_masked[8363];
  assign N5478 = N5477 | data_masked[8491];
  assign N5477 = N5476 | data_masked[8619];
  assign N5476 = N5475 | data_masked[8747];
  assign N5475 = N5474 | data_masked[8875];
  assign N5474 = N5473 | data_masked[9003];
  assign N5473 = N5472 | data_masked[9131];
  assign N5472 = N5471 | data_masked[9259];
  assign N5471 = N5470 | data_masked[9387];
  assign N5470 = N5469 | data_masked[9515];
  assign N5469 = N5468 | data_masked[9643];
  assign N5468 = N5467 | data_masked[9771];
  assign N5467 = N5466 | data_masked[9899];
  assign N5466 = N5465 | data_masked[10027];
  assign N5465 = N5464 | data_masked[10155];
  assign N5464 = N5463 | data_masked[10283];
  assign N5463 = N5462 | data_masked[10411];
  assign N5462 = N5461 | data_masked[10539];
  assign N5461 = N5460 | data_masked[10667];
  assign N5460 = N5459 | data_masked[10795];
  assign N5459 = N5458 | data_masked[10923];
  assign N5458 = N5457 | data_masked[11051];
  assign N5457 = N5456 | data_masked[11179];
  assign N5456 = N5455 | data_masked[11307];
  assign N5455 = N5454 | data_masked[11435];
  assign N5454 = N5453 | data_masked[11563];
  assign N5453 = N5452 | data_masked[11691];
  assign N5452 = N5451 | data_masked[11819];
  assign N5451 = N5450 | data_masked[11947];
  assign N5450 = N5449 | data_masked[12075];
  assign N5449 = N5448 | data_masked[12203];
  assign N5448 = N5447 | data_masked[12331];
  assign N5447 = N5446 | data_masked[12459];
  assign N5446 = N5445 | data_masked[12587];
  assign N5445 = N5444 | data_masked[12715];
  assign N5444 = N5443 | data_masked[12843];
  assign N5443 = N5442 | data_masked[12971];
  assign N5442 = N5441 | data_masked[13099];
  assign N5441 = N5440 | data_masked[13227];
  assign N5440 = N5439 | data_masked[13355];
  assign N5439 = N5438 | data_masked[13483];
  assign N5438 = N5437 | data_masked[13611];
  assign N5437 = N5436 | data_masked[13739];
  assign N5436 = N5435 | data_masked[13867];
  assign N5435 = N5434 | data_masked[13995];
  assign N5434 = N5433 | data_masked[14123];
  assign N5433 = N5432 | data_masked[14251];
  assign N5432 = N5431 | data_masked[14379];
  assign N5431 = N5430 | data_masked[14507];
  assign N5430 = N5429 | data_masked[14635];
  assign N5429 = N5428 | data_masked[14763];
  assign N5428 = N5427 | data_masked[14891];
  assign N5427 = N5426 | data_masked[15019];
  assign N5426 = N5425 | data_masked[15147];
  assign N5425 = N5424 | data_masked[15275];
  assign N5424 = N5423 | data_masked[15403];
  assign N5423 = N5422 | data_masked[15531];
  assign N5422 = N5421 | data_masked[15659];
  assign N5421 = N5420 | data_masked[15787];
  assign N5420 = N5419 | data_masked[15915];
  assign N5419 = N5418 | data_masked[16043];
  assign N5418 = data_masked[16299] | data_masked[16171];
  assign data_o[44] = N5669 | data_masked[44];
  assign N5669 = N5668 | data_masked[172];
  assign N5668 = N5667 | data_masked[300];
  assign N5667 = N5666 | data_masked[428];
  assign N5666 = N5665 | data_masked[556];
  assign N5665 = N5664 | data_masked[684];
  assign N5664 = N5663 | data_masked[812];
  assign N5663 = N5662 | data_masked[940];
  assign N5662 = N5661 | data_masked[1068];
  assign N5661 = N5660 | data_masked[1196];
  assign N5660 = N5659 | data_masked[1324];
  assign N5659 = N5658 | data_masked[1452];
  assign N5658 = N5657 | data_masked[1580];
  assign N5657 = N5656 | data_masked[1708];
  assign N5656 = N5655 | data_masked[1836];
  assign N5655 = N5654 | data_masked[1964];
  assign N5654 = N5653 | data_masked[2092];
  assign N5653 = N5652 | data_masked[2220];
  assign N5652 = N5651 | data_masked[2348];
  assign N5651 = N5650 | data_masked[2476];
  assign N5650 = N5649 | data_masked[2604];
  assign N5649 = N5648 | data_masked[2732];
  assign N5648 = N5647 | data_masked[2860];
  assign N5647 = N5646 | data_masked[2988];
  assign N5646 = N5645 | data_masked[3116];
  assign N5645 = N5644 | data_masked[3244];
  assign N5644 = N5643 | data_masked[3372];
  assign N5643 = N5642 | data_masked[3500];
  assign N5642 = N5641 | data_masked[3628];
  assign N5641 = N5640 | data_masked[3756];
  assign N5640 = N5639 | data_masked[3884];
  assign N5639 = N5638 | data_masked[4012];
  assign N5638 = N5637 | data_masked[4140];
  assign N5637 = N5636 | data_masked[4268];
  assign N5636 = N5635 | data_masked[4396];
  assign N5635 = N5634 | data_masked[4524];
  assign N5634 = N5633 | data_masked[4652];
  assign N5633 = N5632 | data_masked[4780];
  assign N5632 = N5631 | data_masked[4908];
  assign N5631 = N5630 | data_masked[5036];
  assign N5630 = N5629 | data_masked[5164];
  assign N5629 = N5628 | data_masked[5292];
  assign N5628 = N5627 | data_masked[5420];
  assign N5627 = N5626 | data_masked[5548];
  assign N5626 = N5625 | data_masked[5676];
  assign N5625 = N5624 | data_masked[5804];
  assign N5624 = N5623 | data_masked[5932];
  assign N5623 = N5622 | data_masked[6060];
  assign N5622 = N5621 | data_masked[6188];
  assign N5621 = N5620 | data_masked[6316];
  assign N5620 = N5619 | data_masked[6444];
  assign N5619 = N5618 | data_masked[6572];
  assign N5618 = N5617 | data_masked[6700];
  assign N5617 = N5616 | data_masked[6828];
  assign N5616 = N5615 | data_masked[6956];
  assign N5615 = N5614 | data_masked[7084];
  assign N5614 = N5613 | data_masked[7212];
  assign N5613 = N5612 | data_masked[7340];
  assign N5612 = N5611 | data_masked[7468];
  assign N5611 = N5610 | data_masked[7596];
  assign N5610 = N5609 | data_masked[7724];
  assign N5609 = N5608 | data_masked[7852];
  assign N5608 = N5607 | data_masked[7980];
  assign N5607 = N5606 | data_masked[8108];
  assign N5606 = N5605 | data_masked[8236];
  assign N5605 = N5604 | data_masked[8364];
  assign N5604 = N5603 | data_masked[8492];
  assign N5603 = N5602 | data_masked[8620];
  assign N5602 = N5601 | data_masked[8748];
  assign N5601 = N5600 | data_masked[8876];
  assign N5600 = N5599 | data_masked[9004];
  assign N5599 = N5598 | data_masked[9132];
  assign N5598 = N5597 | data_masked[9260];
  assign N5597 = N5596 | data_masked[9388];
  assign N5596 = N5595 | data_masked[9516];
  assign N5595 = N5594 | data_masked[9644];
  assign N5594 = N5593 | data_masked[9772];
  assign N5593 = N5592 | data_masked[9900];
  assign N5592 = N5591 | data_masked[10028];
  assign N5591 = N5590 | data_masked[10156];
  assign N5590 = N5589 | data_masked[10284];
  assign N5589 = N5588 | data_masked[10412];
  assign N5588 = N5587 | data_masked[10540];
  assign N5587 = N5586 | data_masked[10668];
  assign N5586 = N5585 | data_masked[10796];
  assign N5585 = N5584 | data_masked[10924];
  assign N5584 = N5583 | data_masked[11052];
  assign N5583 = N5582 | data_masked[11180];
  assign N5582 = N5581 | data_masked[11308];
  assign N5581 = N5580 | data_masked[11436];
  assign N5580 = N5579 | data_masked[11564];
  assign N5579 = N5578 | data_masked[11692];
  assign N5578 = N5577 | data_masked[11820];
  assign N5577 = N5576 | data_masked[11948];
  assign N5576 = N5575 | data_masked[12076];
  assign N5575 = N5574 | data_masked[12204];
  assign N5574 = N5573 | data_masked[12332];
  assign N5573 = N5572 | data_masked[12460];
  assign N5572 = N5571 | data_masked[12588];
  assign N5571 = N5570 | data_masked[12716];
  assign N5570 = N5569 | data_masked[12844];
  assign N5569 = N5568 | data_masked[12972];
  assign N5568 = N5567 | data_masked[13100];
  assign N5567 = N5566 | data_masked[13228];
  assign N5566 = N5565 | data_masked[13356];
  assign N5565 = N5564 | data_masked[13484];
  assign N5564 = N5563 | data_masked[13612];
  assign N5563 = N5562 | data_masked[13740];
  assign N5562 = N5561 | data_masked[13868];
  assign N5561 = N5560 | data_masked[13996];
  assign N5560 = N5559 | data_masked[14124];
  assign N5559 = N5558 | data_masked[14252];
  assign N5558 = N5557 | data_masked[14380];
  assign N5557 = N5556 | data_masked[14508];
  assign N5556 = N5555 | data_masked[14636];
  assign N5555 = N5554 | data_masked[14764];
  assign N5554 = N5553 | data_masked[14892];
  assign N5553 = N5552 | data_masked[15020];
  assign N5552 = N5551 | data_masked[15148];
  assign N5551 = N5550 | data_masked[15276];
  assign N5550 = N5549 | data_masked[15404];
  assign N5549 = N5548 | data_masked[15532];
  assign N5548 = N5547 | data_masked[15660];
  assign N5547 = N5546 | data_masked[15788];
  assign N5546 = N5545 | data_masked[15916];
  assign N5545 = N5544 | data_masked[16044];
  assign N5544 = data_masked[16300] | data_masked[16172];
  assign data_o[45] = N5795 | data_masked[45];
  assign N5795 = N5794 | data_masked[173];
  assign N5794 = N5793 | data_masked[301];
  assign N5793 = N5792 | data_masked[429];
  assign N5792 = N5791 | data_masked[557];
  assign N5791 = N5790 | data_masked[685];
  assign N5790 = N5789 | data_masked[813];
  assign N5789 = N5788 | data_masked[941];
  assign N5788 = N5787 | data_masked[1069];
  assign N5787 = N5786 | data_masked[1197];
  assign N5786 = N5785 | data_masked[1325];
  assign N5785 = N5784 | data_masked[1453];
  assign N5784 = N5783 | data_masked[1581];
  assign N5783 = N5782 | data_masked[1709];
  assign N5782 = N5781 | data_masked[1837];
  assign N5781 = N5780 | data_masked[1965];
  assign N5780 = N5779 | data_masked[2093];
  assign N5779 = N5778 | data_masked[2221];
  assign N5778 = N5777 | data_masked[2349];
  assign N5777 = N5776 | data_masked[2477];
  assign N5776 = N5775 | data_masked[2605];
  assign N5775 = N5774 | data_masked[2733];
  assign N5774 = N5773 | data_masked[2861];
  assign N5773 = N5772 | data_masked[2989];
  assign N5772 = N5771 | data_masked[3117];
  assign N5771 = N5770 | data_masked[3245];
  assign N5770 = N5769 | data_masked[3373];
  assign N5769 = N5768 | data_masked[3501];
  assign N5768 = N5767 | data_masked[3629];
  assign N5767 = N5766 | data_masked[3757];
  assign N5766 = N5765 | data_masked[3885];
  assign N5765 = N5764 | data_masked[4013];
  assign N5764 = N5763 | data_masked[4141];
  assign N5763 = N5762 | data_masked[4269];
  assign N5762 = N5761 | data_masked[4397];
  assign N5761 = N5760 | data_masked[4525];
  assign N5760 = N5759 | data_masked[4653];
  assign N5759 = N5758 | data_masked[4781];
  assign N5758 = N5757 | data_masked[4909];
  assign N5757 = N5756 | data_masked[5037];
  assign N5756 = N5755 | data_masked[5165];
  assign N5755 = N5754 | data_masked[5293];
  assign N5754 = N5753 | data_masked[5421];
  assign N5753 = N5752 | data_masked[5549];
  assign N5752 = N5751 | data_masked[5677];
  assign N5751 = N5750 | data_masked[5805];
  assign N5750 = N5749 | data_masked[5933];
  assign N5749 = N5748 | data_masked[6061];
  assign N5748 = N5747 | data_masked[6189];
  assign N5747 = N5746 | data_masked[6317];
  assign N5746 = N5745 | data_masked[6445];
  assign N5745 = N5744 | data_masked[6573];
  assign N5744 = N5743 | data_masked[6701];
  assign N5743 = N5742 | data_masked[6829];
  assign N5742 = N5741 | data_masked[6957];
  assign N5741 = N5740 | data_masked[7085];
  assign N5740 = N5739 | data_masked[7213];
  assign N5739 = N5738 | data_masked[7341];
  assign N5738 = N5737 | data_masked[7469];
  assign N5737 = N5736 | data_masked[7597];
  assign N5736 = N5735 | data_masked[7725];
  assign N5735 = N5734 | data_masked[7853];
  assign N5734 = N5733 | data_masked[7981];
  assign N5733 = N5732 | data_masked[8109];
  assign N5732 = N5731 | data_masked[8237];
  assign N5731 = N5730 | data_masked[8365];
  assign N5730 = N5729 | data_masked[8493];
  assign N5729 = N5728 | data_masked[8621];
  assign N5728 = N5727 | data_masked[8749];
  assign N5727 = N5726 | data_masked[8877];
  assign N5726 = N5725 | data_masked[9005];
  assign N5725 = N5724 | data_masked[9133];
  assign N5724 = N5723 | data_masked[9261];
  assign N5723 = N5722 | data_masked[9389];
  assign N5722 = N5721 | data_masked[9517];
  assign N5721 = N5720 | data_masked[9645];
  assign N5720 = N5719 | data_masked[9773];
  assign N5719 = N5718 | data_masked[9901];
  assign N5718 = N5717 | data_masked[10029];
  assign N5717 = N5716 | data_masked[10157];
  assign N5716 = N5715 | data_masked[10285];
  assign N5715 = N5714 | data_masked[10413];
  assign N5714 = N5713 | data_masked[10541];
  assign N5713 = N5712 | data_masked[10669];
  assign N5712 = N5711 | data_masked[10797];
  assign N5711 = N5710 | data_masked[10925];
  assign N5710 = N5709 | data_masked[11053];
  assign N5709 = N5708 | data_masked[11181];
  assign N5708 = N5707 | data_masked[11309];
  assign N5707 = N5706 | data_masked[11437];
  assign N5706 = N5705 | data_masked[11565];
  assign N5705 = N5704 | data_masked[11693];
  assign N5704 = N5703 | data_masked[11821];
  assign N5703 = N5702 | data_masked[11949];
  assign N5702 = N5701 | data_masked[12077];
  assign N5701 = N5700 | data_masked[12205];
  assign N5700 = N5699 | data_masked[12333];
  assign N5699 = N5698 | data_masked[12461];
  assign N5698 = N5697 | data_masked[12589];
  assign N5697 = N5696 | data_masked[12717];
  assign N5696 = N5695 | data_masked[12845];
  assign N5695 = N5694 | data_masked[12973];
  assign N5694 = N5693 | data_masked[13101];
  assign N5693 = N5692 | data_masked[13229];
  assign N5692 = N5691 | data_masked[13357];
  assign N5691 = N5690 | data_masked[13485];
  assign N5690 = N5689 | data_masked[13613];
  assign N5689 = N5688 | data_masked[13741];
  assign N5688 = N5687 | data_masked[13869];
  assign N5687 = N5686 | data_masked[13997];
  assign N5686 = N5685 | data_masked[14125];
  assign N5685 = N5684 | data_masked[14253];
  assign N5684 = N5683 | data_masked[14381];
  assign N5683 = N5682 | data_masked[14509];
  assign N5682 = N5681 | data_masked[14637];
  assign N5681 = N5680 | data_masked[14765];
  assign N5680 = N5679 | data_masked[14893];
  assign N5679 = N5678 | data_masked[15021];
  assign N5678 = N5677 | data_masked[15149];
  assign N5677 = N5676 | data_masked[15277];
  assign N5676 = N5675 | data_masked[15405];
  assign N5675 = N5674 | data_masked[15533];
  assign N5674 = N5673 | data_masked[15661];
  assign N5673 = N5672 | data_masked[15789];
  assign N5672 = N5671 | data_masked[15917];
  assign N5671 = N5670 | data_masked[16045];
  assign N5670 = data_masked[16301] | data_masked[16173];
  assign data_o[46] = N5921 | data_masked[46];
  assign N5921 = N5920 | data_masked[174];
  assign N5920 = N5919 | data_masked[302];
  assign N5919 = N5918 | data_masked[430];
  assign N5918 = N5917 | data_masked[558];
  assign N5917 = N5916 | data_masked[686];
  assign N5916 = N5915 | data_masked[814];
  assign N5915 = N5914 | data_masked[942];
  assign N5914 = N5913 | data_masked[1070];
  assign N5913 = N5912 | data_masked[1198];
  assign N5912 = N5911 | data_masked[1326];
  assign N5911 = N5910 | data_masked[1454];
  assign N5910 = N5909 | data_masked[1582];
  assign N5909 = N5908 | data_masked[1710];
  assign N5908 = N5907 | data_masked[1838];
  assign N5907 = N5906 | data_masked[1966];
  assign N5906 = N5905 | data_masked[2094];
  assign N5905 = N5904 | data_masked[2222];
  assign N5904 = N5903 | data_masked[2350];
  assign N5903 = N5902 | data_masked[2478];
  assign N5902 = N5901 | data_masked[2606];
  assign N5901 = N5900 | data_masked[2734];
  assign N5900 = N5899 | data_masked[2862];
  assign N5899 = N5898 | data_masked[2990];
  assign N5898 = N5897 | data_masked[3118];
  assign N5897 = N5896 | data_masked[3246];
  assign N5896 = N5895 | data_masked[3374];
  assign N5895 = N5894 | data_masked[3502];
  assign N5894 = N5893 | data_masked[3630];
  assign N5893 = N5892 | data_masked[3758];
  assign N5892 = N5891 | data_masked[3886];
  assign N5891 = N5890 | data_masked[4014];
  assign N5890 = N5889 | data_masked[4142];
  assign N5889 = N5888 | data_masked[4270];
  assign N5888 = N5887 | data_masked[4398];
  assign N5887 = N5886 | data_masked[4526];
  assign N5886 = N5885 | data_masked[4654];
  assign N5885 = N5884 | data_masked[4782];
  assign N5884 = N5883 | data_masked[4910];
  assign N5883 = N5882 | data_masked[5038];
  assign N5882 = N5881 | data_masked[5166];
  assign N5881 = N5880 | data_masked[5294];
  assign N5880 = N5879 | data_masked[5422];
  assign N5879 = N5878 | data_masked[5550];
  assign N5878 = N5877 | data_masked[5678];
  assign N5877 = N5876 | data_masked[5806];
  assign N5876 = N5875 | data_masked[5934];
  assign N5875 = N5874 | data_masked[6062];
  assign N5874 = N5873 | data_masked[6190];
  assign N5873 = N5872 | data_masked[6318];
  assign N5872 = N5871 | data_masked[6446];
  assign N5871 = N5870 | data_masked[6574];
  assign N5870 = N5869 | data_masked[6702];
  assign N5869 = N5868 | data_masked[6830];
  assign N5868 = N5867 | data_masked[6958];
  assign N5867 = N5866 | data_masked[7086];
  assign N5866 = N5865 | data_masked[7214];
  assign N5865 = N5864 | data_masked[7342];
  assign N5864 = N5863 | data_masked[7470];
  assign N5863 = N5862 | data_masked[7598];
  assign N5862 = N5861 | data_masked[7726];
  assign N5861 = N5860 | data_masked[7854];
  assign N5860 = N5859 | data_masked[7982];
  assign N5859 = N5858 | data_masked[8110];
  assign N5858 = N5857 | data_masked[8238];
  assign N5857 = N5856 | data_masked[8366];
  assign N5856 = N5855 | data_masked[8494];
  assign N5855 = N5854 | data_masked[8622];
  assign N5854 = N5853 | data_masked[8750];
  assign N5853 = N5852 | data_masked[8878];
  assign N5852 = N5851 | data_masked[9006];
  assign N5851 = N5850 | data_masked[9134];
  assign N5850 = N5849 | data_masked[9262];
  assign N5849 = N5848 | data_masked[9390];
  assign N5848 = N5847 | data_masked[9518];
  assign N5847 = N5846 | data_masked[9646];
  assign N5846 = N5845 | data_masked[9774];
  assign N5845 = N5844 | data_masked[9902];
  assign N5844 = N5843 | data_masked[10030];
  assign N5843 = N5842 | data_masked[10158];
  assign N5842 = N5841 | data_masked[10286];
  assign N5841 = N5840 | data_masked[10414];
  assign N5840 = N5839 | data_masked[10542];
  assign N5839 = N5838 | data_masked[10670];
  assign N5838 = N5837 | data_masked[10798];
  assign N5837 = N5836 | data_masked[10926];
  assign N5836 = N5835 | data_masked[11054];
  assign N5835 = N5834 | data_masked[11182];
  assign N5834 = N5833 | data_masked[11310];
  assign N5833 = N5832 | data_masked[11438];
  assign N5832 = N5831 | data_masked[11566];
  assign N5831 = N5830 | data_masked[11694];
  assign N5830 = N5829 | data_masked[11822];
  assign N5829 = N5828 | data_masked[11950];
  assign N5828 = N5827 | data_masked[12078];
  assign N5827 = N5826 | data_masked[12206];
  assign N5826 = N5825 | data_masked[12334];
  assign N5825 = N5824 | data_masked[12462];
  assign N5824 = N5823 | data_masked[12590];
  assign N5823 = N5822 | data_masked[12718];
  assign N5822 = N5821 | data_masked[12846];
  assign N5821 = N5820 | data_masked[12974];
  assign N5820 = N5819 | data_masked[13102];
  assign N5819 = N5818 | data_masked[13230];
  assign N5818 = N5817 | data_masked[13358];
  assign N5817 = N5816 | data_masked[13486];
  assign N5816 = N5815 | data_masked[13614];
  assign N5815 = N5814 | data_masked[13742];
  assign N5814 = N5813 | data_masked[13870];
  assign N5813 = N5812 | data_masked[13998];
  assign N5812 = N5811 | data_masked[14126];
  assign N5811 = N5810 | data_masked[14254];
  assign N5810 = N5809 | data_masked[14382];
  assign N5809 = N5808 | data_masked[14510];
  assign N5808 = N5807 | data_masked[14638];
  assign N5807 = N5806 | data_masked[14766];
  assign N5806 = N5805 | data_masked[14894];
  assign N5805 = N5804 | data_masked[15022];
  assign N5804 = N5803 | data_masked[15150];
  assign N5803 = N5802 | data_masked[15278];
  assign N5802 = N5801 | data_masked[15406];
  assign N5801 = N5800 | data_masked[15534];
  assign N5800 = N5799 | data_masked[15662];
  assign N5799 = N5798 | data_masked[15790];
  assign N5798 = N5797 | data_masked[15918];
  assign N5797 = N5796 | data_masked[16046];
  assign N5796 = data_masked[16302] | data_masked[16174];
  assign data_o[47] = N6047 | data_masked[47];
  assign N6047 = N6046 | data_masked[175];
  assign N6046 = N6045 | data_masked[303];
  assign N6045 = N6044 | data_masked[431];
  assign N6044 = N6043 | data_masked[559];
  assign N6043 = N6042 | data_masked[687];
  assign N6042 = N6041 | data_masked[815];
  assign N6041 = N6040 | data_masked[943];
  assign N6040 = N6039 | data_masked[1071];
  assign N6039 = N6038 | data_masked[1199];
  assign N6038 = N6037 | data_masked[1327];
  assign N6037 = N6036 | data_masked[1455];
  assign N6036 = N6035 | data_masked[1583];
  assign N6035 = N6034 | data_masked[1711];
  assign N6034 = N6033 | data_masked[1839];
  assign N6033 = N6032 | data_masked[1967];
  assign N6032 = N6031 | data_masked[2095];
  assign N6031 = N6030 | data_masked[2223];
  assign N6030 = N6029 | data_masked[2351];
  assign N6029 = N6028 | data_masked[2479];
  assign N6028 = N6027 | data_masked[2607];
  assign N6027 = N6026 | data_masked[2735];
  assign N6026 = N6025 | data_masked[2863];
  assign N6025 = N6024 | data_masked[2991];
  assign N6024 = N6023 | data_masked[3119];
  assign N6023 = N6022 | data_masked[3247];
  assign N6022 = N6021 | data_masked[3375];
  assign N6021 = N6020 | data_masked[3503];
  assign N6020 = N6019 | data_masked[3631];
  assign N6019 = N6018 | data_masked[3759];
  assign N6018 = N6017 | data_masked[3887];
  assign N6017 = N6016 | data_masked[4015];
  assign N6016 = N6015 | data_masked[4143];
  assign N6015 = N6014 | data_masked[4271];
  assign N6014 = N6013 | data_masked[4399];
  assign N6013 = N6012 | data_masked[4527];
  assign N6012 = N6011 | data_masked[4655];
  assign N6011 = N6010 | data_masked[4783];
  assign N6010 = N6009 | data_masked[4911];
  assign N6009 = N6008 | data_masked[5039];
  assign N6008 = N6007 | data_masked[5167];
  assign N6007 = N6006 | data_masked[5295];
  assign N6006 = N6005 | data_masked[5423];
  assign N6005 = N6004 | data_masked[5551];
  assign N6004 = N6003 | data_masked[5679];
  assign N6003 = N6002 | data_masked[5807];
  assign N6002 = N6001 | data_masked[5935];
  assign N6001 = N6000 | data_masked[6063];
  assign N6000 = N5999 | data_masked[6191];
  assign N5999 = N5998 | data_masked[6319];
  assign N5998 = N5997 | data_masked[6447];
  assign N5997 = N5996 | data_masked[6575];
  assign N5996 = N5995 | data_masked[6703];
  assign N5995 = N5994 | data_masked[6831];
  assign N5994 = N5993 | data_masked[6959];
  assign N5993 = N5992 | data_masked[7087];
  assign N5992 = N5991 | data_masked[7215];
  assign N5991 = N5990 | data_masked[7343];
  assign N5990 = N5989 | data_masked[7471];
  assign N5989 = N5988 | data_masked[7599];
  assign N5988 = N5987 | data_masked[7727];
  assign N5987 = N5986 | data_masked[7855];
  assign N5986 = N5985 | data_masked[7983];
  assign N5985 = N5984 | data_masked[8111];
  assign N5984 = N5983 | data_masked[8239];
  assign N5983 = N5982 | data_masked[8367];
  assign N5982 = N5981 | data_masked[8495];
  assign N5981 = N5980 | data_masked[8623];
  assign N5980 = N5979 | data_masked[8751];
  assign N5979 = N5978 | data_masked[8879];
  assign N5978 = N5977 | data_masked[9007];
  assign N5977 = N5976 | data_masked[9135];
  assign N5976 = N5975 | data_masked[9263];
  assign N5975 = N5974 | data_masked[9391];
  assign N5974 = N5973 | data_masked[9519];
  assign N5973 = N5972 | data_masked[9647];
  assign N5972 = N5971 | data_masked[9775];
  assign N5971 = N5970 | data_masked[9903];
  assign N5970 = N5969 | data_masked[10031];
  assign N5969 = N5968 | data_masked[10159];
  assign N5968 = N5967 | data_masked[10287];
  assign N5967 = N5966 | data_masked[10415];
  assign N5966 = N5965 | data_masked[10543];
  assign N5965 = N5964 | data_masked[10671];
  assign N5964 = N5963 | data_masked[10799];
  assign N5963 = N5962 | data_masked[10927];
  assign N5962 = N5961 | data_masked[11055];
  assign N5961 = N5960 | data_masked[11183];
  assign N5960 = N5959 | data_masked[11311];
  assign N5959 = N5958 | data_masked[11439];
  assign N5958 = N5957 | data_masked[11567];
  assign N5957 = N5956 | data_masked[11695];
  assign N5956 = N5955 | data_masked[11823];
  assign N5955 = N5954 | data_masked[11951];
  assign N5954 = N5953 | data_masked[12079];
  assign N5953 = N5952 | data_masked[12207];
  assign N5952 = N5951 | data_masked[12335];
  assign N5951 = N5950 | data_masked[12463];
  assign N5950 = N5949 | data_masked[12591];
  assign N5949 = N5948 | data_masked[12719];
  assign N5948 = N5947 | data_masked[12847];
  assign N5947 = N5946 | data_masked[12975];
  assign N5946 = N5945 | data_masked[13103];
  assign N5945 = N5944 | data_masked[13231];
  assign N5944 = N5943 | data_masked[13359];
  assign N5943 = N5942 | data_masked[13487];
  assign N5942 = N5941 | data_masked[13615];
  assign N5941 = N5940 | data_masked[13743];
  assign N5940 = N5939 | data_masked[13871];
  assign N5939 = N5938 | data_masked[13999];
  assign N5938 = N5937 | data_masked[14127];
  assign N5937 = N5936 | data_masked[14255];
  assign N5936 = N5935 | data_masked[14383];
  assign N5935 = N5934 | data_masked[14511];
  assign N5934 = N5933 | data_masked[14639];
  assign N5933 = N5932 | data_masked[14767];
  assign N5932 = N5931 | data_masked[14895];
  assign N5931 = N5930 | data_masked[15023];
  assign N5930 = N5929 | data_masked[15151];
  assign N5929 = N5928 | data_masked[15279];
  assign N5928 = N5927 | data_masked[15407];
  assign N5927 = N5926 | data_masked[15535];
  assign N5926 = N5925 | data_masked[15663];
  assign N5925 = N5924 | data_masked[15791];
  assign N5924 = N5923 | data_masked[15919];
  assign N5923 = N5922 | data_masked[16047];
  assign N5922 = data_masked[16303] | data_masked[16175];
  assign data_o[48] = N6173 | data_masked[48];
  assign N6173 = N6172 | data_masked[176];
  assign N6172 = N6171 | data_masked[304];
  assign N6171 = N6170 | data_masked[432];
  assign N6170 = N6169 | data_masked[560];
  assign N6169 = N6168 | data_masked[688];
  assign N6168 = N6167 | data_masked[816];
  assign N6167 = N6166 | data_masked[944];
  assign N6166 = N6165 | data_masked[1072];
  assign N6165 = N6164 | data_masked[1200];
  assign N6164 = N6163 | data_masked[1328];
  assign N6163 = N6162 | data_masked[1456];
  assign N6162 = N6161 | data_masked[1584];
  assign N6161 = N6160 | data_masked[1712];
  assign N6160 = N6159 | data_masked[1840];
  assign N6159 = N6158 | data_masked[1968];
  assign N6158 = N6157 | data_masked[2096];
  assign N6157 = N6156 | data_masked[2224];
  assign N6156 = N6155 | data_masked[2352];
  assign N6155 = N6154 | data_masked[2480];
  assign N6154 = N6153 | data_masked[2608];
  assign N6153 = N6152 | data_masked[2736];
  assign N6152 = N6151 | data_masked[2864];
  assign N6151 = N6150 | data_masked[2992];
  assign N6150 = N6149 | data_masked[3120];
  assign N6149 = N6148 | data_masked[3248];
  assign N6148 = N6147 | data_masked[3376];
  assign N6147 = N6146 | data_masked[3504];
  assign N6146 = N6145 | data_masked[3632];
  assign N6145 = N6144 | data_masked[3760];
  assign N6144 = N6143 | data_masked[3888];
  assign N6143 = N6142 | data_masked[4016];
  assign N6142 = N6141 | data_masked[4144];
  assign N6141 = N6140 | data_masked[4272];
  assign N6140 = N6139 | data_masked[4400];
  assign N6139 = N6138 | data_masked[4528];
  assign N6138 = N6137 | data_masked[4656];
  assign N6137 = N6136 | data_masked[4784];
  assign N6136 = N6135 | data_masked[4912];
  assign N6135 = N6134 | data_masked[5040];
  assign N6134 = N6133 | data_masked[5168];
  assign N6133 = N6132 | data_masked[5296];
  assign N6132 = N6131 | data_masked[5424];
  assign N6131 = N6130 | data_masked[5552];
  assign N6130 = N6129 | data_masked[5680];
  assign N6129 = N6128 | data_masked[5808];
  assign N6128 = N6127 | data_masked[5936];
  assign N6127 = N6126 | data_masked[6064];
  assign N6126 = N6125 | data_masked[6192];
  assign N6125 = N6124 | data_masked[6320];
  assign N6124 = N6123 | data_masked[6448];
  assign N6123 = N6122 | data_masked[6576];
  assign N6122 = N6121 | data_masked[6704];
  assign N6121 = N6120 | data_masked[6832];
  assign N6120 = N6119 | data_masked[6960];
  assign N6119 = N6118 | data_masked[7088];
  assign N6118 = N6117 | data_masked[7216];
  assign N6117 = N6116 | data_masked[7344];
  assign N6116 = N6115 | data_masked[7472];
  assign N6115 = N6114 | data_masked[7600];
  assign N6114 = N6113 | data_masked[7728];
  assign N6113 = N6112 | data_masked[7856];
  assign N6112 = N6111 | data_masked[7984];
  assign N6111 = N6110 | data_masked[8112];
  assign N6110 = N6109 | data_masked[8240];
  assign N6109 = N6108 | data_masked[8368];
  assign N6108 = N6107 | data_masked[8496];
  assign N6107 = N6106 | data_masked[8624];
  assign N6106 = N6105 | data_masked[8752];
  assign N6105 = N6104 | data_masked[8880];
  assign N6104 = N6103 | data_masked[9008];
  assign N6103 = N6102 | data_masked[9136];
  assign N6102 = N6101 | data_masked[9264];
  assign N6101 = N6100 | data_masked[9392];
  assign N6100 = N6099 | data_masked[9520];
  assign N6099 = N6098 | data_masked[9648];
  assign N6098 = N6097 | data_masked[9776];
  assign N6097 = N6096 | data_masked[9904];
  assign N6096 = N6095 | data_masked[10032];
  assign N6095 = N6094 | data_masked[10160];
  assign N6094 = N6093 | data_masked[10288];
  assign N6093 = N6092 | data_masked[10416];
  assign N6092 = N6091 | data_masked[10544];
  assign N6091 = N6090 | data_masked[10672];
  assign N6090 = N6089 | data_masked[10800];
  assign N6089 = N6088 | data_masked[10928];
  assign N6088 = N6087 | data_masked[11056];
  assign N6087 = N6086 | data_masked[11184];
  assign N6086 = N6085 | data_masked[11312];
  assign N6085 = N6084 | data_masked[11440];
  assign N6084 = N6083 | data_masked[11568];
  assign N6083 = N6082 | data_masked[11696];
  assign N6082 = N6081 | data_masked[11824];
  assign N6081 = N6080 | data_masked[11952];
  assign N6080 = N6079 | data_masked[12080];
  assign N6079 = N6078 | data_masked[12208];
  assign N6078 = N6077 | data_masked[12336];
  assign N6077 = N6076 | data_masked[12464];
  assign N6076 = N6075 | data_masked[12592];
  assign N6075 = N6074 | data_masked[12720];
  assign N6074 = N6073 | data_masked[12848];
  assign N6073 = N6072 | data_masked[12976];
  assign N6072 = N6071 | data_masked[13104];
  assign N6071 = N6070 | data_masked[13232];
  assign N6070 = N6069 | data_masked[13360];
  assign N6069 = N6068 | data_masked[13488];
  assign N6068 = N6067 | data_masked[13616];
  assign N6067 = N6066 | data_masked[13744];
  assign N6066 = N6065 | data_masked[13872];
  assign N6065 = N6064 | data_masked[14000];
  assign N6064 = N6063 | data_masked[14128];
  assign N6063 = N6062 | data_masked[14256];
  assign N6062 = N6061 | data_masked[14384];
  assign N6061 = N6060 | data_masked[14512];
  assign N6060 = N6059 | data_masked[14640];
  assign N6059 = N6058 | data_masked[14768];
  assign N6058 = N6057 | data_masked[14896];
  assign N6057 = N6056 | data_masked[15024];
  assign N6056 = N6055 | data_masked[15152];
  assign N6055 = N6054 | data_masked[15280];
  assign N6054 = N6053 | data_masked[15408];
  assign N6053 = N6052 | data_masked[15536];
  assign N6052 = N6051 | data_masked[15664];
  assign N6051 = N6050 | data_masked[15792];
  assign N6050 = N6049 | data_masked[15920];
  assign N6049 = N6048 | data_masked[16048];
  assign N6048 = data_masked[16304] | data_masked[16176];
  assign data_o[49] = N6299 | data_masked[49];
  assign N6299 = N6298 | data_masked[177];
  assign N6298 = N6297 | data_masked[305];
  assign N6297 = N6296 | data_masked[433];
  assign N6296 = N6295 | data_masked[561];
  assign N6295 = N6294 | data_masked[689];
  assign N6294 = N6293 | data_masked[817];
  assign N6293 = N6292 | data_masked[945];
  assign N6292 = N6291 | data_masked[1073];
  assign N6291 = N6290 | data_masked[1201];
  assign N6290 = N6289 | data_masked[1329];
  assign N6289 = N6288 | data_masked[1457];
  assign N6288 = N6287 | data_masked[1585];
  assign N6287 = N6286 | data_masked[1713];
  assign N6286 = N6285 | data_masked[1841];
  assign N6285 = N6284 | data_masked[1969];
  assign N6284 = N6283 | data_masked[2097];
  assign N6283 = N6282 | data_masked[2225];
  assign N6282 = N6281 | data_masked[2353];
  assign N6281 = N6280 | data_masked[2481];
  assign N6280 = N6279 | data_masked[2609];
  assign N6279 = N6278 | data_masked[2737];
  assign N6278 = N6277 | data_masked[2865];
  assign N6277 = N6276 | data_masked[2993];
  assign N6276 = N6275 | data_masked[3121];
  assign N6275 = N6274 | data_masked[3249];
  assign N6274 = N6273 | data_masked[3377];
  assign N6273 = N6272 | data_masked[3505];
  assign N6272 = N6271 | data_masked[3633];
  assign N6271 = N6270 | data_masked[3761];
  assign N6270 = N6269 | data_masked[3889];
  assign N6269 = N6268 | data_masked[4017];
  assign N6268 = N6267 | data_masked[4145];
  assign N6267 = N6266 | data_masked[4273];
  assign N6266 = N6265 | data_masked[4401];
  assign N6265 = N6264 | data_masked[4529];
  assign N6264 = N6263 | data_masked[4657];
  assign N6263 = N6262 | data_masked[4785];
  assign N6262 = N6261 | data_masked[4913];
  assign N6261 = N6260 | data_masked[5041];
  assign N6260 = N6259 | data_masked[5169];
  assign N6259 = N6258 | data_masked[5297];
  assign N6258 = N6257 | data_masked[5425];
  assign N6257 = N6256 | data_masked[5553];
  assign N6256 = N6255 | data_masked[5681];
  assign N6255 = N6254 | data_masked[5809];
  assign N6254 = N6253 | data_masked[5937];
  assign N6253 = N6252 | data_masked[6065];
  assign N6252 = N6251 | data_masked[6193];
  assign N6251 = N6250 | data_masked[6321];
  assign N6250 = N6249 | data_masked[6449];
  assign N6249 = N6248 | data_masked[6577];
  assign N6248 = N6247 | data_masked[6705];
  assign N6247 = N6246 | data_masked[6833];
  assign N6246 = N6245 | data_masked[6961];
  assign N6245 = N6244 | data_masked[7089];
  assign N6244 = N6243 | data_masked[7217];
  assign N6243 = N6242 | data_masked[7345];
  assign N6242 = N6241 | data_masked[7473];
  assign N6241 = N6240 | data_masked[7601];
  assign N6240 = N6239 | data_masked[7729];
  assign N6239 = N6238 | data_masked[7857];
  assign N6238 = N6237 | data_masked[7985];
  assign N6237 = N6236 | data_masked[8113];
  assign N6236 = N6235 | data_masked[8241];
  assign N6235 = N6234 | data_masked[8369];
  assign N6234 = N6233 | data_masked[8497];
  assign N6233 = N6232 | data_masked[8625];
  assign N6232 = N6231 | data_masked[8753];
  assign N6231 = N6230 | data_masked[8881];
  assign N6230 = N6229 | data_masked[9009];
  assign N6229 = N6228 | data_masked[9137];
  assign N6228 = N6227 | data_masked[9265];
  assign N6227 = N6226 | data_masked[9393];
  assign N6226 = N6225 | data_masked[9521];
  assign N6225 = N6224 | data_masked[9649];
  assign N6224 = N6223 | data_masked[9777];
  assign N6223 = N6222 | data_masked[9905];
  assign N6222 = N6221 | data_masked[10033];
  assign N6221 = N6220 | data_masked[10161];
  assign N6220 = N6219 | data_masked[10289];
  assign N6219 = N6218 | data_masked[10417];
  assign N6218 = N6217 | data_masked[10545];
  assign N6217 = N6216 | data_masked[10673];
  assign N6216 = N6215 | data_masked[10801];
  assign N6215 = N6214 | data_masked[10929];
  assign N6214 = N6213 | data_masked[11057];
  assign N6213 = N6212 | data_masked[11185];
  assign N6212 = N6211 | data_masked[11313];
  assign N6211 = N6210 | data_masked[11441];
  assign N6210 = N6209 | data_masked[11569];
  assign N6209 = N6208 | data_masked[11697];
  assign N6208 = N6207 | data_masked[11825];
  assign N6207 = N6206 | data_masked[11953];
  assign N6206 = N6205 | data_masked[12081];
  assign N6205 = N6204 | data_masked[12209];
  assign N6204 = N6203 | data_masked[12337];
  assign N6203 = N6202 | data_masked[12465];
  assign N6202 = N6201 | data_masked[12593];
  assign N6201 = N6200 | data_masked[12721];
  assign N6200 = N6199 | data_masked[12849];
  assign N6199 = N6198 | data_masked[12977];
  assign N6198 = N6197 | data_masked[13105];
  assign N6197 = N6196 | data_masked[13233];
  assign N6196 = N6195 | data_masked[13361];
  assign N6195 = N6194 | data_masked[13489];
  assign N6194 = N6193 | data_masked[13617];
  assign N6193 = N6192 | data_masked[13745];
  assign N6192 = N6191 | data_masked[13873];
  assign N6191 = N6190 | data_masked[14001];
  assign N6190 = N6189 | data_masked[14129];
  assign N6189 = N6188 | data_masked[14257];
  assign N6188 = N6187 | data_masked[14385];
  assign N6187 = N6186 | data_masked[14513];
  assign N6186 = N6185 | data_masked[14641];
  assign N6185 = N6184 | data_masked[14769];
  assign N6184 = N6183 | data_masked[14897];
  assign N6183 = N6182 | data_masked[15025];
  assign N6182 = N6181 | data_masked[15153];
  assign N6181 = N6180 | data_masked[15281];
  assign N6180 = N6179 | data_masked[15409];
  assign N6179 = N6178 | data_masked[15537];
  assign N6178 = N6177 | data_masked[15665];
  assign N6177 = N6176 | data_masked[15793];
  assign N6176 = N6175 | data_masked[15921];
  assign N6175 = N6174 | data_masked[16049];
  assign N6174 = data_masked[16305] | data_masked[16177];
  assign data_o[50] = N6425 | data_masked[50];
  assign N6425 = N6424 | data_masked[178];
  assign N6424 = N6423 | data_masked[306];
  assign N6423 = N6422 | data_masked[434];
  assign N6422 = N6421 | data_masked[562];
  assign N6421 = N6420 | data_masked[690];
  assign N6420 = N6419 | data_masked[818];
  assign N6419 = N6418 | data_masked[946];
  assign N6418 = N6417 | data_masked[1074];
  assign N6417 = N6416 | data_masked[1202];
  assign N6416 = N6415 | data_masked[1330];
  assign N6415 = N6414 | data_masked[1458];
  assign N6414 = N6413 | data_masked[1586];
  assign N6413 = N6412 | data_masked[1714];
  assign N6412 = N6411 | data_masked[1842];
  assign N6411 = N6410 | data_masked[1970];
  assign N6410 = N6409 | data_masked[2098];
  assign N6409 = N6408 | data_masked[2226];
  assign N6408 = N6407 | data_masked[2354];
  assign N6407 = N6406 | data_masked[2482];
  assign N6406 = N6405 | data_masked[2610];
  assign N6405 = N6404 | data_masked[2738];
  assign N6404 = N6403 | data_masked[2866];
  assign N6403 = N6402 | data_masked[2994];
  assign N6402 = N6401 | data_masked[3122];
  assign N6401 = N6400 | data_masked[3250];
  assign N6400 = N6399 | data_masked[3378];
  assign N6399 = N6398 | data_masked[3506];
  assign N6398 = N6397 | data_masked[3634];
  assign N6397 = N6396 | data_masked[3762];
  assign N6396 = N6395 | data_masked[3890];
  assign N6395 = N6394 | data_masked[4018];
  assign N6394 = N6393 | data_masked[4146];
  assign N6393 = N6392 | data_masked[4274];
  assign N6392 = N6391 | data_masked[4402];
  assign N6391 = N6390 | data_masked[4530];
  assign N6390 = N6389 | data_masked[4658];
  assign N6389 = N6388 | data_masked[4786];
  assign N6388 = N6387 | data_masked[4914];
  assign N6387 = N6386 | data_masked[5042];
  assign N6386 = N6385 | data_masked[5170];
  assign N6385 = N6384 | data_masked[5298];
  assign N6384 = N6383 | data_masked[5426];
  assign N6383 = N6382 | data_masked[5554];
  assign N6382 = N6381 | data_masked[5682];
  assign N6381 = N6380 | data_masked[5810];
  assign N6380 = N6379 | data_masked[5938];
  assign N6379 = N6378 | data_masked[6066];
  assign N6378 = N6377 | data_masked[6194];
  assign N6377 = N6376 | data_masked[6322];
  assign N6376 = N6375 | data_masked[6450];
  assign N6375 = N6374 | data_masked[6578];
  assign N6374 = N6373 | data_masked[6706];
  assign N6373 = N6372 | data_masked[6834];
  assign N6372 = N6371 | data_masked[6962];
  assign N6371 = N6370 | data_masked[7090];
  assign N6370 = N6369 | data_masked[7218];
  assign N6369 = N6368 | data_masked[7346];
  assign N6368 = N6367 | data_masked[7474];
  assign N6367 = N6366 | data_masked[7602];
  assign N6366 = N6365 | data_masked[7730];
  assign N6365 = N6364 | data_masked[7858];
  assign N6364 = N6363 | data_masked[7986];
  assign N6363 = N6362 | data_masked[8114];
  assign N6362 = N6361 | data_masked[8242];
  assign N6361 = N6360 | data_masked[8370];
  assign N6360 = N6359 | data_masked[8498];
  assign N6359 = N6358 | data_masked[8626];
  assign N6358 = N6357 | data_masked[8754];
  assign N6357 = N6356 | data_masked[8882];
  assign N6356 = N6355 | data_masked[9010];
  assign N6355 = N6354 | data_masked[9138];
  assign N6354 = N6353 | data_masked[9266];
  assign N6353 = N6352 | data_masked[9394];
  assign N6352 = N6351 | data_masked[9522];
  assign N6351 = N6350 | data_masked[9650];
  assign N6350 = N6349 | data_masked[9778];
  assign N6349 = N6348 | data_masked[9906];
  assign N6348 = N6347 | data_masked[10034];
  assign N6347 = N6346 | data_masked[10162];
  assign N6346 = N6345 | data_masked[10290];
  assign N6345 = N6344 | data_masked[10418];
  assign N6344 = N6343 | data_masked[10546];
  assign N6343 = N6342 | data_masked[10674];
  assign N6342 = N6341 | data_masked[10802];
  assign N6341 = N6340 | data_masked[10930];
  assign N6340 = N6339 | data_masked[11058];
  assign N6339 = N6338 | data_masked[11186];
  assign N6338 = N6337 | data_masked[11314];
  assign N6337 = N6336 | data_masked[11442];
  assign N6336 = N6335 | data_masked[11570];
  assign N6335 = N6334 | data_masked[11698];
  assign N6334 = N6333 | data_masked[11826];
  assign N6333 = N6332 | data_masked[11954];
  assign N6332 = N6331 | data_masked[12082];
  assign N6331 = N6330 | data_masked[12210];
  assign N6330 = N6329 | data_masked[12338];
  assign N6329 = N6328 | data_masked[12466];
  assign N6328 = N6327 | data_masked[12594];
  assign N6327 = N6326 | data_masked[12722];
  assign N6326 = N6325 | data_masked[12850];
  assign N6325 = N6324 | data_masked[12978];
  assign N6324 = N6323 | data_masked[13106];
  assign N6323 = N6322 | data_masked[13234];
  assign N6322 = N6321 | data_masked[13362];
  assign N6321 = N6320 | data_masked[13490];
  assign N6320 = N6319 | data_masked[13618];
  assign N6319 = N6318 | data_masked[13746];
  assign N6318 = N6317 | data_masked[13874];
  assign N6317 = N6316 | data_masked[14002];
  assign N6316 = N6315 | data_masked[14130];
  assign N6315 = N6314 | data_masked[14258];
  assign N6314 = N6313 | data_masked[14386];
  assign N6313 = N6312 | data_masked[14514];
  assign N6312 = N6311 | data_masked[14642];
  assign N6311 = N6310 | data_masked[14770];
  assign N6310 = N6309 | data_masked[14898];
  assign N6309 = N6308 | data_masked[15026];
  assign N6308 = N6307 | data_masked[15154];
  assign N6307 = N6306 | data_masked[15282];
  assign N6306 = N6305 | data_masked[15410];
  assign N6305 = N6304 | data_masked[15538];
  assign N6304 = N6303 | data_masked[15666];
  assign N6303 = N6302 | data_masked[15794];
  assign N6302 = N6301 | data_masked[15922];
  assign N6301 = N6300 | data_masked[16050];
  assign N6300 = data_masked[16306] | data_masked[16178];
  assign data_o[51] = N6551 | data_masked[51];
  assign N6551 = N6550 | data_masked[179];
  assign N6550 = N6549 | data_masked[307];
  assign N6549 = N6548 | data_masked[435];
  assign N6548 = N6547 | data_masked[563];
  assign N6547 = N6546 | data_masked[691];
  assign N6546 = N6545 | data_masked[819];
  assign N6545 = N6544 | data_masked[947];
  assign N6544 = N6543 | data_masked[1075];
  assign N6543 = N6542 | data_masked[1203];
  assign N6542 = N6541 | data_masked[1331];
  assign N6541 = N6540 | data_masked[1459];
  assign N6540 = N6539 | data_masked[1587];
  assign N6539 = N6538 | data_masked[1715];
  assign N6538 = N6537 | data_masked[1843];
  assign N6537 = N6536 | data_masked[1971];
  assign N6536 = N6535 | data_masked[2099];
  assign N6535 = N6534 | data_masked[2227];
  assign N6534 = N6533 | data_masked[2355];
  assign N6533 = N6532 | data_masked[2483];
  assign N6532 = N6531 | data_masked[2611];
  assign N6531 = N6530 | data_masked[2739];
  assign N6530 = N6529 | data_masked[2867];
  assign N6529 = N6528 | data_masked[2995];
  assign N6528 = N6527 | data_masked[3123];
  assign N6527 = N6526 | data_masked[3251];
  assign N6526 = N6525 | data_masked[3379];
  assign N6525 = N6524 | data_masked[3507];
  assign N6524 = N6523 | data_masked[3635];
  assign N6523 = N6522 | data_masked[3763];
  assign N6522 = N6521 | data_masked[3891];
  assign N6521 = N6520 | data_masked[4019];
  assign N6520 = N6519 | data_masked[4147];
  assign N6519 = N6518 | data_masked[4275];
  assign N6518 = N6517 | data_masked[4403];
  assign N6517 = N6516 | data_masked[4531];
  assign N6516 = N6515 | data_masked[4659];
  assign N6515 = N6514 | data_masked[4787];
  assign N6514 = N6513 | data_masked[4915];
  assign N6513 = N6512 | data_masked[5043];
  assign N6512 = N6511 | data_masked[5171];
  assign N6511 = N6510 | data_masked[5299];
  assign N6510 = N6509 | data_masked[5427];
  assign N6509 = N6508 | data_masked[5555];
  assign N6508 = N6507 | data_masked[5683];
  assign N6507 = N6506 | data_masked[5811];
  assign N6506 = N6505 | data_masked[5939];
  assign N6505 = N6504 | data_masked[6067];
  assign N6504 = N6503 | data_masked[6195];
  assign N6503 = N6502 | data_masked[6323];
  assign N6502 = N6501 | data_masked[6451];
  assign N6501 = N6500 | data_masked[6579];
  assign N6500 = N6499 | data_masked[6707];
  assign N6499 = N6498 | data_masked[6835];
  assign N6498 = N6497 | data_masked[6963];
  assign N6497 = N6496 | data_masked[7091];
  assign N6496 = N6495 | data_masked[7219];
  assign N6495 = N6494 | data_masked[7347];
  assign N6494 = N6493 | data_masked[7475];
  assign N6493 = N6492 | data_masked[7603];
  assign N6492 = N6491 | data_masked[7731];
  assign N6491 = N6490 | data_masked[7859];
  assign N6490 = N6489 | data_masked[7987];
  assign N6489 = N6488 | data_masked[8115];
  assign N6488 = N6487 | data_masked[8243];
  assign N6487 = N6486 | data_masked[8371];
  assign N6486 = N6485 | data_masked[8499];
  assign N6485 = N6484 | data_masked[8627];
  assign N6484 = N6483 | data_masked[8755];
  assign N6483 = N6482 | data_masked[8883];
  assign N6482 = N6481 | data_masked[9011];
  assign N6481 = N6480 | data_masked[9139];
  assign N6480 = N6479 | data_masked[9267];
  assign N6479 = N6478 | data_masked[9395];
  assign N6478 = N6477 | data_masked[9523];
  assign N6477 = N6476 | data_masked[9651];
  assign N6476 = N6475 | data_masked[9779];
  assign N6475 = N6474 | data_masked[9907];
  assign N6474 = N6473 | data_masked[10035];
  assign N6473 = N6472 | data_masked[10163];
  assign N6472 = N6471 | data_masked[10291];
  assign N6471 = N6470 | data_masked[10419];
  assign N6470 = N6469 | data_masked[10547];
  assign N6469 = N6468 | data_masked[10675];
  assign N6468 = N6467 | data_masked[10803];
  assign N6467 = N6466 | data_masked[10931];
  assign N6466 = N6465 | data_masked[11059];
  assign N6465 = N6464 | data_masked[11187];
  assign N6464 = N6463 | data_masked[11315];
  assign N6463 = N6462 | data_masked[11443];
  assign N6462 = N6461 | data_masked[11571];
  assign N6461 = N6460 | data_masked[11699];
  assign N6460 = N6459 | data_masked[11827];
  assign N6459 = N6458 | data_masked[11955];
  assign N6458 = N6457 | data_masked[12083];
  assign N6457 = N6456 | data_masked[12211];
  assign N6456 = N6455 | data_masked[12339];
  assign N6455 = N6454 | data_masked[12467];
  assign N6454 = N6453 | data_masked[12595];
  assign N6453 = N6452 | data_masked[12723];
  assign N6452 = N6451 | data_masked[12851];
  assign N6451 = N6450 | data_masked[12979];
  assign N6450 = N6449 | data_masked[13107];
  assign N6449 = N6448 | data_masked[13235];
  assign N6448 = N6447 | data_masked[13363];
  assign N6447 = N6446 | data_masked[13491];
  assign N6446 = N6445 | data_masked[13619];
  assign N6445 = N6444 | data_masked[13747];
  assign N6444 = N6443 | data_masked[13875];
  assign N6443 = N6442 | data_masked[14003];
  assign N6442 = N6441 | data_masked[14131];
  assign N6441 = N6440 | data_masked[14259];
  assign N6440 = N6439 | data_masked[14387];
  assign N6439 = N6438 | data_masked[14515];
  assign N6438 = N6437 | data_masked[14643];
  assign N6437 = N6436 | data_masked[14771];
  assign N6436 = N6435 | data_masked[14899];
  assign N6435 = N6434 | data_masked[15027];
  assign N6434 = N6433 | data_masked[15155];
  assign N6433 = N6432 | data_masked[15283];
  assign N6432 = N6431 | data_masked[15411];
  assign N6431 = N6430 | data_masked[15539];
  assign N6430 = N6429 | data_masked[15667];
  assign N6429 = N6428 | data_masked[15795];
  assign N6428 = N6427 | data_masked[15923];
  assign N6427 = N6426 | data_masked[16051];
  assign N6426 = data_masked[16307] | data_masked[16179];
  assign data_o[52] = N6677 | data_masked[52];
  assign N6677 = N6676 | data_masked[180];
  assign N6676 = N6675 | data_masked[308];
  assign N6675 = N6674 | data_masked[436];
  assign N6674 = N6673 | data_masked[564];
  assign N6673 = N6672 | data_masked[692];
  assign N6672 = N6671 | data_masked[820];
  assign N6671 = N6670 | data_masked[948];
  assign N6670 = N6669 | data_masked[1076];
  assign N6669 = N6668 | data_masked[1204];
  assign N6668 = N6667 | data_masked[1332];
  assign N6667 = N6666 | data_masked[1460];
  assign N6666 = N6665 | data_masked[1588];
  assign N6665 = N6664 | data_masked[1716];
  assign N6664 = N6663 | data_masked[1844];
  assign N6663 = N6662 | data_masked[1972];
  assign N6662 = N6661 | data_masked[2100];
  assign N6661 = N6660 | data_masked[2228];
  assign N6660 = N6659 | data_masked[2356];
  assign N6659 = N6658 | data_masked[2484];
  assign N6658 = N6657 | data_masked[2612];
  assign N6657 = N6656 | data_masked[2740];
  assign N6656 = N6655 | data_masked[2868];
  assign N6655 = N6654 | data_masked[2996];
  assign N6654 = N6653 | data_masked[3124];
  assign N6653 = N6652 | data_masked[3252];
  assign N6652 = N6651 | data_masked[3380];
  assign N6651 = N6650 | data_masked[3508];
  assign N6650 = N6649 | data_masked[3636];
  assign N6649 = N6648 | data_masked[3764];
  assign N6648 = N6647 | data_masked[3892];
  assign N6647 = N6646 | data_masked[4020];
  assign N6646 = N6645 | data_masked[4148];
  assign N6645 = N6644 | data_masked[4276];
  assign N6644 = N6643 | data_masked[4404];
  assign N6643 = N6642 | data_masked[4532];
  assign N6642 = N6641 | data_masked[4660];
  assign N6641 = N6640 | data_masked[4788];
  assign N6640 = N6639 | data_masked[4916];
  assign N6639 = N6638 | data_masked[5044];
  assign N6638 = N6637 | data_masked[5172];
  assign N6637 = N6636 | data_masked[5300];
  assign N6636 = N6635 | data_masked[5428];
  assign N6635 = N6634 | data_masked[5556];
  assign N6634 = N6633 | data_masked[5684];
  assign N6633 = N6632 | data_masked[5812];
  assign N6632 = N6631 | data_masked[5940];
  assign N6631 = N6630 | data_masked[6068];
  assign N6630 = N6629 | data_masked[6196];
  assign N6629 = N6628 | data_masked[6324];
  assign N6628 = N6627 | data_masked[6452];
  assign N6627 = N6626 | data_masked[6580];
  assign N6626 = N6625 | data_masked[6708];
  assign N6625 = N6624 | data_masked[6836];
  assign N6624 = N6623 | data_masked[6964];
  assign N6623 = N6622 | data_masked[7092];
  assign N6622 = N6621 | data_masked[7220];
  assign N6621 = N6620 | data_masked[7348];
  assign N6620 = N6619 | data_masked[7476];
  assign N6619 = N6618 | data_masked[7604];
  assign N6618 = N6617 | data_masked[7732];
  assign N6617 = N6616 | data_masked[7860];
  assign N6616 = N6615 | data_masked[7988];
  assign N6615 = N6614 | data_masked[8116];
  assign N6614 = N6613 | data_masked[8244];
  assign N6613 = N6612 | data_masked[8372];
  assign N6612 = N6611 | data_masked[8500];
  assign N6611 = N6610 | data_masked[8628];
  assign N6610 = N6609 | data_masked[8756];
  assign N6609 = N6608 | data_masked[8884];
  assign N6608 = N6607 | data_masked[9012];
  assign N6607 = N6606 | data_masked[9140];
  assign N6606 = N6605 | data_masked[9268];
  assign N6605 = N6604 | data_masked[9396];
  assign N6604 = N6603 | data_masked[9524];
  assign N6603 = N6602 | data_masked[9652];
  assign N6602 = N6601 | data_masked[9780];
  assign N6601 = N6600 | data_masked[9908];
  assign N6600 = N6599 | data_masked[10036];
  assign N6599 = N6598 | data_masked[10164];
  assign N6598 = N6597 | data_masked[10292];
  assign N6597 = N6596 | data_masked[10420];
  assign N6596 = N6595 | data_masked[10548];
  assign N6595 = N6594 | data_masked[10676];
  assign N6594 = N6593 | data_masked[10804];
  assign N6593 = N6592 | data_masked[10932];
  assign N6592 = N6591 | data_masked[11060];
  assign N6591 = N6590 | data_masked[11188];
  assign N6590 = N6589 | data_masked[11316];
  assign N6589 = N6588 | data_masked[11444];
  assign N6588 = N6587 | data_masked[11572];
  assign N6587 = N6586 | data_masked[11700];
  assign N6586 = N6585 | data_masked[11828];
  assign N6585 = N6584 | data_masked[11956];
  assign N6584 = N6583 | data_masked[12084];
  assign N6583 = N6582 | data_masked[12212];
  assign N6582 = N6581 | data_masked[12340];
  assign N6581 = N6580 | data_masked[12468];
  assign N6580 = N6579 | data_masked[12596];
  assign N6579 = N6578 | data_masked[12724];
  assign N6578 = N6577 | data_masked[12852];
  assign N6577 = N6576 | data_masked[12980];
  assign N6576 = N6575 | data_masked[13108];
  assign N6575 = N6574 | data_masked[13236];
  assign N6574 = N6573 | data_masked[13364];
  assign N6573 = N6572 | data_masked[13492];
  assign N6572 = N6571 | data_masked[13620];
  assign N6571 = N6570 | data_masked[13748];
  assign N6570 = N6569 | data_masked[13876];
  assign N6569 = N6568 | data_masked[14004];
  assign N6568 = N6567 | data_masked[14132];
  assign N6567 = N6566 | data_masked[14260];
  assign N6566 = N6565 | data_masked[14388];
  assign N6565 = N6564 | data_masked[14516];
  assign N6564 = N6563 | data_masked[14644];
  assign N6563 = N6562 | data_masked[14772];
  assign N6562 = N6561 | data_masked[14900];
  assign N6561 = N6560 | data_masked[15028];
  assign N6560 = N6559 | data_masked[15156];
  assign N6559 = N6558 | data_masked[15284];
  assign N6558 = N6557 | data_masked[15412];
  assign N6557 = N6556 | data_masked[15540];
  assign N6556 = N6555 | data_masked[15668];
  assign N6555 = N6554 | data_masked[15796];
  assign N6554 = N6553 | data_masked[15924];
  assign N6553 = N6552 | data_masked[16052];
  assign N6552 = data_masked[16308] | data_masked[16180];
  assign data_o[53] = N6803 | data_masked[53];
  assign N6803 = N6802 | data_masked[181];
  assign N6802 = N6801 | data_masked[309];
  assign N6801 = N6800 | data_masked[437];
  assign N6800 = N6799 | data_masked[565];
  assign N6799 = N6798 | data_masked[693];
  assign N6798 = N6797 | data_masked[821];
  assign N6797 = N6796 | data_masked[949];
  assign N6796 = N6795 | data_masked[1077];
  assign N6795 = N6794 | data_masked[1205];
  assign N6794 = N6793 | data_masked[1333];
  assign N6793 = N6792 | data_masked[1461];
  assign N6792 = N6791 | data_masked[1589];
  assign N6791 = N6790 | data_masked[1717];
  assign N6790 = N6789 | data_masked[1845];
  assign N6789 = N6788 | data_masked[1973];
  assign N6788 = N6787 | data_masked[2101];
  assign N6787 = N6786 | data_masked[2229];
  assign N6786 = N6785 | data_masked[2357];
  assign N6785 = N6784 | data_masked[2485];
  assign N6784 = N6783 | data_masked[2613];
  assign N6783 = N6782 | data_masked[2741];
  assign N6782 = N6781 | data_masked[2869];
  assign N6781 = N6780 | data_masked[2997];
  assign N6780 = N6779 | data_masked[3125];
  assign N6779 = N6778 | data_masked[3253];
  assign N6778 = N6777 | data_masked[3381];
  assign N6777 = N6776 | data_masked[3509];
  assign N6776 = N6775 | data_masked[3637];
  assign N6775 = N6774 | data_masked[3765];
  assign N6774 = N6773 | data_masked[3893];
  assign N6773 = N6772 | data_masked[4021];
  assign N6772 = N6771 | data_masked[4149];
  assign N6771 = N6770 | data_masked[4277];
  assign N6770 = N6769 | data_masked[4405];
  assign N6769 = N6768 | data_masked[4533];
  assign N6768 = N6767 | data_masked[4661];
  assign N6767 = N6766 | data_masked[4789];
  assign N6766 = N6765 | data_masked[4917];
  assign N6765 = N6764 | data_masked[5045];
  assign N6764 = N6763 | data_masked[5173];
  assign N6763 = N6762 | data_masked[5301];
  assign N6762 = N6761 | data_masked[5429];
  assign N6761 = N6760 | data_masked[5557];
  assign N6760 = N6759 | data_masked[5685];
  assign N6759 = N6758 | data_masked[5813];
  assign N6758 = N6757 | data_masked[5941];
  assign N6757 = N6756 | data_masked[6069];
  assign N6756 = N6755 | data_masked[6197];
  assign N6755 = N6754 | data_masked[6325];
  assign N6754 = N6753 | data_masked[6453];
  assign N6753 = N6752 | data_masked[6581];
  assign N6752 = N6751 | data_masked[6709];
  assign N6751 = N6750 | data_masked[6837];
  assign N6750 = N6749 | data_masked[6965];
  assign N6749 = N6748 | data_masked[7093];
  assign N6748 = N6747 | data_masked[7221];
  assign N6747 = N6746 | data_masked[7349];
  assign N6746 = N6745 | data_masked[7477];
  assign N6745 = N6744 | data_masked[7605];
  assign N6744 = N6743 | data_masked[7733];
  assign N6743 = N6742 | data_masked[7861];
  assign N6742 = N6741 | data_masked[7989];
  assign N6741 = N6740 | data_masked[8117];
  assign N6740 = N6739 | data_masked[8245];
  assign N6739 = N6738 | data_masked[8373];
  assign N6738 = N6737 | data_masked[8501];
  assign N6737 = N6736 | data_masked[8629];
  assign N6736 = N6735 | data_masked[8757];
  assign N6735 = N6734 | data_masked[8885];
  assign N6734 = N6733 | data_masked[9013];
  assign N6733 = N6732 | data_masked[9141];
  assign N6732 = N6731 | data_masked[9269];
  assign N6731 = N6730 | data_masked[9397];
  assign N6730 = N6729 | data_masked[9525];
  assign N6729 = N6728 | data_masked[9653];
  assign N6728 = N6727 | data_masked[9781];
  assign N6727 = N6726 | data_masked[9909];
  assign N6726 = N6725 | data_masked[10037];
  assign N6725 = N6724 | data_masked[10165];
  assign N6724 = N6723 | data_masked[10293];
  assign N6723 = N6722 | data_masked[10421];
  assign N6722 = N6721 | data_masked[10549];
  assign N6721 = N6720 | data_masked[10677];
  assign N6720 = N6719 | data_masked[10805];
  assign N6719 = N6718 | data_masked[10933];
  assign N6718 = N6717 | data_masked[11061];
  assign N6717 = N6716 | data_masked[11189];
  assign N6716 = N6715 | data_masked[11317];
  assign N6715 = N6714 | data_masked[11445];
  assign N6714 = N6713 | data_masked[11573];
  assign N6713 = N6712 | data_masked[11701];
  assign N6712 = N6711 | data_masked[11829];
  assign N6711 = N6710 | data_masked[11957];
  assign N6710 = N6709 | data_masked[12085];
  assign N6709 = N6708 | data_masked[12213];
  assign N6708 = N6707 | data_masked[12341];
  assign N6707 = N6706 | data_masked[12469];
  assign N6706 = N6705 | data_masked[12597];
  assign N6705 = N6704 | data_masked[12725];
  assign N6704 = N6703 | data_masked[12853];
  assign N6703 = N6702 | data_masked[12981];
  assign N6702 = N6701 | data_masked[13109];
  assign N6701 = N6700 | data_masked[13237];
  assign N6700 = N6699 | data_masked[13365];
  assign N6699 = N6698 | data_masked[13493];
  assign N6698 = N6697 | data_masked[13621];
  assign N6697 = N6696 | data_masked[13749];
  assign N6696 = N6695 | data_masked[13877];
  assign N6695 = N6694 | data_masked[14005];
  assign N6694 = N6693 | data_masked[14133];
  assign N6693 = N6692 | data_masked[14261];
  assign N6692 = N6691 | data_masked[14389];
  assign N6691 = N6690 | data_masked[14517];
  assign N6690 = N6689 | data_masked[14645];
  assign N6689 = N6688 | data_masked[14773];
  assign N6688 = N6687 | data_masked[14901];
  assign N6687 = N6686 | data_masked[15029];
  assign N6686 = N6685 | data_masked[15157];
  assign N6685 = N6684 | data_masked[15285];
  assign N6684 = N6683 | data_masked[15413];
  assign N6683 = N6682 | data_masked[15541];
  assign N6682 = N6681 | data_masked[15669];
  assign N6681 = N6680 | data_masked[15797];
  assign N6680 = N6679 | data_masked[15925];
  assign N6679 = N6678 | data_masked[16053];
  assign N6678 = data_masked[16309] | data_masked[16181];
  assign data_o[54] = N6929 | data_masked[54];
  assign N6929 = N6928 | data_masked[182];
  assign N6928 = N6927 | data_masked[310];
  assign N6927 = N6926 | data_masked[438];
  assign N6926 = N6925 | data_masked[566];
  assign N6925 = N6924 | data_masked[694];
  assign N6924 = N6923 | data_masked[822];
  assign N6923 = N6922 | data_masked[950];
  assign N6922 = N6921 | data_masked[1078];
  assign N6921 = N6920 | data_masked[1206];
  assign N6920 = N6919 | data_masked[1334];
  assign N6919 = N6918 | data_masked[1462];
  assign N6918 = N6917 | data_masked[1590];
  assign N6917 = N6916 | data_masked[1718];
  assign N6916 = N6915 | data_masked[1846];
  assign N6915 = N6914 | data_masked[1974];
  assign N6914 = N6913 | data_masked[2102];
  assign N6913 = N6912 | data_masked[2230];
  assign N6912 = N6911 | data_masked[2358];
  assign N6911 = N6910 | data_masked[2486];
  assign N6910 = N6909 | data_masked[2614];
  assign N6909 = N6908 | data_masked[2742];
  assign N6908 = N6907 | data_masked[2870];
  assign N6907 = N6906 | data_masked[2998];
  assign N6906 = N6905 | data_masked[3126];
  assign N6905 = N6904 | data_masked[3254];
  assign N6904 = N6903 | data_masked[3382];
  assign N6903 = N6902 | data_masked[3510];
  assign N6902 = N6901 | data_masked[3638];
  assign N6901 = N6900 | data_masked[3766];
  assign N6900 = N6899 | data_masked[3894];
  assign N6899 = N6898 | data_masked[4022];
  assign N6898 = N6897 | data_masked[4150];
  assign N6897 = N6896 | data_masked[4278];
  assign N6896 = N6895 | data_masked[4406];
  assign N6895 = N6894 | data_masked[4534];
  assign N6894 = N6893 | data_masked[4662];
  assign N6893 = N6892 | data_masked[4790];
  assign N6892 = N6891 | data_masked[4918];
  assign N6891 = N6890 | data_masked[5046];
  assign N6890 = N6889 | data_masked[5174];
  assign N6889 = N6888 | data_masked[5302];
  assign N6888 = N6887 | data_masked[5430];
  assign N6887 = N6886 | data_masked[5558];
  assign N6886 = N6885 | data_masked[5686];
  assign N6885 = N6884 | data_masked[5814];
  assign N6884 = N6883 | data_masked[5942];
  assign N6883 = N6882 | data_masked[6070];
  assign N6882 = N6881 | data_masked[6198];
  assign N6881 = N6880 | data_masked[6326];
  assign N6880 = N6879 | data_masked[6454];
  assign N6879 = N6878 | data_masked[6582];
  assign N6878 = N6877 | data_masked[6710];
  assign N6877 = N6876 | data_masked[6838];
  assign N6876 = N6875 | data_masked[6966];
  assign N6875 = N6874 | data_masked[7094];
  assign N6874 = N6873 | data_masked[7222];
  assign N6873 = N6872 | data_masked[7350];
  assign N6872 = N6871 | data_masked[7478];
  assign N6871 = N6870 | data_masked[7606];
  assign N6870 = N6869 | data_masked[7734];
  assign N6869 = N6868 | data_masked[7862];
  assign N6868 = N6867 | data_masked[7990];
  assign N6867 = N6866 | data_masked[8118];
  assign N6866 = N6865 | data_masked[8246];
  assign N6865 = N6864 | data_masked[8374];
  assign N6864 = N6863 | data_masked[8502];
  assign N6863 = N6862 | data_masked[8630];
  assign N6862 = N6861 | data_masked[8758];
  assign N6861 = N6860 | data_masked[8886];
  assign N6860 = N6859 | data_masked[9014];
  assign N6859 = N6858 | data_masked[9142];
  assign N6858 = N6857 | data_masked[9270];
  assign N6857 = N6856 | data_masked[9398];
  assign N6856 = N6855 | data_masked[9526];
  assign N6855 = N6854 | data_masked[9654];
  assign N6854 = N6853 | data_masked[9782];
  assign N6853 = N6852 | data_masked[9910];
  assign N6852 = N6851 | data_masked[10038];
  assign N6851 = N6850 | data_masked[10166];
  assign N6850 = N6849 | data_masked[10294];
  assign N6849 = N6848 | data_masked[10422];
  assign N6848 = N6847 | data_masked[10550];
  assign N6847 = N6846 | data_masked[10678];
  assign N6846 = N6845 | data_masked[10806];
  assign N6845 = N6844 | data_masked[10934];
  assign N6844 = N6843 | data_masked[11062];
  assign N6843 = N6842 | data_masked[11190];
  assign N6842 = N6841 | data_masked[11318];
  assign N6841 = N6840 | data_masked[11446];
  assign N6840 = N6839 | data_masked[11574];
  assign N6839 = N6838 | data_masked[11702];
  assign N6838 = N6837 | data_masked[11830];
  assign N6837 = N6836 | data_masked[11958];
  assign N6836 = N6835 | data_masked[12086];
  assign N6835 = N6834 | data_masked[12214];
  assign N6834 = N6833 | data_masked[12342];
  assign N6833 = N6832 | data_masked[12470];
  assign N6832 = N6831 | data_masked[12598];
  assign N6831 = N6830 | data_masked[12726];
  assign N6830 = N6829 | data_masked[12854];
  assign N6829 = N6828 | data_masked[12982];
  assign N6828 = N6827 | data_masked[13110];
  assign N6827 = N6826 | data_masked[13238];
  assign N6826 = N6825 | data_masked[13366];
  assign N6825 = N6824 | data_masked[13494];
  assign N6824 = N6823 | data_masked[13622];
  assign N6823 = N6822 | data_masked[13750];
  assign N6822 = N6821 | data_masked[13878];
  assign N6821 = N6820 | data_masked[14006];
  assign N6820 = N6819 | data_masked[14134];
  assign N6819 = N6818 | data_masked[14262];
  assign N6818 = N6817 | data_masked[14390];
  assign N6817 = N6816 | data_masked[14518];
  assign N6816 = N6815 | data_masked[14646];
  assign N6815 = N6814 | data_masked[14774];
  assign N6814 = N6813 | data_masked[14902];
  assign N6813 = N6812 | data_masked[15030];
  assign N6812 = N6811 | data_masked[15158];
  assign N6811 = N6810 | data_masked[15286];
  assign N6810 = N6809 | data_masked[15414];
  assign N6809 = N6808 | data_masked[15542];
  assign N6808 = N6807 | data_masked[15670];
  assign N6807 = N6806 | data_masked[15798];
  assign N6806 = N6805 | data_masked[15926];
  assign N6805 = N6804 | data_masked[16054];
  assign N6804 = data_masked[16310] | data_masked[16182];
  assign data_o[55] = N7055 | data_masked[55];
  assign N7055 = N7054 | data_masked[183];
  assign N7054 = N7053 | data_masked[311];
  assign N7053 = N7052 | data_masked[439];
  assign N7052 = N7051 | data_masked[567];
  assign N7051 = N7050 | data_masked[695];
  assign N7050 = N7049 | data_masked[823];
  assign N7049 = N7048 | data_masked[951];
  assign N7048 = N7047 | data_masked[1079];
  assign N7047 = N7046 | data_masked[1207];
  assign N7046 = N7045 | data_masked[1335];
  assign N7045 = N7044 | data_masked[1463];
  assign N7044 = N7043 | data_masked[1591];
  assign N7043 = N7042 | data_masked[1719];
  assign N7042 = N7041 | data_masked[1847];
  assign N7041 = N7040 | data_masked[1975];
  assign N7040 = N7039 | data_masked[2103];
  assign N7039 = N7038 | data_masked[2231];
  assign N7038 = N7037 | data_masked[2359];
  assign N7037 = N7036 | data_masked[2487];
  assign N7036 = N7035 | data_masked[2615];
  assign N7035 = N7034 | data_masked[2743];
  assign N7034 = N7033 | data_masked[2871];
  assign N7033 = N7032 | data_masked[2999];
  assign N7032 = N7031 | data_masked[3127];
  assign N7031 = N7030 | data_masked[3255];
  assign N7030 = N7029 | data_masked[3383];
  assign N7029 = N7028 | data_masked[3511];
  assign N7028 = N7027 | data_masked[3639];
  assign N7027 = N7026 | data_masked[3767];
  assign N7026 = N7025 | data_masked[3895];
  assign N7025 = N7024 | data_masked[4023];
  assign N7024 = N7023 | data_masked[4151];
  assign N7023 = N7022 | data_masked[4279];
  assign N7022 = N7021 | data_masked[4407];
  assign N7021 = N7020 | data_masked[4535];
  assign N7020 = N7019 | data_masked[4663];
  assign N7019 = N7018 | data_masked[4791];
  assign N7018 = N7017 | data_masked[4919];
  assign N7017 = N7016 | data_masked[5047];
  assign N7016 = N7015 | data_masked[5175];
  assign N7015 = N7014 | data_masked[5303];
  assign N7014 = N7013 | data_masked[5431];
  assign N7013 = N7012 | data_masked[5559];
  assign N7012 = N7011 | data_masked[5687];
  assign N7011 = N7010 | data_masked[5815];
  assign N7010 = N7009 | data_masked[5943];
  assign N7009 = N7008 | data_masked[6071];
  assign N7008 = N7007 | data_masked[6199];
  assign N7007 = N7006 | data_masked[6327];
  assign N7006 = N7005 | data_masked[6455];
  assign N7005 = N7004 | data_masked[6583];
  assign N7004 = N7003 | data_masked[6711];
  assign N7003 = N7002 | data_masked[6839];
  assign N7002 = N7001 | data_masked[6967];
  assign N7001 = N7000 | data_masked[7095];
  assign N7000 = N6999 | data_masked[7223];
  assign N6999 = N6998 | data_masked[7351];
  assign N6998 = N6997 | data_masked[7479];
  assign N6997 = N6996 | data_masked[7607];
  assign N6996 = N6995 | data_masked[7735];
  assign N6995 = N6994 | data_masked[7863];
  assign N6994 = N6993 | data_masked[7991];
  assign N6993 = N6992 | data_masked[8119];
  assign N6992 = N6991 | data_masked[8247];
  assign N6991 = N6990 | data_masked[8375];
  assign N6990 = N6989 | data_masked[8503];
  assign N6989 = N6988 | data_masked[8631];
  assign N6988 = N6987 | data_masked[8759];
  assign N6987 = N6986 | data_masked[8887];
  assign N6986 = N6985 | data_masked[9015];
  assign N6985 = N6984 | data_masked[9143];
  assign N6984 = N6983 | data_masked[9271];
  assign N6983 = N6982 | data_masked[9399];
  assign N6982 = N6981 | data_masked[9527];
  assign N6981 = N6980 | data_masked[9655];
  assign N6980 = N6979 | data_masked[9783];
  assign N6979 = N6978 | data_masked[9911];
  assign N6978 = N6977 | data_masked[10039];
  assign N6977 = N6976 | data_masked[10167];
  assign N6976 = N6975 | data_masked[10295];
  assign N6975 = N6974 | data_masked[10423];
  assign N6974 = N6973 | data_masked[10551];
  assign N6973 = N6972 | data_masked[10679];
  assign N6972 = N6971 | data_masked[10807];
  assign N6971 = N6970 | data_masked[10935];
  assign N6970 = N6969 | data_masked[11063];
  assign N6969 = N6968 | data_masked[11191];
  assign N6968 = N6967 | data_masked[11319];
  assign N6967 = N6966 | data_masked[11447];
  assign N6966 = N6965 | data_masked[11575];
  assign N6965 = N6964 | data_masked[11703];
  assign N6964 = N6963 | data_masked[11831];
  assign N6963 = N6962 | data_masked[11959];
  assign N6962 = N6961 | data_masked[12087];
  assign N6961 = N6960 | data_masked[12215];
  assign N6960 = N6959 | data_masked[12343];
  assign N6959 = N6958 | data_masked[12471];
  assign N6958 = N6957 | data_masked[12599];
  assign N6957 = N6956 | data_masked[12727];
  assign N6956 = N6955 | data_masked[12855];
  assign N6955 = N6954 | data_masked[12983];
  assign N6954 = N6953 | data_masked[13111];
  assign N6953 = N6952 | data_masked[13239];
  assign N6952 = N6951 | data_masked[13367];
  assign N6951 = N6950 | data_masked[13495];
  assign N6950 = N6949 | data_masked[13623];
  assign N6949 = N6948 | data_masked[13751];
  assign N6948 = N6947 | data_masked[13879];
  assign N6947 = N6946 | data_masked[14007];
  assign N6946 = N6945 | data_masked[14135];
  assign N6945 = N6944 | data_masked[14263];
  assign N6944 = N6943 | data_masked[14391];
  assign N6943 = N6942 | data_masked[14519];
  assign N6942 = N6941 | data_masked[14647];
  assign N6941 = N6940 | data_masked[14775];
  assign N6940 = N6939 | data_masked[14903];
  assign N6939 = N6938 | data_masked[15031];
  assign N6938 = N6937 | data_masked[15159];
  assign N6937 = N6936 | data_masked[15287];
  assign N6936 = N6935 | data_masked[15415];
  assign N6935 = N6934 | data_masked[15543];
  assign N6934 = N6933 | data_masked[15671];
  assign N6933 = N6932 | data_masked[15799];
  assign N6932 = N6931 | data_masked[15927];
  assign N6931 = N6930 | data_masked[16055];
  assign N6930 = data_masked[16311] | data_masked[16183];
  assign data_o[56] = N7181 | data_masked[56];
  assign N7181 = N7180 | data_masked[184];
  assign N7180 = N7179 | data_masked[312];
  assign N7179 = N7178 | data_masked[440];
  assign N7178 = N7177 | data_masked[568];
  assign N7177 = N7176 | data_masked[696];
  assign N7176 = N7175 | data_masked[824];
  assign N7175 = N7174 | data_masked[952];
  assign N7174 = N7173 | data_masked[1080];
  assign N7173 = N7172 | data_masked[1208];
  assign N7172 = N7171 | data_masked[1336];
  assign N7171 = N7170 | data_masked[1464];
  assign N7170 = N7169 | data_masked[1592];
  assign N7169 = N7168 | data_masked[1720];
  assign N7168 = N7167 | data_masked[1848];
  assign N7167 = N7166 | data_masked[1976];
  assign N7166 = N7165 | data_masked[2104];
  assign N7165 = N7164 | data_masked[2232];
  assign N7164 = N7163 | data_masked[2360];
  assign N7163 = N7162 | data_masked[2488];
  assign N7162 = N7161 | data_masked[2616];
  assign N7161 = N7160 | data_masked[2744];
  assign N7160 = N7159 | data_masked[2872];
  assign N7159 = N7158 | data_masked[3000];
  assign N7158 = N7157 | data_masked[3128];
  assign N7157 = N7156 | data_masked[3256];
  assign N7156 = N7155 | data_masked[3384];
  assign N7155 = N7154 | data_masked[3512];
  assign N7154 = N7153 | data_masked[3640];
  assign N7153 = N7152 | data_masked[3768];
  assign N7152 = N7151 | data_masked[3896];
  assign N7151 = N7150 | data_masked[4024];
  assign N7150 = N7149 | data_masked[4152];
  assign N7149 = N7148 | data_masked[4280];
  assign N7148 = N7147 | data_masked[4408];
  assign N7147 = N7146 | data_masked[4536];
  assign N7146 = N7145 | data_masked[4664];
  assign N7145 = N7144 | data_masked[4792];
  assign N7144 = N7143 | data_masked[4920];
  assign N7143 = N7142 | data_masked[5048];
  assign N7142 = N7141 | data_masked[5176];
  assign N7141 = N7140 | data_masked[5304];
  assign N7140 = N7139 | data_masked[5432];
  assign N7139 = N7138 | data_masked[5560];
  assign N7138 = N7137 | data_masked[5688];
  assign N7137 = N7136 | data_masked[5816];
  assign N7136 = N7135 | data_masked[5944];
  assign N7135 = N7134 | data_masked[6072];
  assign N7134 = N7133 | data_masked[6200];
  assign N7133 = N7132 | data_masked[6328];
  assign N7132 = N7131 | data_masked[6456];
  assign N7131 = N7130 | data_masked[6584];
  assign N7130 = N7129 | data_masked[6712];
  assign N7129 = N7128 | data_masked[6840];
  assign N7128 = N7127 | data_masked[6968];
  assign N7127 = N7126 | data_masked[7096];
  assign N7126 = N7125 | data_masked[7224];
  assign N7125 = N7124 | data_masked[7352];
  assign N7124 = N7123 | data_masked[7480];
  assign N7123 = N7122 | data_masked[7608];
  assign N7122 = N7121 | data_masked[7736];
  assign N7121 = N7120 | data_masked[7864];
  assign N7120 = N7119 | data_masked[7992];
  assign N7119 = N7118 | data_masked[8120];
  assign N7118 = N7117 | data_masked[8248];
  assign N7117 = N7116 | data_masked[8376];
  assign N7116 = N7115 | data_masked[8504];
  assign N7115 = N7114 | data_masked[8632];
  assign N7114 = N7113 | data_masked[8760];
  assign N7113 = N7112 | data_masked[8888];
  assign N7112 = N7111 | data_masked[9016];
  assign N7111 = N7110 | data_masked[9144];
  assign N7110 = N7109 | data_masked[9272];
  assign N7109 = N7108 | data_masked[9400];
  assign N7108 = N7107 | data_masked[9528];
  assign N7107 = N7106 | data_masked[9656];
  assign N7106 = N7105 | data_masked[9784];
  assign N7105 = N7104 | data_masked[9912];
  assign N7104 = N7103 | data_masked[10040];
  assign N7103 = N7102 | data_masked[10168];
  assign N7102 = N7101 | data_masked[10296];
  assign N7101 = N7100 | data_masked[10424];
  assign N7100 = N7099 | data_masked[10552];
  assign N7099 = N7098 | data_masked[10680];
  assign N7098 = N7097 | data_masked[10808];
  assign N7097 = N7096 | data_masked[10936];
  assign N7096 = N7095 | data_masked[11064];
  assign N7095 = N7094 | data_masked[11192];
  assign N7094 = N7093 | data_masked[11320];
  assign N7093 = N7092 | data_masked[11448];
  assign N7092 = N7091 | data_masked[11576];
  assign N7091 = N7090 | data_masked[11704];
  assign N7090 = N7089 | data_masked[11832];
  assign N7089 = N7088 | data_masked[11960];
  assign N7088 = N7087 | data_masked[12088];
  assign N7087 = N7086 | data_masked[12216];
  assign N7086 = N7085 | data_masked[12344];
  assign N7085 = N7084 | data_masked[12472];
  assign N7084 = N7083 | data_masked[12600];
  assign N7083 = N7082 | data_masked[12728];
  assign N7082 = N7081 | data_masked[12856];
  assign N7081 = N7080 | data_masked[12984];
  assign N7080 = N7079 | data_masked[13112];
  assign N7079 = N7078 | data_masked[13240];
  assign N7078 = N7077 | data_masked[13368];
  assign N7077 = N7076 | data_masked[13496];
  assign N7076 = N7075 | data_masked[13624];
  assign N7075 = N7074 | data_masked[13752];
  assign N7074 = N7073 | data_masked[13880];
  assign N7073 = N7072 | data_masked[14008];
  assign N7072 = N7071 | data_masked[14136];
  assign N7071 = N7070 | data_masked[14264];
  assign N7070 = N7069 | data_masked[14392];
  assign N7069 = N7068 | data_masked[14520];
  assign N7068 = N7067 | data_masked[14648];
  assign N7067 = N7066 | data_masked[14776];
  assign N7066 = N7065 | data_masked[14904];
  assign N7065 = N7064 | data_masked[15032];
  assign N7064 = N7063 | data_masked[15160];
  assign N7063 = N7062 | data_masked[15288];
  assign N7062 = N7061 | data_masked[15416];
  assign N7061 = N7060 | data_masked[15544];
  assign N7060 = N7059 | data_masked[15672];
  assign N7059 = N7058 | data_masked[15800];
  assign N7058 = N7057 | data_masked[15928];
  assign N7057 = N7056 | data_masked[16056];
  assign N7056 = data_masked[16312] | data_masked[16184];
  assign data_o[57] = N7307 | data_masked[57];
  assign N7307 = N7306 | data_masked[185];
  assign N7306 = N7305 | data_masked[313];
  assign N7305 = N7304 | data_masked[441];
  assign N7304 = N7303 | data_masked[569];
  assign N7303 = N7302 | data_masked[697];
  assign N7302 = N7301 | data_masked[825];
  assign N7301 = N7300 | data_masked[953];
  assign N7300 = N7299 | data_masked[1081];
  assign N7299 = N7298 | data_masked[1209];
  assign N7298 = N7297 | data_masked[1337];
  assign N7297 = N7296 | data_masked[1465];
  assign N7296 = N7295 | data_masked[1593];
  assign N7295 = N7294 | data_masked[1721];
  assign N7294 = N7293 | data_masked[1849];
  assign N7293 = N7292 | data_masked[1977];
  assign N7292 = N7291 | data_masked[2105];
  assign N7291 = N7290 | data_masked[2233];
  assign N7290 = N7289 | data_masked[2361];
  assign N7289 = N7288 | data_masked[2489];
  assign N7288 = N7287 | data_masked[2617];
  assign N7287 = N7286 | data_masked[2745];
  assign N7286 = N7285 | data_masked[2873];
  assign N7285 = N7284 | data_masked[3001];
  assign N7284 = N7283 | data_masked[3129];
  assign N7283 = N7282 | data_masked[3257];
  assign N7282 = N7281 | data_masked[3385];
  assign N7281 = N7280 | data_masked[3513];
  assign N7280 = N7279 | data_masked[3641];
  assign N7279 = N7278 | data_masked[3769];
  assign N7278 = N7277 | data_masked[3897];
  assign N7277 = N7276 | data_masked[4025];
  assign N7276 = N7275 | data_masked[4153];
  assign N7275 = N7274 | data_masked[4281];
  assign N7274 = N7273 | data_masked[4409];
  assign N7273 = N7272 | data_masked[4537];
  assign N7272 = N7271 | data_masked[4665];
  assign N7271 = N7270 | data_masked[4793];
  assign N7270 = N7269 | data_masked[4921];
  assign N7269 = N7268 | data_masked[5049];
  assign N7268 = N7267 | data_masked[5177];
  assign N7267 = N7266 | data_masked[5305];
  assign N7266 = N7265 | data_masked[5433];
  assign N7265 = N7264 | data_masked[5561];
  assign N7264 = N7263 | data_masked[5689];
  assign N7263 = N7262 | data_masked[5817];
  assign N7262 = N7261 | data_masked[5945];
  assign N7261 = N7260 | data_masked[6073];
  assign N7260 = N7259 | data_masked[6201];
  assign N7259 = N7258 | data_masked[6329];
  assign N7258 = N7257 | data_masked[6457];
  assign N7257 = N7256 | data_masked[6585];
  assign N7256 = N7255 | data_masked[6713];
  assign N7255 = N7254 | data_masked[6841];
  assign N7254 = N7253 | data_masked[6969];
  assign N7253 = N7252 | data_masked[7097];
  assign N7252 = N7251 | data_masked[7225];
  assign N7251 = N7250 | data_masked[7353];
  assign N7250 = N7249 | data_masked[7481];
  assign N7249 = N7248 | data_masked[7609];
  assign N7248 = N7247 | data_masked[7737];
  assign N7247 = N7246 | data_masked[7865];
  assign N7246 = N7245 | data_masked[7993];
  assign N7245 = N7244 | data_masked[8121];
  assign N7244 = N7243 | data_masked[8249];
  assign N7243 = N7242 | data_masked[8377];
  assign N7242 = N7241 | data_masked[8505];
  assign N7241 = N7240 | data_masked[8633];
  assign N7240 = N7239 | data_masked[8761];
  assign N7239 = N7238 | data_masked[8889];
  assign N7238 = N7237 | data_masked[9017];
  assign N7237 = N7236 | data_masked[9145];
  assign N7236 = N7235 | data_masked[9273];
  assign N7235 = N7234 | data_masked[9401];
  assign N7234 = N7233 | data_masked[9529];
  assign N7233 = N7232 | data_masked[9657];
  assign N7232 = N7231 | data_masked[9785];
  assign N7231 = N7230 | data_masked[9913];
  assign N7230 = N7229 | data_masked[10041];
  assign N7229 = N7228 | data_masked[10169];
  assign N7228 = N7227 | data_masked[10297];
  assign N7227 = N7226 | data_masked[10425];
  assign N7226 = N7225 | data_masked[10553];
  assign N7225 = N7224 | data_masked[10681];
  assign N7224 = N7223 | data_masked[10809];
  assign N7223 = N7222 | data_masked[10937];
  assign N7222 = N7221 | data_masked[11065];
  assign N7221 = N7220 | data_masked[11193];
  assign N7220 = N7219 | data_masked[11321];
  assign N7219 = N7218 | data_masked[11449];
  assign N7218 = N7217 | data_masked[11577];
  assign N7217 = N7216 | data_masked[11705];
  assign N7216 = N7215 | data_masked[11833];
  assign N7215 = N7214 | data_masked[11961];
  assign N7214 = N7213 | data_masked[12089];
  assign N7213 = N7212 | data_masked[12217];
  assign N7212 = N7211 | data_masked[12345];
  assign N7211 = N7210 | data_masked[12473];
  assign N7210 = N7209 | data_masked[12601];
  assign N7209 = N7208 | data_masked[12729];
  assign N7208 = N7207 | data_masked[12857];
  assign N7207 = N7206 | data_masked[12985];
  assign N7206 = N7205 | data_masked[13113];
  assign N7205 = N7204 | data_masked[13241];
  assign N7204 = N7203 | data_masked[13369];
  assign N7203 = N7202 | data_masked[13497];
  assign N7202 = N7201 | data_masked[13625];
  assign N7201 = N7200 | data_masked[13753];
  assign N7200 = N7199 | data_masked[13881];
  assign N7199 = N7198 | data_masked[14009];
  assign N7198 = N7197 | data_masked[14137];
  assign N7197 = N7196 | data_masked[14265];
  assign N7196 = N7195 | data_masked[14393];
  assign N7195 = N7194 | data_masked[14521];
  assign N7194 = N7193 | data_masked[14649];
  assign N7193 = N7192 | data_masked[14777];
  assign N7192 = N7191 | data_masked[14905];
  assign N7191 = N7190 | data_masked[15033];
  assign N7190 = N7189 | data_masked[15161];
  assign N7189 = N7188 | data_masked[15289];
  assign N7188 = N7187 | data_masked[15417];
  assign N7187 = N7186 | data_masked[15545];
  assign N7186 = N7185 | data_masked[15673];
  assign N7185 = N7184 | data_masked[15801];
  assign N7184 = N7183 | data_masked[15929];
  assign N7183 = N7182 | data_masked[16057];
  assign N7182 = data_masked[16313] | data_masked[16185];
  assign data_o[58] = N7433 | data_masked[58];
  assign N7433 = N7432 | data_masked[186];
  assign N7432 = N7431 | data_masked[314];
  assign N7431 = N7430 | data_masked[442];
  assign N7430 = N7429 | data_masked[570];
  assign N7429 = N7428 | data_masked[698];
  assign N7428 = N7427 | data_masked[826];
  assign N7427 = N7426 | data_masked[954];
  assign N7426 = N7425 | data_masked[1082];
  assign N7425 = N7424 | data_masked[1210];
  assign N7424 = N7423 | data_masked[1338];
  assign N7423 = N7422 | data_masked[1466];
  assign N7422 = N7421 | data_masked[1594];
  assign N7421 = N7420 | data_masked[1722];
  assign N7420 = N7419 | data_masked[1850];
  assign N7419 = N7418 | data_masked[1978];
  assign N7418 = N7417 | data_masked[2106];
  assign N7417 = N7416 | data_masked[2234];
  assign N7416 = N7415 | data_masked[2362];
  assign N7415 = N7414 | data_masked[2490];
  assign N7414 = N7413 | data_masked[2618];
  assign N7413 = N7412 | data_masked[2746];
  assign N7412 = N7411 | data_masked[2874];
  assign N7411 = N7410 | data_masked[3002];
  assign N7410 = N7409 | data_masked[3130];
  assign N7409 = N7408 | data_masked[3258];
  assign N7408 = N7407 | data_masked[3386];
  assign N7407 = N7406 | data_masked[3514];
  assign N7406 = N7405 | data_masked[3642];
  assign N7405 = N7404 | data_masked[3770];
  assign N7404 = N7403 | data_masked[3898];
  assign N7403 = N7402 | data_masked[4026];
  assign N7402 = N7401 | data_masked[4154];
  assign N7401 = N7400 | data_masked[4282];
  assign N7400 = N7399 | data_masked[4410];
  assign N7399 = N7398 | data_masked[4538];
  assign N7398 = N7397 | data_masked[4666];
  assign N7397 = N7396 | data_masked[4794];
  assign N7396 = N7395 | data_masked[4922];
  assign N7395 = N7394 | data_masked[5050];
  assign N7394 = N7393 | data_masked[5178];
  assign N7393 = N7392 | data_masked[5306];
  assign N7392 = N7391 | data_masked[5434];
  assign N7391 = N7390 | data_masked[5562];
  assign N7390 = N7389 | data_masked[5690];
  assign N7389 = N7388 | data_masked[5818];
  assign N7388 = N7387 | data_masked[5946];
  assign N7387 = N7386 | data_masked[6074];
  assign N7386 = N7385 | data_masked[6202];
  assign N7385 = N7384 | data_masked[6330];
  assign N7384 = N7383 | data_masked[6458];
  assign N7383 = N7382 | data_masked[6586];
  assign N7382 = N7381 | data_masked[6714];
  assign N7381 = N7380 | data_masked[6842];
  assign N7380 = N7379 | data_masked[6970];
  assign N7379 = N7378 | data_masked[7098];
  assign N7378 = N7377 | data_masked[7226];
  assign N7377 = N7376 | data_masked[7354];
  assign N7376 = N7375 | data_masked[7482];
  assign N7375 = N7374 | data_masked[7610];
  assign N7374 = N7373 | data_masked[7738];
  assign N7373 = N7372 | data_masked[7866];
  assign N7372 = N7371 | data_masked[7994];
  assign N7371 = N7370 | data_masked[8122];
  assign N7370 = N7369 | data_masked[8250];
  assign N7369 = N7368 | data_masked[8378];
  assign N7368 = N7367 | data_masked[8506];
  assign N7367 = N7366 | data_masked[8634];
  assign N7366 = N7365 | data_masked[8762];
  assign N7365 = N7364 | data_masked[8890];
  assign N7364 = N7363 | data_masked[9018];
  assign N7363 = N7362 | data_masked[9146];
  assign N7362 = N7361 | data_masked[9274];
  assign N7361 = N7360 | data_masked[9402];
  assign N7360 = N7359 | data_masked[9530];
  assign N7359 = N7358 | data_masked[9658];
  assign N7358 = N7357 | data_masked[9786];
  assign N7357 = N7356 | data_masked[9914];
  assign N7356 = N7355 | data_masked[10042];
  assign N7355 = N7354 | data_masked[10170];
  assign N7354 = N7353 | data_masked[10298];
  assign N7353 = N7352 | data_masked[10426];
  assign N7352 = N7351 | data_masked[10554];
  assign N7351 = N7350 | data_masked[10682];
  assign N7350 = N7349 | data_masked[10810];
  assign N7349 = N7348 | data_masked[10938];
  assign N7348 = N7347 | data_masked[11066];
  assign N7347 = N7346 | data_masked[11194];
  assign N7346 = N7345 | data_masked[11322];
  assign N7345 = N7344 | data_masked[11450];
  assign N7344 = N7343 | data_masked[11578];
  assign N7343 = N7342 | data_masked[11706];
  assign N7342 = N7341 | data_masked[11834];
  assign N7341 = N7340 | data_masked[11962];
  assign N7340 = N7339 | data_masked[12090];
  assign N7339 = N7338 | data_masked[12218];
  assign N7338 = N7337 | data_masked[12346];
  assign N7337 = N7336 | data_masked[12474];
  assign N7336 = N7335 | data_masked[12602];
  assign N7335 = N7334 | data_masked[12730];
  assign N7334 = N7333 | data_masked[12858];
  assign N7333 = N7332 | data_masked[12986];
  assign N7332 = N7331 | data_masked[13114];
  assign N7331 = N7330 | data_masked[13242];
  assign N7330 = N7329 | data_masked[13370];
  assign N7329 = N7328 | data_masked[13498];
  assign N7328 = N7327 | data_masked[13626];
  assign N7327 = N7326 | data_masked[13754];
  assign N7326 = N7325 | data_masked[13882];
  assign N7325 = N7324 | data_masked[14010];
  assign N7324 = N7323 | data_masked[14138];
  assign N7323 = N7322 | data_masked[14266];
  assign N7322 = N7321 | data_masked[14394];
  assign N7321 = N7320 | data_masked[14522];
  assign N7320 = N7319 | data_masked[14650];
  assign N7319 = N7318 | data_masked[14778];
  assign N7318 = N7317 | data_masked[14906];
  assign N7317 = N7316 | data_masked[15034];
  assign N7316 = N7315 | data_masked[15162];
  assign N7315 = N7314 | data_masked[15290];
  assign N7314 = N7313 | data_masked[15418];
  assign N7313 = N7312 | data_masked[15546];
  assign N7312 = N7311 | data_masked[15674];
  assign N7311 = N7310 | data_masked[15802];
  assign N7310 = N7309 | data_masked[15930];
  assign N7309 = N7308 | data_masked[16058];
  assign N7308 = data_masked[16314] | data_masked[16186];
  assign data_o[59] = N7559 | data_masked[59];
  assign N7559 = N7558 | data_masked[187];
  assign N7558 = N7557 | data_masked[315];
  assign N7557 = N7556 | data_masked[443];
  assign N7556 = N7555 | data_masked[571];
  assign N7555 = N7554 | data_masked[699];
  assign N7554 = N7553 | data_masked[827];
  assign N7553 = N7552 | data_masked[955];
  assign N7552 = N7551 | data_masked[1083];
  assign N7551 = N7550 | data_masked[1211];
  assign N7550 = N7549 | data_masked[1339];
  assign N7549 = N7548 | data_masked[1467];
  assign N7548 = N7547 | data_masked[1595];
  assign N7547 = N7546 | data_masked[1723];
  assign N7546 = N7545 | data_masked[1851];
  assign N7545 = N7544 | data_masked[1979];
  assign N7544 = N7543 | data_masked[2107];
  assign N7543 = N7542 | data_masked[2235];
  assign N7542 = N7541 | data_masked[2363];
  assign N7541 = N7540 | data_masked[2491];
  assign N7540 = N7539 | data_masked[2619];
  assign N7539 = N7538 | data_masked[2747];
  assign N7538 = N7537 | data_masked[2875];
  assign N7537 = N7536 | data_masked[3003];
  assign N7536 = N7535 | data_masked[3131];
  assign N7535 = N7534 | data_masked[3259];
  assign N7534 = N7533 | data_masked[3387];
  assign N7533 = N7532 | data_masked[3515];
  assign N7532 = N7531 | data_masked[3643];
  assign N7531 = N7530 | data_masked[3771];
  assign N7530 = N7529 | data_masked[3899];
  assign N7529 = N7528 | data_masked[4027];
  assign N7528 = N7527 | data_masked[4155];
  assign N7527 = N7526 | data_masked[4283];
  assign N7526 = N7525 | data_masked[4411];
  assign N7525 = N7524 | data_masked[4539];
  assign N7524 = N7523 | data_masked[4667];
  assign N7523 = N7522 | data_masked[4795];
  assign N7522 = N7521 | data_masked[4923];
  assign N7521 = N7520 | data_masked[5051];
  assign N7520 = N7519 | data_masked[5179];
  assign N7519 = N7518 | data_masked[5307];
  assign N7518 = N7517 | data_masked[5435];
  assign N7517 = N7516 | data_masked[5563];
  assign N7516 = N7515 | data_masked[5691];
  assign N7515 = N7514 | data_masked[5819];
  assign N7514 = N7513 | data_masked[5947];
  assign N7513 = N7512 | data_masked[6075];
  assign N7512 = N7511 | data_masked[6203];
  assign N7511 = N7510 | data_masked[6331];
  assign N7510 = N7509 | data_masked[6459];
  assign N7509 = N7508 | data_masked[6587];
  assign N7508 = N7507 | data_masked[6715];
  assign N7507 = N7506 | data_masked[6843];
  assign N7506 = N7505 | data_masked[6971];
  assign N7505 = N7504 | data_masked[7099];
  assign N7504 = N7503 | data_masked[7227];
  assign N7503 = N7502 | data_masked[7355];
  assign N7502 = N7501 | data_masked[7483];
  assign N7501 = N7500 | data_masked[7611];
  assign N7500 = N7499 | data_masked[7739];
  assign N7499 = N7498 | data_masked[7867];
  assign N7498 = N7497 | data_masked[7995];
  assign N7497 = N7496 | data_masked[8123];
  assign N7496 = N7495 | data_masked[8251];
  assign N7495 = N7494 | data_masked[8379];
  assign N7494 = N7493 | data_masked[8507];
  assign N7493 = N7492 | data_masked[8635];
  assign N7492 = N7491 | data_masked[8763];
  assign N7491 = N7490 | data_masked[8891];
  assign N7490 = N7489 | data_masked[9019];
  assign N7489 = N7488 | data_masked[9147];
  assign N7488 = N7487 | data_masked[9275];
  assign N7487 = N7486 | data_masked[9403];
  assign N7486 = N7485 | data_masked[9531];
  assign N7485 = N7484 | data_masked[9659];
  assign N7484 = N7483 | data_masked[9787];
  assign N7483 = N7482 | data_masked[9915];
  assign N7482 = N7481 | data_masked[10043];
  assign N7481 = N7480 | data_masked[10171];
  assign N7480 = N7479 | data_masked[10299];
  assign N7479 = N7478 | data_masked[10427];
  assign N7478 = N7477 | data_masked[10555];
  assign N7477 = N7476 | data_masked[10683];
  assign N7476 = N7475 | data_masked[10811];
  assign N7475 = N7474 | data_masked[10939];
  assign N7474 = N7473 | data_masked[11067];
  assign N7473 = N7472 | data_masked[11195];
  assign N7472 = N7471 | data_masked[11323];
  assign N7471 = N7470 | data_masked[11451];
  assign N7470 = N7469 | data_masked[11579];
  assign N7469 = N7468 | data_masked[11707];
  assign N7468 = N7467 | data_masked[11835];
  assign N7467 = N7466 | data_masked[11963];
  assign N7466 = N7465 | data_masked[12091];
  assign N7465 = N7464 | data_masked[12219];
  assign N7464 = N7463 | data_masked[12347];
  assign N7463 = N7462 | data_masked[12475];
  assign N7462 = N7461 | data_masked[12603];
  assign N7461 = N7460 | data_masked[12731];
  assign N7460 = N7459 | data_masked[12859];
  assign N7459 = N7458 | data_masked[12987];
  assign N7458 = N7457 | data_masked[13115];
  assign N7457 = N7456 | data_masked[13243];
  assign N7456 = N7455 | data_masked[13371];
  assign N7455 = N7454 | data_masked[13499];
  assign N7454 = N7453 | data_masked[13627];
  assign N7453 = N7452 | data_masked[13755];
  assign N7452 = N7451 | data_masked[13883];
  assign N7451 = N7450 | data_masked[14011];
  assign N7450 = N7449 | data_masked[14139];
  assign N7449 = N7448 | data_masked[14267];
  assign N7448 = N7447 | data_masked[14395];
  assign N7447 = N7446 | data_masked[14523];
  assign N7446 = N7445 | data_masked[14651];
  assign N7445 = N7444 | data_masked[14779];
  assign N7444 = N7443 | data_masked[14907];
  assign N7443 = N7442 | data_masked[15035];
  assign N7442 = N7441 | data_masked[15163];
  assign N7441 = N7440 | data_masked[15291];
  assign N7440 = N7439 | data_masked[15419];
  assign N7439 = N7438 | data_masked[15547];
  assign N7438 = N7437 | data_masked[15675];
  assign N7437 = N7436 | data_masked[15803];
  assign N7436 = N7435 | data_masked[15931];
  assign N7435 = N7434 | data_masked[16059];
  assign N7434 = data_masked[16315] | data_masked[16187];
  assign data_o[60] = N7685 | data_masked[60];
  assign N7685 = N7684 | data_masked[188];
  assign N7684 = N7683 | data_masked[316];
  assign N7683 = N7682 | data_masked[444];
  assign N7682 = N7681 | data_masked[572];
  assign N7681 = N7680 | data_masked[700];
  assign N7680 = N7679 | data_masked[828];
  assign N7679 = N7678 | data_masked[956];
  assign N7678 = N7677 | data_masked[1084];
  assign N7677 = N7676 | data_masked[1212];
  assign N7676 = N7675 | data_masked[1340];
  assign N7675 = N7674 | data_masked[1468];
  assign N7674 = N7673 | data_masked[1596];
  assign N7673 = N7672 | data_masked[1724];
  assign N7672 = N7671 | data_masked[1852];
  assign N7671 = N7670 | data_masked[1980];
  assign N7670 = N7669 | data_masked[2108];
  assign N7669 = N7668 | data_masked[2236];
  assign N7668 = N7667 | data_masked[2364];
  assign N7667 = N7666 | data_masked[2492];
  assign N7666 = N7665 | data_masked[2620];
  assign N7665 = N7664 | data_masked[2748];
  assign N7664 = N7663 | data_masked[2876];
  assign N7663 = N7662 | data_masked[3004];
  assign N7662 = N7661 | data_masked[3132];
  assign N7661 = N7660 | data_masked[3260];
  assign N7660 = N7659 | data_masked[3388];
  assign N7659 = N7658 | data_masked[3516];
  assign N7658 = N7657 | data_masked[3644];
  assign N7657 = N7656 | data_masked[3772];
  assign N7656 = N7655 | data_masked[3900];
  assign N7655 = N7654 | data_masked[4028];
  assign N7654 = N7653 | data_masked[4156];
  assign N7653 = N7652 | data_masked[4284];
  assign N7652 = N7651 | data_masked[4412];
  assign N7651 = N7650 | data_masked[4540];
  assign N7650 = N7649 | data_masked[4668];
  assign N7649 = N7648 | data_masked[4796];
  assign N7648 = N7647 | data_masked[4924];
  assign N7647 = N7646 | data_masked[5052];
  assign N7646 = N7645 | data_masked[5180];
  assign N7645 = N7644 | data_masked[5308];
  assign N7644 = N7643 | data_masked[5436];
  assign N7643 = N7642 | data_masked[5564];
  assign N7642 = N7641 | data_masked[5692];
  assign N7641 = N7640 | data_masked[5820];
  assign N7640 = N7639 | data_masked[5948];
  assign N7639 = N7638 | data_masked[6076];
  assign N7638 = N7637 | data_masked[6204];
  assign N7637 = N7636 | data_masked[6332];
  assign N7636 = N7635 | data_masked[6460];
  assign N7635 = N7634 | data_masked[6588];
  assign N7634 = N7633 | data_masked[6716];
  assign N7633 = N7632 | data_masked[6844];
  assign N7632 = N7631 | data_masked[6972];
  assign N7631 = N7630 | data_masked[7100];
  assign N7630 = N7629 | data_masked[7228];
  assign N7629 = N7628 | data_masked[7356];
  assign N7628 = N7627 | data_masked[7484];
  assign N7627 = N7626 | data_masked[7612];
  assign N7626 = N7625 | data_masked[7740];
  assign N7625 = N7624 | data_masked[7868];
  assign N7624 = N7623 | data_masked[7996];
  assign N7623 = N7622 | data_masked[8124];
  assign N7622 = N7621 | data_masked[8252];
  assign N7621 = N7620 | data_masked[8380];
  assign N7620 = N7619 | data_masked[8508];
  assign N7619 = N7618 | data_masked[8636];
  assign N7618 = N7617 | data_masked[8764];
  assign N7617 = N7616 | data_masked[8892];
  assign N7616 = N7615 | data_masked[9020];
  assign N7615 = N7614 | data_masked[9148];
  assign N7614 = N7613 | data_masked[9276];
  assign N7613 = N7612 | data_masked[9404];
  assign N7612 = N7611 | data_masked[9532];
  assign N7611 = N7610 | data_masked[9660];
  assign N7610 = N7609 | data_masked[9788];
  assign N7609 = N7608 | data_masked[9916];
  assign N7608 = N7607 | data_masked[10044];
  assign N7607 = N7606 | data_masked[10172];
  assign N7606 = N7605 | data_masked[10300];
  assign N7605 = N7604 | data_masked[10428];
  assign N7604 = N7603 | data_masked[10556];
  assign N7603 = N7602 | data_masked[10684];
  assign N7602 = N7601 | data_masked[10812];
  assign N7601 = N7600 | data_masked[10940];
  assign N7600 = N7599 | data_masked[11068];
  assign N7599 = N7598 | data_masked[11196];
  assign N7598 = N7597 | data_masked[11324];
  assign N7597 = N7596 | data_masked[11452];
  assign N7596 = N7595 | data_masked[11580];
  assign N7595 = N7594 | data_masked[11708];
  assign N7594 = N7593 | data_masked[11836];
  assign N7593 = N7592 | data_masked[11964];
  assign N7592 = N7591 | data_masked[12092];
  assign N7591 = N7590 | data_masked[12220];
  assign N7590 = N7589 | data_masked[12348];
  assign N7589 = N7588 | data_masked[12476];
  assign N7588 = N7587 | data_masked[12604];
  assign N7587 = N7586 | data_masked[12732];
  assign N7586 = N7585 | data_masked[12860];
  assign N7585 = N7584 | data_masked[12988];
  assign N7584 = N7583 | data_masked[13116];
  assign N7583 = N7582 | data_masked[13244];
  assign N7582 = N7581 | data_masked[13372];
  assign N7581 = N7580 | data_masked[13500];
  assign N7580 = N7579 | data_masked[13628];
  assign N7579 = N7578 | data_masked[13756];
  assign N7578 = N7577 | data_masked[13884];
  assign N7577 = N7576 | data_masked[14012];
  assign N7576 = N7575 | data_masked[14140];
  assign N7575 = N7574 | data_masked[14268];
  assign N7574 = N7573 | data_masked[14396];
  assign N7573 = N7572 | data_masked[14524];
  assign N7572 = N7571 | data_masked[14652];
  assign N7571 = N7570 | data_masked[14780];
  assign N7570 = N7569 | data_masked[14908];
  assign N7569 = N7568 | data_masked[15036];
  assign N7568 = N7567 | data_masked[15164];
  assign N7567 = N7566 | data_masked[15292];
  assign N7566 = N7565 | data_masked[15420];
  assign N7565 = N7564 | data_masked[15548];
  assign N7564 = N7563 | data_masked[15676];
  assign N7563 = N7562 | data_masked[15804];
  assign N7562 = N7561 | data_masked[15932];
  assign N7561 = N7560 | data_masked[16060];
  assign N7560 = data_masked[16316] | data_masked[16188];
  assign data_o[61] = N7811 | data_masked[61];
  assign N7811 = N7810 | data_masked[189];
  assign N7810 = N7809 | data_masked[317];
  assign N7809 = N7808 | data_masked[445];
  assign N7808 = N7807 | data_masked[573];
  assign N7807 = N7806 | data_masked[701];
  assign N7806 = N7805 | data_masked[829];
  assign N7805 = N7804 | data_masked[957];
  assign N7804 = N7803 | data_masked[1085];
  assign N7803 = N7802 | data_masked[1213];
  assign N7802 = N7801 | data_masked[1341];
  assign N7801 = N7800 | data_masked[1469];
  assign N7800 = N7799 | data_masked[1597];
  assign N7799 = N7798 | data_masked[1725];
  assign N7798 = N7797 | data_masked[1853];
  assign N7797 = N7796 | data_masked[1981];
  assign N7796 = N7795 | data_masked[2109];
  assign N7795 = N7794 | data_masked[2237];
  assign N7794 = N7793 | data_masked[2365];
  assign N7793 = N7792 | data_masked[2493];
  assign N7792 = N7791 | data_masked[2621];
  assign N7791 = N7790 | data_masked[2749];
  assign N7790 = N7789 | data_masked[2877];
  assign N7789 = N7788 | data_masked[3005];
  assign N7788 = N7787 | data_masked[3133];
  assign N7787 = N7786 | data_masked[3261];
  assign N7786 = N7785 | data_masked[3389];
  assign N7785 = N7784 | data_masked[3517];
  assign N7784 = N7783 | data_masked[3645];
  assign N7783 = N7782 | data_masked[3773];
  assign N7782 = N7781 | data_masked[3901];
  assign N7781 = N7780 | data_masked[4029];
  assign N7780 = N7779 | data_masked[4157];
  assign N7779 = N7778 | data_masked[4285];
  assign N7778 = N7777 | data_masked[4413];
  assign N7777 = N7776 | data_masked[4541];
  assign N7776 = N7775 | data_masked[4669];
  assign N7775 = N7774 | data_masked[4797];
  assign N7774 = N7773 | data_masked[4925];
  assign N7773 = N7772 | data_masked[5053];
  assign N7772 = N7771 | data_masked[5181];
  assign N7771 = N7770 | data_masked[5309];
  assign N7770 = N7769 | data_masked[5437];
  assign N7769 = N7768 | data_masked[5565];
  assign N7768 = N7767 | data_masked[5693];
  assign N7767 = N7766 | data_masked[5821];
  assign N7766 = N7765 | data_masked[5949];
  assign N7765 = N7764 | data_masked[6077];
  assign N7764 = N7763 | data_masked[6205];
  assign N7763 = N7762 | data_masked[6333];
  assign N7762 = N7761 | data_masked[6461];
  assign N7761 = N7760 | data_masked[6589];
  assign N7760 = N7759 | data_masked[6717];
  assign N7759 = N7758 | data_masked[6845];
  assign N7758 = N7757 | data_masked[6973];
  assign N7757 = N7756 | data_masked[7101];
  assign N7756 = N7755 | data_masked[7229];
  assign N7755 = N7754 | data_masked[7357];
  assign N7754 = N7753 | data_masked[7485];
  assign N7753 = N7752 | data_masked[7613];
  assign N7752 = N7751 | data_masked[7741];
  assign N7751 = N7750 | data_masked[7869];
  assign N7750 = N7749 | data_masked[7997];
  assign N7749 = N7748 | data_masked[8125];
  assign N7748 = N7747 | data_masked[8253];
  assign N7747 = N7746 | data_masked[8381];
  assign N7746 = N7745 | data_masked[8509];
  assign N7745 = N7744 | data_masked[8637];
  assign N7744 = N7743 | data_masked[8765];
  assign N7743 = N7742 | data_masked[8893];
  assign N7742 = N7741 | data_masked[9021];
  assign N7741 = N7740 | data_masked[9149];
  assign N7740 = N7739 | data_masked[9277];
  assign N7739 = N7738 | data_masked[9405];
  assign N7738 = N7737 | data_masked[9533];
  assign N7737 = N7736 | data_masked[9661];
  assign N7736 = N7735 | data_masked[9789];
  assign N7735 = N7734 | data_masked[9917];
  assign N7734 = N7733 | data_masked[10045];
  assign N7733 = N7732 | data_masked[10173];
  assign N7732 = N7731 | data_masked[10301];
  assign N7731 = N7730 | data_masked[10429];
  assign N7730 = N7729 | data_masked[10557];
  assign N7729 = N7728 | data_masked[10685];
  assign N7728 = N7727 | data_masked[10813];
  assign N7727 = N7726 | data_masked[10941];
  assign N7726 = N7725 | data_masked[11069];
  assign N7725 = N7724 | data_masked[11197];
  assign N7724 = N7723 | data_masked[11325];
  assign N7723 = N7722 | data_masked[11453];
  assign N7722 = N7721 | data_masked[11581];
  assign N7721 = N7720 | data_masked[11709];
  assign N7720 = N7719 | data_masked[11837];
  assign N7719 = N7718 | data_masked[11965];
  assign N7718 = N7717 | data_masked[12093];
  assign N7717 = N7716 | data_masked[12221];
  assign N7716 = N7715 | data_masked[12349];
  assign N7715 = N7714 | data_masked[12477];
  assign N7714 = N7713 | data_masked[12605];
  assign N7713 = N7712 | data_masked[12733];
  assign N7712 = N7711 | data_masked[12861];
  assign N7711 = N7710 | data_masked[12989];
  assign N7710 = N7709 | data_masked[13117];
  assign N7709 = N7708 | data_masked[13245];
  assign N7708 = N7707 | data_masked[13373];
  assign N7707 = N7706 | data_masked[13501];
  assign N7706 = N7705 | data_masked[13629];
  assign N7705 = N7704 | data_masked[13757];
  assign N7704 = N7703 | data_masked[13885];
  assign N7703 = N7702 | data_masked[14013];
  assign N7702 = N7701 | data_masked[14141];
  assign N7701 = N7700 | data_masked[14269];
  assign N7700 = N7699 | data_masked[14397];
  assign N7699 = N7698 | data_masked[14525];
  assign N7698 = N7697 | data_masked[14653];
  assign N7697 = N7696 | data_masked[14781];
  assign N7696 = N7695 | data_masked[14909];
  assign N7695 = N7694 | data_masked[15037];
  assign N7694 = N7693 | data_masked[15165];
  assign N7693 = N7692 | data_masked[15293];
  assign N7692 = N7691 | data_masked[15421];
  assign N7691 = N7690 | data_masked[15549];
  assign N7690 = N7689 | data_masked[15677];
  assign N7689 = N7688 | data_masked[15805];
  assign N7688 = N7687 | data_masked[15933];
  assign N7687 = N7686 | data_masked[16061];
  assign N7686 = data_masked[16317] | data_masked[16189];
  assign data_o[62] = N7937 | data_masked[62];
  assign N7937 = N7936 | data_masked[190];
  assign N7936 = N7935 | data_masked[318];
  assign N7935 = N7934 | data_masked[446];
  assign N7934 = N7933 | data_masked[574];
  assign N7933 = N7932 | data_masked[702];
  assign N7932 = N7931 | data_masked[830];
  assign N7931 = N7930 | data_masked[958];
  assign N7930 = N7929 | data_masked[1086];
  assign N7929 = N7928 | data_masked[1214];
  assign N7928 = N7927 | data_masked[1342];
  assign N7927 = N7926 | data_masked[1470];
  assign N7926 = N7925 | data_masked[1598];
  assign N7925 = N7924 | data_masked[1726];
  assign N7924 = N7923 | data_masked[1854];
  assign N7923 = N7922 | data_masked[1982];
  assign N7922 = N7921 | data_masked[2110];
  assign N7921 = N7920 | data_masked[2238];
  assign N7920 = N7919 | data_masked[2366];
  assign N7919 = N7918 | data_masked[2494];
  assign N7918 = N7917 | data_masked[2622];
  assign N7917 = N7916 | data_masked[2750];
  assign N7916 = N7915 | data_masked[2878];
  assign N7915 = N7914 | data_masked[3006];
  assign N7914 = N7913 | data_masked[3134];
  assign N7913 = N7912 | data_masked[3262];
  assign N7912 = N7911 | data_masked[3390];
  assign N7911 = N7910 | data_masked[3518];
  assign N7910 = N7909 | data_masked[3646];
  assign N7909 = N7908 | data_masked[3774];
  assign N7908 = N7907 | data_masked[3902];
  assign N7907 = N7906 | data_masked[4030];
  assign N7906 = N7905 | data_masked[4158];
  assign N7905 = N7904 | data_masked[4286];
  assign N7904 = N7903 | data_masked[4414];
  assign N7903 = N7902 | data_masked[4542];
  assign N7902 = N7901 | data_masked[4670];
  assign N7901 = N7900 | data_masked[4798];
  assign N7900 = N7899 | data_masked[4926];
  assign N7899 = N7898 | data_masked[5054];
  assign N7898 = N7897 | data_masked[5182];
  assign N7897 = N7896 | data_masked[5310];
  assign N7896 = N7895 | data_masked[5438];
  assign N7895 = N7894 | data_masked[5566];
  assign N7894 = N7893 | data_masked[5694];
  assign N7893 = N7892 | data_masked[5822];
  assign N7892 = N7891 | data_masked[5950];
  assign N7891 = N7890 | data_masked[6078];
  assign N7890 = N7889 | data_masked[6206];
  assign N7889 = N7888 | data_masked[6334];
  assign N7888 = N7887 | data_masked[6462];
  assign N7887 = N7886 | data_masked[6590];
  assign N7886 = N7885 | data_masked[6718];
  assign N7885 = N7884 | data_masked[6846];
  assign N7884 = N7883 | data_masked[6974];
  assign N7883 = N7882 | data_masked[7102];
  assign N7882 = N7881 | data_masked[7230];
  assign N7881 = N7880 | data_masked[7358];
  assign N7880 = N7879 | data_masked[7486];
  assign N7879 = N7878 | data_masked[7614];
  assign N7878 = N7877 | data_masked[7742];
  assign N7877 = N7876 | data_masked[7870];
  assign N7876 = N7875 | data_masked[7998];
  assign N7875 = N7874 | data_masked[8126];
  assign N7874 = N7873 | data_masked[8254];
  assign N7873 = N7872 | data_masked[8382];
  assign N7872 = N7871 | data_masked[8510];
  assign N7871 = N7870 | data_masked[8638];
  assign N7870 = N7869 | data_masked[8766];
  assign N7869 = N7868 | data_masked[8894];
  assign N7868 = N7867 | data_masked[9022];
  assign N7867 = N7866 | data_masked[9150];
  assign N7866 = N7865 | data_masked[9278];
  assign N7865 = N7864 | data_masked[9406];
  assign N7864 = N7863 | data_masked[9534];
  assign N7863 = N7862 | data_masked[9662];
  assign N7862 = N7861 | data_masked[9790];
  assign N7861 = N7860 | data_masked[9918];
  assign N7860 = N7859 | data_masked[10046];
  assign N7859 = N7858 | data_masked[10174];
  assign N7858 = N7857 | data_masked[10302];
  assign N7857 = N7856 | data_masked[10430];
  assign N7856 = N7855 | data_masked[10558];
  assign N7855 = N7854 | data_masked[10686];
  assign N7854 = N7853 | data_masked[10814];
  assign N7853 = N7852 | data_masked[10942];
  assign N7852 = N7851 | data_masked[11070];
  assign N7851 = N7850 | data_masked[11198];
  assign N7850 = N7849 | data_masked[11326];
  assign N7849 = N7848 | data_masked[11454];
  assign N7848 = N7847 | data_masked[11582];
  assign N7847 = N7846 | data_masked[11710];
  assign N7846 = N7845 | data_masked[11838];
  assign N7845 = N7844 | data_masked[11966];
  assign N7844 = N7843 | data_masked[12094];
  assign N7843 = N7842 | data_masked[12222];
  assign N7842 = N7841 | data_masked[12350];
  assign N7841 = N7840 | data_masked[12478];
  assign N7840 = N7839 | data_masked[12606];
  assign N7839 = N7838 | data_masked[12734];
  assign N7838 = N7837 | data_masked[12862];
  assign N7837 = N7836 | data_masked[12990];
  assign N7836 = N7835 | data_masked[13118];
  assign N7835 = N7834 | data_masked[13246];
  assign N7834 = N7833 | data_masked[13374];
  assign N7833 = N7832 | data_masked[13502];
  assign N7832 = N7831 | data_masked[13630];
  assign N7831 = N7830 | data_masked[13758];
  assign N7830 = N7829 | data_masked[13886];
  assign N7829 = N7828 | data_masked[14014];
  assign N7828 = N7827 | data_masked[14142];
  assign N7827 = N7826 | data_masked[14270];
  assign N7826 = N7825 | data_masked[14398];
  assign N7825 = N7824 | data_masked[14526];
  assign N7824 = N7823 | data_masked[14654];
  assign N7823 = N7822 | data_masked[14782];
  assign N7822 = N7821 | data_masked[14910];
  assign N7821 = N7820 | data_masked[15038];
  assign N7820 = N7819 | data_masked[15166];
  assign N7819 = N7818 | data_masked[15294];
  assign N7818 = N7817 | data_masked[15422];
  assign N7817 = N7816 | data_masked[15550];
  assign N7816 = N7815 | data_masked[15678];
  assign N7815 = N7814 | data_masked[15806];
  assign N7814 = N7813 | data_masked[15934];
  assign N7813 = N7812 | data_masked[16062];
  assign N7812 = data_masked[16318] | data_masked[16190];
  assign data_o[63] = N8063 | data_masked[63];
  assign N8063 = N8062 | data_masked[191];
  assign N8062 = N8061 | data_masked[319];
  assign N8061 = N8060 | data_masked[447];
  assign N8060 = N8059 | data_masked[575];
  assign N8059 = N8058 | data_masked[703];
  assign N8058 = N8057 | data_masked[831];
  assign N8057 = N8056 | data_masked[959];
  assign N8056 = N8055 | data_masked[1087];
  assign N8055 = N8054 | data_masked[1215];
  assign N8054 = N8053 | data_masked[1343];
  assign N8053 = N8052 | data_masked[1471];
  assign N8052 = N8051 | data_masked[1599];
  assign N8051 = N8050 | data_masked[1727];
  assign N8050 = N8049 | data_masked[1855];
  assign N8049 = N8048 | data_masked[1983];
  assign N8048 = N8047 | data_masked[2111];
  assign N8047 = N8046 | data_masked[2239];
  assign N8046 = N8045 | data_masked[2367];
  assign N8045 = N8044 | data_masked[2495];
  assign N8044 = N8043 | data_masked[2623];
  assign N8043 = N8042 | data_masked[2751];
  assign N8042 = N8041 | data_masked[2879];
  assign N8041 = N8040 | data_masked[3007];
  assign N8040 = N8039 | data_masked[3135];
  assign N8039 = N8038 | data_masked[3263];
  assign N8038 = N8037 | data_masked[3391];
  assign N8037 = N8036 | data_masked[3519];
  assign N8036 = N8035 | data_masked[3647];
  assign N8035 = N8034 | data_masked[3775];
  assign N8034 = N8033 | data_masked[3903];
  assign N8033 = N8032 | data_masked[4031];
  assign N8032 = N8031 | data_masked[4159];
  assign N8031 = N8030 | data_masked[4287];
  assign N8030 = N8029 | data_masked[4415];
  assign N8029 = N8028 | data_masked[4543];
  assign N8028 = N8027 | data_masked[4671];
  assign N8027 = N8026 | data_masked[4799];
  assign N8026 = N8025 | data_masked[4927];
  assign N8025 = N8024 | data_masked[5055];
  assign N8024 = N8023 | data_masked[5183];
  assign N8023 = N8022 | data_masked[5311];
  assign N8022 = N8021 | data_masked[5439];
  assign N8021 = N8020 | data_masked[5567];
  assign N8020 = N8019 | data_masked[5695];
  assign N8019 = N8018 | data_masked[5823];
  assign N8018 = N8017 | data_masked[5951];
  assign N8017 = N8016 | data_masked[6079];
  assign N8016 = N8015 | data_masked[6207];
  assign N8015 = N8014 | data_masked[6335];
  assign N8014 = N8013 | data_masked[6463];
  assign N8013 = N8012 | data_masked[6591];
  assign N8012 = N8011 | data_masked[6719];
  assign N8011 = N8010 | data_masked[6847];
  assign N8010 = N8009 | data_masked[6975];
  assign N8009 = N8008 | data_masked[7103];
  assign N8008 = N8007 | data_masked[7231];
  assign N8007 = N8006 | data_masked[7359];
  assign N8006 = N8005 | data_masked[7487];
  assign N8005 = N8004 | data_masked[7615];
  assign N8004 = N8003 | data_masked[7743];
  assign N8003 = N8002 | data_masked[7871];
  assign N8002 = N8001 | data_masked[7999];
  assign N8001 = N8000 | data_masked[8127];
  assign N8000 = N7999 | data_masked[8255];
  assign N7999 = N7998 | data_masked[8383];
  assign N7998 = N7997 | data_masked[8511];
  assign N7997 = N7996 | data_masked[8639];
  assign N7996 = N7995 | data_masked[8767];
  assign N7995 = N7994 | data_masked[8895];
  assign N7994 = N7993 | data_masked[9023];
  assign N7993 = N7992 | data_masked[9151];
  assign N7992 = N7991 | data_masked[9279];
  assign N7991 = N7990 | data_masked[9407];
  assign N7990 = N7989 | data_masked[9535];
  assign N7989 = N7988 | data_masked[9663];
  assign N7988 = N7987 | data_masked[9791];
  assign N7987 = N7986 | data_masked[9919];
  assign N7986 = N7985 | data_masked[10047];
  assign N7985 = N7984 | data_masked[10175];
  assign N7984 = N7983 | data_masked[10303];
  assign N7983 = N7982 | data_masked[10431];
  assign N7982 = N7981 | data_masked[10559];
  assign N7981 = N7980 | data_masked[10687];
  assign N7980 = N7979 | data_masked[10815];
  assign N7979 = N7978 | data_masked[10943];
  assign N7978 = N7977 | data_masked[11071];
  assign N7977 = N7976 | data_masked[11199];
  assign N7976 = N7975 | data_masked[11327];
  assign N7975 = N7974 | data_masked[11455];
  assign N7974 = N7973 | data_masked[11583];
  assign N7973 = N7972 | data_masked[11711];
  assign N7972 = N7971 | data_masked[11839];
  assign N7971 = N7970 | data_masked[11967];
  assign N7970 = N7969 | data_masked[12095];
  assign N7969 = N7968 | data_masked[12223];
  assign N7968 = N7967 | data_masked[12351];
  assign N7967 = N7966 | data_masked[12479];
  assign N7966 = N7965 | data_masked[12607];
  assign N7965 = N7964 | data_masked[12735];
  assign N7964 = N7963 | data_masked[12863];
  assign N7963 = N7962 | data_masked[12991];
  assign N7962 = N7961 | data_masked[13119];
  assign N7961 = N7960 | data_masked[13247];
  assign N7960 = N7959 | data_masked[13375];
  assign N7959 = N7958 | data_masked[13503];
  assign N7958 = N7957 | data_masked[13631];
  assign N7957 = N7956 | data_masked[13759];
  assign N7956 = N7955 | data_masked[13887];
  assign N7955 = N7954 | data_masked[14015];
  assign N7954 = N7953 | data_masked[14143];
  assign N7953 = N7952 | data_masked[14271];
  assign N7952 = N7951 | data_masked[14399];
  assign N7951 = N7950 | data_masked[14527];
  assign N7950 = N7949 | data_masked[14655];
  assign N7949 = N7948 | data_masked[14783];
  assign N7948 = N7947 | data_masked[14911];
  assign N7947 = N7946 | data_masked[15039];
  assign N7946 = N7945 | data_masked[15167];
  assign N7945 = N7944 | data_masked[15295];
  assign N7944 = N7943 | data_masked[15423];
  assign N7943 = N7942 | data_masked[15551];
  assign N7942 = N7941 | data_masked[15679];
  assign N7941 = N7940 | data_masked[15807];
  assign N7940 = N7939 | data_masked[15935];
  assign N7939 = N7938 | data_masked[16063];
  assign N7938 = data_masked[16319] | data_masked[16191];
  assign data_o[64] = N8189 | data_masked[64];
  assign N8189 = N8188 | data_masked[192];
  assign N8188 = N8187 | data_masked[320];
  assign N8187 = N8186 | data_masked[448];
  assign N8186 = N8185 | data_masked[576];
  assign N8185 = N8184 | data_masked[704];
  assign N8184 = N8183 | data_masked[832];
  assign N8183 = N8182 | data_masked[960];
  assign N8182 = N8181 | data_masked[1088];
  assign N8181 = N8180 | data_masked[1216];
  assign N8180 = N8179 | data_masked[1344];
  assign N8179 = N8178 | data_masked[1472];
  assign N8178 = N8177 | data_masked[1600];
  assign N8177 = N8176 | data_masked[1728];
  assign N8176 = N8175 | data_masked[1856];
  assign N8175 = N8174 | data_masked[1984];
  assign N8174 = N8173 | data_masked[2112];
  assign N8173 = N8172 | data_masked[2240];
  assign N8172 = N8171 | data_masked[2368];
  assign N8171 = N8170 | data_masked[2496];
  assign N8170 = N8169 | data_masked[2624];
  assign N8169 = N8168 | data_masked[2752];
  assign N8168 = N8167 | data_masked[2880];
  assign N8167 = N8166 | data_masked[3008];
  assign N8166 = N8165 | data_masked[3136];
  assign N8165 = N8164 | data_masked[3264];
  assign N8164 = N8163 | data_masked[3392];
  assign N8163 = N8162 | data_masked[3520];
  assign N8162 = N8161 | data_masked[3648];
  assign N8161 = N8160 | data_masked[3776];
  assign N8160 = N8159 | data_masked[3904];
  assign N8159 = N8158 | data_masked[4032];
  assign N8158 = N8157 | data_masked[4160];
  assign N8157 = N8156 | data_masked[4288];
  assign N8156 = N8155 | data_masked[4416];
  assign N8155 = N8154 | data_masked[4544];
  assign N8154 = N8153 | data_masked[4672];
  assign N8153 = N8152 | data_masked[4800];
  assign N8152 = N8151 | data_masked[4928];
  assign N8151 = N8150 | data_masked[5056];
  assign N8150 = N8149 | data_masked[5184];
  assign N8149 = N8148 | data_masked[5312];
  assign N8148 = N8147 | data_masked[5440];
  assign N8147 = N8146 | data_masked[5568];
  assign N8146 = N8145 | data_masked[5696];
  assign N8145 = N8144 | data_masked[5824];
  assign N8144 = N8143 | data_masked[5952];
  assign N8143 = N8142 | data_masked[6080];
  assign N8142 = N8141 | data_masked[6208];
  assign N8141 = N8140 | data_masked[6336];
  assign N8140 = N8139 | data_masked[6464];
  assign N8139 = N8138 | data_masked[6592];
  assign N8138 = N8137 | data_masked[6720];
  assign N8137 = N8136 | data_masked[6848];
  assign N8136 = N8135 | data_masked[6976];
  assign N8135 = N8134 | data_masked[7104];
  assign N8134 = N8133 | data_masked[7232];
  assign N8133 = N8132 | data_masked[7360];
  assign N8132 = N8131 | data_masked[7488];
  assign N8131 = N8130 | data_masked[7616];
  assign N8130 = N8129 | data_masked[7744];
  assign N8129 = N8128 | data_masked[7872];
  assign N8128 = N8127 | data_masked[8000];
  assign N8127 = N8126 | data_masked[8128];
  assign N8126 = N8125 | data_masked[8256];
  assign N8125 = N8124 | data_masked[8384];
  assign N8124 = N8123 | data_masked[8512];
  assign N8123 = N8122 | data_masked[8640];
  assign N8122 = N8121 | data_masked[8768];
  assign N8121 = N8120 | data_masked[8896];
  assign N8120 = N8119 | data_masked[9024];
  assign N8119 = N8118 | data_masked[9152];
  assign N8118 = N8117 | data_masked[9280];
  assign N8117 = N8116 | data_masked[9408];
  assign N8116 = N8115 | data_masked[9536];
  assign N8115 = N8114 | data_masked[9664];
  assign N8114 = N8113 | data_masked[9792];
  assign N8113 = N8112 | data_masked[9920];
  assign N8112 = N8111 | data_masked[10048];
  assign N8111 = N8110 | data_masked[10176];
  assign N8110 = N8109 | data_masked[10304];
  assign N8109 = N8108 | data_masked[10432];
  assign N8108 = N8107 | data_masked[10560];
  assign N8107 = N8106 | data_masked[10688];
  assign N8106 = N8105 | data_masked[10816];
  assign N8105 = N8104 | data_masked[10944];
  assign N8104 = N8103 | data_masked[11072];
  assign N8103 = N8102 | data_masked[11200];
  assign N8102 = N8101 | data_masked[11328];
  assign N8101 = N8100 | data_masked[11456];
  assign N8100 = N8099 | data_masked[11584];
  assign N8099 = N8098 | data_masked[11712];
  assign N8098 = N8097 | data_masked[11840];
  assign N8097 = N8096 | data_masked[11968];
  assign N8096 = N8095 | data_masked[12096];
  assign N8095 = N8094 | data_masked[12224];
  assign N8094 = N8093 | data_masked[12352];
  assign N8093 = N8092 | data_masked[12480];
  assign N8092 = N8091 | data_masked[12608];
  assign N8091 = N8090 | data_masked[12736];
  assign N8090 = N8089 | data_masked[12864];
  assign N8089 = N8088 | data_masked[12992];
  assign N8088 = N8087 | data_masked[13120];
  assign N8087 = N8086 | data_masked[13248];
  assign N8086 = N8085 | data_masked[13376];
  assign N8085 = N8084 | data_masked[13504];
  assign N8084 = N8083 | data_masked[13632];
  assign N8083 = N8082 | data_masked[13760];
  assign N8082 = N8081 | data_masked[13888];
  assign N8081 = N8080 | data_masked[14016];
  assign N8080 = N8079 | data_masked[14144];
  assign N8079 = N8078 | data_masked[14272];
  assign N8078 = N8077 | data_masked[14400];
  assign N8077 = N8076 | data_masked[14528];
  assign N8076 = N8075 | data_masked[14656];
  assign N8075 = N8074 | data_masked[14784];
  assign N8074 = N8073 | data_masked[14912];
  assign N8073 = N8072 | data_masked[15040];
  assign N8072 = N8071 | data_masked[15168];
  assign N8071 = N8070 | data_masked[15296];
  assign N8070 = N8069 | data_masked[15424];
  assign N8069 = N8068 | data_masked[15552];
  assign N8068 = N8067 | data_masked[15680];
  assign N8067 = N8066 | data_masked[15808];
  assign N8066 = N8065 | data_masked[15936];
  assign N8065 = N8064 | data_masked[16064];
  assign N8064 = data_masked[16320] | data_masked[16192];
  assign data_o[65] = N8315 | data_masked[65];
  assign N8315 = N8314 | data_masked[193];
  assign N8314 = N8313 | data_masked[321];
  assign N8313 = N8312 | data_masked[449];
  assign N8312 = N8311 | data_masked[577];
  assign N8311 = N8310 | data_masked[705];
  assign N8310 = N8309 | data_masked[833];
  assign N8309 = N8308 | data_masked[961];
  assign N8308 = N8307 | data_masked[1089];
  assign N8307 = N8306 | data_masked[1217];
  assign N8306 = N8305 | data_masked[1345];
  assign N8305 = N8304 | data_masked[1473];
  assign N8304 = N8303 | data_masked[1601];
  assign N8303 = N8302 | data_masked[1729];
  assign N8302 = N8301 | data_masked[1857];
  assign N8301 = N8300 | data_masked[1985];
  assign N8300 = N8299 | data_masked[2113];
  assign N8299 = N8298 | data_masked[2241];
  assign N8298 = N8297 | data_masked[2369];
  assign N8297 = N8296 | data_masked[2497];
  assign N8296 = N8295 | data_masked[2625];
  assign N8295 = N8294 | data_masked[2753];
  assign N8294 = N8293 | data_masked[2881];
  assign N8293 = N8292 | data_masked[3009];
  assign N8292 = N8291 | data_masked[3137];
  assign N8291 = N8290 | data_masked[3265];
  assign N8290 = N8289 | data_masked[3393];
  assign N8289 = N8288 | data_masked[3521];
  assign N8288 = N8287 | data_masked[3649];
  assign N8287 = N8286 | data_masked[3777];
  assign N8286 = N8285 | data_masked[3905];
  assign N8285 = N8284 | data_masked[4033];
  assign N8284 = N8283 | data_masked[4161];
  assign N8283 = N8282 | data_masked[4289];
  assign N8282 = N8281 | data_masked[4417];
  assign N8281 = N8280 | data_masked[4545];
  assign N8280 = N8279 | data_masked[4673];
  assign N8279 = N8278 | data_masked[4801];
  assign N8278 = N8277 | data_masked[4929];
  assign N8277 = N8276 | data_masked[5057];
  assign N8276 = N8275 | data_masked[5185];
  assign N8275 = N8274 | data_masked[5313];
  assign N8274 = N8273 | data_masked[5441];
  assign N8273 = N8272 | data_masked[5569];
  assign N8272 = N8271 | data_masked[5697];
  assign N8271 = N8270 | data_masked[5825];
  assign N8270 = N8269 | data_masked[5953];
  assign N8269 = N8268 | data_masked[6081];
  assign N8268 = N8267 | data_masked[6209];
  assign N8267 = N8266 | data_masked[6337];
  assign N8266 = N8265 | data_masked[6465];
  assign N8265 = N8264 | data_masked[6593];
  assign N8264 = N8263 | data_masked[6721];
  assign N8263 = N8262 | data_masked[6849];
  assign N8262 = N8261 | data_masked[6977];
  assign N8261 = N8260 | data_masked[7105];
  assign N8260 = N8259 | data_masked[7233];
  assign N8259 = N8258 | data_masked[7361];
  assign N8258 = N8257 | data_masked[7489];
  assign N8257 = N8256 | data_masked[7617];
  assign N8256 = N8255 | data_masked[7745];
  assign N8255 = N8254 | data_masked[7873];
  assign N8254 = N8253 | data_masked[8001];
  assign N8253 = N8252 | data_masked[8129];
  assign N8252 = N8251 | data_masked[8257];
  assign N8251 = N8250 | data_masked[8385];
  assign N8250 = N8249 | data_masked[8513];
  assign N8249 = N8248 | data_masked[8641];
  assign N8248 = N8247 | data_masked[8769];
  assign N8247 = N8246 | data_masked[8897];
  assign N8246 = N8245 | data_masked[9025];
  assign N8245 = N8244 | data_masked[9153];
  assign N8244 = N8243 | data_masked[9281];
  assign N8243 = N8242 | data_masked[9409];
  assign N8242 = N8241 | data_masked[9537];
  assign N8241 = N8240 | data_masked[9665];
  assign N8240 = N8239 | data_masked[9793];
  assign N8239 = N8238 | data_masked[9921];
  assign N8238 = N8237 | data_masked[10049];
  assign N8237 = N8236 | data_masked[10177];
  assign N8236 = N8235 | data_masked[10305];
  assign N8235 = N8234 | data_masked[10433];
  assign N8234 = N8233 | data_masked[10561];
  assign N8233 = N8232 | data_masked[10689];
  assign N8232 = N8231 | data_masked[10817];
  assign N8231 = N8230 | data_masked[10945];
  assign N8230 = N8229 | data_masked[11073];
  assign N8229 = N8228 | data_masked[11201];
  assign N8228 = N8227 | data_masked[11329];
  assign N8227 = N8226 | data_masked[11457];
  assign N8226 = N8225 | data_masked[11585];
  assign N8225 = N8224 | data_masked[11713];
  assign N8224 = N8223 | data_masked[11841];
  assign N8223 = N8222 | data_masked[11969];
  assign N8222 = N8221 | data_masked[12097];
  assign N8221 = N8220 | data_masked[12225];
  assign N8220 = N8219 | data_masked[12353];
  assign N8219 = N8218 | data_masked[12481];
  assign N8218 = N8217 | data_masked[12609];
  assign N8217 = N8216 | data_masked[12737];
  assign N8216 = N8215 | data_masked[12865];
  assign N8215 = N8214 | data_masked[12993];
  assign N8214 = N8213 | data_masked[13121];
  assign N8213 = N8212 | data_masked[13249];
  assign N8212 = N8211 | data_masked[13377];
  assign N8211 = N8210 | data_masked[13505];
  assign N8210 = N8209 | data_masked[13633];
  assign N8209 = N8208 | data_masked[13761];
  assign N8208 = N8207 | data_masked[13889];
  assign N8207 = N8206 | data_masked[14017];
  assign N8206 = N8205 | data_masked[14145];
  assign N8205 = N8204 | data_masked[14273];
  assign N8204 = N8203 | data_masked[14401];
  assign N8203 = N8202 | data_masked[14529];
  assign N8202 = N8201 | data_masked[14657];
  assign N8201 = N8200 | data_masked[14785];
  assign N8200 = N8199 | data_masked[14913];
  assign N8199 = N8198 | data_masked[15041];
  assign N8198 = N8197 | data_masked[15169];
  assign N8197 = N8196 | data_masked[15297];
  assign N8196 = N8195 | data_masked[15425];
  assign N8195 = N8194 | data_masked[15553];
  assign N8194 = N8193 | data_masked[15681];
  assign N8193 = N8192 | data_masked[15809];
  assign N8192 = N8191 | data_masked[15937];
  assign N8191 = N8190 | data_masked[16065];
  assign N8190 = data_masked[16321] | data_masked[16193];
  assign data_o[66] = N8441 | data_masked[66];
  assign N8441 = N8440 | data_masked[194];
  assign N8440 = N8439 | data_masked[322];
  assign N8439 = N8438 | data_masked[450];
  assign N8438 = N8437 | data_masked[578];
  assign N8437 = N8436 | data_masked[706];
  assign N8436 = N8435 | data_masked[834];
  assign N8435 = N8434 | data_masked[962];
  assign N8434 = N8433 | data_masked[1090];
  assign N8433 = N8432 | data_masked[1218];
  assign N8432 = N8431 | data_masked[1346];
  assign N8431 = N8430 | data_masked[1474];
  assign N8430 = N8429 | data_masked[1602];
  assign N8429 = N8428 | data_masked[1730];
  assign N8428 = N8427 | data_masked[1858];
  assign N8427 = N8426 | data_masked[1986];
  assign N8426 = N8425 | data_masked[2114];
  assign N8425 = N8424 | data_masked[2242];
  assign N8424 = N8423 | data_masked[2370];
  assign N8423 = N8422 | data_masked[2498];
  assign N8422 = N8421 | data_masked[2626];
  assign N8421 = N8420 | data_masked[2754];
  assign N8420 = N8419 | data_masked[2882];
  assign N8419 = N8418 | data_masked[3010];
  assign N8418 = N8417 | data_masked[3138];
  assign N8417 = N8416 | data_masked[3266];
  assign N8416 = N8415 | data_masked[3394];
  assign N8415 = N8414 | data_masked[3522];
  assign N8414 = N8413 | data_masked[3650];
  assign N8413 = N8412 | data_masked[3778];
  assign N8412 = N8411 | data_masked[3906];
  assign N8411 = N8410 | data_masked[4034];
  assign N8410 = N8409 | data_masked[4162];
  assign N8409 = N8408 | data_masked[4290];
  assign N8408 = N8407 | data_masked[4418];
  assign N8407 = N8406 | data_masked[4546];
  assign N8406 = N8405 | data_masked[4674];
  assign N8405 = N8404 | data_masked[4802];
  assign N8404 = N8403 | data_masked[4930];
  assign N8403 = N8402 | data_masked[5058];
  assign N8402 = N8401 | data_masked[5186];
  assign N8401 = N8400 | data_masked[5314];
  assign N8400 = N8399 | data_masked[5442];
  assign N8399 = N8398 | data_masked[5570];
  assign N8398 = N8397 | data_masked[5698];
  assign N8397 = N8396 | data_masked[5826];
  assign N8396 = N8395 | data_masked[5954];
  assign N8395 = N8394 | data_masked[6082];
  assign N8394 = N8393 | data_masked[6210];
  assign N8393 = N8392 | data_masked[6338];
  assign N8392 = N8391 | data_masked[6466];
  assign N8391 = N8390 | data_masked[6594];
  assign N8390 = N8389 | data_masked[6722];
  assign N8389 = N8388 | data_masked[6850];
  assign N8388 = N8387 | data_masked[6978];
  assign N8387 = N8386 | data_masked[7106];
  assign N8386 = N8385 | data_masked[7234];
  assign N8385 = N8384 | data_masked[7362];
  assign N8384 = N8383 | data_masked[7490];
  assign N8383 = N8382 | data_masked[7618];
  assign N8382 = N8381 | data_masked[7746];
  assign N8381 = N8380 | data_masked[7874];
  assign N8380 = N8379 | data_masked[8002];
  assign N8379 = N8378 | data_masked[8130];
  assign N8378 = N8377 | data_masked[8258];
  assign N8377 = N8376 | data_masked[8386];
  assign N8376 = N8375 | data_masked[8514];
  assign N8375 = N8374 | data_masked[8642];
  assign N8374 = N8373 | data_masked[8770];
  assign N8373 = N8372 | data_masked[8898];
  assign N8372 = N8371 | data_masked[9026];
  assign N8371 = N8370 | data_masked[9154];
  assign N8370 = N8369 | data_masked[9282];
  assign N8369 = N8368 | data_masked[9410];
  assign N8368 = N8367 | data_masked[9538];
  assign N8367 = N8366 | data_masked[9666];
  assign N8366 = N8365 | data_masked[9794];
  assign N8365 = N8364 | data_masked[9922];
  assign N8364 = N8363 | data_masked[10050];
  assign N8363 = N8362 | data_masked[10178];
  assign N8362 = N8361 | data_masked[10306];
  assign N8361 = N8360 | data_masked[10434];
  assign N8360 = N8359 | data_masked[10562];
  assign N8359 = N8358 | data_masked[10690];
  assign N8358 = N8357 | data_masked[10818];
  assign N8357 = N8356 | data_masked[10946];
  assign N8356 = N8355 | data_masked[11074];
  assign N8355 = N8354 | data_masked[11202];
  assign N8354 = N8353 | data_masked[11330];
  assign N8353 = N8352 | data_masked[11458];
  assign N8352 = N8351 | data_masked[11586];
  assign N8351 = N8350 | data_masked[11714];
  assign N8350 = N8349 | data_masked[11842];
  assign N8349 = N8348 | data_masked[11970];
  assign N8348 = N8347 | data_masked[12098];
  assign N8347 = N8346 | data_masked[12226];
  assign N8346 = N8345 | data_masked[12354];
  assign N8345 = N8344 | data_masked[12482];
  assign N8344 = N8343 | data_masked[12610];
  assign N8343 = N8342 | data_masked[12738];
  assign N8342 = N8341 | data_masked[12866];
  assign N8341 = N8340 | data_masked[12994];
  assign N8340 = N8339 | data_masked[13122];
  assign N8339 = N8338 | data_masked[13250];
  assign N8338 = N8337 | data_masked[13378];
  assign N8337 = N8336 | data_masked[13506];
  assign N8336 = N8335 | data_masked[13634];
  assign N8335 = N8334 | data_masked[13762];
  assign N8334 = N8333 | data_masked[13890];
  assign N8333 = N8332 | data_masked[14018];
  assign N8332 = N8331 | data_masked[14146];
  assign N8331 = N8330 | data_masked[14274];
  assign N8330 = N8329 | data_masked[14402];
  assign N8329 = N8328 | data_masked[14530];
  assign N8328 = N8327 | data_masked[14658];
  assign N8327 = N8326 | data_masked[14786];
  assign N8326 = N8325 | data_masked[14914];
  assign N8325 = N8324 | data_masked[15042];
  assign N8324 = N8323 | data_masked[15170];
  assign N8323 = N8322 | data_masked[15298];
  assign N8322 = N8321 | data_masked[15426];
  assign N8321 = N8320 | data_masked[15554];
  assign N8320 = N8319 | data_masked[15682];
  assign N8319 = N8318 | data_masked[15810];
  assign N8318 = N8317 | data_masked[15938];
  assign N8317 = N8316 | data_masked[16066];
  assign N8316 = data_masked[16322] | data_masked[16194];
  assign data_o[67] = N8567 | data_masked[67];
  assign N8567 = N8566 | data_masked[195];
  assign N8566 = N8565 | data_masked[323];
  assign N8565 = N8564 | data_masked[451];
  assign N8564 = N8563 | data_masked[579];
  assign N8563 = N8562 | data_masked[707];
  assign N8562 = N8561 | data_masked[835];
  assign N8561 = N8560 | data_masked[963];
  assign N8560 = N8559 | data_masked[1091];
  assign N8559 = N8558 | data_masked[1219];
  assign N8558 = N8557 | data_masked[1347];
  assign N8557 = N8556 | data_masked[1475];
  assign N8556 = N8555 | data_masked[1603];
  assign N8555 = N8554 | data_masked[1731];
  assign N8554 = N8553 | data_masked[1859];
  assign N8553 = N8552 | data_masked[1987];
  assign N8552 = N8551 | data_masked[2115];
  assign N8551 = N8550 | data_masked[2243];
  assign N8550 = N8549 | data_masked[2371];
  assign N8549 = N8548 | data_masked[2499];
  assign N8548 = N8547 | data_masked[2627];
  assign N8547 = N8546 | data_masked[2755];
  assign N8546 = N8545 | data_masked[2883];
  assign N8545 = N8544 | data_masked[3011];
  assign N8544 = N8543 | data_masked[3139];
  assign N8543 = N8542 | data_masked[3267];
  assign N8542 = N8541 | data_masked[3395];
  assign N8541 = N8540 | data_masked[3523];
  assign N8540 = N8539 | data_masked[3651];
  assign N8539 = N8538 | data_masked[3779];
  assign N8538 = N8537 | data_masked[3907];
  assign N8537 = N8536 | data_masked[4035];
  assign N8536 = N8535 | data_masked[4163];
  assign N8535 = N8534 | data_masked[4291];
  assign N8534 = N8533 | data_masked[4419];
  assign N8533 = N8532 | data_masked[4547];
  assign N8532 = N8531 | data_masked[4675];
  assign N8531 = N8530 | data_masked[4803];
  assign N8530 = N8529 | data_masked[4931];
  assign N8529 = N8528 | data_masked[5059];
  assign N8528 = N8527 | data_masked[5187];
  assign N8527 = N8526 | data_masked[5315];
  assign N8526 = N8525 | data_masked[5443];
  assign N8525 = N8524 | data_masked[5571];
  assign N8524 = N8523 | data_masked[5699];
  assign N8523 = N8522 | data_masked[5827];
  assign N8522 = N8521 | data_masked[5955];
  assign N8521 = N8520 | data_masked[6083];
  assign N8520 = N8519 | data_masked[6211];
  assign N8519 = N8518 | data_masked[6339];
  assign N8518 = N8517 | data_masked[6467];
  assign N8517 = N8516 | data_masked[6595];
  assign N8516 = N8515 | data_masked[6723];
  assign N8515 = N8514 | data_masked[6851];
  assign N8514 = N8513 | data_masked[6979];
  assign N8513 = N8512 | data_masked[7107];
  assign N8512 = N8511 | data_masked[7235];
  assign N8511 = N8510 | data_masked[7363];
  assign N8510 = N8509 | data_masked[7491];
  assign N8509 = N8508 | data_masked[7619];
  assign N8508 = N8507 | data_masked[7747];
  assign N8507 = N8506 | data_masked[7875];
  assign N8506 = N8505 | data_masked[8003];
  assign N8505 = N8504 | data_masked[8131];
  assign N8504 = N8503 | data_masked[8259];
  assign N8503 = N8502 | data_masked[8387];
  assign N8502 = N8501 | data_masked[8515];
  assign N8501 = N8500 | data_masked[8643];
  assign N8500 = N8499 | data_masked[8771];
  assign N8499 = N8498 | data_masked[8899];
  assign N8498 = N8497 | data_masked[9027];
  assign N8497 = N8496 | data_masked[9155];
  assign N8496 = N8495 | data_masked[9283];
  assign N8495 = N8494 | data_masked[9411];
  assign N8494 = N8493 | data_masked[9539];
  assign N8493 = N8492 | data_masked[9667];
  assign N8492 = N8491 | data_masked[9795];
  assign N8491 = N8490 | data_masked[9923];
  assign N8490 = N8489 | data_masked[10051];
  assign N8489 = N8488 | data_masked[10179];
  assign N8488 = N8487 | data_masked[10307];
  assign N8487 = N8486 | data_masked[10435];
  assign N8486 = N8485 | data_masked[10563];
  assign N8485 = N8484 | data_masked[10691];
  assign N8484 = N8483 | data_masked[10819];
  assign N8483 = N8482 | data_masked[10947];
  assign N8482 = N8481 | data_masked[11075];
  assign N8481 = N8480 | data_masked[11203];
  assign N8480 = N8479 | data_masked[11331];
  assign N8479 = N8478 | data_masked[11459];
  assign N8478 = N8477 | data_masked[11587];
  assign N8477 = N8476 | data_masked[11715];
  assign N8476 = N8475 | data_masked[11843];
  assign N8475 = N8474 | data_masked[11971];
  assign N8474 = N8473 | data_masked[12099];
  assign N8473 = N8472 | data_masked[12227];
  assign N8472 = N8471 | data_masked[12355];
  assign N8471 = N8470 | data_masked[12483];
  assign N8470 = N8469 | data_masked[12611];
  assign N8469 = N8468 | data_masked[12739];
  assign N8468 = N8467 | data_masked[12867];
  assign N8467 = N8466 | data_masked[12995];
  assign N8466 = N8465 | data_masked[13123];
  assign N8465 = N8464 | data_masked[13251];
  assign N8464 = N8463 | data_masked[13379];
  assign N8463 = N8462 | data_masked[13507];
  assign N8462 = N8461 | data_masked[13635];
  assign N8461 = N8460 | data_masked[13763];
  assign N8460 = N8459 | data_masked[13891];
  assign N8459 = N8458 | data_masked[14019];
  assign N8458 = N8457 | data_masked[14147];
  assign N8457 = N8456 | data_masked[14275];
  assign N8456 = N8455 | data_masked[14403];
  assign N8455 = N8454 | data_masked[14531];
  assign N8454 = N8453 | data_masked[14659];
  assign N8453 = N8452 | data_masked[14787];
  assign N8452 = N8451 | data_masked[14915];
  assign N8451 = N8450 | data_masked[15043];
  assign N8450 = N8449 | data_masked[15171];
  assign N8449 = N8448 | data_masked[15299];
  assign N8448 = N8447 | data_masked[15427];
  assign N8447 = N8446 | data_masked[15555];
  assign N8446 = N8445 | data_masked[15683];
  assign N8445 = N8444 | data_masked[15811];
  assign N8444 = N8443 | data_masked[15939];
  assign N8443 = N8442 | data_masked[16067];
  assign N8442 = data_masked[16323] | data_masked[16195];
  assign data_o[68] = N8693 | data_masked[68];
  assign N8693 = N8692 | data_masked[196];
  assign N8692 = N8691 | data_masked[324];
  assign N8691 = N8690 | data_masked[452];
  assign N8690 = N8689 | data_masked[580];
  assign N8689 = N8688 | data_masked[708];
  assign N8688 = N8687 | data_masked[836];
  assign N8687 = N8686 | data_masked[964];
  assign N8686 = N8685 | data_masked[1092];
  assign N8685 = N8684 | data_masked[1220];
  assign N8684 = N8683 | data_masked[1348];
  assign N8683 = N8682 | data_masked[1476];
  assign N8682 = N8681 | data_masked[1604];
  assign N8681 = N8680 | data_masked[1732];
  assign N8680 = N8679 | data_masked[1860];
  assign N8679 = N8678 | data_masked[1988];
  assign N8678 = N8677 | data_masked[2116];
  assign N8677 = N8676 | data_masked[2244];
  assign N8676 = N8675 | data_masked[2372];
  assign N8675 = N8674 | data_masked[2500];
  assign N8674 = N8673 | data_masked[2628];
  assign N8673 = N8672 | data_masked[2756];
  assign N8672 = N8671 | data_masked[2884];
  assign N8671 = N8670 | data_masked[3012];
  assign N8670 = N8669 | data_masked[3140];
  assign N8669 = N8668 | data_masked[3268];
  assign N8668 = N8667 | data_masked[3396];
  assign N8667 = N8666 | data_masked[3524];
  assign N8666 = N8665 | data_masked[3652];
  assign N8665 = N8664 | data_masked[3780];
  assign N8664 = N8663 | data_masked[3908];
  assign N8663 = N8662 | data_masked[4036];
  assign N8662 = N8661 | data_masked[4164];
  assign N8661 = N8660 | data_masked[4292];
  assign N8660 = N8659 | data_masked[4420];
  assign N8659 = N8658 | data_masked[4548];
  assign N8658 = N8657 | data_masked[4676];
  assign N8657 = N8656 | data_masked[4804];
  assign N8656 = N8655 | data_masked[4932];
  assign N8655 = N8654 | data_masked[5060];
  assign N8654 = N8653 | data_masked[5188];
  assign N8653 = N8652 | data_masked[5316];
  assign N8652 = N8651 | data_masked[5444];
  assign N8651 = N8650 | data_masked[5572];
  assign N8650 = N8649 | data_masked[5700];
  assign N8649 = N8648 | data_masked[5828];
  assign N8648 = N8647 | data_masked[5956];
  assign N8647 = N8646 | data_masked[6084];
  assign N8646 = N8645 | data_masked[6212];
  assign N8645 = N8644 | data_masked[6340];
  assign N8644 = N8643 | data_masked[6468];
  assign N8643 = N8642 | data_masked[6596];
  assign N8642 = N8641 | data_masked[6724];
  assign N8641 = N8640 | data_masked[6852];
  assign N8640 = N8639 | data_masked[6980];
  assign N8639 = N8638 | data_masked[7108];
  assign N8638 = N8637 | data_masked[7236];
  assign N8637 = N8636 | data_masked[7364];
  assign N8636 = N8635 | data_masked[7492];
  assign N8635 = N8634 | data_masked[7620];
  assign N8634 = N8633 | data_masked[7748];
  assign N8633 = N8632 | data_masked[7876];
  assign N8632 = N8631 | data_masked[8004];
  assign N8631 = N8630 | data_masked[8132];
  assign N8630 = N8629 | data_masked[8260];
  assign N8629 = N8628 | data_masked[8388];
  assign N8628 = N8627 | data_masked[8516];
  assign N8627 = N8626 | data_masked[8644];
  assign N8626 = N8625 | data_masked[8772];
  assign N8625 = N8624 | data_masked[8900];
  assign N8624 = N8623 | data_masked[9028];
  assign N8623 = N8622 | data_masked[9156];
  assign N8622 = N8621 | data_masked[9284];
  assign N8621 = N8620 | data_masked[9412];
  assign N8620 = N8619 | data_masked[9540];
  assign N8619 = N8618 | data_masked[9668];
  assign N8618 = N8617 | data_masked[9796];
  assign N8617 = N8616 | data_masked[9924];
  assign N8616 = N8615 | data_masked[10052];
  assign N8615 = N8614 | data_masked[10180];
  assign N8614 = N8613 | data_masked[10308];
  assign N8613 = N8612 | data_masked[10436];
  assign N8612 = N8611 | data_masked[10564];
  assign N8611 = N8610 | data_masked[10692];
  assign N8610 = N8609 | data_masked[10820];
  assign N8609 = N8608 | data_masked[10948];
  assign N8608 = N8607 | data_masked[11076];
  assign N8607 = N8606 | data_masked[11204];
  assign N8606 = N8605 | data_masked[11332];
  assign N8605 = N8604 | data_masked[11460];
  assign N8604 = N8603 | data_masked[11588];
  assign N8603 = N8602 | data_masked[11716];
  assign N8602 = N8601 | data_masked[11844];
  assign N8601 = N8600 | data_masked[11972];
  assign N8600 = N8599 | data_masked[12100];
  assign N8599 = N8598 | data_masked[12228];
  assign N8598 = N8597 | data_masked[12356];
  assign N8597 = N8596 | data_masked[12484];
  assign N8596 = N8595 | data_masked[12612];
  assign N8595 = N8594 | data_masked[12740];
  assign N8594 = N8593 | data_masked[12868];
  assign N8593 = N8592 | data_masked[12996];
  assign N8592 = N8591 | data_masked[13124];
  assign N8591 = N8590 | data_masked[13252];
  assign N8590 = N8589 | data_masked[13380];
  assign N8589 = N8588 | data_masked[13508];
  assign N8588 = N8587 | data_masked[13636];
  assign N8587 = N8586 | data_masked[13764];
  assign N8586 = N8585 | data_masked[13892];
  assign N8585 = N8584 | data_masked[14020];
  assign N8584 = N8583 | data_masked[14148];
  assign N8583 = N8582 | data_masked[14276];
  assign N8582 = N8581 | data_masked[14404];
  assign N8581 = N8580 | data_masked[14532];
  assign N8580 = N8579 | data_masked[14660];
  assign N8579 = N8578 | data_masked[14788];
  assign N8578 = N8577 | data_masked[14916];
  assign N8577 = N8576 | data_masked[15044];
  assign N8576 = N8575 | data_masked[15172];
  assign N8575 = N8574 | data_masked[15300];
  assign N8574 = N8573 | data_masked[15428];
  assign N8573 = N8572 | data_masked[15556];
  assign N8572 = N8571 | data_masked[15684];
  assign N8571 = N8570 | data_masked[15812];
  assign N8570 = N8569 | data_masked[15940];
  assign N8569 = N8568 | data_masked[16068];
  assign N8568 = data_masked[16324] | data_masked[16196];
  assign data_o[69] = N8819 | data_masked[69];
  assign N8819 = N8818 | data_masked[197];
  assign N8818 = N8817 | data_masked[325];
  assign N8817 = N8816 | data_masked[453];
  assign N8816 = N8815 | data_masked[581];
  assign N8815 = N8814 | data_masked[709];
  assign N8814 = N8813 | data_masked[837];
  assign N8813 = N8812 | data_masked[965];
  assign N8812 = N8811 | data_masked[1093];
  assign N8811 = N8810 | data_masked[1221];
  assign N8810 = N8809 | data_masked[1349];
  assign N8809 = N8808 | data_masked[1477];
  assign N8808 = N8807 | data_masked[1605];
  assign N8807 = N8806 | data_masked[1733];
  assign N8806 = N8805 | data_masked[1861];
  assign N8805 = N8804 | data_masked[1989];
  assign N8804 = N8803 | data_masked[2117];
  assign N8803 = N8802 | data_masked[2245];
  assign N8802 = N8801 | data_masked[2373];
  assign N8801 = N8800 | data_masked[2501];
  assign N8800 = N8799 | data_masked[2629];
  assign N8799 = N8798 | data_masked[2757];
  assign N8798 = N8797 | data_masked[2885];
  assign N8797 = N8796 | data_masked[3013];
  assign N8796 = N8795 | data_masked[3141];
  assign N8795 = N8794 | data_masked[3269];
  assign N8794 = N8793 | data_masked[3397];
  assign N8793 = N8792 | data_masked[3525];
  assign N8792 = N8791 | data_masked[3653];
  assign N8791 = N8790 | data_masked[3781];
  assign N8790 = N8789 | data_masked[3909];
  assign N8789 = N8788 | data_masked[4037];
  assign N8788 = N8787 | data_masked[4165];
  assign N8787 = N8786 | data_masked[4293];
  assign N8786 = N8785 | data_masked[4421];
  assign N8785 = N8784 | data_masked[4549];
  assign N8784 = N8783 | data_masked[4677];
  assign N8783 = N8782 | data_masked[4805];
  assign N8782 = N8781 | data_masked[4933];
  assign N8781 = N8780 | data_masked[5061];
  assign N8780 = N8779 | data_masked[5189];
  assign N8779 = N8778 | data_masked[5317];
  assign N8778 = N8777 | data_masked[5445];
  assign N8777 = N8776 | data_masked[5573];
  assign N8776 = N8775 | data_masked[5701];
  assign N8775 = N8774 | data_masked[5829];
  assign N8774 = N8773 | data_masked[5957];
  assign N8773 = N8772 | data_masked[6085];
  assign N8772 = N8771 | data_masked[6213];
  assign N8771 = N8770 | data_masked[6341];
  assign N8770 = N8769 | data_masked[6469];
  assign N8769 = N8768 | data_masked[6597];
  assign N8768 = N8767 | data_masked[6725];
  assign N8767 = N8766 | data_masked[6853];
  assign N8766 = N8765 | data_masked[6981];
  assign N8765 = N8764 | data_masked[7109];
  assign N8764 = N8763 | data_masked[7237];
  assign N8763 = N8762 | data_masked[7365];
  assign N8762 = N8761 | data_masked[7493];
  assign N8761 = N8760 | data_masked[7621];
  assign N8760 = N8759 | data_masked[7749];
  assign N8759 = N8758 | data_masked[7877];
  assign N8758 = N8757 | data_masked[8005];
  assign N8757 = N8756 | data_masked[8133];
  assign N8756 = N8755 | data_masked[8261];
  assign N8755 = N8754 | data_masked[8389];
  assign N8754 = N8753 | data_masked[8517];
  assign N8753 = N8752 | data_masked[8645];
  assign N8752 = N8751 | data_masked[8773];
  assign N8751 = N8750 | data_masked[8901];
  assign N8750 = N8749 | data_masked[9029];
  assign N8749 = N8748 | data_masked[9157];
  assign N8748 = N8747 | data_masked[9285];
  assign N8747 = N8746 | data_masked[9413];
  assign N8746 = N8745 | data_masked[9541];
  assign N8745 = N8744 | data_masked[9669];
  assign N8744 = N8743 | data_masked[9797];
  assign N8743 = N8742 | data_masked[9925];
  assign N8742 = N8741 | data_masked[10053];
  assign N8741 = N8740 | data_masked[10181];
  assign N8740 = N8739 | data_masked[10309];
  assign N8739 = N8738 | data_masked[10437];
  assign N8738 = N8737 | data_masked[10565];
  assign N8737 = N8736 | data_masked[10693];
  assign N8736 = N8735 | data_masked[10821];
  assign N8735 = N8734 | data_masked[10949];
  assign N8734 = N8733 | data_masked[11077];
  assign N8733 = N8732 | data_masked[11205];
  assign N8732 = N8731 | data_masked[11333];
  assign N8731 = N8730 | data_masked[11461];
  assign N8730 = N8729 | data_masked[11589];
  assign N8729 = N8728 | data_masked[11717];
  assign N8728 = N8727 | data_masked[11845];
  assign N8727 = N8726 | data_masked[11973];
  assign N8726 = N8725 | data_masked[12101];
  assign N8725 = N8724 | data_masked[12229];
  assign N8724 = N8723 | data_masked[12357];
  assign N8723 = N8722 | data_masked[12485];
  assign N8722 = N8721 | data_masked[12613];
  assign N8721 = N8720 | data_masked[12741];
  assign N8720 = N8719 | data_masked[12869];
  assign N8719 = N8718 | data_masked[12997];
  assign N8718 = N8717 | data_masked[13125];
  assign N8717 = N8716 | data_masked[13253];
  assign N8716 = N8715 | data_masked[13381];
  assign N8715 = N8714 | data_masked[13509];
  assign N8714 = N8713 | data_masked[13637];
  assign N8713 = N8712 | data_masked[13765];
  assign N8712 = N8711 | data_masked[13893];
  assign N8711 = N8710 | data_masked[14021];
  assign N8710 = N8709 | data_masked[14149];
  assign N8709 = N8708 | data_masked[14277];
  assign N8708 = N8707 | data_masked[14405];
  assign N8707 = N8706 | data_masked[14533];
  assign N8706 = N8705 | data_masked[14661];
  assign N8705 = N8704 | data_masked[14789];
  assign N8704 = N8703 | data_masked[14917];
  assign N8703 = N8702 | data_masked[15045];
  assign N8702 = N8701 | data_masked[15173];
  assign N8701 = N8700 | data_masked[15301];
  assign N8700 = N8699 | data_masked[15429];
  assign N8699 = N8698 | data_masked[15557];
  assign N8698 = N8697 | data_masked[15685];
  assign N8697 = N8696 | data_masked[15813];
  assign N8696 = N8695 | data_masked[15941];
  assign N8695 = N8694 | data_masked[16069];
  assign N8694 = data_masked[16325] | data_masked[16197];
  assign data_o[70] = N8945 | data_masked[70];
  assign N8945 = N8944 | data_masked[198];
  assign N8944 = N8943 | data_masked[326];
  assign N8943 = N8942 | data_masked[454];
  assign N8942 = N8941 | data_masked[582];
  assign N8941 = N8940 | data_masked[710];
  assign N8940 = N8939 | data_masked[838];
  assign N8939 = N8938 | data_masked[966];
  assign N8938 = N8937 | data_masked[1094];
  assign N8937 = N8936 | data_masked[1222];
  assign N8936 = N8935 | data_masked[1350];
  assign N8935 = N8934 | data_masked[1478];
  assign N8934 = N8933 | data_masked[1606];
  assign N8933 = N8932 | data_masked[1734];
  assign N8932 = N8931 | data_masked[1862];
  assign N8931 = N8930 | data_masked[1990];
  assign N8930 = N8929 | data_masked[2118];
  assign N8929 = N8928 | data_masked[2246];
  assign N8928 = N8927 | data_masked[2374];
  assign N8927 = N8926 | data_masked[2502];
  assign N8926 = N8925 | data_masked[2630];
  assign N8925 = N8924 | data_masked[2758];
  assign N8924 = N8923 | data_masked[2886];
  assign N8923 = N8922 | data_masked[3014];
  assign N8922 = N8921 | data_masked[3142];
  assign N8921 = N8920 | data_masked[3270];
  assign N8920 = N8919 | data_masked[3398];
  assign N8919 = N8918 | data_masked[3526];
  assign N8918 = N8917 | data_masked[3654];
  assign N8917 = N8916 | data_masked[3782];
  assign N8916 = N8915 | data_masked[3910];
  assign N8915 = N8914 | data_masked[4038];
  assign N8914 = N8913 | data_masked[4166];
  assign N8913 = N8912 | data_masked[4294];
  assign N8912 = N8911 | data_masked[4422];
  assign N8911 = N8910 | data_masked[4550];
  assign N8910 = N8909 | data_masked[4678];
  assign N8909 = N8908 | data_masked[4806];
  assign N8908 = N8907 | data_masked[4934];
  assign N8907 = N8906 | data_masked[5062];
  assign N8906 = N8905 | data_masked[5190];
  assign N8905 = N8904 | data_masked[5318];
  assign N8904 = N8903 | data_masked[5446];
  assign N8903 = N8902 | data_masked[5574];
  assign N8902 = N8901 | data_masked[5702];
  assign N8901 = N8900 | data_masked[5830];
  assign N8900 = N8899 | data_masked[5958];
  assign N8899 = N8898 | data_masked[6086];
  assign N8898 = N8897 | data_masked[6214];
  assign N8897 = N8896 | data_masked[6342];
  assign N8896 = N8895 | data_masked[6470];
  assign N8895 = N8894 | data_masked[6598];
  assign N8894 = N8893 | data_masked[6726];
  assign N8893 = N8892 | data_masked[6854];
  assign N8892 = N8891 | data_masked[6982];
  assign N8891 = N8890 | data_masked[7110];
  assign N8890 = N8889 | data_masked[7238];
  assign N8889 = N8888 | data_masked[7366];
  assign N8888 = N8887 | data_masked[7494];
  assign N8887 = N8886 | data_masked[7622];
  assign N8886 = N8885 | data_masked[7750];
  assign N8885 = N8884 | data_masked[7878];
  assign N8884 = N8883 | data_masked[8006];
  assign N8883 = N8882 | data_masked[8134];
  assign N8882 = N8881 | data_masked[8262];
  assign N8881 = N8880 | data_masked[8390];
  assign N8880 = N8879 | data_masked[8518];
  assign N8879 = N8878 | data_masked[8646];
  assign N8878 = N8877 | data_masked[8774];
  assign N8877 = N8876 | data_masked[8902];
  assign N8876 = N8875 | data_masked[9030];
  assign N8875 = N8874 | data_masked[9158];
  assign N8874 = N8873 | data_masked[9286];
  assign N8873 = N8872 | data_masked[9414];
  assign N8872 = N8871 | data_masked[9542];
  assign N8871 = N8870 | data_masked[9670];
  assign N8870 = N8869 | data_masked[9798];
  assign N8869 = N8868 | data_masked[9926];
  assign N8868 = N8867 | data_masked[10054];
  assign N8867 = N8866 | data_masked[10182];
  assign N8866 = N8865 | data_masked[10310];
  assign N8865 = N8864 | data_masked[10438];
  assign N8864 = N8863 | data_masked[10566];
  assign N8863 = N8862 | data_masked[10694];
  assign N8862 = N8861 | data_masked[10822];
  assign N8861 = N8860 | data_masked[10950];
  assign N8860 = N8859 | data_masked[11078];
  assign N8859 = N8858 | data_masked[11206];
  assign N8858 = N8857 | data_masked[11334];
  assign N8857 = N8856 | data_masked[11462];
  assign N8856 = N8855 | data_masked[11590];
  assign N8855 = N8854 | data_masked[11718];
  assign N8854 = N8853 | data_masked[11846];
  assign N8853 = N8852 | data_masked[11974];
  assign N8852 = N8851 | data_masked[12102];
  assign N8851 = N8850 | data_masked[12230];
  assign N8850 = N8849 | data_masked[12358];
  assign N8849 = N8848 | data_masked[12486];
  assign N8848 = N8847 | data_masked[12614];
  assign N8847 = N8846 | data_masked[12742];
  assign N8846 = N8845 | data_masked[12870];
  assign N8845 = N8844 | data_masked[12998];
  assign N8844 = N8843 | data_masked[13126];
  assign N8843 = N8842 | data_masked[13254];
  assign N8842 = N8841 | data_masked[13382];
  assign N8841 = N8840 | data_masked[13510];
  assign N8840 = N8839 | data_masked[13638];
  assign N8839 = N8838 | data_masked[13766];
  assign N8838 = N8837 | data_masked[13894];
  assign N8837 = N8836 | data_masked[14022];
  assign N8836 = N8835 | data_masked[14150];
  assign N8835 = N8834 | data_masked[14278];
  assign N8834 = N8833 | data_masked[14406];
  assign N8833 = N8832 | data_masked[14534];
  assign N8832 = N8831 | data_masked[14662];
  assign N8831 = N8830 | data_masked[14790];
  assign N8830 = N8829 | data_masked[14918];
  assign N8829 = N8828 | data_masked[15046];
  assign N8828 = N8827 | data_masked[15174];
  assign N8827 = N8826 | data_masked[15302];
  assign N8826 = N8825 | data_masked[15430];
  assign N8825 = N8824 | data_masked[15558];
  assign N8824 = N8823 | data_masked[15686];
  assign N8823 = N8822 | data_masked[15814];
  assign N8822 = N8821 | data_masked[15942];
  assign N8821 = N8820 | data_masked[16070];
  assign N8820 = data_masked[16326] | data_masked[16198];
  assign data_o[71] = N9071 | data_masked[71];
  assign N9071 = N9070 | data_masked[199];
  assign N9070 = N9069 | data_masked[327];
  assign N9069 = N9068 | data_masked[455];
  assign N9068 = N9067 | data_masked[583];
  assign N9067 = N9066 | data_masked[711];
  assign N9066 = N9065 | data_masked[839];
  assign N9065 = N9064 | data_masked[967];
  assign N9064 = N9063 | data_masked[1095];
  assign N9063 = N9062 | data_masked[1223];
  assign N9062 = N9061 | data_masked[1351];
  assign N9061 = N9060 | data_masked[1479];
  assign N9060 = N9059 | data_masked[1607];
  assign N9059 = N9058 | data_masked[1735];
  assign N9058 = N9057 | data_masked[1863];
  assign N9057 = N9056 | data_masked[1991];
  assign N9056 = N9055 | data_masked[2119];
  assign N9055 = N9054 | data_masked[2247];
  assign N9054 = N9053 | data_masked[2375];
  assign N9053 = N9052 | data_masked[2503];
  assign N9052 = N9051 | data_masked[2631];
  assign N9051 = N9050 | data_masked[2759];
  assign N9050 = N9049 | data_masked[2887];
  assign N9049 = N9048 | data_masked[3015];
  assign N9048 = N9047 | data_masked[3143];
  assign N9047 = N9046 | data_masked[3271];
  assign N9046 = N9045 | data_masked[3399];
  assign N9045 = N9044 | data_masked[3527];
  assign N9044 = N9043 | data_masked[3655];
  assign N9043 = N9042 | data_masked[3783];
  assign N9042 = N9041 | data_masked[3911];
  assign N9041 = N9040 | data_masked[4039];
  assign N9040 = N9039 | data_masked[4167];
  assign N9039 = N9038 | data_masked[4295];
  assign N9038 = N9037 | data_masked[4423];
  assign N9037 = N9036 | data_masked[4551];
  assign N9036 = N9035 | data_masked[4679];
  assign N9035 = N9034 | data_masked[4807];
  assign N9034 = N9033 | data_masked[4935];
  assign N9033 = N9032 | data_masked[5063];
  assign N9032 = N9031 | data_masked[5191];
  assign N9031 = N9030 | data_masked[5319];
  assign N9030 = N9029 | data_masked[5447];
  assign N9029 = N9028 | data_masked[5575];
  assign N9028 = N9027 | data_masked[5703];
  assign N9027 = N9026 | data_masked[5831];
  assign N9026 = N9025 | data_masked[5959];
  assign N9025 = N9024 | data_masked[6087];
  assign N9024 = N9023 | data_masked[6215];
  assign N9023 = N9022 | data_masked[6343];
  assign N9022 = N9021 | data_masked[6471];
  assign N9021 = N9020 | data_masked[6599];
  assign N9020 = N9019 | data_masked[6727];
  assign N9019 = N9018 | data_masked[6855];
  assign N9018 = N9017 | data_masked[6983];
  assign N9017 = N9016 | data_masked[7111];
  assign N9016 = N9015 | data_masked[7239];
  assign N9015 = N9014 | data_masked[7367];
  assign N9014 = N9013 | data_masked[7495];
  assign N9013 = N9012 | data_masked[7623];
  assign N9012 = N9011 | data_masked[7751];
  assign N9011 = N9010 | data_masked[7879];
  assign N9010 = N9009 | data_masked[8007];
  assign N9009 = N9008 | data_masked[8135];
  assign N9008 = N9007 | data_masked[8263];
  assign N9007 = N9006 | data_masked[8391];
  assign N9006 = N9005 | data_masked[8519];
  assign N9005 = N9004 | data_masked[8647];
  assign N9004 = N9003 | data_masked[8775];
  assign N9003 = N9002 | data_masked[8903];
  assign N9002 = N9001 | data_masked[9031];
  assign N9001 = N9000 | data_masked[9159];
  assign N9000 = N8999 | data_masked[9287];
  assign N8999 = N8998 | data_masked[9415];
  assign N8998 = N8997 | data_masked[9543];
  assign N8997 = N8996 | data_masked[9671];
  assign N8996 = N8995 | data_masked[9799];
  assign N8995 = N8994 | data_masked[9927];
  assign N8994 = N8993 | data_masked[10055];
  assign N8993 = N8992 | data_masked[10183];
  assign N8992 = N8991 | data_masked[10311];
  assign N8991 = N8990 | data_masked[10439];
  assign N8990 = N8989 | data_masked[10567];
  assign N8989 = N8988 | data_masked[10695];
  assign N8988 = N8987 | data_masked[10823];
  assign N8987 = N8986 | data_masked[10951];
  assign N8986 = N8985 | data_masked[11079];
  assign N8985 = N8984 | data_masked[11207];
  assign N8984 = N8983 | data_masked[11335];
  assign N8983 = N8982 | data_masked[11463];
  assign N8982 = N8981 | data_masked[11591];
  assign N8981 = N8980 | data_masked[11719];
  assign N8980 = N8979 | data_masked[11847];
  assign N8979 = N8978 | data_masked[11975];
  assign N8978 = N8977 | data_masked[12103];
  assign N8977 = N8976 | data_masked[12231];
  assign N8976 = N8975 | data_masked[12359];
  assign N8975 = N8974 | data_masked[12487];
  assign N8974 = N8973 | data_masked[12615];
  assign N8973 = N8972 | data_masked[12743];
  assign N8972 = N8971 | data_masked[12871];
  assign N8971 = N8970 | data_masked[12999];
  assign N8970 = N8969 | data_masked[13127];
  assign N8969 = N8968 | data_masked[13255];
  assign N8968 = N8967 | data_masked[13383];
  assign N8967 = N8966 | data_masked[13511];
  assign N8966 = N8965 | data_masked[13639];
  assign N8965 = N8964 | data_masked[13767];
  assign N8964 = N8963 | data_masked[13895];
  assign N8963 = N8962 | data_masked[14023];
  assign N8962 = N8961 | data_masked[14151];
  assign N8961 = N8960 | data_masked[14279];
  assign N8960 = N8959 | data_masked[14407];
  assign N8959 = N8958 | data_masked[14535];
  assign N8958 = N8957 | data_masked[14663];
  assign N8957 = N8956 | data_masked[14791];
  assign N8956 = N8955 | data_masked[14919];
  assign N8955 = N8954 | data_masked[15047];
  assign N8954 = N8953 | data_masked[15175];
  assign N8953 = N8952 | data_masked[15303];
  assign N8952 = N8951 | data_masked[15431];
  assign N8951 = N8950 | data_masked[15559];
  assign N8950 = N8949 | data_masked[15687];
  assign N8949 = N8948 | data_masked[15815];
  assign N8948 = N8947 | data_masked[15943];
  assign N8947 = N8946 | data_masked[16071];
  assign N8946 = data_masked[16327] | data_masked[16199];
  assign data_o[72] = N9197 | data_masked[72];
  assign N9197 = N9196 | data_masked[200];
  assign N9196 = N9195 | data_masked[328];
  assign N9195 = N9194 | data_masked[456];
  assign N9194 = N9193 | data_masked[584];
  assign N9193 = N9192 | data_masked[712];
  assign N9192 = N9191 | data_masked[840];
  assign N9191 = N9190 | data_masked[968];
  assign N9190 = N9189 | data_masked[1096];
  assign N9189 = N9188 | data_masked[1224];
  assign N9188 = N9187 | data_masked[1352];
  assign N9187 = N9186 | data_masked[1480];
  assign N9186 = N9185 | data_masked[1608];
  assign N9185 = N9184 | data_masked[1736];
  assign N9184 = N9183 | data_masked[1864];
  assign N9183 = N9182 | data_masked[1992];
  assign N9182 = N9181 | data_masked[2120];
  assign N9181 = N9180 | data_masked[2248];
  assign N9180 = N9179 | data_masked[2376];
  assign N9179 = N9178 | data_masked[2504];
  assign N9178 = N9177 | data_masked[2632];
  assign N9177 = N9176 | data_masked[2760];
  assign N9176 = N9175 | data_masked[2888];
  assign N9175 = N9174 | data_masked[3016];
  assign N9174 = N9173 | data_masked[3144];
  assign N9173 = N9172 | data_masked[3272];
  assign N9172 = N9171 | data_masked[3400];
  assign N9171 = N9170 | data_masked[3528];
  assign N9170 = N9169 | data_masked[3656];
  assign N9169 = N9168 | data_masked[3784];
  assign N9168 = N9167 | data_masked[3912];
  assign N9167 = N9166 | data_masked[4040];
  assign N9166 = N9165 | data_masked[4168];
  assign N9165 = N9164 | data_masked[4296];
  assign N9164 = N9163 | data_masked[4424];
  assign N9163 = N9162 | data_masked[4552];
  assign N9162 = N9161 | data_masked[4680];
  assign N9161 = N9160 | data_masked[4808];
  assign N9160 = N9159 | data_masked[4936];
  assign N9159 = N9158 | data_masked[5064];
  assign N9158 = N9157 | data_masked[5192];
  assign N9157 = N9156 | data_masked[5320];
  assign N9156 = N9155 | data_masked[5448];
  assign N9155 = N9154 | data_masked[5576];
  assign N9154 = N9153 | data_masked[5704];
  assign N9153 = N9152 | data_masked[5832];
  assign N9152 = N9151 | data_masked[5960];
  assign N9151 = N9150 | data_masked[6088];
  assign N9150 = N9149 | data_masked[6216];
  assign N9149 = N9148 | data_masked[6344];
  assign N9148 = N9147 | data_masked[6472];
  assign N9147 = N9146 | data_masked[6600];
  assign N9146 = N9145 | data_masked[6728];
  assign N9145 = N9144 | data_masked[6856];
  assign N9144 = N9143 | data_masked[6984];
  assign N9143 = N9142 | data_masked[7112];
  assign N9142 = N9141 | data_masked[7240];
  assign N9141 = N9140 | data_masked[7368];
  assign N9140 = N9139 | data_masked[7496];
  assign N9139 = N9138 | data_masked[7624];
  assign N9138 = N9137 | data_masked[7752];
  assign N9137 = N9136 | data_masked[7880];
  assign N9136 = N9135 | data_masked[8008];
  assign N9135 = N9134 | data_masked[8136];
  assign N9134 = N9133 | data_masked[8264];
  assign N9133 = N9132 | data_masked[8392];
  assign N9132 = N9131 | data_masked[8520];
  assign N9131 = N9130 | data_masked[8648];
  assign N9130 = N9129 | data_masked[8776];
  assign N9129 = N9128 | data_masked[8904];
  assign N9128 = N9127 | data_masked[9032];
  assign N9127 = N9126 | data_masked[9160];
  assign N9126 = N9125 | data_masked[9288];
  assign N9125 = N9124 | data_masked[9416];
  assign N9124 = N9123 | data_masked[9544];
  assign N9123 = N9122 | data_masked[9672];
  assign N9122 = N9121 | data_masked[9800];
  assign N9121 = N9120 | data_masked[9928];
  assign N9120 = N9119 | data_masked[10056];
  assign N9119 = N9118 | data_masked[10184];
  assign N9118 = N9117 | data_masked[10312];
  assign N9117 = N9116 | data_masked[10440];
  assign N9116 = N9115 | data_masked[10568];
  assign N9115 = N9114 | data_masked[10696];
  assign N9114 = N9113 | data_masked[10824];
  assign N9113 = N9112 | data_masked[10952];
  assign N9112 = N9111 | data_masked[11080];
  assign N9111 = N9110 | data_masked[11208];
  assign N9110 = N9109 | data_masked[11336];
  assign N9109 = N9108 | data_masked[11464];
  assign N9108 = N9107 | data_masked[11592];
  assign N9107 = N9106 | data_masked[11720];
  assign N9106 = N9105 | data_masked[11848];
  assign N9105 = N9104 | data_masked[11976];
  assign N9104 = N9103 | data_masked[12104];
  assign N9103 = N9102 | data_masked[12232];
  assign N9102 = N9101 | data_masked[12360];
  assign N9101 = N9100 | data_masked[12488];
  assign N9100 = N9099 | data_masked[12616];
  assign N9099 = N9098 | data_masked[12744];
  assign N9098 = N9097 | data_masked[12872];
  assign N9097 = N9096 | data_masked[13000];
  assign N9096 = N9095 | data_masked[13128];
  assign N9095 = N9094 | data_masked[13256];
  assign N9094 = N9093 | data_masked[13384];
  assign N9093 = N9092 | data_masked[13512];
  assign N9092 = N9091 | data_masked[13640];
  assign N9091 = N9090 | data_masked[13768];
  assign N9090 = N9089 | data_masked[13896];
  assign N9089 = N9088 | data_masked[14024];
  assign N9088 = N9087 | data_masked[14152];
  assign N9087 = N9086 | data_masked[14280];
  assign N9086 = N9085 | data_masked[14408];
  assign N9085 = N9084 | data_masked[14536];
  assign N9084 = N9083 | data_masked[14664];
  assign N9083 = N9082 | data_masked[14792];
  assign N9082 = N9081 | data_masked[14920];
  assign N9081 = N9080 | data_masked[15048];
  assign N9080 = N9079 | data_masked[15176];
  assign N9079 = N9078 | data_masked[15304];
  assign N9078 = N9077 | data_masked[15432];
  assign N9077 = N9076 | data_masked[15560];
  assign N9076 = N9075 | data_masked[15688];
  assign N9075 = N9074 | data_masked[15816];
  assign N9074 = N9073 | data_masked[15944];
  assign N9073 = N9072 | data_masked[16072];
  assign N9072 = data_masked[16328] | data_masked[16200];
  assign data_o[73] = N9323 | data_masked[73];
  assign N9323 = N9322 | data_masked[201];
  assign N9322 = N9321 | data_masked[329];
  assign N9321 = N9320 | data_masked[457];
  assign N9320 = N9319 | data_masked[585];
  assign N9319 = N9318 | data_masked[713];
  assign N9318 = N9317 | data_masked[841];
  assign N9317 = N9316 | data_masked[969];
  assign N9316 = N9315 | data_masked[1097];
  assign N9315 = N9314 | data_masked[1225];
  assign N9314 = N9313 | data_masked[1353];
  assign N9313 = N9312 | data_masked[1481];
  assign N9312 = N9311 | data_masked[1609];
  assign N9311 = N9310 | data_masked[1737];
  assign N9310 = N9309 | data_masked[1865];
  assign N9309 = N9308 | data_masked[1993];
  assign N9308 = N9307 | data_masked[2121];
  assign N9307 = N9306 | data_masked[2249];
  assign N9306 = N9305 | data_masked[2377];
  assign N9305 = N9304 | data_masked[2505];
  assign N9304 = N9303 | data_masked[2633];
  assign N9303 = N9302 | data_masked[2761];
  assign N9302 = N9301 | data_masked[2889];
  assign N9301 = N9300 | data_masked[3017];
  assign N9300 = N9299 | data_masked[3145];
  assign N9299 = N9298 | data_masked[3273];
  assign N9298 = N9297 | data_masked[3401];
  assign N9297 = N9296 | data_masked[3529];
  assign N9296 = N9295 | data_masked[3657];
  assign N9295 = N9294 | data_masked[3785];
  assign N9294 = N9293 | data_masked[3913];
  assign N9293 = N9292 | data_masked[4041];
  assign N9292 = N9291 | data_masked[4169];
  assign N9291 = N9290 | data_masked[4297];
  assign N9290 = N9289 | data_masked[4425];
  assign N9289 = N9288 | data_masked[4553];
  assign N9288 = N9287 | data_masked[4681];
  assign N9287 = N9286 | data_masked[4809];
  assign N9286 = N9285 | data_masked[4937];
  assign N9285 = N9284 | data_masked[5065];
  assign N9284 = N9283 | data_masked[5193];
  assign N9283 = N9282 | data_masked[5321];
  assign N9282 = N9281 | data_masked[5449];
  assign N9281 = N9280 | data_masked[5577];
  assign N9280 = N9279 | data_masked[5705];
  assign N9279 = N9278 | data_masked[5833];
  assign N9278 = N9277 | data_masked[5961];
  assign N9277 = N9276 | data_masked[6089];
  assign N9276 = N9275 | data_masked[6217];
  assign N9275 = N9274 | data_masked[6345];
  assign N9274 = N9273 | data_masked[6473];
  assign N9273 = N9272 | data_masked[6601];
  assign N9272 = N9271 | data_masked[6729];
  assign N9271 = N9270 | data_masked[6857];
  assign N9270 = N9269 | data_masked[6985];
  assign N9269 = N9268 | data_masked[7113];
  assign N9268 = N9267 | data_masked[7241];
  assign N9267 = N9266 | data_masked[7369];
  assign N9266 = N9265 | data_masked[7497];
  assign N9265 = N9264 | data_masked[7625];
  assign N9264 = N9263 | data_masked[7753];
  assign N9263 = N9262 | data_masked[7881];
  assign N9262 = N9261 | data_masked[8009];
  assign N9261 = N9260 | data_masked[8137];
  assign N9260 = N9259 | data_masked[8265];
  assign N9259 = N9258 | data_masked[8393];
  assign N9258 = N9257 | data_masked[8521];
  assign N9257 = N9256 | data_masked[8649];
  assign N9256 = N9255 | data_masked[8777];
  assign N9255 = N9254 | data_masked[8905];
  assign N9254 = N9253 | data_masked[9033];
  assign N9253 = N9252 | data_masked[9161];
  assign N9252 = N9251 | data_masked[9289];
  assign N9251 = N9250 | data_masked[9417];
  assign N9250 = N9249 | data_masked[9545];
  assign N9249 = N9248 | data_masked[9673];
  assign N9248 = N9247 | data_masked[9801];
  assign N9247 = N9246 | data_masked[9929];
  assign N9246 = N9245 | data_masked[10057];
  assign N9245 = N9244 | data_masked[10185];
  assign N9244 = N9243 | data_masked[10313];
  assign N9243 = N9242 | data_masked[10441];
  assign N9242 = N9241 | data_masked[10569];
  assign N9241 = N9240 | data_masked[10697];
  assign N9240 = N9239 | data_masked[10825];
  assign N9239 = N9238 | data_masked[10953];
  assign N9238 = N9237 | data_masked[11081];
  assign N9237 = N9236 | data_masked[11209];
  assign N9236 = N9235 | data_masked[11337];
  assign N9235 = N9234 | data_masked[11465];
  assign N9234 = N9233 | data_masked[11593];
  assign N9233 = N9232 | data_masked[11721];
  assign N9232 = N9231 | data_masked[11849];
  assign N9231 = N9230 | data_masked[11977];
  assign N9230 = N9229 | data_masked[12105];
  assign N9229 = N9228 | data_masked[12233];
  assign N9228 = N9227 | data_masked[12361];
  assign N9227 = N9226 | data_masked[12489];
  assign N9226 = N9225 | data_masked[12617];
  assign N9225 = N9224 | data_masked[12745];
  assign N9224 = N9223 | data_masked[12873];
  assign N9223 = N9222 | data_masked[13001];
  assign N9222 = N9221 | data_masked[13129];
  assign N9221 = N9220 | data_masked[13257];
  assign N9220 = N9219 | data_masked[13385];
  assign N9219 = N9218 | data_masked[13513];
  assign N9218 = N9217 | data_masked[13641];
  assign N9217 = N9216 | data_masked[13769];
  assign N9216 = N9215 | data_masked[13897];
  assign N9215 = N9214 | data_masked[14025];
  assign N9214 = N9213 | data_masked[14153];
  assign N9213 = N9212 | data_masked[14281];
  assign N9212 = N9211 | data_masked[14409];
  assign N9211 = N9210 | data_masked[14537];
  assign N9210 = N9209 | data_masked[14665];
  assign N9209 = N9208 | data_masked[14793];
  assign N9208 = N9207 | data_masked[14921];
  assign N9207 = N9206 | data_masked[15049];
  assign N9206 = N9205 | data_masked[15177];
  assign N9205 = N9204 | data_masked[15305];
  assign N9204 = N9203 | data_masked[15433];
  assign N9203 = N9202 | data_masked[15561];
  assign N9202 = N9201 | data_masked[15689];
  assign N9201 = N9200 | data_masked[15817];
  assign N9200 = N9199 | data_masked[15945];
  assign N9199 = N9198 | data_masked[16073];
  assign N9198 = data_masked[16329] | data_masked[16201];
  assign data_o[74] = N9449 | data_masked[74];
  assign N9449 = N9448 | data_masked[202];
  assign N9448 = N9447 | data_masked[330];
  assign N9447 = N9446 | data_masked[458];
  assign N9446 = N9445 | data_masked[586];
  assign N9445 = N9444 | data_masked[714];
  assign N9444 = N9443 | data_masked[842];
  assign N9443 = N9442 | data_masked[970];
  assign N9442 = N9441 | data_masked[1098];
  assign N9441 = N9440 | data_masked[1226];
  assign N9440 = N9439 | data_masked[1354];
  assign N9439 = N9438 | data_masked[1482];
  assign N9438 = N9437 | data_masked[1610];
  assign N9437 = N9436 | data_masked[1738];
  assign N9436 = N9435 | data_masked[1866];
  assign N9435 = N9434 | data_masked[1994];
  assign N9434 = N9433 | data_masked[2122];
  assign N9433 = N9432 | data_masked[2250];
  assign N9432 = N9431 | data_masked[2378];
  assign N9431 = N9430 | data_masked[2506];
  assign N9430 = N9429 | data_masked[2634];
  assign N9429 = N9428 | data_masked[2762];
  assign N9428 = N9427 | data_masked[2890];
  assign N9427 = N9426 | data_masked[3018];
  assign N9426 = N9425 | data_masked[3146];
  assign N9425 = N9424 | data_masked[3274];
  assign N9424 = N9423 | data_masked[3402];
  assign N9423 = N9422 | data_masked[3530];
  assign N9422 = N9421 | data_masked[3658];
  assign N9421 = N9420 | data_masked[3786];
  assign N9420 = N9419 | data_masked[3914];
  assign N9419 = N9418 | data_masked[4042];
  assign N9418 = N9417 | data_masked[4170];
  assign N9417 = N9416 | data_masked[4298];
  assign N9416 = N9415 | data_masked[4426];
  assign N9415 = N9414 | data_masked[4554];
  assign N9414 = N9413 | data_masked[4682];
  assign N9413 = N9412 | data_masked[4810];
  assign N9412 = N9411 | data_masked[4938];
  assign N9411 = N9410 | data_masked[5066];
  assign N9410 = N9409 | data_masked[5194];
  assign N9409 = N9408 | data_masked[5322];
  assign N9408 = N9407 | data_masked[5450];
  assign N9407 = N9406 | data_masked[5578];
  assign N9406 = N9405 | data_masked[5706];
  assign N9405 = N9404 | data_masked[5834];
  assign N9404 = N9403 | data_masked[5962];
  assign N9403 = N9402 | data_masked[6090];
  assign N9402 = N9401 | data_masked[6218];
  assign N9401 = N9400 | data_masked[6346];
  assign N9400 = N9399 | data_masked[6474];
  assign N9399 = N9398 | data_masked[6602];
  assign N9398 = N9397 | data_masked[6730];
  assign N9397 = N9396 | data_masked[6858];
  assign N9396 = N9395 | data_masked[6986];
  assign N9395 = N9394 | data_masked[7114];
  assign N9394 = N9393 | data_masked[7242];
  assign N9393 = N9392 | data_masked[7370];
  assign N9392 = N9391 | data_masked[7498];
  assign N9391 = N9390 | data_masked[7626];
  assign N9390 = N9389 | data_masked[7754];
  assign N9389 = N9388 | data_masked[7882];
  assign N9388 = N9387 | data_masked[8010];
  assign N9387 = N9386 | data_masked[8138];
  assign N9386 = N9385 | data_masked[8266];
  assign N9385 = N9384 | data_masked[8394];
  assign N9384 = N9383 | data_masked[8522];
  assign N9383 = N9382 | data_masked[8650];
  assign N9382 = N9381 | data_masked[8778];
  assign N9381 = N9380 | data_masked[8906];
  assign N9380 = N9379 | data_masked[9034];
  assign N9379 = N9378 | data_masked[9162];
  assign N9378 = N9377 | data_masked[9290];
  assign N9377 = N9376 | data_masked[9418];
  assign N9376 = N9375 | data_masked[9546];
  assign N9375 = N9374 | data_masked[9674];
  assign N9374 = N9373 | data_masked[9802];
  assign N9373 = N9372 | data_masked[9930];
  assign N9372 = N9371 | data_masked[10058];
  assign N9371 = N9370 | data_masked[10186];
  assign N9370 = N9369 | data_masked[10314];
  assign N9369 = N9368 | data_masked[10442];
  assign N9368 = N9367 | data_masked[10570];
  assign N9367 = N9366 | data_masked[10698];
  assign N9366 = N9365 | data_masked[10826];
  assign N9365 = N9364 | data_masked[10954];
  assign N9364 = N9363 | data_masked[11082];
  assign N9363 = N9362 | data_masked[11210];
  assign N9362 = N9361 | data_masked[11338];
  assign N9361 = N9360 | data_masked[11466];
  assign N9360 = N9359 | data_masked[11594];
  assign N9359 = N9358 | data_masked[11722];
  assign N9358 = N9357 | data_masked[11850];
  assign N9357 = N9356 | data_masked[11978];
  assign N9356 = N9355 | data_masked[12106];
  assign N9355 = N9354 | data_masked[12234];
  assign N9354 = N9353 | data_masked[12362];
  assign N9353 = N9352 | data_masked[12490];
  assign N9352 = N9351 | data_masked[12618];
  assign N9351 = N9350 | data_masked[12746];
  assign N9350 = N9349 | data_masked[12874];
  assign N9349 = N9348 | data_masked[13002];
  assign N9348 = N9347 | data_masked[13130];
  assign N9347 = N9346 | data_masked[13258];
  assign N9346 = N9345 | data_masked[13386];
  assign N9345 = N9344 | data_masked[13514];
  assign N9344 = N9343 | data_masked[13642];
  assign N9343 = N9342 | data_masked[13770];
  assign N9342 = N9341 | data_masked[13898];
  assign N9341 = N9340 | data_masked[14026];
  assign N9340 = N9339 | data_masked[14154];
  assign N9339 = N9338 | data_masked[14282];
  assign N9338 = N9337 | data_masked[14410];
  assign N9337 = N9336 | data_masked[14538];
  assign N9336 = N9335 | data_masked[14666];
  assign N9335 = N9334 | data_masked[14794];
  assign N9334 = N9333 | data_masked[14922];
  assign N9333 = N9332 | data_masked[15050];
  assign N9332 = N9331 | data_masked[15178];
  assign N9331 = N9330 | data_masked[15306];
  assign N9330 = N9329 | data_masked[15434];
  assign N9329 = N9328 | data_masked[15562];
  assign N9328 = N9327 | data_masked[15690];
  assign N9327 = N9326 | data_masked[15818];
  assign N9326 = N9325 | data_masked[15946];
  assign N9325 = N9324 | data_masked[16074];
  assign N9324 = data_masked[16330] | data_masked[16202];
  assign data_o[75] = N9575 | data_masked[75];
  assign N9575 = N9574 | data_masked[203];
  assign N9574 = N9573 | data_masked[331];
  assign N9573 = N9572 | data_masked[459];
  assign N9572 = N9571 | data_masked[587];
  assign N9571 = N9570 | data_masked[715];
  assign N9570 = N9569 | data_masked[843];
  assign N9569 = N9568 | data_masked[971];
  assign N9568 = N9567 | data_masked[1099];
  assign N9567 = N9566 | data_masked[1227];
  assign N9566 = N9565 | data_masked[1355];
  assign N9565 = N9564 | data_masked[1483];
  assign N9564 = N9563 | data_masked[1611];
  assign N9563 = N9562 | data_masked[1739];
  assign N9562 = N9561 | data_masked[1867];
  assign N9561 = N9560 | data_masked[1995];
  assign N9560 = N9559 | data_masked[2123];
  assign N9559 = N9558 | data_masked[2251];
  assign N9558 = N9557 | data_masked[2379];
  assign N9557 = N9556 | data_masked[2507];
  assign N9556 = N9555 | data_masked[2635];
  assign N9555 = N9554 | data_masked[2763];
  assign N9554 = N9553 | data_masked[2891];
  assign N9553 = N9552 | data_masked[3019];
  assign N9552 = N9551 | data_masked[3147];
  assign N9551 = N9550 | data_masked[3275];
  assign N9550 = N9549 | data_masked[3403];
  assign N9549 = N9548 | data_masked[3531];
  assign N9548 = N9547 | data_masked[3659];
  assign N9547 = N9546 | data_masked[3787];
  assign N9546 = N9545 | data_masked[3915];
  assign N9545 = N9544 | data_masked[4043];
  assign N9544 = N9543 | data_masked[4171];
  assign N9543 = N9542 | data_masked[4299];
  assign N9542 = N9541 | data_masked[4427];
  assign N9541 = N9540 | data_masked[4555];
  assign N9540 = N9539 | data_masked[4683];
  assign N9539 = N9538 | data_masked[4811];
  assign N9538 = N9537 | data_masked[4939];
  assign N9537 = N9536 | data_masked[5067];
  assign N9536 = N9535 | data_masked[5195];
  assign N9535 = N9534 | data_masked[5323];
  assign N9534 = N9533 | data_masked[5451];
  assign N9533 = N9532 | data_masked[5579];
  assign N9532 = N9531 | data_masked[5707];
  assign N9531 = N9530 | data_masked[5835];
  assign N9530 = N9529 | data_masked[5963];
  assign N9529 = N9528 | data_masked[6091];
  assign N9528 = N9527 | data_masked[6219];
  assign N9527 = N9526 | data_masked[6347];
  assign N9526 = N9525 | data_masked[6475];
  assign N9525 = N9524 | data_masked[6603];
  assign N9524 = N9523 | data_masked[6731];
  assign N9523 = N9522 | data_masked[6859];
  assign N9522 = N9521 | data_masked[6987];
  assign N9521 = N9520 | data_masked[7115];
  assign N9520 = N9519 | data_masked[7243];
  assign N9519 = N9518 | data_masked[7371];
  assign N9518 = N9517 | data_masked[7499];
  assign N9517 = N9516 | data_masked[7627];
  assign N9516 = N9515 | data_masked[7755];
  assign N9515 = N9514 | data_masked[7883];
  assign N9514 = N9513 | data_masked[8011];
  assign N9513 = N9512 | data_masked[8139];
  assign N9512 = N9511 | data_masked[8267];
  assign N9511 = N9510 | data_masked[8395];
  assign N9510 = N9509 | data_masked[8523];
  assign N9509 = N9508 | data_masked[8651];
  assign N9508 = N9507 | data_masked[8779];
  assign N9507 = N9506 | data_masked[8907];
  assign N9506 = N9505 | data_masked[9035];
  assign N9505 = N9504 | data_masked[9163];
  assign N9504 = N9503 | data_masked[9291];
  assign N9503 = N9502 | data_masked[9419];
  assign N9502 = N9501 | data_masked[9547];
  assign N9501 = N9500 | data_masked[9675];
  assign N9500 = N9499 | data_masked[9803];
  assign N9499 = N9498 | data_masked[9931];
  assign N9498 = N9497 | data_masked[10059];
  assign N9497 = N9496 | data_masked[10187];
  assign N9496 = N9495 | data_masked[10315];
  assign N9495 = N9494 | data_masked[10443];
  assign N9494 = N9493 | data_masked[10571];
  assign N9493 = N9492 | data_masked[10699];
  assign N9492 = N9491 | data_masked[10827];
  assign N9491 = N9490 | data_masked[10955];
  assign N9490 = N9489 | data_masked[11083];
  assign N9489 = N9488 | data_masked[11211];
  assign N9488 = N9487 | data_masked[11339];
  assign N9487 = N9486 | data_masked[11467];
  assign N9486 = N9485 | data_masked[11595];
  assign N9485 = N9484 | data_masked[11723];
  assign N9484 = N9483 | data_masked[11851];
  assign N9483 = N9482 | data_masked[11979];
  assign N9482 = N9481 | data_masked[12107];
  assign N9481 = N9480 | data_masked[12235];
  assign N9480 = N9479 | data_masked[12363];
  assign N9479 = N9478 | data_masked[12491];
  assign N9478 = N9477 | data_masked[12619];
  assign N9477 = N9476 | data_masked[12747];
  assign N9476 = N9475 | data_masked[12875];
  assign N9475 = N9474 | data_masked[13003];
  assign N9474 = N9473 | data_masked[13131];
  assign N9473 = N9472 | data_masked[13259];
  assign N9472 = N9471 | data_masked[13387];
  assign N9471 = N9470 | data_masked[13515];
  assign N9470 = N9469 | data_masked[13643];
  assign N9469 = N9468 | data_masked[13771];
  assign N9468 = N9467 | data_masked[13899];
  assign N9467 = N9466 | data_masked[14027];
  assign N9466 = N9465 | data_masked[14155];
  assign N9465 = N9464 | data_masked[14283];
  assign N9464 = N9463 | data_masked[14411];
  assign N9463 = N9462 | data_masked[14539];
  assign N9462 = N9461 | data_masked[14667];
  assign N9461 = N9460 | data_masked[14795];
  assign N9460 = N9459 | data_masked[14923];
  assign N9459 = N9458 | data_masked[15051];
  assign N9458 = N9457 | data_masked[15179];
  assign N9457 = N9456 | data_masked[15307];
  assign N9456 = N9455 | data_masked[15435];
  assign N9455 = N9454 | data_masked[15563];
  assign N9454 = N9453 | data_masked[15691];
  assign N9453 = N9452 | data_masked[15819];
  assign N9452 = N9451 | data_masked[15947];
  assign N9451 = N9450 | data_masked[16075];
  assign N9450 = data_masked[16331] | data_masked[16203];
  assign data_o[76] = N9701 | data_masked[76];
  assign N9701 = N9700 | data_masked[204];
  assign N9700 = N9699 | data_masked[332];
  assign N9699 = N9698 | data_masked[460];
  assign N9698 = N9697 | data_masked[588];
  assign N9697 = N9696 | data_masked[716];
  assign N9696 = N9695 | data_masked[844];
  assign N9695 = N9694 | data_masked[972];
  assign N9694 = N9693 | data_masked[1100];
  assign N9693 = N9692 | data_masked[1228];
  assign N9692 = N9691 | data_masked[1356];
  assign N9691 = N9690 | data_masked[1484];
  assign N9690 = N9689 | data_masked[1612];
  assign N9689 = N9688 | data_masked[1740];
  assign N9688 = N9687 | data_masked[1868];
  assign N9687 = N9686 | data_masked[1996];
  assign N9686 = N9685 | data_masked[2124];
  assign N9685 = N9684 | data_masked[2252];
  assign N9684 = N9683 | data_masked[2380];
  assign N9683 = N9682 | data_masked[2508];
  assign N9682 = N9681 | data_masked[2636];
  assign N9681 = N9680 | data_masked[2764];
  assign N9680 = N9679 | data_masked[2892];
  assign N9679 = N9678 | data_masked[3020];
  assign N9678 = N9677 | data_masked[3148];
  assign N9677 = N9676 | data_masked[3276];
  assign N9676 = N9675 | data_masked[3404];
  assign N9675 = N9674 | data_masked[3532];
  assign N9674 = N9673 | data_masked[3660];
  assign N9673 = N9672 | data_masked[3788];
  assign N9672 = N9671 | data_masked[3916];
  assign N9671 = N9670 | data_masked[4044];
  assign N9670 = N9669 | data_masked[4172];
  assign N9669 = N9668 | data_masked[4300];
  assign N9668 = N9667 | data_masked[4428];
  assign N9667 = N9666 | data_masked[4556];
  assign N9666 = N9665 | data_masked[4684];
  assign N9665 = N9664 | data_masked[4812];
  assign N9664 = N9663 | data_masked[4940];
  assign N9663 = N9662 | data_masked[5068];
  assign N9662 = N9661 | data_masked[5196];
  assign N9661 = N9660 | data_masked[5324];
  assign N9660 = N9659 | data_masked[5452];
  assign N9659 = N9658 | data_masked[5580];
  assign N9658 = N9657 | data_masked[5708];
  assign N9657 = N9656 | data_masked[5836];
  assign N9656 = N9655 | data_masked[5964];
  assign N9655 = N9654 | data_masked[6092];
  assign N9654 = N9653 | data_masked[6220];
  assign N9653 = N9652 | data_masked[6348];
  assign N9652 = N9651 | data_masked[6476];
  assign N9651 = N9650 | data_masked[6604];
  assign N9650 = N9649 | data_masked[6732];
  assign N9649 = N9648 | data_masked[6860];
  assign N9648 = N9647 | data_masked[6988];
  assign N9647 = N9646 | data_masked[7116];
  assign N9646 = N9645 | data_masked[7244];
  assign N9645 = N9644 | data_masked[7372];
  assign N9644 = N9643 | data_masked[7500];
  assign N9643 = N9642 | data_masked[7628];
  assign N9642 = N9641 | data_masked[7756];
  assign N9641 = N9640 | data_masked[7884];
  assign N9640 = N9639 | data_masked[8012];
  assign N9639 = N9638 | data_masked[8140];
  assign N9638 = N9637 | data_masked[8268];
  assign N9637 = N9636 | data_masked[8396];
  assign N9636 = N9635 | data_masked[8524];
  assign N9635 = N9634 | data_masked[8652];
  assign N9634 = N9633 | data_masked[8780];
  assign N9633 = N9632 | data_masked[8908];
  assign N9632 = N9631 | data_masked[9036];
  assign N9631 = N9630 | data_masked[9164];
  assign N9630 = N9629 | data_masked[9292];
  assign N9629 = N9628 | data_masked[9420];
  assign N9628 = N9627 | data_masked[9548];
  assign N9627 = N9626 | data_masked[9676];
  assign N9626 = N9625 | data_masked[9804];
  assign N9625 = N9624 | data_masked[9932];
  assign N9624 = N9623 | data_masked[10060];
  assign N9623 = N9622 | data_masked[10188];
  assign N9622 = N9621 | data_masked[10316];
  assign N9621 = N9620 | data_masked[10444];
  assign N9620 = N9619 | data_masked[10572];
  assign N9619 = N9618 | data_masked[10700];
  assign N9618 = N9617 | data_masked[10828];
  assign N9617 = N9616 | data_masked[10956];
  assign N9616 = N9615 | data_masked[11084];
  assign N9615 = N9614 | data_masked[11212];
  assign N9614 = N9613 | data_masked[11340];
  assign N9613 = N9612 | data_masked[11468];
  assign N9612 = N9611 | data_masked[11596];
  assign N9611 = N9610 | data_masked[11724];
  assign N9610 = N9609 | data_masked[11852];
  assign N9609 = N9608 | data_masked[11980];
  assign N9608 = N9607 | data_masked[12108];
  assign N9607 = N9606 | data_masked[12236];
  assign N9606 = N9605 | data_masked[12364];
  assign N9605 = N9604 | data_masked[12492];
  assign N9604 = N9603 | data_masked[12620];
  assign N9603 = N9602 | data_masked[12748];
  assign N9602 = N9601 | data_masked[12876];
  assign N9601 = N9600 | data_masked[13004];
  assign N9600 = N9599 | data_masked[13132];
  assign N9599 = N9598 | data_masked[13260];
  assign N9598 = N9597 | data_masked[13388];
  assign N9597 = N9596 | data_masked[13516];
  assign N9596 = N9595 | data_masked[13644];
  assign N9595 = N9594 | data_masked[13772];
  assign N9594 = N9593 | data_masked[13900];
  assign N9593 = N9592 | data_masked[14028];
  assign N9592 = N9591 | data_masked[14156];
  assign N9591 = N9590 | data_masked[14284];
  assign N9590 = N9589 | data_masked[14412];
  assign N9589 = N9588 | data_masked[14540];
  assign N9588 = N9587 | data_masked[14668];
  assign N9587 = N9586 | data_masked[14796];
  assign N9586 = N9585 | data_masked[14924];
  assign N9585 = N9584 | data_masked[15052];
  assign N9584 = N9583 | data_masked[15180];
  assign N9583 = N9582 | data_masked[15308];
  assign N9582 = N9581 | data_masked[15436];
  assign N9581 = N9580 | data_masked[15564];
  assign N9580 = N9579 | data_masked[15692];
  assign N9579 = N9578 | data_masked[15820];
  assign N9578 = N9577 | data_masked[15948];
  assign N9577 = N9576 | data_masked[16076];
  assign N9576 = data_masked[16332] | data_masked[16204];
  assign data_o[77] = N9827 | data_masked[77];
  assign N9827 = N9826 | data_masked[205];
  assign N9826 = N9825 | data_masked[333];
  assign N9825 = N9824 | data_masked[461];
  assign N9824 = N9823 | data_masked[589];
  assign N9823 = N9822 | data_masked[717];
  assign N9822 = N9821 | data_masked[845];
  assign N9821 = N9820 | data_masked[973];
  assign N9820 = N9819 | data_masked[1101];
  assign N9819 = N9818 | data_masked[1229];
  assign N9818 = N9817 | data_masked[1357];
  assign N9817 = N9816 | data_masked[1485];
  assign N9816 = N9815 | data_masked[1613];
  assign N9815 = N9814 | data_masked[1741];
  assign N9814 = N9813 | data_masked[1869];
  assign N9813 = N9812 | data_masked[1997];
  assign N9812 = N9811 | data_masked[2125];
  assign N9811 = N9810 | data_masked[2253];
  assign N9810 = N9809 | data_masked[2381];
  assign N9809 = N9808 | data_masked[2509];
  assign N9808 = N9807 | data_masked[2637];
  assign N9807 = N9806 | data_masked[2765];
  assign N9806 = N9805 | data_masked[2893];
  assign N9805 = N9804 | data_masked[3021];
  assign N9804 = N9803 | data_masked[3149];
  assign N9803 = N9802 | data_masked[3277];
  assign N9802 = N9801 | data_masked[3405];
  assign N9801 = N9800 | data_masked[3533];
  assign N9800 = N9799 | data_masked[3661];
  assign N9799 = N9798 | data_masked[3789];
  assign N9798 = N9797 | data_masked[3917];
  assign N9797 = N9796 | data_masked[4045];
  assign N9796 = N9795 | data_masked[4173];
  assign N9795 = N9794 | data_masked[4301];
  assign N9794 = N9793 | data_masked[4429];
  assign N9793 = N9792 | data_masked[4557];
  assign N9792 = N9791 | data_masked[4685];
  assign N9791 = N9790 | data_masked[4813];
  assign N9790 = N9789 | data_masked[4941];
  assign N9789 = N9788 | data_masked[5069];
  assign N9788 = N9787 | data_masked[5197];
  assign N9787 = N9786 | data_masked[5325];
  assign N9786 = N9785 | data_masked[5453];
  assign N9785 = N9784 | data_masked[5581];
  assign N9784 = N9783 | data_masked[5709];
  assign N9783 = N9782 | data_masked[5837];
  assign N9782 = N9781 | data_masked[5965];
  assign N9781 = N9780 | data_masked[6093];
  assign N9780 = N9779 | data_masked[6221];
  assign N9779 = N9778 | data_masked[6349];
  assign N9778 = N9777 | data_masked[6477];
  assign N9777 = N9776 | data_masked[6605];
  assign N9776 = N9775 | data_masked[6733];
  assign N9775 = N9774 | data_masked[6861];
  assign N9774 = N9773 | data_masked[6989];
  assign N9773 = N9772 | data_masked[7117];
  assign N9772 = N9771 | data_masked[7245];
  assign N9771 = N9770 | data_masked[7373];
  assign N9770 = N9769 | data_masked[7501];
  assign N9769 = N9768 | data_masked[7629];
  assign N9768 = N9767 | data_masked[7757];
  assign N9767 = N9766 | data_masked[7885];
  assign N9766 = N9765 | data_masked[8013];
  assign N9765 = N9764 | data_masked[8141];
  assign N9764 = N9763 | data_masked[8269];
  assign N9763 = N9762 | data_masked[8397];
  assign N9762 = N9761 | data_masked[8525];
  assign N9761 = N9760 | data_masked[8653];
  assign N9760 = N9759 | data_masked[8781];
  assign N9759 = N9758 | data_masked[8909];
  assign N9758 = N9757 | data_masked[9037];
  assign N9757 = N9756 | data_masked[9165];
  assign N9756 = N9755 | data_masked[9293];
  assign N9755 = N9754 | data_masked[9421];
  assign N9754 = N9753 | data_masked[9549];
  assign N9753 = N9752 | data_masked[9677];
  assign N9752 = N9751 | data_masked[9805];
  assign N9751 = N9750 | data_masked[9933];
  assign N9750 = N9749 | data_masked[10061];
  assign N9749 = N9748 | data_masked[10189];
  assign N9748 = N9747 | data_masked[10317];
  assign N9747 = N9746 | data_masked[10445];
  assign N9746 = N9745 | data_masked[10573];
  assign N9745 = N9744 | data_masked[10701];
  assign N9744 = N9743 | data_masked[10829];
  assign N9743 = N9742 | data_masked[10957];
  assign N9742 = N9741 | data_masked[11085];
  assign N9741 = N9740 | data_masked[11213];
  assign N9740 = N9739 | data_masked[11341];
  assign N9739 = N9738 | data_masked[11469];
  assign N9738 = N9737 | data_masked[11597];
  assign N9737 = N9736 | data_masked[11725];
  assign N9736 = N9735 | data_masked[11853];
  assign N9735 = N9734 | data_masked[11981];
  assign N9734 = N9733 | data_masked[12109];
  assign N9733 = N9732 | data_masked[12237];
  assign N9732 = N9731 | data_masked[12365];
  assign N9731 = N9730 | data_masked[12493];
  assign N9730 = N9729 | data_masked[12621];
  assign N9729 = N9728 | data_masked[12749];
  assign N9728 = N9727 | data_masked[12877];
  assign N9727 = N9726 | data_masked[13005];
  assign N9726 = N9725 | data_masked[13133];
  assign N9725 = N9724 | data_masked[13261];
  assign N9724 = N9723 | data_masked[13389];
  assign N9723 = N9722 | data_masked[13517];
  assign N9722 = N9721 | data_masked[13645];
  assign N9721 = N9720 | data_masked[13773];
  assign N9720 = N9719 | data_masked[13901];
  assign N9719 = N9718 | data_masked[14029];
  assign N9718 = N9717 | data_masked[14157];
  assign N9717 = N9716 | data_masked[14285];
  assign N9716 = N9715 | data_masked[14413];
  assign N9715 = N9714 | data_masked[14541];
  assign N9714 = N9713 | data_masked[14669];
  assign N9713 = N9712 | data_masked[14797];
  assign N9712 = N9711 | data_masked[14925];
  assign N9711 = N9710 | data_masked[15053];
  assign N9710 = N9709 | data_masked[15181];
  assign N9709 = N9708 | data_masked[15309];
  assign N9708 = N9707 | data_masked[15437];
  assign N9707 = N9706 | data_masked[15565];
  assign N9706 = N9705 | data_masked[15693];
  assign N9705 = N9704 | data_masked[15821];
  assign N9704 = N9703 | data_masked[15949];
  assign N9703 = N9702 | data_masked[16077];
  assign N9702 = data_masked[16333] | data_masked[16205];
  assign data_o[78] = N9953 | data_masked[78];
  assign N9953 = N9952 | data_masked[206];
  assign N9952 = N9951 | data_masked[334];
  assign N9951 = N9950 | data_masked[462];
  assign N9950 = N9949 | data_masked[590];
  assign N9949 = N9948 | data_masked[718];
  assign N9948 = N9947 | data_masked[846];
  assign N9947 = N9946 | data_masked[974];
  assign N9946 = N9945 | data_masked[1102];
  assign N9945 = N9944 | data_masked[1230];
  assign N9944 = N9943 | data_masked[1358];
  assign N9943 = N9942 | data_masked[1486];
  assign N9942 = N9941 | data_masked[1614];
  assign N9941 = N9940 | data_masked[1742];
  assign N9940 = N9939 | data_masked[1870];
  assign N9939 = N9938 | data_masked[1998];
  assign N9938 = N9937 | data_masked[2126];
  assign N9937 = N9936 | data_masked[2254];
  assign N9936 = N9935 | data_masked[2382];
  assign N9935 = N9934 | data_masked[2510];
  assign N9934 = N9933 | data_masked[2638];
  assign N9933 = N9932 | data_masked[2766];
  assign N9932 = N9931 | data_masked[2894];
  assign N9931 = N9930 | data_masked[3022];
  assign N9930 = N9929 | data_masked[3150];
  assign N9929 = N9928 | data_masked[3278];
  assign N9928 = N9927 | data_masked[3406];
  assign N9927 = N9926 | data_masked[3534];
  assign N9926 = N9925 | data_masked[3662];
  assign N9925 = N9924 | data_masked[3790];
  assign N9924 = N9923 | data_masked[3918];
  assign N9923 = N9922 | data_masked[4046];
  assign N9922 = N9921 | data_masked[4174];
  assign N9921 = N9920 | data_masked[4302];
  assign N9920 = N9919 | data_masked[4430];
  assign N9919 = N9918 | data_masked[4558];
  assign N9918 = N9917 | data_masked[4686];
  assign N9917 = N9916 | data_masked[4814];
  assign N9916 = N9915 | data_masked[4942];
  assign N9915 = N9914 | data_masked[5070];
  assign N9914 = N9913 | data_masked[5198];
  assign N9913 = N9912 | data_masked[5326];
  assign N9912 = N9911 | data_masked[5454];
  assign N9911 = N9910 | data_masked[5582];
  assign N9910 = N9909 | data_masked[5710];
  assign N9909 = N9908 | data_masked[5838];
  assign N9908 = N9907 | data_masked[5966];
  assign N9907 = N9906 | data_masked[6094];
  assign N9906 = N9905 | data_masked[6222];
  assign N9905 = N9904 | data_masked[6350];
  assign N9904 = N9903 | data_masked[6478];
  assign N9903 = N9902 | data_masked[6606];
  assign N9902 = N9901 | data_masked[6734];
  assign N9901 = N9900 | data_masked[6862];
  assign N9900 = N9899 | data_masked[6990];
  assign N9899 = N9898 | data_masked[7118];
  assign N9898 = N9897 | data_masked[7246];
  assign N9897 = N9896 | data_masked[7374];
  assign N9896 = N9895 | data_masked[7502];
  assign N9895 = N9894 | data_masked[7630];
  assign N9894 = N9893 | data_masked[7758];
  assign N9893 = N9892 | data_masked[7886];
  assign N9892 = N9891 | data_masked[8014];
  assign N9891 = N9890 | data_masked[8142];
  assign N9890 = N9889 | data_masked[8270];
  assign N9889 = N9888 | data_masked[8398];
  assign N9888 = N9887 | data_masked[8526];
  assign N9887 = N9886 | data_masked[8654];
  assign N9886 = N9885 | data_masked[8782];
  assign N9885 = N9884 | data_masked[8910];
  assign N9884 = N9883 | data_masked[9038];
  assign N9883 = N9882 | data_masked[9166];
  assign N9882 = N9881 | data_masked[9294];
  assign N9881 = N9880 | data_masked[9422];
  assign N9880 = N9879 | data_masked[9550];
  assign N9879 = N9878 | data_masked[9678];
  assign N9878 = N9877 | data_masked[9806];
  assign N9877 = N9876 | data_masked[9934];
  assign N9876 = N9875 | data_masked[10062];
  assign N9875 = N9874 | data_masked[10190];
  assign N9874 = N9873 | data_masked[10318];
  assign N9873 = N9872 | data_masked[10446];
  assign N9872 = N9871 | data_masked[10574];
  assign N9871 = N9870 | data_masked[10702];
  assign N9870 = N9869 | data_masked[10830];
  assign N9869 = N9868 | data_masked[10958];
  assign N9868 = N9867 | data_masked[11086];
  assign N9867 = N9866 | data_masked[11214];
  assign N9866 = N9865 | data_masked[11342];
  assign N9865 = N9864 | data_masked[11470];
  assign N9864 = N9863 | data_masked[11598];
  assign N9863 = N9862 | data_masked[11726];
  assign N9862 = N9861 | data_masked[11854];
  assign N9861 = N9860 | data_masked[11982];
  assign N9860 = N9859 | data_masked[12110];
  assign N9859 = N9858 | data_masked[12238];
  assign N9858 = N9857 | data_masked[12366];
  assign N9857 = N9856 | data_masked[12494];
  assign N9856 = N9855 | data_masked[12622];
  assign N9855 = N9854 | data_masked[12750];
  assign N9854 = N9853 | data_masked[12878];
  assign N9853 = N9852 | data_masked[13006];
  assign N9852 = N9851 | data_masked[13134];
  assign N9851 = N9850 | data_masked[13262];
  assign N9850 = N9849 | data_masked[13390];
  assign N9849 = N9848 | data_masked[13518];
  assign N9848 = N9847 | data_masked[13646];
  assign N9847 = N9846 | data_masked[13774];
  assign N9846 = N9845 | data_masked[13902];
  assign N9845 = N9844 | data_masked[14030];
  assign N9844 = N9843 | data_masked[14158];
  assign N9843 = N9842 | data_masked[14286];
  assign N9842 = N9841 | data_masked[14414];
  assign N9841 = N9840 | data_masked[14542];
  assign N9840 = N9839 | data_masked[14670];
  assign N9839 = N9838 | data_masked[14798];
  assign N9838 = N9837 | data_masked[14926];
  assign N9837 = N9836 | data_masked[15054];
  assign N9836 = N9835 | data_masked[15182];
  assign N9835 = N9834 | data_masked[15310];
  assign N9834 = N9833 | data_masked[15438];
  assign N9833 = N9832 | data_masked[15566];
  assign N9832 = N9831 | data_masked[15694];
  assign N9831 = N9830 | data_masked[15822];
  assign N9830 = N9829 | data_masked[15950];
  assign N9829 = N9828 | data_masked[16078];
  assign N9828 = data_masked[16334] | data_masked[16206];
  assign data_o[79] = N10079 | data_masked[79];
  assign N10079 = N10078 | data_masked[207];
  assign N10078 = N10077 | data_masked[335];
  assign N10077 = N10076 | data_masked[463];
  assign N10076 = N10075 | data_masked[591];
  assign N10075 = N10074 | data_masked[719];
  assign N10074 = N10073 | data_masked[847];
  assign N10073 = N10072 | data_masked[975];
  assign N10072 = N10071 | data_masked[1103];
  assign N10071 = N10070 | data_masked[1231];
  assign N10070 = N10069 | data_masked[1359];
  assign N10069 = N10068 | data_masked[1487];
  assign N10068 = N10067 | data_masked[1615];
  assign N10067 = N10066 | data_masked[1743];
  assign N10066 = N10065 | data_masked[1871];
  assign N10065 = N10064 | data_masked[1999];
  assign N10064 = N10063 | data_masked[2127];
  assign N10063 = N10062 | data_masked[2255];
  assign N10062 = N10061 | data_masked[2383];
  assign N10061 = N10060 | data_masked[2511];
  assign N10060 = N10059 | data_masked[2639];
  assign N10059 = N10058 | data_masked[2767];
  assign N10058 = N10057 | data_masked[2895];
  assign N10057 = N10056 | data_masked[3023];
  assign N10056 = N10055 | data_masked[3151];
  assign N10055 = N10054 | data_masked[3279];
  assign N10054 = N10053 | data_masked[3407];
  assign N10053 = N10052 | data_masked[3535];
  assign N10052 = N10051 | data_masked[3663];
  assign N10051 = N10050 | data_masked[3791];
  assign N10050 = N10049 | data_masked[3919];
  assign N10049 = N10048 | data_masked[4047];
  assign N10048 = N10047 | data_masked[4175];
  assign N10047 = N10046 | data_masked[4303];
  assign N10046 = N10045 | data_masked[4431];
  assign N10045 = N10044 | data_masked[4559];
  assign N10044 = N10043 | data_masked[4687];
  assign N10043 = N10042 | data_masked[4815];
  assign N10042 = N10041 | data_masked[4943];
  assign N10041 = N10040 | data_masked[5071];
  assign N10040 = N10039 | data_masked[5199];
  assign N10039 = N10038 | data_masked[5327];
  assign N10038 = N10037 | data_masked[5455];
  assign N10037 = N10036 | data_masked[5583];
  assign N10036 = N10035 | data_masked[5711];
  assign N10035 = N10034 | data_masked[5839];
  assign N10034 = N10033 | data_masked[5967];
  assign N10033 = N10032 | data_masked[6095];
  assign N10032 = N10031 | data_masked[6223];
  assign N10031 = N10030 | data_masked[6351];
  assign N10030 = N10029 | data_masked[6479];
  assign N10029 = N10028 | data_masked[6607];
  assign N10028 = N10027 | data_masked[6735];
  assign N10027 = N10026 | data_masked[6863];
  assign N10026 = N10025 | data_masked[6991];
  assign N10025 = N10024 | data_masked[7119];
  assign N10024 = N10023 | data_masked[7247];
  assign N10023 = N10022 | data_masked[7375];
  assign N10022 = N10021 | data_masked[7503];
  assign N10021 = N10020 | data_masked[7631];
  assign N10020 = N10019 | data_masked[7759];
  assign N10019 = N10018 | data_masked[7887];
  assign N10018 = N10017 | data_masked[8015];
  assign N10017 = N10016 | data_masked[8143];
  assign N10016 = N10015 | data_masked[8271];
  assign N10015 = N10014 | data_masked[8399];
  assign N10014 = N10013 | data_masked[8527];
  assign N10013 = N10012 | data_masked[8655];
  assign N10012 = N10011 | data_masked[8783];
  assign N10011 = N10010 | data_masked[8911];
  assign N10010 = N10009 | data_masked[9039];
  assign N10009 = N10008 | data_masked[9167];
  assign N10008 = N10007 | data_masked[9295];
  assign N10007 = N10006 | data_masked[9423];
  assign N10006 = N10005 | data_masked[9551];
  assign N10005 = N10004 | data_masked[9679];
  assign N10004 = N10003 | data_masked[9807];
  assign N10003 = N10002 | data_masked[9935];
  assign N10002 = N10001 | data_masked[10063];
  assign N10001 = N10000 | data_masked[10191];
  assign N10000 = N9999 | data_masked[10319];
  assign N9999 = N9998 | data_masked[10447];
  assign N9998 = N9997 | data_masked[10575];
  assign N9997 = N9996 | data_masked[10703];
  assign N9996 = N9995 | data_masked[10831];
  assign N9995 = N9994 | data_masked[10959];
  assign N9994 = N9993 | data_masked[11087];
  assign N9993 = N9992 | data_masked[11215];
  assign N9992 = N9991 | data_masked[11343];
  assign N9991 = N9990 | data_masked[11471];
  assign N9990 = N9989 | data_masked[11599];
  assign N9989 = N9988 | data_masked[11727];
  assign N9988 = N9987 | data_masked[11855];
  assign N9987 = N9986 | data_masked[11983];
  assign N9986 = N9985 | data_masked[12111];
  assign N9985 = N9984 | data_masked[12239];
  assign N9984 = N9983 | data_masked[12367];
  assign N9983 = N9982 | data_masked[12495];
  assign N9982 = N9981 | data_masked[12623];
  assign N9981 = N9980 | data_masked[12751];
  assign N9980 = N9979 | data_masked[12879];
  assign N9979 = N9978 | data_masked[13007];
  assign N9978 = N9977 | data_masked[13135];
  assign N9977 = N9976 | data_masked[13263];
  assign N9976 = N9975 | data_masked[13391];
  assign N9975 = N9974 | data_masked[13519];
  assign N9974 = N9973 | data_masked[13647];
  assign N9973 = N9972 | data_masked[13775];
  assign N9972 = N9971 | data_masked[13903];
  assign N9971 = N9970 | data_masked[14031];
  assign N9970 = N9969 | data_masked[14159];
  assign N9969 = N9968 | data_masked[14287];
  assign N9968 = N9967 | data_masked[14415];
  assign N9967 = N9966 | data_masked[14543];
  assign N9966 = N9965 | data_masked[14671];
  assign N9965 = N9964 | data_masked[14799];
  assign N9964 = N9963 | data_masked[14927];
  assign N9963 = N9962 | data_masked[15055];
  assign N9962 = N9961 | data_masked[15183];
  assign N9961 = N9960 | data_masked[15311];
  assign N9960 = N9959 | data_masked[15439];
  assign N9959 = N9958 | data_masked[15567];
  assign N9958 = N9957 | data_masked[15695];
  assign N9957 = N9956 | data_masked[15823];
  assign N9956 = N9955 | data_masked[15951];
  assign N9955 = N9954 | data_masked[16079];
  assign N9954 = data_masked[16335] | data_masked[16207];
  assign data_o[80] = N10205 | data_masked[80];
  assign N10205 = N10204 | data_masked[208];
  assign N10204 = N10203 | data_masked[336];
  assign N10203 = N10202 | data_masked[464];
  assign N10202 = N10201 | data_masked[592];
  assign N10201 = N10200 | data_masked[720];
  assign N10200 = N10199 | data_masked[848];
  assign N10199 = N10198 | data_masked[976];
  assign N10198 = N10197 | data_masked[1104];
  assign N10197 = N10196 | data_masked[1232];
  assign N10196 = N10195 | data_masked[1360];
  assign N10195 = N10194 | data_masked[1488];
  assign N10194 = N10193 | data_masked[1616];
  assign N10193 = N10192 | data_masked[1744];
  assign N10192 = N10191 | data_masked[1872];
  assign N10191 = N10190 | data_masked[2000];
  assign N10190 = N10189 | data_masked[2128];
  assign N10189 = N10188 | data_masked[2256];
  assign N10188 = N10187 | data_masked[2384];
  assign N10187 = N10186 | data_masked[2512];
  assign N10186 = N10185 | data_masked[2640];
  assign N10185 = N10184 | data_masked[2768];
  assign N10184 = N10183 | data_masked[2896];
  assign N10183 = N10182 | data_masked[3024];
  assign N10182 = N10181 | data_masked[3152];
  assign N10181 = N10180 | data_masked[3280];
  assign N10180 = N10179 | data_masked[3408];
  assign N10179 = N10178 | data_masked[3536];
  assign N10178 = N10177 | data_masked[3664];
  assign N10177 = N10176 | data_masked[3792];
  assign N10176 = N10175 | data_masked[3920];
  assign N10175 = N10174 | data_masked[4048];
  assign N10174 = N10173 | data_masked[4176];
  assign N10173 = N10172 | data_masked[4304];
  assign N10172 = N10171 | data_masked[4432];
  assign N10171 = N10170 | data_masked[4560];
  assign N10170 = N10169 | data_masked[4688];
  assign N10169 = N10168 | data_masked[4816];
  assign N10168 = N10167 | data_masked[4944];
  assign N10167 = N10166 | data_masked[5072];
  assign N10166 = N10165 | data_masked[5200];
  assign N10165 = N10164 | data_masked[5328];
  assign N10164 = N10163 | data_masked[5456];
  assign N10163 = N10162 | data_masked[5584];
  assign N10162 = N10161 | data_masked[5712];
  assign N10161 = N10160 | data_masked[5840];
  assign N10160 = N10159 | data_masked[5968];
  assign N10159 = N10158 | data_masked[6096];
  assign N10158 = N10157 | data_masked[6224];
  assign N10157 = N10156 | data_masked[6352];
  assign N10156 = N10155 | data_masked[6480];
  assign N10155 = N10154 | data_masked[6608];
  assign N10154 = N10153 | data_masked[6736];
  assign N10153 = N10152 | data_masked[6864];
  assign N10152 = N10151 | data_masked[6992];
  assign N10151 = N10150 | data_masked[7120];
  assign N10150 = N10149 | data_masked[7248];
  assign N10149 = N10148 | data_masked[7376];
  assign N10148 = N10147 | data_masked[7504];
  assign N10147 = N10146 | data_masked[7632];
  assign N10146 = N10145 | data_masked[7760];
  assign N10145 = N10144 | data_masked[7888];
  assign N10144 = N10143 | data_masked[8016];
  assign N10143 = N10142 | data_masked[8144];
  assign N10142 = N10141 | data_masked[8272];
  assign N10141 = N10140 | data_masked[8400];
  assign N10140 = N10139 | data_masked[8528];
  assign N10139 = N10138 | data_masked[8656];
  assign N10138 = N10137 | data_masked[8784];
  assign N10137 = N10136 | data_masked[8912];
  assign N10136 = N10135 | data_masked[9040];
  assign N10135 = N10134 | data_masked[9168];
  assign N10134 = N10133 | data_masked[9296];
  assign N10133 = N10132 | data_masked[9424];
  assign N10132 = N10131 | data_masked[9552];
  assign N10131 = N10130 | data_masked[9680];
  assign N10130 = N10129 | data_masked[9808];
  assign N10129 = N10128 | data_masked[9936];
  assign N10128 = N10127 | data_masked[10064];
  assign N10127 = N10126 | data_masked[10192];
  assign N10126 = N10125 | data_masked[10320];
  assign N10125 = N10124 | data_masked[10448];
  assign N10124 = N10123 | data_masked[10576];
  assign N10123 = N10122 | data_masked[10704];
  assign N10122 = N10121 | data_masked[10832];
  assign N10121 = N10120 | data_masked[10960];
  assign N10120 = N10119 | data_masked[11088];
  assign N10119 = N10118 | data_masked[11216];
  assign N10118 = N10117 | data_masked[11344];
  assign N10117 = N10116 | data_masked[11472];
  assign N10116 = N10115 | data_masked[11600];
  assign N10115 = N10114 | data_masked[11728];
  assign N10114 = N10113 | data_masked[11856];
  assign N10113 = N10112 | data_masked[11984];
  assign N10112 = N10111 | data_masked[12112];
  assign N10111 = N10110 | data_masked[12240];
  assign N10110 = N10109 | data_masked[12368];
  assign N10109 = N10108 | data_masked[12496];
  assign N10108 = N10107 | data_masked[12624];
  assign N10107 = N10106 | data_masked[12752];
  assign N10106 = N10105 | data_masked[12880];
  assign N10105 = N10104 | data_masked[13008];
  assign N10104 = N10103 | data_masked[13136];
  assign N10103 = N10102 | data_masked[13264];
  assign N10102 = N10101 | data_masked[13392];
  assign N10101 = N10100 | data_masked[13520];
  assign N10100 = N10099 | data_masked[13648];
  assign N10099 = N10098 | data_masked[13776];
  assign N10098 = N10097 | data_masked[13904];
  assign N10097 = N10096 | data_masked[14032];
  assign N10096 = N10095 | data_masked[14160];
  assign N10095 = N10094 | data_masked[14288];
  assign N10094 = N10093 | data_masked[14416];
  assign N10093 = N10092 | data_masked[14544];
  assign N10092 = N10091 | data_masked[14672];
  assign N10091 = N10090 | data_masked[14800];
  assign N10090 = N10089 | data_masked[14928];
  assign N10089 = N10088 | data_masked[15056];
  assign N10088 = N10087 | data_masked[15184];
  assign N10087 = N10086 | data_masked[15312];
  assign N10086 = N10085 | data_masked[15440];
  assign N10085 = N10084 | data_masked[15568];
  assign N10084 = N10083 | data_masked[15696];
  assign N10083 = N10082 | data_masked[15824];
  assign N10082 = N10081 | data_masked[15952];
  assign N10081 = N10080 | data_masked[16080];
  assign N10080 = data_masked[16336] | data_masked[16208];
  assign data_o[81] = N10331 | data_masked[81];
  assign N10331 = N10330 | data_masked[209];
  assign N10330 = N10329 | data_masked[337];
  assign N10329 = N10328 | data_masked[465];
  assign N10328 = N10327 | data_masked[593];
  assign N10327 = N10326 | data_masked[721];
  assign N10326 = N10325 | data_masked[849];
  assign N10325 = N10324 | data_masked[977];
  assign N10324 = N10323 | data_masked[1105];
  assign N10323 = N10322 | data_masked[1233];
  assign N10322 = N10321 | data_masked[1361];
  assign N10321 = N10320 | data_masked[1489];
  assign N10320 = N10319 | data_masked[1617];
  assign N10319 = N10318 | data_masked[1745];
  assign N10318 = N10317 | data_masked[1873];
  assign N10317 = N10316 | data_masked[2001];
  assign N10316 = N10315 | data_masked[2129];
  assign N10315 = N10314 | data_masked[2257];
  assign N10314 = N10313 | data_masked[2385];
  assign N10313 = N10312 | data_masked[2513];
  assign N10312 = N10311 | data_masked[2641];
  assign N10311 = N10310 | data_masked[2769];
  assign N10310 = N10309 | data_masked[2897];
  assign N10309 = N10308 | data_masked[3025];
  assign N10308 = N10307 | data_masked[3153];
  assign N10307 = N10306 | data_masked[3281];
  assign N10306 = N10305 | data_masked[3409];
  assign N10305 = N10304 | data_masked[3537];
  assign N10304 = N10303 | data_masked[3665];
  assign N10303 = N10302 | data_masked[3793];
  assign N10302 = N10301 | data_masked[3921];
  assign N10301 = N10300 | data_masked[4049];
  assign N10300 = N10299 | data_masked[4177];
  assign N10299 = N10298 | data_masked[4305];
  assign N10298 = N10297 | data_masked[4433];
  assign N10297 = N10296 | data_masked[4561];
  assign N10296 = N10295 | data_masked[4689];
  assign N10295 = N10294 | data_masked[4817];
  assign N10294 = N10293 | data_masked[4945];
  assign N10293 = N10292 | data_masked[5073];
  assign N10292 = N10291 | data_masked[5201];
  assign N10291 = N10290 | data_masked[5329];
  assign N10290 = N10289 | data_masked[5457];
  assign N10289 = N10288 | data_masked[5585];
  assign N10288 = N10287 | data_masked[5713];
  assign N10287 = N10286 | data_masked[5841];
  assign N10286 = N10285 | data_masked[5969];
  assign N10285 = N10284 | data_masked[6097];
  assign N10284 = N10283 | data_masked[6225];
  assign N10283 = N10282 | data_masked[6353];
  assign N10282 = N10281 | data_masked[6481];
  assign N10281 = N10280 | data_masked[6609];
  assign N10280 = N10279 | data_masked[6737];
  assign N10279 = N10278 | data_masked[6865];
  assign N10278 = N10277 | data_masked[6993];
  assign N10277 = N10276 | data_masked[7121];
  assign N10276 = N10275 | data_masked[7249];
  assign N10275 = N10274 | data_masked[7377];
  assign N10274 = N10273 | data_masked[7505];
  assign N10273 = N10272 | data_masked[7633];
  assign N10272 = N10271 | data_masked[7761];
  assign N10271 = N10270 | data_masked[7889];
  assign N10270 = N10269 | data_masked[8017];
  assign N10269 = N10268 | data_masked[8145];
  assign N10268 = N10267 | data_masked[8273];
  assign N10267 = N10266 | data_masked[8401];
  assign N10266 = N10265 | data_masked[8529];
  assign N10265 = N10264 | data_masked[8657];
  assign N10264 = N10263 | data_masked[8785];
  assign N10263 = N10262 | data_masked[8913];
  assign N10262 = N10261 | data_masked[9041];
  assign N10261 = N10260 | data_masked[9169];
  assign N10260 = N10259 | data_masked[9297];
  assign N10259 = N10258 | data_masked[9425];
  assign N10258 = N10257 | data_masked[9553];
  assign N10257 = N10256 | data_masked[9681];
  assign N10256 = N10255 | data_masked[9809];
  assign N10255 = N10254 | data_masked[9937];
  assign N10254 = N10253 | data_masked[10065];
  assign N10253 = N10252 | data_masked[10193];
  assign N10252 = N10251 | data_masked[10321];
  assign N10251 = N10250 | data_masked[10449];
  assign N10250 = N10249 | data_masked[10577];
  assign N10249 = N10248 | data_masked[10705];
  assign N10248 = N10247 | data_masked[10833];
  assign N10247 = N10246 | data_masked[10961];
  assign N10246 = N10245 | data_masked[11089];
  assign N10245 = N10244 | data_masked[11217];
  assign N10244 = N10243 | data_masked[11345];
  assign N10243 = N10242 | data_masked[11473];
  assign N10242 = N10241 | data_masked[11601];
  assign N10241 = N10240 | data_masked[11729];
  assign N10240 = N10239 | data_masked[11857];
  assign N10239 = N10238 | data_masked[11985];
  assign N10238 = N10237 | data_masked[12113];
  assign N10237 = N10236 | data_masked[12241];
  assign N10236 = N10235 | data_masked[12369];
  assign N10235 = N10234 | data_masked[12497];
  assign N10234 = N10233 | data_masked[12625];
  assign N10233 = N10232 | data_masked[12753];
  assign N10232 = N10231 | data_masked[12881];
  assign N10231 = N10230 | data_masked[13009];
  assign N10230 = N10229 | data_masked[13137];
  assign N10229 = N10228 | data_masked[13265];
  assign N10228 = N10227 | data_masked[13393];
  assign N10227 = N10226 | data_masked[13521];
  assign N10226 = N10225 | data_masked[13649];
  assign N10225 = N10224 | data_masked[13777];
  assign N10224 = N10223 | data_masked[13905];
  assign N10223 = N10222 | data_masked[14033];
  assign N10222 = N10221 | data_masked[14161];
  assign N10221 = N10220 | data_masked[14289];
  assign N10220 = N10219 | data_masked[14417];
  assign N10219 = N10218 | data_masked[14545];
  assign N10218 = N10217 | data_masked[14673];
  assign N10217 = N10216 | data_masked[14801];
  assign N10216 = N10215 | data_masked[14929];
  assign N10215 = N10214 | data_masked[15057];
  assign N10214 = N10213 | data_masked[15185];
  assign N10213 = N10212 | data_masked[15313];
  assign N10212 = N10211 | data_masked[15441];
  assign N10211 = N10210 | data_masked[15569];
  assign N10210 = N10209 | data_masked[15697];
  assign N10209 = N10208 | data_masked[15825];
  assign N10208 = N10207 | data_masked[15953];
  assign N10207 = N10206 | data_masked[16081];
  assign N10206 = data_masked[16337] | data_masked[16209];
  assign data_o[82] = N10457 | data_masked[82];
  assign N10457 = N10456 | data_masked[210];
  assign N10456 = N10455 | data_masked[338];
  assign N10455 = N10454 | data_masked[466];
  assign N10454 = N10453 | data_masked[594];
  assign N10453 = N10452 | data_masked[722];
  assign N10452 = N10451 | data_masked[850];
  assign N10451 = N10450 | data_masked[978];
  assign N10450 = N10449 | data_masked[1106];
  assign N10449 = N10448 | data_masked[1234];
  assign N10448 = N10447 | data_masked[1362];
  assign N10447 = N10446 | data_masked[1490];
  assign N10446 = N10445 | data_masked[1618];
  assign N10445 = N10444 | data_masked[1746];
  assign N10444 = N10443 | data_masked[1874];
  assign N10443 = N10442 | data_masked[2002];
  assign N10442 = N10441 | data_masked[2130];
  assign N10441 = N10440 | data_masked[2258];
  assign N10440 = N10439 | data_masked[2386];
  assign N10439 = N10438 | data_masked[2514];
  assign N10438 = N10437 | data_masked[2642];
  assign N10437 = N10436 | data_masked[2770];
  assign N10436 = N10435 | data_masked[2898];
  assign N10435 = N10434 | data_masked[3026];
  assign N10434 = N10433 | data_masked[3154];
  assign N10433 = N10432 | data_masked[3282];
  assign N10432 = N10431 | data_masked[3410];
  assign N10431 = N10430 | data_masked[3538];
  assign N10430 = N10429 | data_masked[3666];
  assign N10429 = N10428 | data_masked[3794];
  assign N10428 = N10427 | data_masked[3922];
  assign N10427 = N10426 | data_masked[4050];
  assign N10426 = N10425 | data_masked[4178];
  assign N10425 = N10424 | data_masked[4306];
  assign N10424 = N10423 | data_masked[4434];
  assign N10423 = N10422 | data_masked[4562];
  assign N10422 = N10421 | data_masked[4690];
  assign N10421 = N10420 | data_masked[4818];
  assign N10420 = N10419 | data_masked[4946];
  assign N10419 = N10418 | data_masked[5074];
  assign N10418 = N10417 | data_masked[5202];
  assign N10417 = N10416 | data_masked[5330];
  assign N10416 = N10415 | data_masked[5458];
  assign N10415 = N10414 | data_masked[5586];
  assign N10414 = N10413 | data_masked[5714];
  assign N10413 = N10412 | data_masked[5842];
  assign N10412 = N10411 | data_masked[5970];
  assign N10411 = N10410 | data_masked[6098];
  assign N10410 = N10409 | data_masked[6226];
  assign N10409 = N10408 | data_masked[6354];
  assign N10408 = N10407 | data_masked[6482];
  assign N10407 = N10406 | data_masked[6610];
  assign N10406 = N10405 | data_masked[6738];
  assign N10405 = N10404 | data_masked[6866];
  assign N10404 = N10403 | data_masked[6994];
  assign N10403 = N10402 | data_masked[7122];
  assign N10402 = N10401 | data_masked[7250];
  assign N10401 = N10400 | data_masked[7378];
  assign N10400 = N10399 | data_masked[7506];
  assign N10399 = N10398 | data_masked[7634];
  assign N10398 = N10397 | data_masked[7762];
  assign N10397 = N10396 | data_masked[7890];
  assign N10396 = N10395 | data_masked[8018];
  assign N10395 = N10394 | data_masked[8146];
  assign N10394 = N10393 | data_masked[8274];
  assign N10393 = N10392 | data_masked[8402];
  assign N10392 = N10391 | data_masked[8530];
  assign N10391 = N10390 | data_masked[8658];
  assign N10390 = N10389 | data_masked[8786];
  assign N10389 = N10388 | data_masked[8914];
  assign N10388 = N10387 | data_masked[9042];
  assign N10387 = N10386 | data_masked[9170];
  assign N10386 = N10385 | data_masked[9298];
  assign N10385 = N10384 | data_masked[9426];
  assign N10384 = N10383 | data_masked[9554];
  assign N10383 = N10382 | data_masked[9682];
  assign N10382 = N10381 | data_masked[9810];
  assign N10381 = N10380 | data_masked[9938];
  assign N10380 = N10379 | data_masked[10066];
  assign N10379 = N10378 | data_masked[10194];
  assign N10378 = N10377 | data_masked[10322];
  assign N10377 = N10376 | data_masked[10450];
  assign N10376 = N10375 | data_masked[10578];
  assign N10375 = N10374 | data_masked[10706];
  assign N10374 = N10373 | data_masked[10834];
  assign N10373 = N10372 | data_masked[10962];
  assign N10372 = N10371 | data_masked[11090];
  assign N10371 = N10370 | data_masked[11218];
  assign N10370 = N10369 | data_masked[11346];
  assign N10369 = N10368 | data_masked[11474];
  assign N10368 = N10367 | data_masked[11602];
  assign N10367 = N10366 | data_masked[11730];
  assign N10366 = N10365 | data_masked[11858];
  assign N10365 = N10364 | data_masked[11986];
  assign N10364 = N10363 | data_masked[12114];
  assign N10363 = N10362 | data_masked[12242];
  assign N10362 = N10361 | data_masked[12370];
  assign N10361 = N10360 | data_masked[12498];
  assign N10360 = N10359 | data_masked[12626];
  assign N10359 = N10358 | data_masked[12754];
  assign N10358 = N10357 | data_masked[12882];
  assign N10357 = N10356 | data_masked[13010];
  assign N10356 = N10355 | data_masked[13138];
  assign N10355 = N10354 | data_masked[13266];
  assign N10354 = N10353 | data_masked[13394];
  assign N10353 = N10352 | data_masked[13522];
  assign N10352 = N10351 | data_masked[13650];
  assign N10351 = N10350 | data_masked[13778];
  assign N10350 = N10349 | data_masked[13906];
  assign N10349 = N10348 | data_masked[14034];
  assign N10348 = N10347 | data_masked[14162];
  assign N10347 = N10346 | data_masked[14290];
  assign N10346 = N10345 | data_masked[14418];
  assign N10345 = N10344 | data_masked[14546];
  assign N10344 = N10343 | data_masked[14674];
  assign N10343 = N10342 | data_masked[14802];
  assign N10342 = N10341 | data_masked[14930];
  assign N10341 = N10340 | data_masked[15058];
  assign N10340 = N10339 | data_masked[15186];
  assign N10339 = N10338 | data_masked[15314];
  assign N10338 = N10337 | data_masked[15442];
  assign N10337 = N10336 | data_masked[15570];
  assign N10336 = N10335 | data_masked[15698];
  assign N10335 = N10334 | data_masked[15826];
  assign N10334 = N10333 | data_masked[15954];
  assign N10333 = N10332 | data_masked[16082];
  assign N10332 = data_masked[16338] | data_masked[16210];
  assign data_o[83] = N10583 | data_masked[83];
  assign N10583 = N10582 | data_masked[211];
  assign N10582 = N10581 | data_masked[339];
  assign N10581 = N10580 | data_masked[467];
  assign N10580 = N10579 | data_masked[595];
  assign N10579 = N10578 | data_masked[723];
  assign N10578 = N10577 | data_masked[851];
  assign N10577 = N10576 | data_masked[979];
  assign N10576 = N10575 | data_masked[1107];
  assign N10575 = N10574 | data_masked[1235];
  assign N10574 = N10573 | data_masked[1363];
  assign N10573 = N10572 | data_masked[1491];
  assign N10572 = N10571 | data_masked[1619];
  assign N10571 = N10570 | data_masked[1747];
  assign N10570 = N10569 | data_masked[1875];
  assign N10569 = N10568 | data_masked[2003];
  assign N10568 = N10567 | data_masked[2131];
  assign N10567 = N10566 | data_masked[2259];
  assign N10566 = N10565 | data_masked[2387];
  assign N10565 = N10564 | data_masked[2515];
  assign N10564 = N10563 | data_masked[2643];
  assign N10563 = N10562 | data_masked[2771];
  assign N10562 = N10561 | data_masked[2899];
  assign N10561 = N10560 | data_masked[3027];
  assign N10560 = N10559 | data_masked[3155];
  assign N10559 = N10558 | data_masked[3283];
  assign N10558 = N10557 | data_masked[3411];
  assign N10557 = N10556 | data_masked[3539];
  assign N10556 = N10555 | data_masked[3667];
  assign N10555 = N10554 | data_masked[3795];
  assign N10554 = N10553 | data_masked[3923];
  assign N10553 = N10552 | data_masked[4051];
  assign N10552 = N10551 | data_masked[4179];
  assign N10551 = N10550 | data_masked[4307];
  assign N10550 = N10549 | data_masked[4435];
  assign N10549 = N10548 | data_masked[4563];
  assign N10548 = N10547 | data_masked[4691];
  assign N10547 = N10546 | data_masked[4819];
  assign N10546 = N10545 | data_masked[4947];
  assign N10545 = N10544 | data_masked[5075];
  assign N10544 = N10543 | data_masked[5203];
  assign N10543 = N10542 | data_masked[5331];
  assign N10542 = N10541 | data_masked[5459];
  assign N10541 = N10540 | data_masked[5587];
  assign N10540 = N10539 | data_masked[5715];
  assign N10539 = N10538 | data_masked[5843];
  assign N10538 = N10537 | data_masked[5971];
  assign N10537 = N10536 | data_masked[6099];
  assign N10536 = N10535 | data_masked[6227];
  assign N10535 = N10534 | data_masked[6355];
  assign N10534 = N10533 | data_masked[6483];
  assign N10533 = N10532 | data_masked[6611];
  assign N10532 = N10531 | data_masked[6739];
  assign N10531 = N10530 | data_masked[6867];
  assign N10530 = N10529 | data_masked[6995];
  assign N10529 = N10528 | data_masked[7123];
  assign N10528 = N10527 | data_masked[7251];
  assign N10527 = N10526 | data_masked[7379];
  assign N10526 = N10525 | data_masked[7507];
  assign N10525 = N10524 | data_masked[7635];
  assign N10524 = N10523 | data_masked[7763];
  assign N10523 = N10522 | data_masked[7891];
  assign N10522 = N10521 | data_masked[8019];
  assign N10521 = N10520 | data_masked[8147];
  assign N10520 = N10519 | data_masked[8275];
  assign N10519 = N10518 | data_masked[8403];
  assign N10518 = N10517 | data_masked[8531];
  assign N10517 = N10516 | data_masked[8659];
  assign N10516 = N10515 | data_masked[8787];
  assign N10515 = N10514 | data_masked[8915];
  assign N10514 = N10513 | data_masked[9043];
  assign N10513 = N10512 | data_masked[9171];
  assign N10512 = N10511 | data_masked[9299];
  assign N10511 = N10510 | data_masked[9427];
  assign N10510 = N10509 | data_masked[9555];
  assign N10509 = N10508 | data_masked[9683];
  assign N10508 = N10507 | data_masked[9811];
  assign N10507 = N10506 | data_masked[9939];
  assign N10506 = N10505 | data_masked[10067];
  assign N10505 = N10504 | data_masked[10195];
  assign N10504 = N10503 | data_masked[10323];
  assign N10503 = N10502 | data_masked[10451];
  assign N10502 = N10501 | data_masked[10579];
  assign N10501 = N10500 | data_masked[10707];
  assign N10500 = N10499 | data_masked[10835];
  assign N10499 = N10498 | data_masked[10963];
  assign N10498 = N10497 | data_masked[11091];
  assign N10497 = N10496 | data_masked[11219];
  assign N10496 = N10495 | data_masked[11347];
  assign N10495 = N10494 | data_masked[11475];
  assign N10494 = N10493 | data_masked[11603];
  assign N10493 = N10492 | data_masked[11731];
  assign N10492 = N10491 | data_masked[11859];
  assign N10491 = N10490 | data_masked[11987];
  assign N10490 = N10489 | data_masked[12115];
  assign N10489 = N10488 | data_masked[12243];
  assign N10488 = N10487 | data_masked[12371];
  assign N10487 = N10486 | data_masked[12499];
  assign N10486 = N10485 | data_masked[12627];
  assign N10485 = N10484 | data_masked[12755];
  assign N10484 = N10483 | data_masked[12883];
  assign N10483 = N10482 | data_masked[13011];
  assign N10482 = N10481 | data_masked[13139];
  assign N10481 = N10480 | data_masked[13267];
  assign N10480 = N10479 | data_masked[13395];
  assign N10479 = N10478 | data_masked[13523];
  assign N10478 = N10477 | data_masked[13651];
  assign N10477 = N10476 | data_masked[13779];
  assign N10476 = N10475 | data_masked[13907];
  assign N10475 = N10474 | data_masked[14035];
  assign N10474 = N10473 | data_masked[14163];
  assign N10473 = N10472 | data_masked[14291];
  assign N10472 = N10471 | data_masked[14419];
  assign N10471 = N10470 | data_masked[14547];
  assign N10470 = N10469 | data_masked[14675];
  assign N10469 = N10468 | data_masked[14803];
  assign N10468 = N10467 | data_masked[14931];
  assign N10467 = N10466 | data_masked[15059];
  assign N10466 = N10465 | data_masked[15187];
  assign N10465 = N10464 | data_masked[15315];
  assign N10464 = N10463 | data_masked[15443];
  assign N10463 = N10462 | data_masked[15571];
  assign N10462 = N10461 | data_masked[15699];
  assign N10461 = N10460 | data_masked[15827];
  assign N10460 = N10459 | data_masked[15955];
  assign N10459 = N10458 | data_masked[16083];
  assign N10458 = data_masked[16339] | data_masked[16211];
  assign data_o[84] = N10709 | data_masked[84];
  assign N10709 = N10708 | data_masked[212];
  assign N10708 = N10707 | data_masked[340];
  assign N10707 = N10706 | data_masked[468];
  assign N10706 = N10705 | data_masked[596];
  assign N10705 = N10704 | data_masked[724];
  assign N10704 = N10703 | data_masked[852];
  assign N10703 = N10702 | data_masked[980];
  assign N10702 = N10701 | data_masked[1108];
  assign N10701 = N10700 | data_masked[1236];
  assign N10700 = N10699 | data_masked[1364];
  assign N10699 = N10698 | data_masked[1492];
  assign N10698 = N10697 | data_masked[1620];
  assign N10697 = N10696 | data_masked[1748];
  assign N10696 = N10695 | data_masked[1876];
  assign N10695 = N10694 | data_masked[2004];
  assign N10694 = N10693 | data_masked[2132];
  assign N10693 = N10692 | data_masked[2260];
  assign N10692 = N10691 | data_masked[2388];
  assign N10691 = N10690 | data_masked[2516];
  assign N10690 = N10689 | data_masked[2644];
  assign N10689 = N10688 | data_masked[2772];
  assign N10688 = N10687 | data_masked[2900];
  assign N10687 = N10686 | data_masked[3028];
  assign N10686 = N10685 | data_masked[3156];
  assign N10685 = N10684 | data_masked[3284];
  assign N10684 = N10683 | data_masked[3412];
  assign N10683 = N10682 | data_masked[3540];
  assign N10682 = N10681 | data_masked[3668];
  assign N10681 = N10680 | data_masked[3796];
  assign N10680 = N10679 | data_masked[3924];
  assign N10679 = N10678 | data_masked[4052];
  assign N10678 = N10677 | data_masked[4180];
  assign N10677 = N10676 | data_masked[4308];
  assign N10676 = N10675 | data_masked[4436];
  assign N10675 = N10674 | data_masked[4564];
  assign N10674 = N10673 | data_masked[4692];
  assign N10673 = N10672 | data_masked[4820];
  assign N10672 = N10671 | data_masked[4948];
  assign N10671 = N10670 | data_masked[5076];
  assign N10670 = N10669 | data_masked[5204];
  assign N10669 = N10668 | data_masked[5332];
  assign N10668 = N10667 | data_masked[5460];
  assign N10667 = N10666 | data_masked[5588];
  assign N10666 = N10665 | data_masked[5716];
  assign N10665 = N10664 | data_masked[5844];
  assign N10664 = N10663 | data_masked[5972];
  assign N10663 = N10662 | data_masked[6100];
  assign N10662 = N10661 | data_masked[6228];
  assign N10661 = N10660 | data_masked[6356];
  assign N10660 = N10659 | data_masked[6484];
  assign N10659 = N10658 | data_masked[6612];
  assign N10658 = N10657 | data_masked[6740];
  assign N10657 = N10656 | data_masked[6868];
  assign N10656 = N10655 | data_masked[6996];
  assign N10655 = N10654 | data_masked[7124];
  assign N10654 = N10653 | data_masked[7252];
  assign N10653 = N10652 | data_masked[7380];
  assign N10652 = N10651 | data_masked[7508];
  assign N10651 = N10650 | data_masked[7636];
  assign N10650 = N10649 | data_masked[7764];
  assign N10649 = N10648 | data_masked[7892];
  assign N10648 = N10647 | data_masked[8020];
  assign N10647 = N10646 | data_masked[8148];
  assign N10646 = N10645 | data_masked[8276];
  assign N10645 = N10644 | data_masked[8404];
  assign N10644 = N10643 | data_masked[8532];
  assign N10643 = N10642 | data_masked[8660];
  assign N10642 = N10641 | data_masked[8788];
  assign N10641 = N10640 | data_masked[8916];
  assign N10640 = N10639 | data_masked[9044];
  assign N10639 = N10638 | data_masked[9172];
  assign N10638 = N10637 | data_masked[9300];
  assign N10637 = N10636 | data_masked[9428];
  assign N10636 = N10635 | data_masked[9556];
  assign N10635 = N10634 | data_masked[9684];
  assign N10634 = N10633 | data_masked[9812];
  assign N10633 = N10632 | data_masked[9940];
  assign N10632 = N10631 | data_masked[10068];
  assign N10631 = N10630 | data_masked[10196];
  assign N10630 = N10629 | data_masked[10324];
  assign N10629 = N10628 | data_masked[10452];
  assign N10628 = N10627 | data_masked[10580];
  assign N10627 = N10626 | data_masked[10708];
  assign N10626 = N10625 | data_masked[10836];
  assign N10625 = N10624 | data_masked[10964];
  assign N10624 = N10623 | data_masked[11092];
  assign N10623 = N10622 | data_masked[11220];
  assign N10622 = N10621 | data_masked[11348];
  assign N10621 = N10620 | data_masked[11476];
  assign N10620 = N10619 | data_masked[11604];
  assign N10619 = N10618 | data_masked[11732];
  assign N10618 = N10617 | data_masked[11860];
  assign N10617 = N10616 | data_masked[11988];
  assign N10616 = N10615 | data_masked[12116];
  assign N10615 = N10614 | data_masked[12244];
  assign N10614 = N10613 | data_masked[12372];
  assign N10613 = N10612 | data_masked[12500];
  assign N10612 = N10611 | data_masked[12628];
  assign N10611 = N10610 | data_masked[12756];
  assign N10610 = N10609 | data_masked[12884];
  assign N10609 = N10608 | data_masked[13012];
  assign N10608 = N10607 | data_masked[13140];
  assign N10607 = N10606 | data_masked[13268];
  assign N10606 = N10605 | data_masked[13396];
  assign N10605 = N10604 | data_masked[13524];
  assign N10604 = N10603 | data_masked[13652];
  assign N10603 = N10602 | data_masked[13780];
  assign N10602 = N10601 | data_masked[13908];
  assign N10601 = N10600 | data_masked[14036];
  assign N10600 = N10599 | data_masked[14164];
  assign N10599 = N10598 | data_masked[14292];
  assign N10598 = N10597 | data_masked[14420];
  assign N10597 = N10596 | data_masked[14548];
  assign N10596 = N10595 | data_masked[14676];
  assign N10595 = N10594 | data_masked[14804];
  assign N10594 = N10593 | data_masked[14932];
  assign N10593 = N10592 | data_masked[15060];
  assign N10592 = N10591 | data_masked[15188];
  assign N10591 = N10590 | data_masked[15316];
  assign N10590 = N10589 | data_masked[15444];
  assign N10589 = N10588 | data_masked[15572];
  assign N10588 = N10587 | data_masked[15700];
  assign N10587 = N10586 | data_masked[15828];
  assign N10586 = N10585 | data_masked[15956];
  assign N10585 = N10584 | data_masked[16084];
  assign N10584 = data_masked[16340] | data_masked[16212];
  assign data_o[85] = N10835 | data_masked[85];
  assign N10835 = N10834 | data_masked[213];
  assign N10834 = N10833 | data_masked[341];
  assign N10833 = N10832 | data_masked[469];
  assign N10832 = N10831 | data_masked[597];
  assign N10831 = N10830 | data_masked[725];
  assign N10830 = N10829 | data_masked[853];
  assign N10829 = N10828 | data_masked[981];
  assign N10828 = N10827 | data_masked[1109];
  assign N10827 = N10826 | data_masked[1237];
  assign N10826 = N10825 | data_masked[1365];
  assign N10825 = N10824 | data_masked[1493];
  assign N10824 = N10823 | data_masked[1621];
  assign N10823 = N10822 | data_masked[1749];
  assign N10822 = N10821 | data_masked[1877];
  assign N10821 = N10820 | data_masked[2005];
  assign N10820 = N10819 | data_masked[2133];
  assign N10819 = N10818 | data_masked[2261];
  assign N10818 = N10817 | data_masked[2389];
  assign N10817 = N10816 | data_masked[2517];
  assign N10816 = N10815 | data_masked[2645];
  assign N10815 = N10814 | data_masked[2773];
  assign N10814 = N10813 | data_masked[2901];
  assign N10813 = N10812 | data_masked[3029];
  assign N10812 = N10811 | data_masked[3157];
  assign N10811 = N10810 | data_masked[3285];
  assign N10810 = N10809 | data_masked[3413];
  assign N10809 = N10808 | data_masked[3541];
  assign N10808 = N10807 | data_masked[3669];
  assign N10807 = N10806 | data_masked[3797];
  assign N10806 = N10805 | data_masked[3925];
  assign N10805 = N10804 | data_masked[4053];
  assign N10804 = N10803 | data_masked[4181];
  assign N10803 = N10802 | data_masked[4309];
  assign N10802 = N10801 | data_masked[4437];
  assign N10801 = N10800 | data_masked[4565];
  assign N10800 = N10799 | data_masked[4693];
  assign N10799 = N10798 | data_masked[4821];
  assign N10798 = N10797 | data_masked[4949];
  assign N10797 = N10796 | data_masked[5077];
  assign N10796 = N10795 | data_masked[5205];
  assign N10795 = N10794 | data_masked[5333];
  assign N10794 = N10793 | data_masked[5461];
  assign N10793 = N10792 | data_masked[5589];
  assign N10792 = N10791 | data_masked[5717];
  assign N10791 = N10790 | data_masked[5845];
  assign N10790 = N10789 | data_masked[5973];
  assign N10789 = N10788 | data_masked[6101];
  assign N10788 = N10787 | data_masked[6229];
  assign N10787 = N10786 | data_masked[6357];
  assign N10786 = N10785 | data_masked[6485];
  assign N10785 = N10784 | data_masked[6613];
  assign N10784 = N10783 | data_masked[6741];
  assign N10783 = N10782 | data_masked[6869];
  assign N10782 = N10781 | data_masked[6997];
  assign N10781 = N10780 | data_masked[7125];
  assign N10780 = N10779 | data_masked[7253];
  assign N10779 = N10778 | data_masked[7381];
  assign N10778 = N10777 | data_masked[7509];
  assign N10777 = N10776 | data_masked[7637];
  assign N10776 = N10775 | data_masked[7765];
  assign N10775 = N10774 | data_masked[7893];
  assign N10774 = N10773 | data_masked[8021];
  assign N10773 = N10772 | data_masked[8149];
  assign N10772 = N10771 | data_masked[8277];
  assign N10771 = N10770 | data_masked[8405];
  assign N10770 = N10769 | data_masked[8533];
  assign N10769 = N10768 | data_masked[8661];
  assign N10768 = N10767 | data_masked[8789];
  assign N10767 = N10766 | data_masked[8917];
  assign N10766 = N10765 | data_masked[9045];
  assign N10765 = N10764 | data_masked[9173];
  assign N10764 = N10763 | data_masked[9301];
  assign N10763 = N10762 | data_masked[9429];
  assign N10762 = N10761 | data_masked[9557];
  assign N10761 = N10760 | data_masked[9685];
  assign N10760 = N10759 | data_masked[9813];
  assign N10759 = N10758 | data_masked[9941];
  assign N10758 = N10757 | data_masked[10069];
  assign N10757 = N10756 | data_masked[10197];
  assign N10756 = N10755 | data_masked[10325];
  assign N10755 = N10754 | data_masked[10453];
  assign N10754 = N10753 | data_masked[10581];
  assign N10753 = N10752 | data_masked[10709];
  assign N10752 = N10751 | data_masked[10837];
  assign N10751 = N10750 | data_masked[10965];
  assign N10750 = N10749 | data_masked[11093];
  assign N10749 = N10748 | data_masked[11221];
  assign N10748 = N10747 | data_masked[11349];
  assign N10747 = N10746 | data_masked[11477];
  assign N10746 = N10745 | data_masked[11605];
  assign N10745 = N10744 | data_masked[11733];
  assign N10744 = N10743 | data_masked[11861];
  assign N10743 = N10742 | data_masked[11989];
  assign N10742 = N10741 | data_masked[12117];
  assign N10741 = N10740 | data_masked[12245];
  assign N10740 = N10739 | data_masked[12373];
  assign N10739 = N10738 | data_masked[12501];
  assign N10738 = N10737 | data_masked[12629];
  assign N10737 = N10736 | data_masked[12757];
  assign N10736 = N10735 | data_masked[12885];
  assign N10735 = N10734 | data_masked[13013];
  assign N10734 = N10733 | data_masked[13141];
  assign N10733 = N10732 | data_masked[13269];
  assign N10732 = N10731 | data_masked[13397];
  assign N10731 = N10730 | data_masked[13525];
  assign N10730 = N10729 | data_masked[13653];
  assign N10729 = N10728 | data_masked[13781];
  assign N10728 = N10727 | data_masked[13909];
  assign N10727 = N10726 | data_masked[14037];
  assign N10726 = N10725 | data_masked[14165];
  assign N10725 = N10724 | data_masked[14293];
  assign N10724 = N10723 | data_masked[14421];
  assign N10723 = N10722 | data_masked[14549];
  assign N10722 = N10721 | data_masked[14677];
  assign N10721 = N10720 | data_masked[14805];
  assign N10720 = N10719 | data_masked[14933];
  assign N10719 = N10718 | data_masked[15061];
  assign N10718 = N10717 | data_masked[15189];
  assign N10717 = N10716 | data_masked[15317];
  assign N10716 = N10715 | data_masked[15445];
  assign N10715 = N10714 | data_masked[15573];
  assign N10714 = N10713 | data_masked[15701];
  assign N10713 = N10712 | data_masked[15829];
  assign N10712 = N10711 | data_masked[15957];
  assign N10711 = N10710 | data_masked[16085];
  assign N10710 = data_masked[16341] | data_masked[16213];
  assign data_o[86] = N10961 | data_masked[86];
  assign N10961 = N10960 | data_masked[214];
  assign N10960 = N10959 | data_masked[342];
  assign N10959 = N10958 | data_masked[470];
  assign N10958 = N10957 | data_masked[598];
  assign N10957 = N10956 | data_masked[726];
  assign N10956 = N10955 | data_masked[854];
  assign N10955 = N10954 | data_masked[982];
  assign N10954 = N10953 | data_masked[1110];
  assign N10953 = N10952 | data_masked[1238];
  assign N10952 = N10951 | data_masked[1366];
  assign N10951 = N10950 | data_masked[1494];
  assign N10950 = N10949 | data_masked[1622];
  assign N10949 = N10948 | data_masked[1750];
  assign N10948 = N10947 | data_masked[1878];
  assign N10947 = N10946 | data_masked[2006];
  assign N10946 = N10945 | data_masked[2134];
  assign N10945 = N10944 | data_masked[2262];
  assign N10944 = N10943 | data_masked[2390];
  assign N10943 = N10942 | data_masked[2518];
  assign N10942 = N10941 | data_masked[2646];
  assign N10941 = N10940 | data_masked[2774];
  assign N10940 = N10939 | data_masked[2902];
  assign N10939 = N10938 | data_masked[3030];
  assign N10938 = N10937 | data_masked[3158];
  assign N10937 = N10936 | data_masked[3286];
  assign N10936 = N10935 | data_masked[3414];
  assign N10935 = N10934 | data_masked[3542];
  assign N10934 = N10933 | data_masked[3670];
  assign N10933 = N10932 | data_masked[3798];
  assign N10932 = N10931 | data_masked[3926];
  assign N10931 = N10930 | data_masked[4054];
  assign N10930 = N10929 | data_masked[4182];
  assign N10929 = N10928 | data_masked[4310];
  assign N10928 = N10927 | data_masked[4438];
  assign N10927 = N10926 | data_masked[4566];
  assign N10926 = N10925 | data_masked[4694];
  assign N10925 = N10924 | data_masked[4822];
  assign N10924 = N10923 | data_masked[4950];
  assign N10923 = N10922 | data_masked[5078];
  assign N10922 = N10921 | data_masked[5206];
  assign N10921 = N10920 | data_masked[5334];
  assign N10920 = N10919 | data_masked[5462];
  assign N10919 = N10918 | data_masked[5590];
  assign N10918 = N10917 | data_masked[5718];
  assign N10917 = N10916 | data_masked[5846];
  assign N10916 = N10915 | data_masked[5974];
  assign N10915 = N10914 | data_masked[6102];
  assign N10914 = N10913 | data_masked[6230];
  assign N10913 = N10912 | data_masked[6358];
  assign N10912 = N10911 | data_masked[6486];
  assign N10911 = N10910 | data_masked[6614];
  assign N10910 = N10909 | data_masked[6742];
  assign N10909 = N10908 | data_masked[6870];
  assign N10908 = N10907 | data_masked[6998];
  assign N10907 = N10906 | data_masked[7126];
  assign N10906 = N10905 | data_masked[7254];
  assign N10905 = N10904 | data_masked[7382];
  assign N10904 = N10903 | data_masked[7510];
  assign N10903 = N10902 | data_masked[7638];
  assign N10902 = N10901 | data_masked[7766];
  assign N10901 = N10900 | data_masked[7894];
  assign N10900 = N10899 | data_masked[8022];
  assign N10899 = N10898 | data_masked[8150];
  assign N10898 = N10897 | data_masked[8278];
  assign N10897 = N10896 | data_masked[8406];
  assign N10896 = N10895 | data_masked[8534];
  assign N10895 = N10894 | data_masked[8662];
  assign N10894 = N10893 | data_masked[8790];
  assign N10893 = N10892 | data_masked[8918];
  assign N10892 = N10891 | data_masked[9046];
  assign N10891 = N10890 | data_masked[9174];
  assign N10890 = N10889 | data_masked[9302];
  assign N10889 = N10888 | data_masked[9430];
  assign N10888 = N10887 | data_masked[9558];
  assign N10887 = N10886 | data_masked[9686];
  assign N10886 = N10885 | data_masked[9814];
  assign N10885 = N10884 | data_masked[9942];
  assign N10884 = N10883 | data_masked[10070];
  assign N10883 = N10882 | data_masked[10198];
  assign N10882 = N10881 | data_masked[10326];
  assign N10881 = N10880 | data_masked[10454];
  assign N10880 = N10879 | data_masked[10582];
  assign N10879 = N10878 | data_masked[10710];
  assign N10878 = N10877 | data_masked[10838];
  assign N10877 = N10876 | data_masked[10966];
  assign N10876 = N10875 | data_masked[11094];
  assign N10875 = N10874 | data_masked[11222];
  assign N10874 = N10873 | data_masked[11350];
  assign N10873 = N10872 | data_masked[11478];
  assign N10872 = N10871 | data_masked[11606];
  assign N10871 = N10870 | data_masked[11734];
  assign N10870 = N10869 | data_masked[11862];
  assign N10869 = N10868 | data_masked[11990];
  assign N10868 = N10867 | data_masked[12118];
  assign N10867 = N10866 | data_masked[12246];
  assign N10866 = N10865 | data_masked[12374];
  assign N10865 = N10864 | data_masked[12502];
  assign N10864 = N10863 | data_masked[12630];
  assign N10863 = N10862 | data_masked[12758];
  assign N10862 = N10861 | data_masked[12886];
  assign N10861 = N10860 | data_masked[13014];
  assign N10860 = N10859 | data_masked[13142];
  assign N10859 = N10858 | data_masked[13270];
  assign N10858 = N10857 | data_masked[13398];
  assign N10857 = N10856 | data_masked[13526];
  assign N10856 = N10855 | data_masked[13654];
  assign N10855 = N10854 | data_masked[13782];
  assign N10854 = N10853 | data_masked[13910];
  assign N10853 = N10852 | data_masked[14038];
  assign N10852 = N10851 | data_masked[14166];
  assign N10851 = N10850 | data_masked[14294];
  assign N10850 = N10849 | data_masked[14422];
  assign N10849 = N10848 | data_masked[14550];
  assign N10848 = N10847 | data_masked[14678];
  assign N10847 = N10846 | data_masked[14806];
  assign N10846 = N10845 | data_masked[14934];
  assign N10845 = N10844 | data_masked[15062];
  assign N10844 = N10843 | data_masked[15190];
  assign N10843 = N10842 | data_masked[15318];
  assign N10842 = N10841 | data_masked[15446];
  assign N10841 = N10840 | data_masked[15574];
  assign N10840 = N10839 | data_masked[15702];
  assign N10839 = N10838 | data_masked[15830];
  assign N10838 = N10837 | data_masked[15958];
  assign N10837 = N10836 | data_masked[16086];
  assign N10836 = data_masked[16342] | data_masked[16214];
  assign data_o[87] = N11087 | data_masked[87];
  assign N11087 = N11086 | data_masked[215];
  assign N11086 = N11085 | data_masked[343];
  assign N11085 = N11084 | data_masked[471];
  assign N11084 = N11083 | data_masked[599];
  assign N11083 = N11082 | data_masked[727];
  assign N11082 = N11081 | data_masked[855];
  assign N11081 = N11080 | data_masked[983];
  assign N11080 = N11079 | data_masked[1111];
  assign N11079 = N11078 | data_masked[1239];
  assign N11078 = N11077 | data_masked[1367];
  assign N11077 = N11076 | data_masked[1495];
  assign N11076 = N11075 | data_masked[1623];
  assign N11075 = N11074 | data_masked[1751];
  assign N11074 = N11073 | data_masked[1879];
  assign N11073 = N11072 | data_masked[2007];
  assign N11072 = N11071 | data_masked[2135];
  assign N11071 = N11070 | data_masked[2263];
  assign N11070 = N11069 | data_masked[2391];
  assign N11069 = N11068 | data_masked[2519];
  assign N11068 = N11067 | data_masked[2647];
  assign N11067 = N11066 | data_masked[2775];
  assign N11066 = N11065 | data_masked[2903];
  assign N11065 = N11064 | data_masked[3031];
  assign N11064 = N11063 | data_masked[3159];
  assign N11063 = N11062 | data_masked[3287];
  assign N11062 = N11061 | data_masked[3415];
  assign N11061 = N11060 | data_masked[3543];
  assign N11060 = N11059 | data_masked[3671];
  assign N11059 = N11058 | data_masked[3799];
  assign N11058 = N11057 | data_masked[3927];
  assign N11057 = N11056 | data_masked[4055];
  assign N11056 = N11055 | data_masked[4183];
  assign N11055 = N11054 | data_masked[4311];
  assign N11054 = N11053 | data_masked[4439];
  assign N11053 = N11052 | data_masked[4567];
  assign N11052 = N11051 | data_masked[4695];
  assign N11051 = N11050 | data_masked[4823];
  assign N11050 = N11049 | data_masked[4951];
  assign N11049 = N11048 | data_masked[5079];
  assign N11048 = N11047 | data_masked[5207];
  assign N11047 = N11046 | data_masked[5335];
  assign N11046 = N11045 | data_masked[5463];
  assign N11045 = N11044 | data_masked[5591];
  assign N11044 = N11043 | data_masked[5719];
  assign N11043 = N11042 | data_masked[5847];
  assign N11042 = N11041 | data_masked[5975];
  assign N11041 = N11040 | data_masked[6103];
  assign N11040 = N11039 | data_masked[6231];
  assign N11039 = N11038 | data_masked[6359];
  assign N11038 = N11037 | data_masked[6487];
  assign N11037 = N11036 | data_masked[6615];
  assign N11036 = N11035 | data_masked[6743];
  assign N11035 = N11034 | data_masked[6871];
  assign N11034 = N11033 | data_masked[6999];
  assign N11033 = N11032 | data_masked[7127];
  assign N11032 = N11031 | data_masked[7255];
  assign N11031 = N11030 | data_masked[7383];
  assign N11030 = N11029 | data_masked[7511];
  assign N11029 = N11028 | data_masked[7639];
  assign N11028 = N11027 | data_masked[7767];
  assign N11027 = N11026 | data_masked[7895];
  assign N11026 = N11025 | data_masked[8023];
  assign N11025 = N11024 | data_masked[8151];
  assign N11024 = N11023 | data_masked[8279];
  assign N11023 = N11022 | data_masked[8407];
  assign N11022 = N11021 | data_masked[8535];
  assign N11021 = N11020 | data_masked[8663];
  assign N11020 = N11019 | data_masked[8791];
  assign N11019 = N11018 | data_masked[8919];
  assign N11018 = N11017 | data_masked[9047];
  assign N11017 = N11016 | data_masked[9175];
  assign N11016 = N11015 | data_masked[9303];
  assign N11015 = N11014 | data_masked[9431];
  assign N11014 = N11013 | data_masked[9559];
  assign N11013 = N11012 | data_masked[9687];
  assign N11012 = N11011 | data_masked[9815];
  assign N11011 = N11010 | data_masked[9943];
  assign N11010 = N11009 | data_masked[10071];
  assign N11009 = N11008 | data_masked[10199];
  assign N11008 = N11007 | data_masked[10327];
  assign N11007 = N11006 | data_masked[10455];
  assign N11006 = N11005 | data_masked[10583];
  assign N11005 = N11004 | data_masked[10711];
  assign N11004 = N11003 | data_masked[10839];
  assign N11003 = N11002 | data_masked[10967];
  assign N11002 = N11001 | data_masked[11095];
  assign N11001 = N11000 | data_masked[11223];
  assign N11000 = N10999 | data_masked[11351];
  assign N10999 = N10998 | data_masked[11479];
  assign N10998 = N10997 | data_masked[11607];
  assign N10997 = N10996 | data_masked[11735];
  assign N10996 = N10995 | data_masked[11863];
  assign N10995 = N10994 | data_masked[11991];
  assign N10994 = N10993 | data_masked[12119];
  assign N10993 = N10992 | data_masked[12247];
  assign N10992 = N10991 | data_masked[12375];
  assign N10991 = N10990 | data_masked[12503];
  assign N10990 = N10989 | data_masked[12631];
  assign N10989 = N10988 | data_masked[12759];
  assign N10988 = N10987 | data_masked[12887];
  assign N10987 = N10986 | data_masked[13015];
  assign N10986 = N10985 | data_masked[13143];
  assign N10985 = N10984 | data_masked[13271];
  assign N10984 = N10983 | data_masked[13399];
  assign N10983 = N10982 | data_masked[13527];
  assign N10982 = N10981 | data_masked[13655];
  assign N10981 = N10980 | data_masked[13783];
  assign N10980 = N10979 | data_masked[13911];
  assign N10979 = N10978 | data_masked[14039];
  assign N10978 = N10977 | data_masked[14167];
  assign N10977 = N10976 | data_masked[14295];
  assign N10976 = N10975 | data_masked[14423];
  assign N10975 = N10974 | data_masked[14551];
  assign N10974 = N10973 | data_masked[14679];
  assign N10973 = N10972 | data_masked[14807];
  assign N10972 = N10971 | data_masked[14935];
  assign N10971 = N10970 | data_masked[15063];
  assign N10970 = N10969 | data_masked[15191];
  assign N10969 = N10968 | data_masked[15319];
  assign N10968 = N10967 | data_masked[15447];
  assign N10967 = N10966 | data_masked[15575];
  assign N10966 = N10965 | data_masked[15703];
  assign N10965 = N10964 | data_masked[15831];
  assign N10964 = N10963 | data_masked[15959];
  assign N10963 = N10962 | data_masked[16087];
  assign N10962 = data_masked[16343] | data_masked[16215];
  assign data_o[88] = N11213 | data_masked[88];
  assign N11213 = N11212 | data_masked[216];
  assign N11212 = N11211 | data_masked[344];
  assign N11211 = N11210 | data_masked[472];
  assign N11210 = N11209 | data_masked[600];
  assign N11209 = N11208 | data_masked[728];
  assign N11208 = N11207 | data_masked[856];
  assign N11207 = N11206 | data_masked[984];
  assign N11206 = N11205 | data_masked[1112];
  assign N11205 = N11204 | data_masked[1240];
  assign N11204 = N11203 | data_masked[1368];
  assign N11203 = N11202 | data_masked[1496];
  assign N11202 = N11201 | data_masked[1624];
  assign N11201 = N11200 | data_masked[1752];
  assign N11200 = N11199 | data_masked[1880];
  assign N11199 = N11198 | data_masked[2008];
  assign N11198 = N11197 | data_masked[2136];
  assign N11197 = N11196 | data_masked[2264];
  assign N11196 = N11195 | data_masked[2392];
  assign N11195 = N11194 | data_masked[2520];
  assign N11194 = N11193 | data_masked[2648];
  assign N11193 = N11192 | data_masked[2776];
  assign N11192 = N11191 | data_masked[2904];
  assign N11191 = N11190 | data_masked[3032];
  assign N11190 = N11189 | data_masked[3160];
  assign N11189 = N11188 | data_masked[3288];
  assign N11188 = N11187 | data_masked[3416];
  assign N11187 = N11186 | data_masked[3544];
  assign N11186 = N11185 | data_masked[3672];
  assign N11185 = N11184 | data_masked[3800];
  assign N11184 = N11183 | data_masked[3928];
  assign N11183 = N11182 | data_masked[4056];
  assign N11182 = N11181 | data_masked[4184];
  assign N11181 = N11180 | data_masked[4312];
  assign N11180 = N11179 | data_masked[4440];
  assign N11179 = N11178 | data_masked[4568];
  assign N11178 = N11177 | data_masked[4696];
  assign N11177 = N11176 | data_masked[4824];
  assign N11176 = N11175 | data_masked[4952];
  assign N11175 = N11174 | data_masked[5080];
  assign N11174 = N11173 | data_masked[5208];
  assign N11173 = N11172 | data_masked[5336];
  assign N11172 = N11171 | data_masked[5464];
  assign N11171 = N11170 | data_masked[5592];
  assign N11170 = N11169 | data_masked[5720];
  assign N11169 = N11168 | data_masked[5848];
  assign N11168 = N11167 | data_masked[5976];
  assign N11167 = N11166 | data_masked[6104];
  assign N11166 = N11165 | data_masked[6232];
  assign N11165 = N11164 | data_masked[6360];
  assign N11164 = N11163 | data_masked[6488];
  assign N11163 = N11162 | data_masked[6616];
  assign N11162 = N11161 | data_masked[6744];
  assign N11161 = N11160 | data_masked[6872];
  assign N11160 = N11159 | data_masked[7000];
  assign N11159 = N11158 | data_masked[7128];
  assign N11158 = N11157 | data_masked[7256];
  assign N11157 = N11156 | data_masked[7384];
  assign N11156 = N11155 | data_masked[7512];
  assign N11155 = N11154 | data_masked[7640];
  assign N11154 = N11153 | data_masked[7768];
  assign N11153 = N11152 | data_masked[7896];
  assign N11152 = N11151 | data_masked[8024];
  assign N11151 = N11150 | data_masked[8152];
  assign N11150 = N11149 | data_masked[8280];
  assign N11149 = N11148 | data_masked[8408];
  assign N11148 = N11147 | data_masked[8536];
  assign N11147 = N11146 | data_masked[8664];
  assign N11146 = N11145 | data_masked[8792];
  assign N11145 = N11144 | data_masked[8920];
  assign N11144 = N11143 | data_masked[9048];
  assign N11143 = N11142 | data_masked[9176];
  assign N11142 = N11141 | data_masked[9304];
  assign N11141 = N11140 | data_masked[9432];
  assign N11140 = N11139 | data_masked[9560];
  assign N11139 = N11138 | data_masked[9688];
  assign N11138 = N11137 | data_masked[9816];
  assign N11137 = N11136 | data_masked[9944];
  assign N11136 = N11135 | data_masked[10072];
  assign N11135 = N11134 | data_masked[10200];
  assign N11134 = N11133 | data_masked[10328];
  assign N11133 = N11132 | data_masked[10456];
  assign N11132 = N11131 | data_masked[10584];
  assign N11131 = N11130 | data_masked[10712];
  assign N11130 = N11129 | data_masked[10840];
  assign N11129 = N11128 | data_masked[10968];
  assign N11128 = N11127 | data_masked[11096];
  assign N11127 = N11126 | data_masked[11224];
  assign N11126 = N11125 | data_masked[11352];
  assign N11125 = N11124 | data_masked[11480];
  assign N11124 = N11123 | data_masked[11608];
  assign N11123 = N11122 | data_masked[11736];
  assign N11122 = N11121 | data_masked[11864];
  assign N11121 = N11120 | data_masked[11992];
  assign N11120 = N11119 | data_masked[12120];
  assign N11119 = N11118 | data_masked[12248];
  assign N11118 = N11117 | data_masked[12376];
  assign N11117 = N11116 | data_masked[12504];
  assign N11116 = N11115 | data_masked[12632];
  assign N11115 = N11114 | data_masked[12760];
  assign N11114 = N11113 | data_masked[12888];
  assign N11113 = N11112 | data_masked[13016];
  assign N11112 = N11111 | data_masked[13144];
  assign N11111 = N11110 | data_masked[13272];
  assign N11110 = N11109 | data_masked[13400];
  assign N11109 = N11108 | data_masked[13528];
  assign N11108 = N11107 | data_masked[13656];
  assign N11107 = N11106 | data_masked[13784];
  assign N11106 = N11105 | data_masked[13912];
  assign N11105 = N11104 | data_masked[14040];
  assign N11104 = N11103 | data_masked[14168];
  assign N11103 = N11102 | data_masked[14296];
  assign N11102 = N11101 | data_masked[14424];
  assign N11101 = N11100 | data_masked[14552];
  assign N11100 = N11099 | data_masked[14680];
  assign N11099 = N11098 | data_masked[14808];
  assign N11098 = N11097 | data_masked[14936];
  assign N11097 = N11096 | data_masked[15064];
  assign N11096 = N11095 | data_masked[15192];
  assign N11095 = N11094 | data_masked[15320];
  assign N11094 = N11093 | data_masked[15448];
  assign N11093 = N11092 | data_masked[15576];
  assign N11092 = N11091 | data_masked[15704];
  assign N11091 = N11090 | data_masked[15832];
  assign N11090 = N11089 | data_masked[15960];
  assign N11089 = N11088 | data_masked[16088];
  assign N11088 = data_masked[16344] | data_masked[16216];
  assign data_o[89] = N11339 | data_masked[89];
  assign N11339 = N11338 | data_masked[217];
  assign N11338 = N11337 | data_masked[345];
  assign N11337 = N11336 | data_masked[473];
  assign N11336 = N11335 | data_masked[601];
  assign N11335 = N11334 | data_masked[729];
  assign N11334 = N11333 | data_masked[857];
  assign N11333 = N11332 | data_masked[985];
  assign N11332 = N11331 | data_masked[1113];
  assign N11331 = N11330 | data_masked[1241];
  assign N11330 = N11329 | data_masked[1369];
  assign N11329 = N11328 | data_masked[1497];
  assign N11328 = N11327 | data_masked[1625];
  assign N11327 = N11326 | data_masked[1753];
  assign N11326 = N11325 | data_masked[1881];
  assign N11325 = N11324 | data_masked[2009];
  assign N11324 = N11323 | data_masked[2137];
  assign N11323 = N11322 | data_masked[2265];
  assign N11322 = N11321 | data_masked[2393];
  assign N11321 = N11320 | data_masked[2521];
  assign N11320 = N11319 | data_masked[2649];
  assign N11319 = N11318 | data_masked[2777];
  assign N11318 = N11317 | data_masked[2905];
  assign N11317 = N11316 | data_masked[3033];
  assign N11316 = N11315 | data_masked[3161];
  assign N11315 = N11314 | data_masked[3289];
  assign N11314 = N11313 | data_masked[3417];
  assign N11313 = N11312 | data_masked[3545];
  assign N11312 = N11311 | data_masked[3673];
  assign N11311 = N11310 | data_masked[3801];
  assign N11310 = N11309 | data_masked[3929];
  assign N11309 = N11308 | data_masked[4057];
  assign N11308 = N11307 | data_masked[4185];
  assign N11307 = N11306 | data_masked[4313];
  assign N11306 = N11305 | data_masked[4441];
  assign N11305 = N11304 | data_masked[4569];
  assign N11304 = N11303 | data_masked[4697];
  assign N11303 = N11302 | data_masked[4825];
  assign N11302 = N11301 | data_masked[4953];
  assign N11301 = N11300 | data_masked[5081];
  assign N11300 = N11299 | data_masked[5209];
  assign N11299 = N11298 | data_masked[5337];
  assign N11298 = N11297 | data_masked[5465];
  assign N11297 = N11296 | data_masked[5593];
  assign N11296 = N11295 | data_masked[5721];
  assign N11295 = N11294 | data_masked[5849];
  assign N11294 = N11293 | data_masked[5977];
  assign N11293 = N11292 | data_masked[6105];
  assign N11292 = N11291 | data_masked[6233];
  assign N11291 = N11290 | data_masked[6361];
  assign N11290 = N11289 | data_masked[6489];
  assign N11289 = N11288 | data_masked[6617];
  assign N11288 = N11287 | data_masked[6745];
  assign N11287 = N11286 | data_masked[6873];
  assign N11286 = N11285 | data_masked[7001];
  assign N11285 = N11284 | data_masked[7129];
  assign N11284 = N11283 | data_masked[7257];
  assign N11283 = N11282 | data_masked[7385];
  assign N11282 = N11281 | data_masked[7513];
  assign N11281 = N11280 | data_masked[7641];
  assign N11280 = N11279 | data_masked[7769];
  assign N11279 = N11278 | data_masked[7897];
  assign N11278 = N11277 | data_masked[8025];
  assign N11277 = N11276 | data_masked[8153];
  assign N11276 = N11275 | data_masked[8281];
  assign N11275 = N11274 | data_masked[8409];
  assign N11274 = N11273 | data_masked[8537];
  assign N11273 = N11272 | data_masked[8665];
  assign N11272 = N11271 | data_masked[8793];
  assign N11271 = N11270 | data_masked[8921];
  assign N11270 = N11269 | data_masked[9049];
  assign N11269 = N11268 | data_masked[9177];
  assign N11268 = N11267 | data_masked[9305];
  assign N11267 = N11266 | data_masked[9433];
  assign N11266 = N11265 | data_masked[9561];
  assign N11265 = N11264 | data_masked[9689];
  assign N11264 = N11263 | data_masked[9817];
  assign N11263 = N11262 | data_masked[9945];
  assign N11262 = N11261 | data_masked[10073];
  assign N11261 = N11260 | data_masked[10201];
  assign N11260 = N11259 | data_masked[10329];
  assign N11259 = N11258 | data_masked[10457];
  assign N11258 = N11257 | data_masked[10585];
  assign N11257 = N11256 | data_masked[10713];
  assign N11256 = N11255 | data_masked[10841];
  assign N11255 = N11254 | data_masked[10969];
  assign N11254 = N11253 | data_masked[11097];
  assign N11253 = N11252 | data_masked[11225];
  assign N11252 = N11251 | data_masked[11353];
  assign N11251 = N11250 | data_masked[11481];
  assign N11250 = N11249 | data_masked[11609];
  assign N11249 = N11248 | data_masked[11737];
  assign N11248 = N11247 | data_masked[11865];
  assign N11247 = N11246 | data_masked[11993];
  assign N11246 = N11245 | data_masked[12121];
  assign N11245 = N11244 | data_masked[12249];
  assign N11244 = N11243 | data_masked[12377];
  assign N11243 = N11242 | data_masked[12505];
  assign N11242 = N11241 | data_masked[12633];
  assign N11241 = N11240 | data_masked[12761];
  assign N11240 = N11239 | data_masked[12889];
  assign N11239 = N11238 | data_masked[13017];
  assign N11238 = N11237 | data_masked[13145];
  assign N11237 = N11236 | data_masked[13273];
  assign N11236 = N11235 | data_masked[13401];
  assign N11235 = N11234 | data_masked[13529];
  assign N11234 = N11233 | data_masked[13657];
  assign N11233 = N11232 | data_masked[13785];
  assign N11232 = N11231 | data_masked[13913];
  assign N11231 = N11230 | data_masked[14041];
  assign N11230 = N11229 | data_masked[14169];
  assign N11229 = N11228 | data_masked[14297];
  assign N11228 = N11227 | data_masked[14425];
  assign N11227 = N11226 | data_masked[14553];
  assign N11226 = N11225 | data_masked[14681];
  assign N11225 = N11224 | data_masked[14809];
  assign N11224 = N11223 | data_masked[14937];
  assign N11223 = N11222 | data_masked[15065];
  assign N11222 = N11221 | data_masked[15193];
  assign N11221 = N11220 | data_masked[15321];
  assign N11220 = N11219 | data_masked[15449];
  assign N11219 = N11218 | data_masked[15577];
  assign N11218 = N11217 | data_masked[15705];
  assign N11217 = N11216 | data_masked[15833];
  assign N11216 = N11215 | data_masked[15961];
  assign N11215 = N11214 | data_masked[16089];
  assign N11214 = data_masked[16345] | data_masked[16217];
  assign data_o[90] = N11465 | data_masked[90];
  assign N11465 = N11464 | data_masked[218];
  assign N11464 = N11463 | data_masked[346];
  assign N11463 = N11462 | data_masked[474];
  assign N11462 = N11461 | data_masked[602];
  assign N11461 = N11460 | data_masked[730];
  assign N11460 = N11459 | data_masked[858];
  assign N11459 = N11458 | data_masked[986];
  assign N11458 = N11457 | data_masked[1114];
  assign N11457 = N11456 | data_masked[1242];
  assign N11456 = N11455 | data_masked[1370];
  assign N11455 = N11454 | data_masked[1498];
  assign N11454 = N11453 | data_masked[1626];
  assign N11453 = N11452 | data_masked[1754];
  assign N11452 = N11451 | data_masked[1882];
  assign N11451 = N11450 | data_masked[2010];
  assign N11450 = N11449 | data_masked[2138];
  assign N11449 = N11448 | data_masked[2266];
  assign N11448 = N11447 | data_masked[2394];
  assign N11447 = N11446 | data_masked[2522];
  assign N11446 = N11445 | data_masked[2650];
  assign N11445 = N11444 | data_masked[2778];
  assign N11444 = N11443 | data_masked[2906];
  assign N11443 = N11442 | data_masked[3034];
  assign N11442 = N11441 | data_masked[3162];
  assign N11441 = N11440 | data_masked[3290];
  assign N11440 = N11439 | data_masked[3418];
  assign N11439 = N11438 | data_masked[3546];
  assign N11438 = N11437 | data_masked[3674];
  assign N11437 = N11436 | data_masked[3802];
  assign N11436 = N11435 | data_masked[3930];
  assign N11435 = N11434 | data_masked[4058];
  assign N11434 = N11433 | data_masked[4186];
  assign N11433 = N11432 | data_masked[4314];
  assign N11432 = N11431 | data_masked[4442];
  assign N11431 = N11430 | data_masked[4570];
  assign N11430 = N11429 | data_masked[4698];
  assign N11429 = N11428 | data_masked[4826];
  assign N11428 = N11427 | data_masked[4954];
  assign N11427 = N11426 | data_masked[5082];
  assign N11426 = N11425 | data_masked[5210];
  assign N11425 = N11424 | data_masked[5338];
  assign N11424 = N11423 | data_masked[5466];
  assign N11423 = N11422 | data_masked[5594];
  assign N11422 = N11421 | data_masked[5722];
  assign N11421 = N11420 | data_masked[5850];
  assign N11420 = N11419 | data_masked[5978];
  assign N11419 = N11418 | data_masked[6106];
  assign N11418 = N11417 | data_masked[6234];
  assign N11417 = N11416 | data_masked[6362];
  assign N11416 = N11415 | data_masked[6490];
  assign N11415 = N11414 | data_masked[6618];
  assign N11414 = N11413 | data_masked[6746];
  assign N11413 = N11412 | data_masked[6874];
  assign N11412 = N11411 | data_masked[7002];
  assign N11411 = N11410 | data_masked[7130];
  assign N11410 = N11409 | data_masked[7258];
  assign N11409 = N11408 | data_masked[7386];
  assign N11408 = N11407 | data_masked[7514];
  assign N11407 = N11406 | data_masked[7642];
  assign N11406 = N11405 | data_masked[7770];
  assign N11405 = N11404 | data_masked[7898];
  assign N11404 = N11403 | data_masked[8026];
  assign N11403 = N11402 | data_masked[8154];
  assign N11402 = N11401 | data_masked[8282];
  assign N11401 = N11400 | data_masked[8410];
  assign N11400 = N11399 | data_masked[8538];
  assign N11399 = N11398 | data_masked[8666];
  assign N11398 = N11397 | data_masked[8794];
  assign N11397 = N11396 | data_masked[8922];
  assign N11396 = N11395 | data_masked[9050];
  assign N11395 = N11394 | data_masked[9178];
  assign N11394 = N11393 | data_masked[9306];
  assign N11393 = N11392 | data_masked[9434];
  assign N11392 = N11391 | data_masked[9562];
  assign N11391 = N11390 | data_masked[9690];
  assign N11390 = N11389 | data_masked[9818];
  assign N11389 = N11388 | data_masked[9946];
  assign N11388 = N11387 | data_masked[10074];
  assign N11387 = N11386 | data_masked[10202];
  assign N11386 = N11385 | data_masked[10330];
  assign N11385 = N11384 | data_masked[10458];
  assign N11384 = N11383 | data_masked[10586];
  assign N11383 = N11382 | data_masked[10714];
  assign N11382 = N11381 | data_masked[10842];
  assign N11381 = N11380 | data_masked[10970];
  assign N11380 = N11379 | data_masked[11098];
  assign N11379 = N11378 | data_masked[11226];
  assign N11378 = N11377 | data_masked[11354];
  assign N11377 = N11376 | data_masked[11482];
  assign N11376 = N11375 | data_masked[11610];
  assign N11375 = N11374 | data_masked[11738];
  assign N11374 = N11373 | data_masked[11866];
  assign N11373 = N11372 | data_masked[11994];
  assign N11372 = N11371 | data_masked[12122];
  assign N11371 = N11370 | data_masked[12250];
  assign N11370 = N11369 | data_masked[12378];
  assign N11369 = N11368 | data_masked[12506];
  assign N11368 = N11367 | data_masked[12634];
  assign N11367 = N11366 | data_masked[12762];
  assign N11366 = N11365 | data_masked[12890];
  assign N11365 = N11364 | data_masked[13018];
  assign N11364 = N11363 | data_masked[13146];
  assign N11363 = N11362 | data_masked[13274];
  assign N11362 = N11361 | data_masked[13402];
  assign N11361 = N11360 | data_masked[13530];
  assign N11360 = N11359 | data_masked[13658];
  assign N11359 = N11358 | data_masked[13786];
  assign N11358 = N11357 | data_masked[13914];
  assign N11357 = N11356 | data_masked[14042];
  assign N11356 = N11355 | data_masked[14170];
  assign N11355 = N11354 | data_masked[14298];
  assign N11354 = N11353 | data_masked[14426];
  assign N11353 = N11352 | data_masked[14554];
  assign N11352 = N11351 | data_masked[14682];
  assign N11351 = N11350 | data_masked[14810];
  assign N11350 = N11349 | data_masked[14938];
  assign N11349 = N11348 | data_masked[15066];
  assign N11348 = N11347 | data_masked[15194];
  assign N11347 = N11346 | data_masked[15322];
  assign N11346 = N11345 | data_masked[15450];
  assign N11345 = N11344 | data_masked[15578];
  assign N11344 = N11343 | data_masked[15706];
  assign N11343 = N11342 | data_masked[15834];
  assign N11342 = N11341 | data_masked[15962];
  assign N11341 = N11340 | data_masked[16090];
  assign N11340 = data_masked[16346] | data_masked[16218];
  assign data_o[91] = N11591 | data_masked[91];
  assign N11591 = N11590 | data_masked[219];
  assign N11590 = N11589 | data_masked[347];
  assign N11589 = N11588 | data_masked[475];
  assign N11588 = N11587 | data_masked[603];
  assign N11587 = N11586 | data_masked[731];
  assign N11586 = N11585 | data_masked[859];
  assign N11585 = N11584 | data_masked[987];
  assign N11584 = N11583 | data_masked[1115];
  assign N11583 = N11582 | data_masked[1243];
  assign N11582 = N11581 | data_masked[1371];
  assign N11581 = N11580 | data_masked[1499];
  assign N11580 = N11579 | data_masked[1627];
  assign N11579 = N11578 | data_masked[1755];
  assign N11578 = N11577 | data_masked[1883];
  assign N11577 = N11576 | data_masked[2011];
  assign N11576 = N11575 | data_masked[2139];
  assign N11575 = N11574 | data_masked[2267];
  assign N11574 = N11573 | data_masked[2395];
  assign N11573 = N11572 | data_masked[2523];
  assign N11572 = N11571 | data_masked[2651];
  assign N11571 = N11570 | data_masked[2779];
  assign N11570 = N11569 | data_masked[2907];
  assign N11569 = N11568 | data_masked[3035];
  assign N11568 = N11567 | data_masked[3163];
  assign N11567 = N11566 | data_masked[3291];
  assign N11566 = N11565 | data_masked[3419];
  assign N11565 = N11564 | data_masked[3547];
  assign N11564 = N11563 | data_masked[3675];
  assign N11563 = N11562 | data_masked[3803];
  assign N11562 = N11561 | data_masked[3931];
  assign N11561 = N11560 | data_masked[4059];
  assign N11560 = N11559 | data_masked[4187];
  assign N11559 = N11558 | data_masked[4315];
  assign N11558 = N11557 | data_masked[4443];
  assign N11557 = N11556 | data_masked[4571];
  assign N11556 = N11555 | data_masked[4699];
  assign N11555 = N11554 | data_masked[4827];
  assign N11554 = N11553 | data_masked[4955];
  assign N11553 = N11552 | data_masked[5083];
  assign N11552 = N11551 | data_masked[5211];
  assign N11551 = N11550 | data_masked[5339];
  assign N11550 = N11549 | data_masked[5467];
  assign N11549 = N11548 | data_masked[5595];
  assign N11548 = N11547 | data_masked[5723];
  assign N11547 = N11546 | data_masked[5851];
  assign N11546 = N11545 | data_masked[5979];
  assign N11545 = N11544 | data_masked[6107];
  assign N11544 = N11543 | data_masked[6235];
  assign N11543 = N11542 | data_masked[6363];
  assign N11542 = N11541 | data_masked[6491];
  assign N11541 = N11540 | data_masked[6619];
  assign N11540 = N11539 | data_masked[6747];
  assign N11539 = N11538 | data_masked[6875];
  assign N11538 = N11537 | data_masked[7003];
  assign N11537 = N11536 | data_masked[7131];
  assign N11536 = N11535 | data_masked[7259];
  assign N11535 = N11534 | data_masked[7387];
  assign N11534 = N11533 | data_masked[7515];
  assign N11533 = N11532 | data_masked[7643];
  assign N11532 = N11531 | data_masked[7771];
  assign N11531 = N11530 | data_masked[7899];
  assign N11530 = N11529 | data_masked[8027];
  assign N11529 = N11528 | data_masked[8155];
  assign N11528 = N11527 | data_masked[8283];
  assign N11527 = N11526 | data_masked[8411];
  assign N11526 = N11525 | data_masked[8539];
  assign N11525 = N11524 | data_masked[8667];
  assign N11524 = N11523 | data_masked[8795];
  assign N11523 = N11522 | data_masked[8923];
  assign N11522 = N11521 | data_masked[9051];
  assign N11521 = N11520 | data_masked[9179];
  assign N11520 = N11519 | data_masked[9307];
  assign N11519 = N11518 | data_masked[9435];
  assign N11518 = N11517 | data_masked[9563];
  assign N11517 = N11516 | data_masked[9691];
  assign N11516 = N11515 | data_masked[9819];
  assign N11515 = N11514 | data_masked[9947];
  assign N11514 = N11513 | data_masked[10075];
  assign N11513 = N11512 | data_masked[10203];
  assign N11512 = N11511 | data_masked[10331];
  assign N11511 = N11510 | data_masked[10459];
  assign N11510 = N11509 | data_masked[10587];
  assign N11509 = N11508 | data_masked[10715];
  assign N11508 = N11507 | data_masked[10843];
  assign N11507 = N11506 | data_masked[10971];
  assign N11506 = N11505 | data_masked[11099];
  assign N11505 = N11504 | data_masked[11227];
  assign N11504 = N11503 | data_masked[11355];
  assign N11503 = N11502 | data_masked[11483];
  assign N11502 = N11501 | data_masked[11611];
  assign N11501 = N11500 | data_masked[11739];
  assign N11500 = N11499 | data_masked[11867];
  assign N11499 = N11498 | data_masked[11995];
  assign N11498 = N11497 | data_masked[12123];
  assign N11497 = N11496 | data_masked[12251];
  assign N11496 = N11495 | data_masked[12379];
  assign N11495 = N11494 | data_masked[12507];
  assign N11494 = N11493 | data_masked[12635];
  assign N11493 = N11492 | data_masked[12763];
  assign N11492 = N11491 | data_masked[12891];
  assign N11491 = N11490 | data_masked[13019];
  assign N11490 = N11489 | data_masked[13147];
  assign N11489 = N11488 | data_masked[13275];
  assign N11488 = N11487 | data_masked[13403];
  assign N11487 = N11486 | data_masked[13531];
  assign N11486 = N11485 | data_masked[13659];
  assign N11485 = N11484 | data_masked[13787];
  assign N11484 = N11483 | data_masked[13915];
  assign N11483 = N11482 | data_masked[14043];
  assign N11482 = N11481 | data_masked[14171];
  assign N11481 = N11480 | data_masked[14299];
  assign N11480 = N11479 | data_masked[14427];
  assign N11479 = N11478 | data_masked[14555];
  assign N11478 = N11477 | data_masked[14683];
  assign N11477 = N11476 | data_masked[14811];
  assign N11476 = N11475 | data_masked[14939];
  assign N11475 = N11474 | data_masked[15067];
  assign N11474 = N11473 | data_masked[15195];
  assign N11473 = N11472 | data_masked[15323];
  assign N11472 = N11471 | data_masked[15451];
  assign N11471 = N11470 | data_masked[15579];
  assign N11470 = N11469 | data_masked[15707];
  assign N11469 = N11468 | data_masked[15835];
  assign N11468 = N11467 | data_masked[15963];
  assign N11467 = N11466 | data_masked[16091];
  assign N11466 = data_masked[16347] | data_masked[16219];
  assign data_o[92] = N11717 | data_masked[92];
  assign N11717 = N11716 | data_masked[220];
  assign N11716 = N11715 | data_masked[348];
  assign N11715 = N11714 | data_masked[476];
  assign N11714 = N11713 | data_masked[604];
  assign N11713 = N11712 | data_masked[732];
  assign N11712 = N11711 | data_masked[860];
  assign N11711 = N11710 | data_masked[988];
  assign N11710 = N11709 | data_masked[1116];
  assign N11709 = N11708 | data_masked[1244];
  assign N11708 = N11707 | data_masked[1372];
  assign N11707 = N11706 | data_masked[1500];
  assign N11706 = N11705 | data_masked[1628];
  assign N11705 = N11704 | data_masked[1756];
  assign N11704 = N11703 | data_masked[1884];
  assign N11703 = N11702 | data_masked[2012];
  assign N11702 = N11701 | data_masked[2140];
  assign N11701 = N11700 | data_masked[2268];
  assign N11700 = N11699 | data_masked[2396];
  assign N11699 = N11698 | data_masked[2524];
  assign N11698 = N11697 | data_masked[2652];
  assign N11697 = N11696 | data_masked[2780];
  assign N11696 = N11695 | data_masked[2908];
  assign N11695 = N11694 | data_masked[3036];
  assign N11694 = N11693 | data_masked[3164];
  assign N11693 = N11692 | data_masked[3292];
  assign N11692 = N11691 | data_masked[3420];
  assign N11691 = N11690 | data_masked[3548];
  assign N11690 = N11689 | data_masked[3676];
  assign N11689 = N11688 | data_masked[3804];
  assign N11688 = N11687 | data_masked[3932];
  assign N11687 = N11686 | data_masked[4060];
  assign N11686 = N11685 | data_masked[4188];
  assign N11685 = N11684 | data_masked[4316];
  assign N11684 = N11683 | data_masked[4444];
  assign N11683 = N11682 | data_masked[4572];
  assign N11682 = N11681 | data_masked[4700];
  assign N11681 = N11680 | data_masked[4828];
  assign N11680 = N11679 | data_masked[4956];
  assign N11679 = N11678 | data_masked[5084];
  assign N11678 = N11677 | data_masked[5212];
  assign N11677 = N11676 | data_masked[5340];
  assign N11676 = N11675 | data_masked[5468];
  assign N11675 = N11674 | data_masked[5596];
  assign N11674 = N11673 | data_masked[5724];
  assign N11673 = N11672 | data_masked[5852];
  assign N11672 = N11671 | data_masked[5980];
  assign N11671 = N11670 | data_masked[6108];
  assign N11670 = N11669 | data_masked[6236];
  assign N11669 = N11668 | data_masked[6364];
  assign N11668 = N11667 | data_masked[6492];
  assign N11667 = N11666 | data_masked[6620];
  assign N11666 = N11665 | data_masked[6748];
  assign N11665 = N11664 | data_masked[6876];
  assign N11664 = N11663 | data_masked[7004];
  assign N11663 = N11662 | data_masked[7132];
  assign N11662 = N11661 | data_masked[7260];
  assign N11661 = N11660 | data_masked[7388];
  assign N11660 = N11659 | data_masked[7516];
  assign N11659 = N11658 | data_masked[7644];
  assign N11658 = N11657 | data_masked[7772];
  assign N11657 = N11656 | data_masked[7900];
  assign N11656 = N11655 | data_masked[8028];
  assign N11655 = N11654 | data_masked[8156];
  assign N11654 = N11653 | data_masked[8284];
  assign N11653 = N11652 | data_masked[8412];
  assign N11652 = N11651 | data_masked[8540];
  assign N11651 = N11650 | data_masked[8668];
  assign N11650 = N11649 | data_masked[8796];
  assign N11649 = N11648 | data_masked[8924];
  assign N11648 = N11647 | data_masked[9052];
  assign N11647 = N11646 | data_masked[9180];
  assign N11646 = N11645 | data_masked[9308];
  assign N11645 = N11644 | data_masked[9436];
  assign N11644 = N11643 | data_masked[9564];
  assign N11643 = N11642 | data_masked[9692];
  assign N11642 = N11641 | data_masked[9820];
  assign N11641 = N11640 | data_masked[9948];
  assign N11640 = N11639 | data_masked[10076];
  assign N11639 = N11638 | data_masked[10204];
  assign N11638 = N11637 | data_masked[10332];
  assign N11637 = N11636 | data_masked[10460];
  assign N11636 = N11635 | data_masked[10588];
  assign N11635 = N11634 | data_masked[10716];
  assign N11634 = N11633 | data_masked[10844];
  assign N11633 = N11632 | data_masked[10972];
  assign N11632 = N11631 | data_masked[11100];
  assign N11631 = N11630 | data_masked[11228];
  assign N11630 = N11629 | data_masked[11356];
  assign N11629 = N11628 | data_masked[11484];
  assign N11628 = N11627 | data_masked[11612];
  assign N11627 = N11626 | data_masked[11740];
  assign N11626 = N11625 | data_masked[11868];
  assign N11625 = N11624 | data_masked[11996];
  assign N11624 = N11623 | data_masked[12124];
  assign N11623 = N11622 | data_masked[12252];
  assign N11622 = N11621 | data_masked[12380];
  assign N11621 = N11620 | data_masked[12508];
  assign N11620 = N11619 | data_masked[12636];
  assign N11619 = N11618 | data_masked[12764];
  assign N11618 = N11617 | data_masked[12892];
  assign N11617 = N11616 | data_masked[13020];
  assign N11616 = N11615 | data_masked[13148];
  assign N11615 = N11614 | data_masked[13276];
  assign N11614 = N11613 | data_masked[13404];
  assign N11613 = N11612 | data_masked[13532];
  assign N11612 = N11611 | data_masked[13660];
  assign N11611 = N11610 | data_masked[13788];
  assign N11610 = N11609 | data_masked[13916];
  assign N11609 = N11608 | data_masked[14044];
  assign N11608 = N11607 | data_masked[14172];
  assign N11607 = N11606 | data_masked[14300];
  assign N11606 = N11605 | data_masked[14428];
  assign N11605 = N11604 | data_masked[14556];
  assign N11604 = N11603 | data_masked[14684];
  assign N11603 = N11602 | data_masked[14812];
  assign N11602 = N11601 | data_masked[14940];
  assign N11601 = N11600 | data_masked[15068];
  assign N11600 = N11599 | data_masked[15196];
  assign N11599 = N11598 | data_masked[15324];
  assign N11598 = N11597 | data_masked[15452];
  assign N11597 = N11596 | data_masked[15580];
  assign N11596 = N11595 | data_masked[15708];
  assign N11595 = N11594 | data_masked[15836];
  assign N11594 = N11593 | data_masked[15964];
  assign N11593 = N11592 | data_masked[16092];
  assign N11592 = data_masked[16348] | data_masked[16220];
  assign data_o[93] = N11843 | data_masked[93];
  assign N11843 = N11842 | data_masked[221];
  assign N11842 = N11841 | data_masked[349];
  assign N11841 = N11840 | data_masked[477];
  assign N11840 = N11839 | data_masked[605];
  assign N11839 = N11838 | data_masked[733];
  assign N11838 = N11837 | data_masked[861];
  assign N11837 = N11836 | data_masked[989];
  assign N11836 = N11835 | data_masked[1117];
  assign N11835 = N11834 | data_masked[1245];
  assign N11834 = N11833 | data_masked[1373];
  assign N11833 = N11832 | data_masked[1501];
  assign N11832 = N11831 | data_masked[1629];
  assign N11831 = N11830 | data_masked[1757];
  assign N11830 = N11829 | data_masked[1885];
  assign N11829 = N11828 | data_masked[2013];
  assign N11828 = N11827 | data_masked[2141];
  assign N11827 = N11826 | data_masked[2269];
  assign N11826 = N11825 | data_masked[2397];
  assign N11825 = N11824 | data_masked[2525];
  assign N11824 = N11823 | data_masked[2653];
  assign N11823 = N11822 | data_masked[2781];
  assign N11822 = N11821 | data_masked[2909];
  assign N11821 = N11820 | data_masked[3037];
  assign N11820 = N11819 | data_masked[3165];
  assign N11819 = N11818 | data_masked[3293];
  assign N11818 = N11817 | data_masked[3421];
  assign N11817 = N11816 | data_masked[3549];
  assign N11816 = N11815 | data_masked[3677];
  assign N11815 = N11814 | data_masked[3805];
  assign N11814 = N11813 | data_masked[3933];
  assign N11813 = N11812 | data_masked[4061];
  assign N11812 = N11811 | data_masked[4189];
  assign N11811 = N11810 | data_masked[4317];
  assign N11810 = N11809 | data_masked[4445];
  assign N11809 = N11808 | data_masked[4573];
  assign N11808 = N11807 | data_masked[4701];
  assign N11807 = N11806 | data_masked[4829];
  assign N11806 = N11805 | data_masked[4957];
  assign N11805 = N11804 | data_masked[5085];
  assign N11804 = N11803 | data_masked[5213];
  assign N11803 = N11802 | data_masked[5341];
  assign N11802 = N11801 | data_masked[5469];
  assign N11801 = N11800 | data_masked[5597];
  assign N11800 = N11799 | data_masked[5725];
  assign N11799 = N11798 | data_masked[5853];
  assign N11798 = N11797 | data_masked[5981];
  assign N11797 = N11796 | data_masked[6109];
  assign N11796 = N11795 | data_masked[6237];
  assign N11795 = N11794 | data_masked[6365];
  assign N11794 = N11793 | data_masked[6493];
  assign N11793 = N11792 | data_masked[6621];
  assign N11792 = N11791 | data_masked[6749];
  assign N11791 = N11790 | data_masked[6877];
  assign N11790 = N11789 | data_masked[7005];
  assign N11789 = N11788 | data_masked[7133];
  assign N11788 = N11787 | data_masked[7261];
  assign N11787 = N11786 | data_masked[7389];
  assign N11786 = N11785 | data_masked[7517];
  assign N11785 = N11784 | data_masked[7645];
  assign N11784 = N11783 | data_masked[7773];
  assign N11783 = N11782 | data_masked[7901];
  assign N11782 = N11781 | data_masked[8029];
  assign N11781 = N11780 | data_masked[8157];
  assign N11780 = N11779 | data_masked[8285];
  assign N11779 = N11778 | data_masked[8413];
  assign N11778 = N11777 | data_masked[8541];
  assign N11777 = N11776 | data_masked[8669];
  assign N11776 = N11775 | data_masked[8797];
  assign N11775 = N11774 | data_masked[8925];
  assign N11774 = N11773 | data_masked[9053];
  assign N11773 = N11772 | data_masked[9181];
  assign N11772 = N11771 | data_masked[9309];
  assign N11771 = N11770 | data_masked[9437];
  assign N11770 = N11769 | data_masked[9565];
  assign N11769 = N11768 | data_masked[9693];
  assign N11768 = N11767 | data_masked[9821];
  assign N11767 = N11766 | data_masked[9949];
  assign N11766 = N11765 | data_masked[10077];
  assign N11765 = N11764 | data_masked[10205];
  assign N11764 = N11763 | data_masked[10333];
  assign N11763 = N11762 | data_masked[10461];
  assign N11762 = N11761 | data_masked[10589];
  assign N11761 = N11760 | data_masked[10717];
  assign N11760 = N11759 | data_masked[10845];
  assign N11759 = N11758 | data_masked[10973];
  assign N11758 = N11757 | data_masked[11101];
  assign N11757 = N11756 | data_masked[11229];
  assign N11756 = N11755 | data_masked[11357];
  assign N11755 = N11754 | data_masked[11485];
  assign N11754 = N11753 | data_masked[11613];
  assign N11753 = N11752 | data_masked[11741];
  assign N11752 = N11751 | data_masked[11869];
  assign N11751 = N11750 | data_masked[11997];
  assign N11750 = N11749 | data_masked[12125];
  assign N11749 = N11748 | data_masked[12253];
  assign N11748 = N11747 | data_masked[12381];
  assign N11747 = N11746 | data_masked[12509];
  assign N11746 = N11745 | data_masked[12637];
  assign N11745 = N11744 | data_masked[12765];
  assign N11744 = N11743 | data_masked[12893];
  assign N11743 = N11742 | data_masked[13021];
  assign N11742 = N11741 | data_masked[13149];
  assign N11741 = N11740 | data_masked[13277];
  assign N11740 = N11739 | data_masked[13405];
  assign N11739 = N11738 | data_masked[13533];
  assign N11738 = N11737 | data_masked[13661];
  assign N11737 = N11736 | data_masked[13789];
  assign N11736 = N11735 | data_masked[13917];
  assign N11735 = N11734 | data_masked[14045];
  assign N11734 = N11733 | data_masked[14173];
  assign N11733 = N11732 | data_masked[14301];
  assign N11732 = N11731 | data_masked[14429];
  assign N11731 = N11730 | data_masked[14557];
  assign N11730 = N11729 | data_masked[14685];
  assign N11729 = N11728 | data_masked[14813];
  assign N11728 = N11727 | data_masked[14941];
  assign N11727 = N11726 | data_masked[15069];
  assign N11726 = N11725 | data_masked[15197];
  assign N11725 = N11724 | data_masked[15325];
  assign N11724 = N11723 | data_masked[15453];
  assign N11723 = N11722 | data_masked[15581];
  assign N11722 = N11721 | data_masked[15709];
  assign N11721 = N11720 | data_masked[15837];
  assign N11720 = N11719 | data_masked[15965];
  assign N11719 = N11718 | data_masked[16093];
  assign N11718 = data_masked[16349] | data_masked[16221];
  assign data_o[94] = N11969 | data_masked[94];
  assign N11969 = N11968 | data_masked[222];
  assign N11968 = N11967 | data_masked[350];
  assign N11967 = N11966 | data_masked[478];
  assign N11966 = N11965 | data_masked[606];
  assign N11965 = N11964 | data_masked[734];
  assign N11964 = N11963 | data_masked[862];
  assign N11963 = N11962 | data_masked[990];
  assign N11962 = N11961 | data_masked[1118];
  assign N11961 = N11960 | data_masked[1246];
  assign N11960 = N11959 | data_masked[1374];
  assign N11959 = N11958 | data_masked[1502];
  assign N11958 = N11957 | data_masked[1630];
  assign N11957 = N11956 | data_masked[1758];
  assign N11956 = N11955 | data_masked[1886];
  assign N11955 = N11954 | data_masked[2014];
  assign N11954 = N11953 | data_masked[2142];
  assign N11953 = N11952 | data_masked[2270];
  assign N11952 = N11951 | data_masked[2398];
  assign N11951 = N11950 | data_masked[2526];
  assign N11950 = N11949 | data_masked[2654];
  assign N11949 = N11948 | data_masked[2782];
  assign N11948 = N11947 | data_masked[2910];
  assign N11947 = N11946 | data_masked[3038];
  assign N11946 = N11945 | data_masked[3166];
  assign N11945 = N11944 | data_masked[3294];
  assign N11944 = N11943 | data_masked[3422];
  assign N11943 = N11942 | data_masked[3550];
  assign N11942 = N11941 | data_masked[3678];
  assign N11941 = N11940 | data_masked[3806];
  assign N11940 = N11939 | data_masked[3934];
  assign N11939 = N11938 | data_masked[4062];
  assign N11938 = N11937 | data_masked[4190];
  assign N11937 = N11936 | data_masked[4318];
  assign N11936 = N11935 | data_masked[4446];
  assign N11935 = N11934 | data_masked[4574];
  assign N11934 = N11933 | data_masked[4702];
  assign N11933 = N11932 | data_masked[4830];
  assign N11932 = N11931 | data_masked[4958];
  assign N11931 = N11930 | data_masked[5086];
  assign N11930 = N11929 | data_masked[5214];
  assign N11929 = N11928 | data_masked[5342];
  assign N11928 = N11927 | data_masked[5470];
  assign N11927 = N11926 | data_masked[5598];
  assign N11926 = N11925 | data_masked[5726];
  assign N11925 = N11924 | data_masked[5854];
  assign N11924 = N11923 | data_masked[5982];
  assign N11923 = N11922 | data_masked[6110];
  assign N11922 = N11921 | data_masked[6238];
  assign N11921 = N11920 | data_masked[6366];
  assign N11920 = N11919 | data_masked[6494];
  assign N11919 = N11918 | data_masked[6622];
  assign N11918 = N11917 | data_masked[6750];
  assign N11917 = N11916 | data_masked[6878];
  assign N11916 = N11915 | data_masked[7006];
  assign N11915 = N11914 | data_masked[7134];
  assign N11914 = N11913 | data_masked[7262];
  assign N11913 = N11912 | data_masked[7390];
  assign N11912 = N11911 | data_masked[7518];
  assign N11911 = N11910 | data_masked[7646];
  assign N11910 = N11909 | data_masked[7774];
  assign N11909 = N11908 | data_masked[7902];
  assign N11908 = N11907 | data_masked[8030];
  assign N11907 = N11906 | data_masked[8158];
  assign N11906 = N11905 | data_masked[8286];
  assign N11905 = N11904 | data_masked[8414];
  assign N11904 = N11903 | data_masked[8542];
  assign N11903 = N11902 | data_masked[8670];
  assign N11902 = N11901 | data_masked[8798];
  assign N11901 = N11900 | data_masked[8926];
  assign N11900 = N11899 | data_masked[9054];
  assign N11899 = N11898 | data_masked[9182];
  assign N11898 = N11897 | data_masked[9310];
  assign N11897 = N11896 | data_masked[9438];
  assign N11896 = N11895 | data_masked[9566];
  assign N11895 = N11894 | data_masked[9694];
  assign N11894 = N11893 | data_masked[9822];
  assign N11893 = N11892 | data_masked[9950];
  assign N11892 = N11891 | data_masked[10078];
  assign N11891 = N11890 | data_masked[10206];
  assign N11890 = N11889 | data_masked[10334];
  assign N11889 = N11888 | data_masked[10462];
  assign N11888 = N11887 | data_masked[10590];
  assign N11887 = N11886 | data_masked[10718];
  assign N11886 = N11885 | data_masked[10846];
  assign N11885 = N11884 | data_masked[10974];
  assign N11884 = N11883 | data_masked[11102];
  assign N11883 = N11882 | data_masked[11230];
  assign N11882 = N11881 | data_masked[11358];
  assign N11881 = N11880 | data_masked[11486];
  assign N11880 = N11879 | data_masked[11614];
  assign N11879 = N11878 | data_masked[11742];
  assign N11878 = N11877 | data_masked[11870];
  assign N11877 = N11876 | data_masked[11998];
  assign N11876 = N11875 | data_masked[12126];
  assign N11875 = N11874 | data_masked[12254];
  assign N11874 = N11873 | data_masked[12382];
  assign N11873 = N11872 | data_masked[12510];
  assign N11872 = N11871 | data_masked[12638];
  assign N11871 = N11870 | data_masked[12766];
  assign N11870 = N11869 | data_masked[12894];
  assign N11869 = N11868 | data_masked[13022];
  assign N11868 = N11867 | data_masked[13150];
  assign N11867 = N11866 | data_masked[13278];
  assign N11866 = N11865 | data_masked[13406];
  assign N11865 = N11864 | data_masked[13534];
  assign N11864 = N11863 | data_masked[13662];
  assign N11863 = N11862 | data_masked[13790];
  assign N11862 = N11861 | data_masked[13918];
  assign N11861 = N11860 | data_masked[14046];
  assign N11860 = N11859 | data_masked[14174];
  assign N11859 = N11858 | data_masked[14302];
  assign N11858 = N11857 | data_masked[14430];
  assign N11857 = N11856 | data_masked[14558];
  assign N11856 = N11855 | data_masked[14686];
  assign N11855 = N11854 | data_masked[14814];
  assign N11854 = N11853 | data_masked[14942];
  assign N11853 = N11852 | data_masked[15070];
  assign N11852 = N11851 | data_masked[15198];
  assign N11851 = N11850 | data_masked[15326];
  assign N11850 = N11849 | data_masked[15454];
  assign N11849 = N11848 | data_masked[15582];
  assign N11848 = N11847 | data_masked[15710];
  assign N11847 = N11846 | data_masked[15838];
  assign N11846 = N11845 | data_masked[15966];
  assign N11845 = N11844 | data_masked[16094];
  assign N11844 = data_masked[16350] | data_masked[16222];
  assign data_o[95] = N12095 | data_masked[95];
  assign N12095 = N12094 | data_masked[223];
  assign N12094 = N12093 | data_masked[351];
  assign N12093 = N12092 | data_masked[479];
  assign N12092 = N12091 | data_masked[607];
  assign N12091 = N12090 | data_masked[735];
  assign N12090 = N12089 | data_masked[863];
  assign N12089 = N12088 | data_masked[991];
  assign N12088 = N12087 | data_masked[1119];
  assign N12087 = N12086 | data_masked[1247];
  assign N12086 = N12085 | data_masked[1375];
  assign N12085 = N12084 | data_masked[1503];
  assign N12084 = N12083 | data_masked[1631];
  assign N12083 = N12082 | data_masked[1759];
  assign N12082 = N12081 | data_masked[1887];
  assign N12081 = N12080 | data_masked[2015];
  assign N12080 = N12079 | data_masked[2143];
  assign N12079 = N12078 | data_masked[2271];
  assign N12078 = N12077 | data_masked[2399];
  assign N12077 = N12076 | data_masked[2527];
  assign N12076 = N12075 | data_masked[2655];
  assign N12075 = N12074 | data_masked[2783];
  assign N12074 = N12073 | data_masked[2911];
  assign N12073 = N12072 | data_masked[3039];
  assign N12072 = N12071 | data_masked[3167];
  assign N12071 = N12070 | data_masked[3295];
  assign N12070 = N12069 | data_masked[3423];
  assign N12069 = N12068 | data_masked[3551];
  assign N12068 = N12067 | data_masked[3679];
  assign N12067 = N12066 | data_masked[3807];
  assign N12066 = N12065 | data_masked[3935];
  assign N12065 = N12064 | data_masked[4063];
  assign N12064 = N12063 | data_masked[4191];
  assign N12063 = N12062 | data_masked[4319];
  assign N12062 = N12061 | data_masked[4447];
  assign N12061 = N12060 | data_masked[4575];
  assign N12060 = N12059 | data_masked[4703];
  assign N12059 = N12058 | data_masked[4831];
  assign N12058 = N12057 | data_masked[4959];
  assign N12057 = N12056 | data_masked[5087];
  assign N12056 = N12055 | data_masked[5215];
  assign N12055 = N12054 | data_masked[5343];
  assign N12054 = N12053 | data_masked[5471];
  assign N12053 = N12052 | data_masked[5599];
  assign N12052 = N12051 | data_masked[5727];
  assign N12051 = N12050 | data_masked[5855];
  assign N12050 = N12049 | data_masked[5983];
  assign N12049 = N12048 | data_masked[6111];
  assign N12048 = N12047 | data_masked[6239];
  assign N12047 = N12046 | data_masked[6367];
  assign N12046 = N12045 | data_masked[6495];
  assign N12045 = N12044 | data_masked[6623];
  assign N12044 = N12043 | data_masked[6751];
  assign N12043 = N12042 | data_masked[6879];
  assign N12042 = N12041 | data_masked[7007];
  assign N12041 = N12040 | data_masked[7135];
  assign N12040 = N12039 | data_masked[7263];
  assign N12039 = N12038 | data_masked[7391];
  assign N12038 = N12037 | data_masked[7519];
  assign N12037 = N12036 | data_masked[7647];
  assign N12036 = N12035 | data_masked[7775];
  assign N12035 = N12034 | data_masked[7903];
  assign N12034 = N12033 | data_masked[8031];
  assign N12033 = N12032 | data_masked[8159];
  assign N12032 = N12031 | data_masked[8287];
  assign N12031 = N12030 | data_masked[8415];
  assign N12030 = N12029 | data_masked[8543];
  assign N12029 = N12028 | data_masked[8671];
  assign N12028 = N12027 | data_masked[8799];
  assign N12027 = N12026 | data_masked[8927];
  assign N12026 = N12025 | data_masked[9055];
  assign N12025 = N12024 | data_masked[9183];
  assign N12024 = N12023 | data_masked[9311];
  assign N12023 = N12022 | data_masked[9439];
  assign N12022 = N12021 | data_masked[9567];
  assign N12021 = N12020 | data_masked[9695];
  assign N12020 = N12019 | data_masked[9823];
  assign N12019 = N12018 | data_masked[9951];
  assign N12018 = N12017 | data_masked[10079];
  assign N12017 = N12016 | data_masked[10207];
  assign N12016 = N12015 | data_masked[10335];
  assign N12015 = N12014 | data_masked[10463];
  assign N12014 = N12013 | data_masked[10591];
  assign N12013 = N12012 | data_masked[10719];
  assign N12012 = N12011 | data_masked[10847];
  assign N12011 = N12010 | data_masked[10975];
  assign N12010 = N12009 | data_masked[11103];
  assign N12009 = N12008 | data_masked[11231];
  assign N12008 = N12007 | data_masked[11359];
  assign N12007 = N12006 | data_masked[11487];
  assign N12006 = N12005 | data_masked[11615];
  assign N12005 = N12004 | data_masked[11743];
  assign N12004 = N12003 | data_masked[11871];
  assign N12003 = N12002 | data_masked[11999];
  assign N12002 = N12001 | data_masked[12127];
  assign N12001 = N12000 | data_masked[12255];
  assign N12000 = N11999 | data_masked[12383];
  assign N11999 = N11998 | data_masked[12511];
  assign N11998 = N11997 | data_masked[12639];
  assign N11997 = N11996 | data_masked[12767];
  assign N11996 = N11995 | data_masked[12895];
  assign N11995 = N11994 | data_masked[13023];
  assign N11994 = N11993 | data_masked[13151];
  assign N11993 = N11992 | data_masked[13279];
  assign N11992 = N11991 | data_masked[13407];
  assign N11991 = N11990 | data_masked[13535];
  assign N11990 = N11989 | data_masked[13663];
  assign N11989 = N11988 | data_masked[13791];
  assign N11988 = N11987 | data_masked[13919];
  assign N11987 = N11986 | data_masked[14047];
  assign N11986 = N11985 | data_masked[14175];
  assign N11985 = N11984 | data_masked[14303];
  assign N11984 = N11983 | data_masked[14431];
  assign N11983 = N11982 | data_masked[14559];
  assign N11982 = N11981 | data_masked[14687];
  assign N11981 = N11980 | data_masked[14815];
  assign N11980 = N11979 | data_masked[14943];
  assign N11979 = N11978 | data_masked[15071];
  assign N11978 = N11977 | data_masked[15199];
  assign N11977 = N11976 | data_masked[15327];
  assign N11976 = N11975 | data_masked[15455];
  assign N11975 = N11974 | data_masked[15583];
  assign N11974 = N11973 | data_masked[15711];
  assign N11973 = N11972 | data_masked[15839];
  assign N11972 = N11971 | data_masked[15967];
  assign N11971 = N11970 | data_masked[16095];
  assign N11970 = data_masked[16351] | data_masked[16223];
  assign data_o[96] = N12221 | data_masked[96];
  assign N12221 = N12220 | data_masked[224];
  assign N12220 = N12219 | data_masked[352];
  assign N12219 = N12218 | data_masked[480];
  assign N12218 = N12217 | data_masked[608];
  assign N12217 = N12216 | data_masked[736];
  assign N12216 = N12215 | data_masked[864];
  assign N12215 = N12214 | data_masked[992];
  assign N12214 = N12213 | data_masked[1120];
  assign N12213 = N12212 | data_masked[1248];
  assign N12212 = N12211 | data_masked[1376];
  assign N12211 = N12210 | data_masked[1504];
  assign N12210 = N12209 | data_masked[1632];
  assign N12209 = N12208 | data_masked[1760];
  assign N12208 = N12207 | data_masked[1888];
  assign N12207 = N12206 | data_masked[2016];
  assign N12206 = N12205 | data_masked[2144];
  assign N12205 = N12204 | data_masked[2272];
  assign N12204 = N12203 | data_masked[2400];
  assign N12203 = N12202 | data_masked[2528];
  assign N12202 = N12201 | data_masked[2656];
  assign N12201 = N12200 | data_masked[2784];
  assign N12200 = N12199 | data_masked[2912];
  assign N12199 = N12198 | data_masked[3040];
  assign N12198 = N12197 | data_masked[3168];
  assign N12197 = N12196 | data_masked[3296];
  assign N12196 = N12195 | data_masked[3424];
  assign N12195 = N12194 | data_masked[3552];
  assign N12194 = N12193 | data_masked[3680];
  assign N12193 = N12192 | data_masked[3808];
  assign N12192 = N12191 | data_masked[3936];
  assign N12191 = N12190 | data_masked[4064];
  assign N12190 = N12189 | data_masked[4192];
  assign N12189 = N12188 | data_masked[4320];
  assign N12188 = N12187 | data_masked[4448];
  assign N12187 = N12186 | data_masked[4576];
  assign N12186 = N12185 | data_masked[4704];
  assign N12185 = N12184 | data_masked[4832];
  assign N12184 = N12183 | data_masked[4960];
  assign N12183 = N12182 | data_masked[5088];
  assign N12182 = N12181 | data_masked[5216];
  assign N12181 = N12180 | data_masked[5344];
  assign N12180 = N12179 | data_masked[5472];
  assign N12179 = N12178 | data_masked[5600];
  assign N12178 = N12177 | data_masked[5728];
  assign N12177 = N12176 | data_masked[5856];
  assign N12176 = N12175 | data_masked[5984];
  assign N12175 = N12174 | data_masked[6112];
  assign N12174 = N12173 | data_masked[6240];
  assign N12173 = N12172 | data_masked[6368];
  assign N12172 = N12171 | data_masked[6496];
  assign N12171 = N12170 | data_masked[6624];
  assign N12170 = N12169 | data_masked[6752];
  assign N12169 = N12168 | data_masked[6880];
  assign N12168 = N12167 | data_masked[7008];
  assign N12167 = N12166 | data_masked[7136];
  assign N12166 = N12165 | data_masked[7264];
  assign N12165 = N12164 | data_masked[7392];
  assign N12164 = N12163 | data_masked[7520];
  assign N12163 = N12162 | data_masked[7648];
  assign N12162 = N12161 | data_masked[7776];
  assign N12161 = N12160 | data_masked[7904];
  assign N12160 = N12159 | data_masked[8032];
  assign N12159 = N12158 | data_masked[8160];
  assign N12158 = N12157 | data_masked[8288];
  assign N12157 = N12156 | data_masked[8416];
  assign N12156 = N12155 | data_masked[8544];
  assign N12155 = N12154 | data_masked[8672];
  assign N12154 = N12153 | data_masked[8800];
  assign N12153 = N12152 | data_masked[8928];
  assign N12152 = N12151 | data_masked[9056];
  assign N12151 = N12150 | data_masked[9184];
  assign N12150 = N12149 | data_masked[9312];
  assign N12149 = N12148 | data_masked[9440];
  assign N12148 = N12147 | data_masked[9568];
  assign N12147 = N12146 | data_masked[9696];
  assign N12146 = N12145 | data_masked[9824];
  assign N12145 = N12144 | data_masked[9952];
  assign N12144 = N12143 | data_masked[10080];
  assign N12143 = N12142 | data_masked[10208];
  assign N12142 = N12141 | data_masked[10336];
  assign N12141 = N12140 | data_masked[10464];
  assign N12140 = N12139 | data_masked[10592];
  assign N12139 = N12138 | data_masked[10720];
  assign N12138 = N12137 | data_masked[10848];
  assign N12137 = N12136 | data_masked[10976];
  assign N12136 = N12135 | data_masked[11104];
  assign N12135 = N12134 | data_masked[11232];
  assign N12134 = N12133 | data_masked[11360];
  assign N12133 = N12132 | data_masked[11488];
  assign N12132 = N12131 | data_masked[11616];
  assign N12131 = N12130 | data_masked[11744];
  assign N12130 = N12129 | data_masked[11872];
  assign N12129 = N12128 | data_masked[12000];
  assign N12128 = N12127 | data_masked[12128];
  assign N12127 = N12126 | data_masked[12256];
  assign N12126 = N12125 | data_masked[12384];
  assign N12125 = N12124 | data_masked[12512];
  assign N12124 = N12123 | data_masked[12640];
  assign N12123 = N12122 | data_masked[12768];
  assign N12122 = N12121 | data_masked[12896];
  assign N12121 = N12120 | data_masked[13024];
  assign N12120 = N12119 | data_masked[13152];
  assign N12119 = N12118 | data_masked[13280];
  assign N12118 = N12117 | data_masked[13408];
  assign N12117 = N12116 | data_masked[13536];
  assign N12116 = N12115 | data_masked[13664];
  assign N12115 = N12114 | data_masked[13792];
  assign N12114 = N12113 | data_masked[13920];
  assign N12113 = N12112 | data_masked[14048];
  assign N12112 = N12111 | data_masked[14176];
  assign N12111 = N12110 | data_masked[14304];
  assign N12110 = N12109 | data_masked[14432];
  assign N12109 = N12108 | data_masked[14560];
  assign N12108 = N12107 | data_masked[14688];
  assign N12107 = N12106 | data_masked[14816];
  assign N12106 = N12105 | data_masked[14944];
  assign N12105 = N12104 | data_masked[15072];
  assign N12104 = N12103 | data_masked[15200];
  assign N12103 = N12102 | data_masked[15328];
  assign N12102 = N12101 | data_masked[15456];
  assign N12101 = N12100 | data_masked[15584];
  assign N12100 = N12099 | data_masked[15712];
  assign N12099 = N12098 | data_masked[15840];
  assign N12098 = N12097 | data_masked[15968];
  assign N12097 = N12096 | data_masked[16096];
  assign N12096 = data_masked[16352] | data_masked[16224];
  assign data_o[97] = N12347 | data_masked[97];
  assign N12347 = N12346 | data_masked[225];
  assign N12346 = N12345 | data_masked[353];
  assign N12345 = N12344 | data_masked[481];
  assign N12344 = N12343 | data_masked[609];
  assign N12343 = N12342 | data_masked[737];
  assign N12342 = N12341 | data_masked[865];
  assign N12341 = N12340 | data_masked[993];
  assign N12340 = N12339 | data_masked[1121];
  assign N12339 = N12338 | data_masked[1249];
  assign N12338 = N12337 | data_masked[1377];
  assign N12337 = N12336 | data_masked[1505];
  assign N12336 = N12335 | data_masked[1633];
  assign N12335 = N12334 | data_masked[1761];
  assign N12334 = N12333 | data_masked[1889];
  assign N12333 = N12332 | data_masked[2017];
  assign N12332 = N12331 | data_masked[2145];
  assign N12331 = N12330 | data_masked[2273];
  assign N12330 = N12329 | data_masked[2401];
  assign N12329 = N12328 | data_masked[2529];
  assign N12328 = N12327 | data_masked[2657];
  assign N12327 = N12326 | data_masked[2785];
  assign N12326 = N12325 | data_masked[2913];
  assign N12325 = N12324 | data_masked[3041];
  assign N12324 = N12323 | data_masked[3169];
  assign N12323 = N12322 | data_masked[3297];
  assign N12322 = N12321 | data_masked[3425];
  assign N12321 = N12320 | data_masked[3553];
  assign N12320 = N12319 | data_masked[3681];
  assign N12319 = N12318 | data_masked[3809];
  assign N12318 = N12317 | data_masked[3937];
  assign N12317 = N12316 | data_masked[4065];
  assign N12316 = N12315 | data_masked[4193];
  assign N12315 = N12314 | data_masked[4321];
  assign N12314 = N12313 | data_masked[4449];
  assign N12313 = N12312 | data_masked[4577];
  assign N12312 = N12311 | data_masked[4705];
  assign N12311 = N12310 | data_masked[4833];
  assign N12310 = N12309 | data_masked[4961];
  assign N12309 = N12308 | data_masked[5089];
  assign N12308 = N12307 | data_masked[5217];
  assign N12307 = N12306 | data_masked[5345];
  assign N12306 = N12305 | data_masked[5473];
  assign N12305 = N12304 | data_masked[5601];
  assign N12304 = N12303 | data_masked[5729];
  assign N12303 = N12302 | data_masked[5857];
  assign N12302 = N12301 | data_masked[5985];
  assign N12301 = N12300 | data_masked[6113];
  assign N12300 = N12299 | data_masked[6241];
  assign N12299 = N12298 | data_masked[6369];
  assign N12298 = N12297 | data_masked[6497];
  assign N12297 = N12296 | data_masked[6625];
  assign N12296 = N12295 | data_masked[6753];
  assign N12295 = N12294 | data_masked[6881];
  assign N12294 = N12293 | data_masked[7009];
  assign N12293 = N12292 | data_masked[7137];
  assign N12292 = N12291 | data_masked[7265];
  assign N12291 = N12290 | data_masked[7393];
  assign N12290 = N12289 | data_masked[7521];
  assign N12289 = N12288 | data_masked[7649];
  assign N12288 = N12287 | data_masked[7777];
  assign N12287 = N12286 | data_masked[7905];
  assign N12286 = N12285 | data_masked[8033];
  assign N12285 = N12284 | data_masked[8161];
  assign N12284 = N12283 | data_masked[8289];
  assign N12283 = N12282 | data_masked[8417];
  assign N12282 = N12281 | data_masked[8545];
  assign N12281 = N12280 | data_masked[8673];
  assign N12280 = N12279 | data_masked[8801];
  assign N12279 = N12278 | data_masked[8929];
  assign N12278 = N12277 | data_masked[9057];
  assign N12277 = N12276 | data_masked[9185];
  assign N12276 = N12275 | data_masked[9313];
  assign N12275 = N12274 | data_masked[9441];
  assign N12274 = N12273 | data_masked[9569];
  assign N12273 = N12272 | data_masked[9697];
  assign N12272 = N12271 | data_masked[9825];
  assign N12271 = N12270 | data_masked[9953];
  assign N12270 = N12269 | data_masked[10081];
  assign N12269 = N12268 | data_masked[10209];
  assign N12268 = N12267 | data_masked[10337];
  assign N12267 = N12266 | data_masked[10465];
  assign N12266 = N12265 | data_masked[10593];
  assign N12265 = N12264 | data_masked[10721];
  assign N12264 = N12263 | data_masked[10849];
  assign N12263 = N12262 | data_masked[10977];
  assign N12262 = N12261 | data_masked[11105];
  assign N12261 = N12260 | data_masked[11233];
  assign N12260 = N12259 | data_masked[11361];
  assign N12259 = N12258 | data_masked[11489];
  assign N12258 = N12257 | data_masked[11617];
  assign N12257 = N12256 | data_masked[11745];
  assign N12256 = N12255 | data_masked[11873];
  assign N12255 = N12254 | data_masked[12001];
  assign N12254 = N12253 | data_masked[12129];
  assign N12253 = N12252 | data_masked[12257];
  assign N12252 = N12251 | data_masked[12385];
  assign N12251 = N12250 | data_masked[12513];
  assign N12250 = N12249 | data_masked[12641];
  assign N12249 = N12248 | data_masked[12769];
  assign N12248 = N12247 | data_masked[12897];
  assign N12247 = N12246 | data_masked[13025];
  assign N12246 = N12245 | data_masked[13153];
  assign N12245 = N12244 | data_masked[13281];
  assign N12244 = N12243 | data_masked[13409];
  assign N12243 = N12242 | data_masked[13537];
  assign N12242 = N12241 | data_masked[13665];
  assign N12241 = N12240 | data_masked[13793];
  assign N12240 = N12239 | data_masked[13921];
  assign N12239 = N12238 | data_masked[14049];
  assign N12238 = N12237 | data_masked[14177];
  assign N12237 = N12236 | data_masked[14305];
  assign N12236 = N12235 | data_masked[14433];
  assign N12235 = N12234 | data_masked[14561];
  assign N12234 = N12233 | data_masked[14689];
  assign N12233 = N12232 | data_masked[14817];
  assign N12232 = N12231 | data_masked[14945];
  assign N12231 = N12230 | data_masked[15073];
  assign N12230 = N12229 | data_masked[15201];
  assign N12229 = N12228 | data_masked[15329];
  assign N12228 = N12227 | data_masked[15457];
  assign N12227 = N12226 | data_masked[15585];
  assign N12226 = N12225 | data_masked[15713];
  assign N12225 = N12224 | data_masked[15841];
  assign N12224 = N12223 | data_masked[15969];
  assign N12223 = N12222 | data_masked[16097];
  assign N12222 = data_masked[16353] | data_masked[16225];
  assign data_o[98] = N12473 | data_masked[98];
  assign N12473 = N12472 | data_masked[226];
  assign N12472 = N12471 | data_masked[354];
  assign N12471 = N12470 | data_masked[482];
  assign N12470 = N12469 | data_masked[610];
  assign N12469 = N12468 | data_masked[738];
  assign N12468 = N12467 | data_masked[866];
  assign N12467 = N12466 | data_masked[994];
  assign N12466 = N12465 | data_masked[1122];
  assign N12465 = N12464 | data_masked[1250];
  assign N12464 = N12463 | data_masked[1378];
  assign N12463 = N12462 | data_masked[1506];
  assign N12462 = N12461 | data_masked[1634];
  assign N12461 = N12460 | data_masked[1762];
  assign N12460 = N12459 | data_masked[1890];
  assign N12459 = N12458 | data_masked[2018];
  assign N12458 = N12457 | data_masked[2146];
  assign N12457 = N12456 | data_masked[2274];
  assign N12456 = N12455 | data_masked[2402];
  assign N12455 = N12454 | data_masked[2530];
  assign N12454 = N12453 | data_masked[2658];
  assign N12453 = N12452 | data_masked[2786];
  assign N12452 = N12451 | data_masked[2914];
  assign N12451 = N12450 | data_masked[3042];
  assign N12450 = N12449 | data_masked[3170];
  assign N12449 = N12448 | data_masked[3298];
  assign N12448 = N12447 | data_masked[3426];
  assign N12447 = N12446 | data_masked[3554];
  assign N12446 = N12445 | data_masked[3682];
  assign N12445 = N12444 | data_masked[3810];
  assign N12444 = N12443 | data_masked[3938];
  assign N12443 = N12442 | data_masked[4066];
  assign N12442 = N12441 | data_masked[4194];
  assign N12441 = N12440 | data_masked[4322];
  assign N12440 = N12439 | data_masked[4450];
  assign N12439 = N12438 | data_masked[4578];
  assign N12438 = N12437 | data_masked[4706];
  assign N12437 = N12436 | data_masked[4834];
  assign N12436 = N12435 | data_masked[4962];
  assign N12435 = N12434 | data_masked[5090];
  assign N12434 = N12433 | data_masked[5218];
  assign N12433 = N12432 | data_masked[5346];
  assign N12432 = N12431 | data_masked[5474];
  assign N12431 = N12430 | data_masked[5602];
  assign N12430 = N12429 | data_masked[5730];
  assign N12429 = N12428 | data_masked[5858];
  assign N12428 = N12427 | data_masked[5986];
  assign N12427 = N12426 | data_masked[6114];
  assign N12426 = N12425 | data_masked[6242];
  assign N12425 = N12424 | data_masked[6370];
  assign N12424 = N12423 | data_masked[6498];
  assign N12423 = N12422 | data_masked[6626];
  assign N12422 = N12421 | data_masked[6754];
  assign N12421 = N12420 | data_masked[6882];
  assign N12420 = N12419 | data_masked[7010];
  assign N12419 = N12418 | data_masked[7138];
  assign N12418 = N12417 | data_masked[7266];
  assign N12417 = N12416 | data_masked[7394];
  assign N12416 = N12415 | data_masked[7522];
  assign N12415 = N12414 | data_masked[7650];
  assign N12414 = N12413 | data_masked[7778];
  assign N12413 = N12412 | data_masked[7906];
  assign N12412 = N12411 | data_masked[8034];
  assign N12411 = N12410 | data_masked[8162];
  assign N12410 = N12409 | data_masked[8290];
  assign N12409 = N12408 | data_masked[8418];
  assign N12408 = N12407 | data_masked[8546];
  assign N12407 = N12406 | data_masked[8674];
  assign N12406 = N12405 | data_masked[8802];
  assign N12405 = N12404 | data_masked[8930];
  assign N12404 = N12403 | data_masked[9058];
  assign N12403 = N12402 | data_masked[9186];
  assign N12402 = N12401 | data_masked[9314];
  assign N12401 = N12400 | data_masked[9442];
  assign N12400 = N12399 | data_masked[9570];
  assign N12399 = N12398 | data_masked[9698];
  assign N12398 = N12397 | data_masked[9826];
  assign N12397 = N12396 | data_masked[9954];
  assign N12396 = N12395 | data_masked[10082];
  assign N12395 = N12394 | data_masked[10210];
  assign N12394 = N12393 | data_masked[10338];
  assign N12393 = N12392 | data_masked[10466];
  assign N12392 = N12391 | data_masked[10594];
  assign N12391 = N12390 | data_masked[10722];
  assign N12390 = N12389 | data_masked[10850];
  assign N12389 = N12388 | data_masked[10978];
  assign N12388 = N12387 | data_masked[11106];
  assign N12387 = N12386 | data_masked[11234];
  assign N12386 = N12385 | data_masked[11362];
  assign N12385 = N12384 | data_masked[11490];
  assign N12384 = N12383 | data_masked[11618];
  assign N12383 = N12382 | data_masked[11746];
  assign N12382 = N12381 | data_masked[11874];
  assign N12381 = N12380 | data_masked[12002];
  assign N12380 = N12379 | data_masked[12130];
  assign N12379 = N12378 | data_masked[12258];
  assign N12378 = N12377 | data_masked[12386];
  assign N12377 = N12376 | data_masked[12514];
  assign N12376 = N12375 | data_masked[12642];
  assign N12375 = N12374 | data_masked[12770];
  assign N12374 = N12373 | data_masked[12898];
  assign N12373 = N12372 | data_masked[13026];
  assign N12372 = N12371 | data_masked[13154];
  assign N12371 = N12370 | data_masked[13282];
  assign N12370 = N12369 | data_masked[13410];
  assign N12369 = N12368 | data_masked[13538];
  assign N12368 = N12367 | data_masked[13666];
  assign N12367 = N12366 | data_masked[13794];
  assign N12366 = N12365 | data_masked[13922];
  assign N12365 = N12364 | data_masked[14050];
  assign N12364 = N12363 | data_masked[14178];
  assign N12363 = N12362 | data_masked[14306];
  assign N12362 = N12361 | data_masked[14434];
  assign N12361 = N12360 | data_masked[14562];
  assign N12360 = N12359 | data_masked[14690];
  assign N12359 = N12358 | data_masked[14818];
  assign N12358 = N12357 | data_masked[14946];
  assign N12357 = N12356 | data_masked[15074];
  assign N12356 = N12355 | data_masked[15202];
  assign N12355 = N12354 | data_masked[15330];
  assign N12354 = N12353 | data_masked[15458];
  assign N12353 = N12352 | data_masked[15586];
  assign N12352 = N12351 | data_masked[15714];
  assign N12351 = N12350 | data_masked[15842];
  assign N12350 = N12349 | data_masked[15970];
  assign N12349 = N12348 | data_masked[16098];
  assign N12348 = data_masked[16354] | data_masked[16226];
  assign data_o[99] = N12599 | data_masked[99];
  assign N12599 = N12598 | data_masked[227];
  assign N12598 = N12597 | data_masked[355];
  assign N12597 = N12596 | data_masked[483];
  assign N12596 = N12595 | data_masked[611];
  assign N12595 = N12594 | data_masked[739];
  assign N12594 = N12593 | data_masked[867];
  assign N12593 = N12592 | data_masked[995];
  assign N12592 = N12591 | data_masked[1123];
  assign N12591 = N12590 | data_masked[1251];
  assign N12590 = N12589 | data_masked[1379];
  assign N12589 = N12588 | data_masked[1507];
  assign N12588 = N12587 | data_masked[1635];
  assign N12587 = N12586 | data_masked[1763];
  assign N12586 = N12585 | data_masked[1891];
  assign N12585 = N12584 | data_masked[2019];
  assign N12584 = N12583 | data_masked[2147];
  assign N12583 = N12582 | data_masked[2275];
  assign N12582 = N12581 | data_masked[2403];
  assign N12581 = N12580 | data_masked[2531];
  assign N12580 = N12579 | data_masked[2659];
  assign N12579 = N12578 | data_masked[2787];
  assign N12578 = N12577 | data_masked[2915];
  assign N12577 = N12576 | data_masked[3043];
  assign N12576 = N12575 | data_masked[3171];
  assign N12575 = N12574 | data_masked[3299];
  assign N12574 = N12573 | data_masked[3427];
  assign N12573 = N12572 | data_masked[3555];
  assign N12572 = N12571 | data_masked[3683];
  assign N12571 = N12570 | data_masked[3811];
  assign N12570 = N12569 | data_masked[3939];
  assign N12569 = N12568 | data_masked[4067];
  assign N12568 = N12567 | data_masked[4195];
  assign N12567 = N12566 | data_masked[4323];
  assign N12566 = N12565 | data_masked[4451];
  assign N12565 = N12564 | data_masked[4579];
  assign N12564 = N12563 | data_masked[4707];
  assign N12563 = N12562 | data_masked[4835];
  assign N12562 = N12561 | data_masked[4963];
  assign N12561 = N12560 | data_masked[5091];
  assign N12560 = N12559 | data_masked[5219];
  assign N12559 = N12558 | data_masked[5347];
  assign N12558 = N12557 | data_masked[5475];
  assign N12557 = N12556 | data_masked[5603];
  assign N12556 = N12555 | data_masked[5731];
  assign N12555 = N12554 | data_masked[5859];
  assign N12554 = N12553 | data_masked[5987];
  assign N12553 = N12552 | data_masked[6115];
  assign N12552 = N12551 | data_masked[6243];
  assign N12551 = N12550 | data_masked[6371];
  assign N12550 = N12549 | data_masked[6499];
  assign N12549 = N12548 | data_masked[6627];
  assign N12548 = N12547 | data_masked[6755];
  assign N12547 = N12546 | data_masked[6883];
  assign N12546 = N12545 | data_masked[7011];
  assign N12545 = N12544 | data_masked[7139];
  assign N12544 = N12543 | data_masked[7267];
  assign N12543 = N12542 | data_masked[7395];
  assign N12542 = N12541 | data_masked[7523];
  assign N12541 = N12540 | data_masked[7651];
  assign N12540 = N12539 | data_masked[7779];
  assign N12539 = N12538 | data_masked[7907];
  assign N12538 = N12537 | data_masked[8035];
  assign N12537 = N12536 | data_masked[8163];
  assign N12536 = N12535 | data_masked[8291];
  assign N12535 = N12534 | data_masked[8419];
  assign N12534 = N12533 | data_masked[8547];
  assign N12533 = N12532 | data_masked[8675];
  assign N12532 = N12531 | data_masked[8803];
  assign N12531 = N12530 | data_masked[8931];
  assign N12530 = N12529 | data_masked[9059];
  assign N12529 = N12528 | data_masked[9187];
  assign N12528 = N12527 | data_masked[9315];
  assign N12527 = N12526 | data_masked[9443];
  assign N12526 = N12525 | data_masked[9571];
  assign N12525 = N12524 | data_masked[9699];
  assign N12524 = N12523 | data_masked[9827];
  assign N12523 = N12522 | data_masked[9955];
  assign N12522 = N12521 | data_masked[10083];
  assign N12521 = N12520 | data_masked[10211];
  assign N12520 = N12519 | data_masked[10339];
  assign N12519 = N12518 | data_masked[10467];
  assign N12518 = N12517 | data_masked[10595];
  assign N12517 = N12516 | data_masked[10723];
  assign N12516 = N12515 | data_masked[10851];
  assign N12515 = N12514 | data_masked[10979];
  assign N12514 = N12513 | data_masked[11107];
  assign N12513 = N12512 | data_masked[11235];
  assign N12512 = N12511 | data_masked[11363];
  assign N12511 = N12510 | data_masked[11491];
  assign N12510 = N12509 | data_masked[11619];
  assign N12509 = N12508 | data_masked[11747];
  assign N12508 = N12507 | data_masked[11875];
  assign N12507 = N12506 | data_masked[12003];
  assign N12506 = N12505 | data_masked[12131];
  assign N12505 = N12504 | data_masked[12259];
  assign N12504 = N12503 | data_masked[12387];
  assign N12503 = N12502 | data_masked[12515];
  assign N12502 = N12501 | data_masked[12643];
  assign N12501 = N12500 | data_masked[12771];
  assign N12500 = N12499 | data_masked[12899];
  assign N12499 = N12498 | data_masked[13027];
  assign N12498 = N12497 | data_masked[13155];
  assign N12497 = N12496 | data_masked[13283];
  assign N12496 = N12495 | data_masked[13411];
  assign N12495 = N12494 | data_masked[13539];
  assign N12494 = N12493 | data_masked[13667];
  assign N12493 = N12492 | data_masked[13795];
  assign N12492 = N12491 | data_masked[13923];
  assign N12491 = N12490 | data_masked[14051];
  assign N12490 = N12489 | data_masked[14179];
  assign N12489 = N12488 | data_masked[14307];
  assign N12488 = N12487 | data_masked[14435];
  assign N12487 = N12486 | data_masked[14563];
  assign N12486 = N12485 | data_masked[14691];
  assign N12485 = N12484 | data_masked[14819];
  assign N12484 = N12483 | data_masked[14947];
  assign N12483 = N12482 | data_masked[15075];
  assign N12482 = N12481 | data_masked[15203];
  assign N12481 = N12480 | data_masked[15331];
  assign N12480 = N12479 | data_masked[15459];
  assign N12479 = N12478 | data_masked[15587];
  assign N12478 = N12477 | data_masked[15715];
  assign N12477 = N12476 | data_masked[15843];
  assign N12476 = N12475 | data_masked[15971];
  assign N12475 = N12474 | data_masked[16099];
  assign N12474 = data_masked[16355] | data_masked[16227];
  assign data_o[100] = N12725 | data_masked[100];
  assign N12725 = N12724 | data_masked[228];
  assign N12724 = N12723 | data_masked[356];
  assign N12723 = N12722 | data_masked[484];
  assign N12722 = N12721 | data_masked[612];
  assign N12721 = N12720 | data_masked[740];
  assign N12720 = N12719 | data_masked[868];
  assign N12719 = N12718 | data_masked[996];
  assign N12718 = N12717 | data_masked[1124];
  assign N12717 = N12716 | data_masked[1252];
  assign N12716 = N12715 | data_masked[1380];
  assign N12715 = N12714 | data_masked[1508];
  assign N12714 = N12713 | data_masked[1636];
  assign N12713 = N12712 | data_masked[1764];
  assign N12712 = N12711 | data_masked[1892];
  assign N12711 = N12710 | data_masked[2020];
  assign N12710 = N12709 | data_masked[2148];
  assign N12709 = N12708 | data_masked[2276];
  assign N12708 = N12707 | data_masked[2404];
  assign N12707 = N12706 | data_masked[2532];
  assign N12706 = N12705 | data_masked[2660];
  assign N12705 = N12704 | data_masked[2788];
  assign N12704 = N12703 | data_masked[2916];
  assign N12703 = N12702 | data_masked[3044];
  assign N12702 = N12701 | data_masked[3172];
  assign N12701 = N12700 | data_masked[3300];
  assign N12700 = N12699 | data_masked[3428];
  assign N12699 = N12698 | data_masked[3556];
  assign N12698 = N12697 | data_masked[3684];
  assign N12697 = N12696 | data_masked[3812];
  assign N12696 = N12695 | data_masked[3940];
  assign N12695 = N12694 | data_masked[4068];
  assign N12694 = N12693 | data_masked[4196];
  assign N12693 = N12692 | data_masked[4324];
  assign N12692 = N12691 | data_masked[4452];
  assign N12691 = N12690 | data_masked[4580];
  assign N12690 = N12689 | data_masked[4708];
  assign N12689 = N12688 | data_masked[4836];
  assign N12688 = N12687 | data_masked[4964];
  assign N12687 = N12686 | data_masked[5092];
  assign N12686 = N12685 | data_masked[5220];
  assign N12685 = N12684 | data_masked[5348];
  assign N12684 = N12683 | data_masked[5476];
  assign N12683 = N12682 | data_masked[5604];
  assign N12682 = N12681 | data_masked[5732];
  assign N12681 = N12680 | data_masked[5860];
  assign N12680 = N12679 | data_masked[5988];
  assign N12679 = N12678 | data_masked[6116];
  assign N12678 = N12677 | data_masked[6244];
  assign N12677 = N12676 | data_masked[6372];
  assign N12676 = N12675 | data_masked[6500];
  assign N12675 = N12674 | data_masked[6628];
  assign N12674 = N12673 | data_masked[6756];
  assign N12673 = N12672 | data_masked[6884];
  assign N12672 = N12671 | data_masked[7012];
  assign N12671 = N12670 | data_masked[7140];
  assign N12670 = N12669 | data_masked[7268];
  assign N12669 = N12668 | data_masked[7396];
  assign N12668 = N12667 | data_masked[7524];
  assign N12667 = N12666 | data_masked[7652];
  assign N12666 = N12665 | data_masked[7780];
  assign N12665 = N12664 | data_masked[7908];
  assign N12664 = N12663 | data_masked[8036];
  assign N12663 = N12662 | data_masked[8164];
  assign N12662 = N12661 | data_masked[8292];
  assign N12661 = N12660 | data_masked[8420];
  assign N12660 = N12659 | data_masked[8548];
  assign N12659 = N12658 | data_masked[8676];
  assign N12658 = N12657 | data_masked[8804];
  assign N12657 = N12656 | data_masked[8932];
  assign N12656 = N12655 | data_masked[9060];
  assign N12655 = N12654 | data_masked[9188];
  assign N12654 = N12653 | data_masked[9316];
  assign N12653 = N12652 | data_masked[9444];
  assign N12652 = N12651 | data_masked[9572];
  assign N12651 = N12650 | data_masked[9700];
  assign N12650 = N12649 | data_masked[9828];
  assign N12649 = N12648 | data_masked[9956];
  assign N12648 = N12647 | data_masked[10084];
  assign N12647 = N12646 | data_masked[10212];
  assign N12646 = N12645 | data_masked[10340];
  assign N12645 = N12644 | data_masked[10468];
  assign N12644 = N12643 | data_masked[10596];
  assign N12643 = N12642 | data_masked[10724];
  assign N12642 = N12641 | data_masked[10852];
  assign N12641 = N12640 | data_masked[10980];
  assign N12640 = N12639 | data_masked[11108];
  assign N12639 = N12638 | data_masked[11236];
  assign N12638 = N12637 | data_masked[11364];
  assign N12637 = N12636 | data_masked[11492];
  assign N12636 = N12635 | data_masked[11620];
  assign N12635 = N12634 | data_masked[11748];
  assign N12634 = N12633 | data_masked[11876];
  assign N12633 = N12632 | data_masked[12004];
  assign N12632 = N12631 | data_masked[12132];
  assign N12631 = N12630 | data_masked[12260];
  assign N12630 = N12629 | data_masked[12388];
  assign N12629 = N12628 | data_masked[12516];
  assign N12628 = N12627 | data_masked[12644];
  assign N12627 = N12626 | data_masked[12772];
  assign N12626 = N12625 | data_masked[12900];
  assign N12625 = N12624 | data_masked[13028];
  assign N12624 = N12623 | data_masked[13156];
  assign N12623 = N12622 | data_masked[13284];
  assign N12622 = N12621 | data_masked[13412];
  assign N12621 = N12620 | data_masked[13540];
  assign N12620 = N12619 | data_masked[13668];
  assign N12619 = N12618 | data_masked[13796];
  assign N12618 = N12617 | data_masked[13924];
  assign N12617 = N12616 | data_masked[14052];
  assign N12616 = N12615 | data_masked[14180];
  assign N12615 = N12614 | data_masked[14308];
  assign N12614 = N12613 | data_masked[14436];
  assign N12613 = N12612 | data_masked[14564];
  assign N12612 = N12611 | data_masked[14692];
  assign N12611 = N12610 | data_masked[14820];
  assign N12610 = N12609 | data_masked[14948];
  assign N12609 = N12608 | data_masked[15076];
  assign N12608 = N12607 | data_masked[15204];
  assign N12607 = N12606 | data_masked[15332];
  assign N12606 = N12605 | data_masked[15460];
  assign N12605 = N12604 | data_masked[15588];
  assign N12604 = N12603 | data_masked[15716];
  assign N12603 = N12602 | data_masked[15844];
  assign N12602 = N12601 | data_masked[15972];
  assign N12601 = N12600 | data_masked[16100];
  assign N12600 = data_masked[16356] | data_masked[16228];
  assign data_o[101] = N12851 | data_masked[101];
  assign N12851 = N12850 | data_masked[229];
  assign N12850 = N12849 | data_masked[357];
  assign N12849 = N12848 | data_masked[485];
  assign N12848 = N12847 | data_masked[613];
  assign N12847 = N12846 | data_masked[741];
  assign N12846 = N12845 | data_masked[869];
  assign N12845 = N12844 | data_masked[997];
  assign N12844 = N12843 | data_masked[1125];
  assign N12843 = N12842 | data_masked[1253];
  assign N12842 = N12841 | data_masked[1381];
  assign N12841 = N12840 | data_masked[1509];
  assign N12840 = N12839 | data_masked[1637];
  assign N12839 = N12838 | data_masked[1765];
  assign N12838 = N12837 | data_masked[1893];
  assign N12837 = N12836 | data_masked[2021];
  assign N12836 = N12835 | data_masked[2149];
  assign N12835 = N12834 | data_masked[2277];
  assign N12834 = N12833 | data_masked[2405];
  assign N12833 = N12832 | data_masked[2533];
  assign N12832 = N12831 | data_masked[2661];
  assign N12831 = N12830 | data_masked[2789];
  assign N12830 = N12829 | data_masked[2917];
  assign N12829 = N12828 | data_masked[3045];
  assign N12828 = N12827 | data_masked[3173];
  assign N12827 = N12826 | data_masked[3301];
  assign N12826 = N12825 | data_masked[3429];
  assign N12825 = N12824 | data_masked[3557];
  assign N12824 = N12823 | data_masked[3685];
  assign N12823 = N12822 | data_masked[3813];
  assign N12822 = N12821 | data_masked[3941];
  assign N12821 = N12820 | data_masked[4069];
  assign N12820 = N12819 | data_masked[4197];
  assign N12819 = N12818 | data_masked[4325];
  assign N12818 = N12817 | data_masked[4453];
  assign N12817 = N12816 | data_masked[4581];
  assign N12816 = N12815 | data_masked[4709];
  assign N12815 = N12814 | data_masked[4837];
  assign N12814 = N12813 | data_masked[4965];
  assign N12813 = N12812 | data_masked[5093];
  assign N12812 = N12811 | data_masked[5221];
  assign N12811 = N12810 | data_masked[5349];
  assign N12810 = N12809 | data_masked[5477];
  assign N12809 = N12808 | data_masked[5605];
  assign N12808 = N12807 | data_masked[5733];
  assign N12807 = N12806 | data_masked[5861];
  assign N12806 = N12805 | data_masked[5989];
  assign N12805 = N12804 | data_masked[6117];
  assign N12804 = N12803 | data_masked[6245];
  assign N12803 = N12802 | data_masked[6373];
  assign N12802 = N12801 | data_masked[6501];
  assign N12801 = N12800 | data_masked[6629];
  assign N12800 = N12799 | data_masked[6757];
  assign N12799 = N12798 | data_masked[6885];
  assign N12798 = N12797 | data_masked[7013];
  assign N12797 = N12796 | data_masked[7141];
  assign N12796 = N12795 | data_masked[7269];
  assign N12795 = N12794 | data_masked[7397];
  assign N12794 = N12793 | data_masked[7525];
  assign N12793 = N12792 | data_masked[7653];
  assign N12792 = N12791 | data_masked[7781];
  assign N12791 = N12790 | data_masked[7909];
  assign N12790 = N12789 | data_masked[8037];
  assign N12789 = N12788 | data_masked[8165];
  assign N12788 = N12787 | data_masked[8293];
  assign N12787 = N12786 | data_masked[8421];
  assign N12786 = N12785 | data_masked[8549];
  assign N12785 = N12784 | data_masked[8677];
  assign N12784 = N12783 | data_masked[8805];
  assign N12783 = N12782 | data_masked[8933];
  assign N12782 = N12781 | data_masked[9061];
  assign N12781 = N12780 | data_masked[9189];
  assign N12780 = N12779 | data_masked[9317];
  assign N12779 = N12778 | data_masked[9445];
  assign N12778 = N12777 | data_masked[9573];
  assign N12777 = N12776 | data_masked[9701];
  assign N12776 = N12775 | data_masked[9829];
  assign N12775 = N12774 | data_masked[9957];
  assign N12774 = N12773 | data_masked[10085];
  assign N12773 = N12772 | data_masked[10213];
  assign N12772 = N12771 | data_masked[10341];
  assign N12771 = N12770 | data_masked[10469];
  assign N12770 = N12769 | data_masked[10597];
  assign N12769 = N12768 | data_masked[10725];
  assign N12768 = N12767 | data_masked[10853];
  assign N12767 = N12766 | data_masked[10981];
  assign N12766 = N12765 | data_masked[11109];
  assign N12765 = N12764 | data_masked[11237];
  assign N12764 = N12763 | data_masked[11365];
  assign N12763 = N12762 | data_masked[11493];
  assign N12762 = N12761 | data_masked[11621];
  assign N12761 = N12760 | data_masked[11749];
  assign N12760 = N12759 | data_masked[11877];
  assign N12759 = N12758 | data_masked[12005];
  assign N12758 = N12757 | data_masked[12133];
  assign N12757 = N12756 | data_masked[12261];
  assign N12756 = N12755 | data_masked[12389];
  assign N12755 = N12754 | data_masked[12517];
  assign N12754 = N12753 | data_masked[12645];
  assign N12753 = N12752 | data_masked[12773];
  assign N12752 = N12751 | data_masked[12901];
  assign N12751 = N12750 | data_masked[13029];
  assign N12750 = N12749 | data_masked[13157];
  assign N12749 = N12748 | data_masked[13285];
  assign N12748 = N12747 | data_masked[13413];
  assign N12747 = N12746 | data_masked[13541];
  assign N12746 = N12745 | data_masked[13669];
  assign N12745 = N12744 | data_masked[13797];
  assign N12744 = N12743 | data_masked[13925];
  assign N12743 = N12742 | data_masked[14053];
  assign N12742 = N12741 | data_masked[14181];
  assign N12741 = N12740 | data_masked[14309];
  assign N12740 = N12739 | data_masked[14437];
  assign N12739 = N12738 | data_masked[14565];
  assign N12738 = N12737 | data_masked[14693];
  assign N12737 = N12736 | data_masked[14821];
  assign N12736 = N12735 | data_masked[14949];
  assign N12735 = N12734 | data_masked[15077];
  assign N12734 = N12733 | data_masked[15205];
  assign N12733 = N12732 | data_masked[15333];
  assign N12732 = N12731 | data_masked[15461];
  assign N12731 = N12730 | data_masked[15589];
  assign N12730 = N12729 | data_masked[15717];
  assign N12729 = N12728 | data_masked[15845];
  assign N12728 = N12727 | data_masked[15973];
  assign N12727 = N12726 | data_masked[16101];
  assign N12726 = data_masked[16357] | data_masked[16229];
  assign data_o[102] = N12977 | data_masked[102];
  assign N12977 = N12976 | data_masked[230];
  assign N12976 = N12975 | data_masked[358];
  assign N12975 = N12974 | data_masked[486];
  assign N12974 = N12973 | data_masked[614];
  assign N12973 = N12972 | data_masked[742];
  assign N12972 = N12971 | data_masked[870];
  assign N12971 = N12970 | data_masked[998];
  assign N12970 = N12969 | data_masked[1126];
  assign N12969 = N12968 | data_masked[1254];
  assign N12968 = N12967 | data_masked[1382];
  assign N12967 = N12966 | data_masked[1510];
  assign N12966 = N12965 | data_masked[1638];
  assign N12965 = N12964 | data_masked[1766];
  assign N12964 = N12963 | data_masked[1894];
  assign N12963 = N12962 | data_masked[2022];
  assign N12962 = N12961 | data_masked[2150];
  assign N12961 = N12960 | data_masked[2278];
  assign N12960 = N12959 | data_masked[2406];
  assign N12959 = N12958 | data_masked[2534];
  assign N12958 = N12957 | data_masked[2662];
  assign N12957 = N12956 | data_masked[2790];
  assign N12956 = N12955 | data_masked[2918];
  assign N12955 = N12954 | data_masked[3046];
  assign N12954 = N12953 | data_masked[3174];
  assign N12953 = N12952 | data_masked[3302];
  assign N12952 = N12951 | data_masked[3430];
  assign N12951 = N12950 | data_masked[3558];
  assign N12950 = N12949 | data_masked[3686];
  assign N12949 = N12948 | data_masked[3814];
  assign N12948 = N12947 | data_masked[3942];
  assign N12947 = N12946 | data_masked[4070];
  assign N12946 = N12945 | data_masked[4198];
  assign N12945 = N12944 | data_masked[4326];
  assign N12944 = N12943 | data_masked[4454];
  assign N12943 = N12942 | data_masked[4582];
  assign N12942 = N12941 | data_masked[4710];
  assign N12941 = N12940 | data_masked[4838];
  assign N12940 = N12939 | data_masked[4966];
  assign N12939 = N12938 | data_masked[5094];
  assign N12938 = N12937 | data_masked[5222];
  assign N12937 = N12936 | data_masked[5350];
  assign N12936 = N12935 | data_masked[5478];
  assign N12935 = N12934 | data_masked[5606];
  assign N12934 = N12933 | data_masked[5734];
  assign N12933 = N12932 | data_masked[5862];
  assign N12932 = N12931 | data_masked[5990];
  assign N12931 = N12930 | data_masked[6118];
  assign N12930 = N12929 | data_masked[6246];
  assign N12929 = N12928 | data_masked[6374];
  assign N12928 = N12927 | data_masked[6502];
  assign N12927 = N12926 | data_masked[6630];
  assign N12926 = N12925 | data_masked[6758];
  assign N12925 = N12924 | data_masked[6886];
  assign N12924 = N12923 | data_masked[7014];
  assign N12923 = N12922 | data_masked[7142];
  assign N12922 = N12921 | data_masked[7270];
  assign N12921 = N12920 | data_masked[7398];
  assign N12920 = N12919 | data_masked[7526];
  assign N12919 = N12918 | data_masked[7654];
  assign N12918 = N12917 | data_masked[7782];
  assign N12917 = N12916 | data_masked[7910];
  assign N12916 = N12915 | data_masked[8038];
  assign N12915 = N12914 | data_masked[8166];
  assign N12914 = N12913 | data_masked[8294];
  assign N12913 = N12912 | data_masked[8422];
  assign N12912 = N12911 | data_masked[8550];
  assign N12911 = N12910 | data_masked[8678];
  assign N12910 = N12909 | data_masked[8806];
  assign N12909 = N12908 | data_masked[8934];
  assign N12908 = N12907 | data_masked[9062];
  assign N12907 = N12906 | data_masked[9190];
  assign N12906 = N12905 | data_masked[9318];
  assign N12905 = N12904 | data_masked[9446];
  assign N12904 = N12903 | data_masked[9574];
  assign N12903 = N12902 | data_masked[9702];
  assign N12902 = N12901 | data_masked[9830];
  assign N12901 = N12900 | data_masked[9958];
  assign N12900 = N12899 | data_masked[10086];
  assign N12899 = N12898 | data_masked[10214];
  assign N12898 = N12897 | data_masked[10342];
  assign N12897 = N12896 | data_masked[10470];
  assign N12896 = N12895 | data_masked[10598];
  assign N12895 = N12894 | data_masked[10726];
  assign N12894 = N12893 | data_masked[10854];
  assign N12893 = N12892 | data_masked[10982];
  assign N12892 = N12891 | data_masked[11110];
  assign N12891 = N12890 | data_masked[11238];
  assign N12890 = N12889 | data_masked[11366];
  assign N12889 = N12888 | data_masked[11494];
  assign N12888 = N12887 | data_masked[11622];
  assign N12887 = N12886 | data_masked[11750];
  assign N12886 = N12885 | data_masked[11878];
  assign N12885 = N12884 | data_masked[12006];
  assign N12884 = N12883 | data_masked[12134];
  assign N12883 = N12882 | data_masked[12262];
  assign N12882 = N12881 | data_masked[12390];
  assign N12881 = N12880 | data_masked[12518];
  assign N12880 = N12879 | data_masked[12646];
  assign N12879 = N12878 | data_masked[12774];
  assign N12878 = N12877 | data_masked[12902];
  assign N12877 = N12876 | data_masked[13030];
  assign N12876 = N12875 | data_masked[13158];
  assign N12875 = N12874 | data_masked[13286];
  assign N12874 = N12873 | data_masked[13414];
  assign N12873 = N12872 | data_masked[13542];
  assign N12872 = N12871 | data_masked[13670];
  assign N12871 = N12870 | data_masked[13798];
  assign N12870 = N12869 | data_masked[13926];
  assign N12869 = N12868 | data_masked[14054];
  assign N12868 = N12867 | data_masked[14182];
  assign N12867 = N12866 | data_masked[14310];
  assign N12866 = N12865 | data_masked[14438];
  assign N12865 = N12864 | data_masked[14566];
  assign N12864 = N12863 | data_masked[14694];
  assign N12863 = N12862 | data_masked[14822];
  assign N12862 = N12861 | data_masked[14950];
  assign N12861 = N12860 | data_masked[15078];
  assign N12860 = N12859 | data_masked[15206];
  assign N12859 = N12858 | data_masked[15334];
  assign N12858 = N12857 | data_masked[15462];
  assign N12857 = N12856 | data_masked[15590];
  assign N12856 = N12855 | data_masked[15718];
  assign N12855 = N12854 | data_masked[15846];
  assign N12854 = N12853 | data_masked[15974];
  assign N12853 = N12852 | data_masked[16102];
  assign N12852 = data_masked[16358] | data_masked[16230];
  assign data_o[103] = N13103 | data_masked[103];
  assign N13103 = N13102 | data_masked[231];
  assign N13102 = N13101 | data_masked[359];
  assign N13101 = N13100 | data_masked[487];
  assign N13100 = N13099 | data_masked[615];
  assign N13099 = N13098 | data_masked[743];
  assign N13098 = N13097 | data_masked[871];
  assign N13097 = N13096 | data_masked[999];
  assign N13096 = N13095 | data_masked[1127];
  assign N13095 = N13094 | data_masked[1255];
  assign N13094 = N13093 | data_masked[1383];
  assign N13093 = N13092 | data_masked[1511];
  assign N13092 = N13091 | data_masked[1639];
  assign N13091 = N13090 | data_masked[1767];
  assign N13090 = N13089 | data_masked[1895];
  assign N13089 = N13088 | data_masked[2023];
  assign N13088 = N13087 | data_masked[2151];
  assign N13087 = N13086 | data_masked[2279];
  assign N13086 = N13085 | data_masked[2407];
  assign N13085 = N13084 | data_masked[2535];
  assign N13084 = N13083 | data_masked[2663];
  assign N13083 = N13082 | data_masked[2791];
  assign N13082 = N13081 | data_masked[2919];
  assign N13081 = N13080 | data_masked[3047];
  assign N13080 = N13079 | data_masked[3175];
  assign N13079 = N13078 | data_masked[3303];
  assign N13078 = N13077 | data_masked[3431];
  assign N13077 = N13076 | data_masked[3559];
  assign N13076 = N13075 | data_masked[3687];
  assign N13075 = N13074 | data_masked[3815];
  assign N13074 = N13073 | data_masked[3943];
  assign N13073 = N13072 | data_masked[4071];
  assign N13072 = N13071 | data_masked[4199];
  assign N13071 = N13070 | data_masked[4327];
  assign N13070 = N13069 | data_masked[4455];
  assign N13069 = N13068 | data_masked[4583];
  assign N13068 = N13067 | data_masked[4711];
  assign N13067 = N13066 | data_masked[4839];
  assign N13066 = N13065 | data_masked[4967];
  assign N13065 = N13064 | data_masked[5095];
  assign N13064 = N13063 | data_masked[5223];
  assign N13063 = N13062 | data_masked[5351];
  assign N13062 = N13061 | data_masked[5479];
  assign N13061 = N13060 | data_masked[5607];
  assign N13060 = N13059 | data_masked[5735];
  assign N13059 = N13058 | data_masked[5863];
  assign N13058 = N13057 | data_masked[5991];
  assign N13057 = N13056 | data_masked[6119];
  assign N13056 = N13055 | data_masked[6247];
  assign N13055 = N13054 | data_masked[6375];
  assign N13054 = N13053 | data_masked[6503];
  assign N13053 = N13052 | data_masked[6631];
  assign N13052 = N13051 | data_masked[6759];
  assign N13051 = N13050 | data_masked[6887];
  assign N13050 = N13049 | data_masked[7015];
  assign N13049 = N13048 | data_masked[7143];
  assign N13048 = N13047 | data_masked[7271];
  assign N13047 = N13046 | data_masked[7399];
  assign N13046 = N13045 | data_masked[7527];
  assign N13045 = N13044 | data_masked[7655];
  assign N13044 = N13043 | data_masked[7783];
  assign N13043 = N13042 | data_masked[7911];
  assign N13042 = N13041 | data_masked[8039];
  assign N13041 = N13040 | data_masked[8167];
  assign N13040 = N13039 | data_masked[8295];
  assign N13039 = N13038 | data_masked[8423];
  assign N13038 = N13037 | data_masked[8551];
  assign N13037 = N13036 | data_masked[8679];
  assign N13036 = N13035 | data_masked[8807];
  assign N13035 = N13034 | data_masked[8935];
  assign N13034 = N13033 | data_masked[9063];
  assign N13033 = N13032 | data_masked[9191];
  assign N13032 = N13031 | data_masked[9319];
  assign N13031 = N13030 | data_masked[9447];
  assign N13030 = N13029 | data_masked[9575];
  assign N13029 = N13028 | data_masked[9703];
  assign N13028 = N13027 | data_masked[9831];
  assign N13027 = N13026 | data_masked[9959];
  assign N13026 = N13025 | data_masked[10087];
  assign N13025 = N13024 | data_masked[10215];
  assign N13024 = N13023 | data_masked[10343];
  assign N13023 = N13022 | data_masked[10471];
  assign N13022 = N13021 | data_masked[10599];
  assign N13021 = N13020 | data_masked[10727];
  assign N13020 = N13019 | data_masked[10855];
  assign N13019 = N13018 | data_masked[10983];
  assign N13018 = N13017 | data_masked[11111];
  assign N13017 = N13016 | data_masked[11239];
  assign N13016 = N13015 | data_masked[11367];
  assign N13015 = N13014 | data_masked[11495];
  assign N13014 = N13013 | data_masked[11623];
  assign N13013 = N13012 | data_masked[11751];
  assign N13012 = N13011 | data_masked[11879];
  assign N13011 = N13010 | data_masked[12007];
  assign N13010 = N13009 | data_masked[12135];
  assign N13009 = N13008 | data_masked[12263];
  assign N13008 = N13007 | data_masked[12391];
  assign N13007 = N13006 | data_masked[12519];
  assign N13006 = N13005 | data_masked[12647];
  assign N13005 = N13004 | data_masked[12775];
  assign N13004 = N13003 | data_masked[12903];
  assign N13003 = N13002 | data_masked[13031];
  assign N13002 = N13001 | data_masked[13159];
  assign N13001 = N13000 | data_masked[13287];
  assign N13000 = N12999 | data_masked[13415];
  assign N12999 = N12998 | data_masked[13543];
  assign N12998 = N12997 | data_masked[13671];
  assign N12997 = N12996 | data_masked[13799];
  assign N12996 = N12995 | data_masked[13927];
  assign N12995 = N12994 | data_masked[14055];
  assign N12994 = N12993 | data_masked[14183];
  assign N12993 = N12992 | data_masked[14311];
  assign N12992 = N12991 | data_masked[14439];
  assign N12991 = N12990 | data_masked[14567];
  assign N12990 = N12989 | data_masked[14695];
  assign N12989 = N12988 | data_masked[14823];
  assign N12988 = N12987 | data_masked[14951];
  assign N12987 = N12986 | data_masked[15079];
  assign N12986 = N12985 | data_masked[15207];
  assign N12985 = N12984 | data_masked[15335];
  assign N12984 = N12983 | data_masked[15463];
  assign N12983 = N12982 | data_masked[15591];
  assign N12982 = N12981 | data_masked[15719];
  assign N12981 = N12980 | data_masked[15847];
  assign N12980 = N12979 | data_masked[15975];
  assign N12979 = N12978 | data_masked[16103];
  assign N12978 = data_masked[16359] | data_masked[16231];
  assign data_o[104] = N13229 | data_masked[104];
  assign N13229 = N13228 | data_masked[232];
  assign N13228 = N13227 | data_masked[360];
  assign N13227 = N13226 | data_masked[488];
  assign N13226 = N13225 | data_masked[616];
  assign N13225 = N13224 | data_masked[744];
  assign N13224 = N13223 | data_masked[872];
  assign N13223 = N13222 | data_masked[1000];
  assign N13222 = N13221 | data_masked[1128];
  assign N13221 = N13220 | data_masked[1256];
  assign N13220 = N13219 | data_masked[1384];
  assign N13219 = N13218 | data_masked[1512];
  assign N13218 = N13217 | data_masked[1640];
  assign N13217 = N13216 | data_masked[1768];
  assign N13216 = N13215 | data_masked[1896];
  assign N13215 = N13214 | data_masked[2024];
  assign N13214 = N13213 | data_masked[2152];
  assign N13213 = N13212 | data_masked[2280];
  assign N13212 = N13211 | data_masked[2408];
  assign N13211 = N13210 | data_masked[2536];
  assign N13210 = N13209 | data_masked[2664];
  assign N13209 = N13208 | data_masked[2792];
  assign N13208 = N13207 | data_masked[2920];
  assign N13207 = N13206 | data_masked[3048];
  assign N13206 = N13205 | data_masked[3176];
  assign N13205 = N13204 | data_masked[3304];
  assign N13204 = N13203 | data_masked[3432];
  assign N13203 = N13202 | data_masked[3560];
  assign N13202 = N13201 | data_masked[3688];
  assign N13201 = N13200 | data_masked[3816];
  assign N13200 = N13199 | data_masked[3944];
  assign N13199 = N13198 | data_masked[4072];
  assign N13198 = N13197 | data_masked[4200];
  assign N13197 = N13196 | data_masked[4328];
  assign N13196 = N13195 | data_masked[4456];
  assign N13195 = N13194 | data_masked[4584];
  assign N13194 = N13193 | data_masked[4712];
  assign N13193 = N13192 | data_masked[4840];
  assign N13192 = N13191 | data_masked[4968];
  assign N13191 = N13190 | data_masked[5096];
  assign N13190 = N13189 | data_masked[5224];
  assign N13189 = N13188 | data_masked[5352];
  assign N13188 = N13187 | data_masked[5480];
  assign N13187 = N13186 | data_masked[5608];
  assign N13186 = N13185 | data_masked[5736];
  assign N13185 = N13184 | data_masked[5864];
  assign N13184 = N13183 | data_masked[5992];
  assign N13183 = N13182 | data_masked[6120];
  assign N13182 = N13181 | data_masked[6248];
  assign N13181 = N13180 | data_masked[6376];
  assign N13180 = N13179 | data_masked[6504];
  assign N13179 = N13178 | data_masked[6632];
  assign N13178 = N13177 | data_masked[6760];
  assign N13177 = N13176 | data_masked[6888];
  assign N13176 = N13175 | data_masked[7016];
  assign N13175 = N13174 | data_masked[7144];
  assign N13174 = N13173 | data_masked[7272];
  assign N13173 = N13172 | data_masked[7400];
  assign N13172 = N13171 | data_masked[7528];
  assign N13171 = N13170 | data_masked[7656];
  assign N13170 = N13169 | data_masked[7784];
  assign N13169 = N13168 | data_masked[7912];
  assign N13168 = N13167 | data_masked[8040];
  assign N13167 = N13166 | data_masked[8168];
  assign N13166 = N13165 | data_masked[8296];
  assign N13165 = N13164 | data_masked[8424];
  assign N13164 = N13163 | data_masked[8552];
  assign N13163 = N13162 | data_masked[8680];
  assign N13162 = N13161 | data_masked[8808];
  assign N13161 = N13160 | data_masked[8936];
  assign N13160 = N13159 | data_masked[9064];
  assign N13159 = N13158 | data_masked[9192];
  assign N13158 = N13157 | data_masked[9320];
  assign N13157 = N13156 | data_masked[9448];
  assign N13156 = N13155 | data_masked[9576];
  assign N13155 = N13154 | data_masked[9704];
  assign N13154 = N13153 | data_masked[9832];
  assign N13153 = N13152 | data_masked[9960];
  assign N13152 = N13151 | data_masked[10088];
  assign N13151 = N13150 | data_masked[10216];
  assign N13150 = N13149 | data_masked[10344];
  assign N13149 = N13148 | data_masked[10472];
  assign N13148 = N13147 | data_masked[10600];
  assign N13147 = N13146 | data_masked[10728];
  assign N13146 = N13145 | data_masked[10856];
  assign N13145 = N13144 | data_masked[10984];
  assign N13144 = N13143 | data_masked[11112];
  assign N13143 = N13142 | data_masked[11240];
  assign N13142 = N13141 | data_masked[11368];
  assign N13141 = N13140 | data_masked[11496];
  assign N13140 = N13139 | data_masked[11624];
  assign N13139 = N13138 | data_masked[11752];
  assign N13138 = N13137 | data_masked[11880];
  assign N13137 = N13136 | data_masked[12008];
  assign N13136 = N13135 | data_masked[12136];
  assign N13135 = N13134 | data_masked[12264];
  assign N13134 = N13133 | data_masked[12392];
  assign N13133 = N13132 | data_masked[12520];
  assign N13132 = N13131 | data_masked[12648];
  assign N13131 = N13130 | data_masked[12776];
  assign N13130 = N13129 | data_masked[12904];
  assign N13129 = N13128 | data_masked[13032];
  assign N13128 = N13127 | data_masked[13160];
  assign N13127 = N13126 | data_masked[13288];
  assign N13126 = N13125 | data_masked[13416];
  assign N13125 = N13124 | data_masked[13544];
  assign N13124 = N13123 | data_masked[13672];
  assign N13123 = N13122 | data_masked[13800];
  assign N13122 = N13121 | data_masked[13928];
  assign N13121 = N13120 | data_masked[14056];
  assign N13120 = N13119 | data_masked[14184];
  assign N13119 = N13118 | data_masked[14312];
  assign N13118 = N13117 | data_masked[14440];
  assign N13117 = N13116 | data_masked[14568];
  assign N13116 = N13115 | data_masked[14696];
  assign N13115 = N13114 | data_masked[14824];
  assign N13114 = N13113 | data_masked[14952];
  assign N13113 = N13112 | data_masked[15080];
  assign N13112 = N13111 | data_masked[15208];
  assign N13111 = N13110 | data_masked[15336];
  assign N13110 = N13109 | data_masked[15464];
  assign N13109 = N13108 | data_masked[15592];
  assign N13108 = N13107 | data_masked[15720];
  assign N13107 = N13106 | data_masked[15848];
  assign N13106 = N13105 | data_masked[15976];
  assign N13105 = N13104 | data_masked[16104];
  assign N13104 = data_masked[16360] | data_masked[16232];
  assign data_o[105] = N13355 | data_masked[105];
  assign N13355 = N13354 | data_masked[233];
  assign N13354 = N13353 | data_masked[361];
  assign N13353 = N13352 | data_masked[489];
  assign N13352 = N13351 | data_masked[617];
  assign N13351 = N13350 | data_masked[745];
  assign N13350 = N13349 | data_masked[873];
  assign N13349 = N13348 | data_masked[1001];
  assign N13348 = N13347 | data_masked[1129];
  assign N13347 = N13346 | data_masked[1257];
  assign N13346 = N13345 | data_masked[1385];
  assign N13345 = N13344 | data_masked[1513];
  assign N13344 = N13343 | data_masked[1641];
  assign N13343 = N13342 | data_masked[1769];
  assign N13342 = N13341 | data_masked[1897];
  assign N13341 = N13340 | data_masked[2025];
  assign N13340 = N13339 | data_masked[2153];
  assign N13339 = N13338 | data_masked[2281];
  assign N13338 = N13337 | data_masked[2409];
  assign N13337 = N13336 | data_masked[2537];
  assign N13336 = N13335 | data_masked[2665];
  assign N13335 = N13334 | data_masked[2793];
  assign N13334 = N13333 | data_masked[2921];
  assign N13333 = N13332 | data_masked[3049];
  assign N13332 = N13331 | data_masked[3177];
  assign N13331 = N13330 | data_masked[3305];
  assign N13330 = N13329 | data_masked[3433];
  assign N13329 = N13328 | data_masked[3561];
  assign N13328 = N13327 | data_masked[3689];
  assign N13327 = N13326 | data_masked[3817];
  assign N13326 = N13325 | data_masked[3945];
  assign N13325 = N13324 | data_masked[4073];
  assign N13324 = N13323 | data_masked[4201];
  assign N13323 = N13322 | data_masked[4329];
  assign N13322 = N13321 | data_masked[4457];
  assign N13321 = N13320 | data_masked[4585];
  assign N13320 = N13319 | data_masked[4713];
  assign N13319 = N13318 | data_masked[4841];
  assign N13318 = N13317 | data_masked[4969];
  assign N13317 = N13316 | data_masked[5097];
  assign N13316 = N13315 | data_masked[5225];
  assign N13315 = N13314 | data_masked[5353];
  assign N13314 = N13313 | data_masked[5481];
  assign N13313 = N13312 | data_masked[5609];
  assign N13312 = N13311 | data_masked[5737];
  assign N13311 = N13310 | data_masked[5865];
  assign N13310 = N13309 | data_masked[5993];
  assign N13309 = N13308 | data_masked[6121];
  assign N13308 = N13307 | data_masked[6249];
  assign N13307 = N13306 | data_masked[6377];
  assign N13306 = N13305 | data_masked[6505];
  assign N13305 = N13304 | data_masked[6633];
  assign N13304 = N13303 | data_masked[6761];
  assign N13303 = N13302 | data_masked[6889];
  assign N13302 = N13301 | data_masked[7017];
  assign N13301 = N13300 | data_masked[7145];
  assign N13300 = N13299 | data_masked[7273];
  assign N13299 = N13298 | data_masked[7401];
  assign N13298 = N13297 | data_masked[7529];
  assign N13297 = N13296 | data_masked[7657];
  assign N13296 = N13295 | data_masked[7785];
  assign N13295 = N13294 | data_masked[7913];
  assign N13294 = N13293 | data_masked[8041];
  assign N13293 = N13292 | data_masked[8169];
  assign N13292 = N13291 | data_masked[8297];
  assign N13291 = N13290 | data_masked[8425];
  assign N13290 = N13289 | data_masked[8553];
  assign N13289 = N13288 | data_masked[8681];
  assign N13288 = N13287 | data_masked[8809];
  assign N13287 = N13286 | data_masked[8937];
  assign N13286 = N13285 | data_masked[9065];
  assign N13285 = N13284 | data_masked[9193];
  assign N13284 = N13283 | data_masked[9321];
  assign N13283 = N13282 | data_masked[9449];
  assign N13282 = N13281 | data_masked[9577];
  assign N13281 = N13280 | data_masked[9705];
  assign N13280 = N13279 | data_masked[9833];
  assign N13279 = N13278 | data_masked[9961];
  assign N13278 = N13277 | data_masked[10089];
  assign N13277 = N13276 | data_masked[10217];
  assign N13276 = N13275 | data_masked[10345];
  assign N13275 = N13274 | data_masked[10473];
  assign N13274 = N13273 | data_masked[10601];
  assign N13273 = N13272 | data_masked[10729];
  assign N13272 = N13271 | data_masked[10857];
  assign N13271 = N13270 | data_masked[10985];
  assign N13270 = N13269 | data_masked[11113];
  assign N13269 = N13268 | data_masked[11241];
  assign N13268 = N13267 | data_masked[11369];
  assign N13267 = N13266 | data_masked[11497];
  assign N13266 = N13265 | data_masked[11625];
  assign N13265 = N13264 | data_masked[11753];
  assign N13264 = N13263 | data_masked[11881];
  assign N13263 = N13262 | data_masked[12009];
  assign N13262 = N13261 | data_masked[12137];
  assign N13261 = N13260 | data_masked[12265];
  assign N13260 = N13259 | data_masked[12393];
  assign N13259 = N13258 | data_masked[12521];
  assign N13258 = N13257 | data_masked[12649];
  assign N13257 = N13256 | data_masked[12777];
  assign N13256 = N13255 | data_masked[12905];
  assign N13255 = N13254 | data_masked[13033];
  assign N13254 = N13253 | data_masked[13161];
  assign N13253 = N13252 | data_masked[13289];
  assign N13252 = N13251 | data_masked[13417];
  assign N13251 = N13250 | data_masked[13545];
  assign N13250 = N13249 | data_masked[13673];
  assign N13249 = N13248 | data_masked[13801];
  assign N13248 = N13247 | data_masked[13929];
  assign N13247 = N13246 | data_masked[14057];
  assign N13246 = N13245 | data_masked[14185];
  assign N13245 = N13244 | data_masked[14313];
  assign N13244 = N13243 | data_masked[14441];
  assign N13243 = N13242 | data_masked[14569];
  assign N13242 = N13241 | data_masked[14697];
  assign N13241 = N13240 | data_masked[14825];
  assign N13240 = N13239 | data_masked[14953];
  assign N13239 = N13238 | data_masked[15081];
  assign N13238 = N13237 | data_masked[15209];
  assign N13237 = N13236 | data_masked[15337];
  assign N13236 = N13235 | data_masked[15465];
  assign N13235 = N13234 | data_masked[15593];
  assign N13234 = N13233 | data_masked[15721];
  assign N13233 = N13232 | data_masked[15849];
  assign N13232 = N13231 | data_masked[15977];
  assign N13231 = N13230 | data_masked[16105];
  assign N13230 = data_masked[16361] | data_masked[16233];
  assign data_o[106] = N13481 | data_masked[106];
  assign N13481 = N13480 | data_masked[234];
  assign N13480 = N13479 | data_masked[362];
  assign N13479 = N13478 | data_masked[490];
  assign N13478 = N13477 | data_masked[618];
  assign N13477 = N13476 | data_masked[746];
  assign N13476 = N13475 | data_masked[874];
  assign N13475 = N13474 | data_masked[1002];
  assign N13474 = N13473 | data_masked[1130];
  assign N13473 = N13472 | data_masked[1258];
  assign N13472 = N13471 | data_masked[1386];
  assign N13471 = N13470 | data_masked[1514];
  assign N13470 = N13469 | data_masked[1642];
  assign N13469 = N13468 | data_masked[1770];
  assign N13468 = N13467 | data_masked[1898];
  assign N13467 = N13466 | data_masked[2026];
  assign N13466 = N13465 | data_masked[2154];
  assign N13465 = N13464 | data_masked[2282];
  assign N13464 = N13463 | data_masked[2410];
  assign N13463 = N13462 | data_masked[2538];
  assign N13462 = N13461 | data_masked[2666];
  assign N13461 = N13460 | data_masked[2794];
  assign N13460 = N13459 | data_masked[2922];
  assign N13459 = N13458 | data_masked[3050];
  assign N13458 = N13457 | data_masked[3178];
  assign N13457 = N13456 | data_masked[3306];
  assign N13456 = N13455 | data_masked[3434];
  assign N13455 = N13454 | data_masked[3562];
  assign N13454 = N13453 | data_masked[3690];
  assign N13453 = N13452 | data_masked[3818];
  assign N13452 = N13451 | data_masked[3946];
  assign N13451 = N13450 | data_masked[4074];
  assign N13450 = N13449 | data_masked[4202];
  assign N13449 = N13448 | data_masked[4330];
  assign N13448 = N13447 | data_masked[4458];
  assign N13447 = N13446 | data_masked[4586];
  assign N13446 = N13445 | data_masked[4714];
  assign N13445 = N13444 | data_masked[4842];
  assign N13444 = N13443 | data_masked[4970];
  assign N13443 = N13442 | data_masked[5098];
  assign N13442 = N13441 | data_masked[5226];
  assign N13441 = N13440 | data_masked[5354];
  assign N13440 = N13439 | data_masked[5482];
  assign N13439 = N13438 | data_masked[5610];
  assign N13438 = N13437 | data_masked[5738];
  assign N13437 = N13436 | data_masked[5866];
  assign N13436 = N13435 | data_masked[5994];
  assign N13435 = N13434 | data_masked[6122];
  assign N13434 = N13433 | data_masked[6250];
  assign N13433 = N13432 | data_masked[6378];
  assign N13432 = N13431 | data_masked[6506];
  assign N13431 = N13430 | data_masked[6634];
  assign N13430 = N13429 | data_masked[6762];
  assign N13429 = N13428 | data_masked[6890];
  assign N13428 = N13427 | data_masked[7018];
  assign N13427 = N13426 | data_masked[7146];
  assign N13426 = N13425 | data_masked[7274];
  assign N13425 = N13424 | data_masked[7402];
  assign N13424 = N13423 | data_masked[7530];
  assign N13423 = N13422 | data_masked[7658];
  assign N13422 = N13421 | data_masked[7786];
  assign N13421 = N13420 | data_masked[7914];
  assign N13420 = N13419 | data_masked[8042];
  assign N13419 = N13418 | data_masked[8170];
  assign N13418 = N13417 | data_masked[8298];
  assign N13417 = N13416 | data_masked[8426];
  assign N13416 = N13415 | data_masked[8554];
  assign N13415 = N13414 | data_masked[8682];
  assign N13414 = N13413 | data_masked[8810];
  assign N13413 = N13412 | data_masked[8938];
  assign N13412 = N13411 | data_masked[9066];
  assign N13411 = N13410 | data_masked[9194];
  assign N13410 = N13409 | data_masked[9322];
  assign N13409 = N13408 | data_masked[9450];
  assign N13408 = N13407 | data_masked[9578];
  assign N13407 = N13406 | data_masked[9706];
  assign N13406 = N13405 | data_masked[9834];
  assign N13405 = N13404 | data_masked[9962];
  assign N13404 = N13403 | data_masked[10090];
  assign N13403 = N13402 | data_masked[10218];
  assign N13402 = N13401 | data_masked[10346];
  assign N13401 = N13400 | data_masked[10474];
  assign N13400 = N13399 | data_masked[10602];
  assign N13399 = N13398 | data_masked[10730];
  assign N13398 = N13397 | data_masked[10858];
  assign N13397 = N13396 | data_masked[10986];
  assign N13396 = N13395 | data_masked[11114];
  assign N13395 = N13394 | data_masked[11242];
  assign N13394 = N13393 | data_masked[11370];
  assign N13393 = N13392 | data_masked[11498];
  assign N13392 = N13391 | data_masked[11626];
  assign N13391 = N13390 | data_masked[11754];
  assign N13390 = N13389 | data_masked[11882];
  assign N13389 = N13388 | data_masked[12010];
  assign N13388 = N13387 | data_masked[12138];
  assign N13387 = N13386 | data_masked[12266];
  assign N13386 = N13385 | data_masked[12394];
  assign N13385 = N13384 | data_masked[12522];
  assign N13384 = N13383 | data_masked[12650];
  assign N13383 = N13382 | data_masked[12778];
  assign N13382 = N13381 | data_masked[12906];
  assign N13381 = N13380 | data_masked[13034];
  assign N13380 = N13379 | data_masked[13162];
  assign N13379 = N13378 | data_masked[13290];
  assign N13378 = N13377 | data_masked[13418];
  assign N13377 = N13376 | data_masked[13546];
  assign N13376 = N13375 | data_masked[13674];
  assign N13375 = N13374 | data_masked[13802];
  assign N13374 = N13373 | data_masked[13930];
  assign N13373 = N13372 | data_masked[14058];
  assign N13372 = N13371 | data_masked[14186];
  assign N13371 = N13370 | data_masked[14314];
  assign N13370 = N13369 | data_masked[14442];
  assign N13369 = N13368 | data_masked[14570];
  assign N13368 = N13367 | data_masked[14698];
  assign N13367 = N13366 | data_masked[14826];
  assign N13366 = N13365 | data_masked[14954];
  assign N13365 = N13364 | data_masked[15082];
  assign N13364 = N13363 | data_masked[15210];
  assign N13363 = N13362 | data_masked[15338];
  assign N13362 = N13361 | data_masked[15466];
  assign N13361 = N13360 | data_masked[15594];
  assign N13360 = N13359 | data_masked[15722];
  assign N13359 = N13358 | data_masked[15850];
  assign N13358 = N13357 | data_masked[15978];
  assign N13357 = N13356 | data_masked[16106];
  assign N13356 = data_masked[16362] | data_masked[16234];
  assign data_o[107] = N13607 | data_masked[107];
  assign N13607 = N13606 | data_masked[235];
  assign N13606 = N13605 | data_masked[363];
  assign N13605 = N13604 | data_masked[491];
  assign N13604 = N13603 | data_masked[619];
  assign N13603 = N13602 | data_masked[747];
  assign N13602 = N13601 | data_masked[875];
  assign N13601 = N13600 | data_masked[1003];
  assign N13600 = N13599 | data_masked[1131];
  assign N13599 = N13598 | data_masked[1259];
  assign N13598 = N13597 | data_masked[1387];
  assign N13597 = N13596 | data_masked[1515];
  assign N13596 = N13595 | data_masked[1643];
  assign N13595 = N13594 | data_masked[1771];
  assign N13594 = N13593 | data_masked[1899];
  assign N13593 = N13592 | data_masked[2027];
  assign N13592 = N13591 | data_masked[2155];
  assign N13591 = N13590 | data_masked[2283];
  assign N13590 = N13589 | data_masked[2411];
  assign N13589 = N13588 | data_masked[2539];
  assign N13588 = N13587 | data_masked[2667];
  assign N13587 = N13586 | data_masked[2795];
  assign N13586 = N13585 | data_masked[2923];
  assign N13585 = N13584 | data_masked[3051];
  assign N13584 = N13583 | data_masked[3179];
  assign N13583 = N13582 | data_masked[3307];
  assign N13582 = N13581 | data_masked[3435];
  assign N13581 = N13580 | data_masked[3563];
  assign N13580 = N13579 | data_masked[3691];
  assign N13579 = N13578 | data_masked[3819];
  assign N13578 = N13577 | data_masked[3947];
  assign N13577 = N13576 | data_masked[4075];
  assign N13576 = N13575 | data_masked[4203];
  assign N13575 = N13574 | data_masked[4331];
  assign N13574 = N13573 | data_masked[4459];
  assign N13573 = N13572 | data_masked[4587];
  assign N13572 = N13571 | data_masked[4715];
  assign N13571 = N13570 | data_masked[4843];
  assign N13570 = N13569 | data_masked[4971];
  assign N13569 = N13568 | data_masked[5099];
  assign N13568 = N13567 | data_masked[5227];
  assign N13567 = N13566 | data_masked[5355];
  assign N13566 = N13565 | data_masked[5483];
  assign N13565 = N13564 | data_masked[5611];
  assign N13564 = N13563 | data_masked[5739];
  assign N13563 = N13562 | data_masked[5867];
  assign N13562 = N13561 | data_masked[5995];
  assign N13561 = N13560 | data_masked[6123];
  assign N13560 = N13559 | data_masked[6251];
  assign N13559 = N13558 | data_masked[6379];
  assign N13558 = N13557 | data_masked[6507];
  assign N13557 = N13556 | data_masked[6635];
  assign N13556 = N13555 | data_masked[6763];
  assign N13555 = N13554 | data_masked[6891];
  assign N13554 = N13553 | data_masked[7019];
  assign N13553 = N13552 | data_masked[7147];
  assign N13552 = N13551 | data_masked[7275];
  assign N13551 = N13550 | data_masked[7403];
  assign N13550 = N13549 | data_masked[7531];
  assign N13549 = N13548 | data_masked[7659];
  assign N13548 = N13547 | data_masked[7787];
  assign N13547 = N13546 | data_masked[7915];
  assign N13546 = N13545 | data_masked[8043];
  assign N13545 = N13544 | data_masked[8171];
  assign N13544 = N13543 | data_masked[8299];
  assign N13543 = N13542 | data_masked[8427];
  assign N13542 = N13541 | data_masked[8555];
  assign N13541 = N13540 | data_masked[8683];
  assign N13540 = N13539 | data_masked[8811];
  assign N13539 = N13538 | data_masked[8939];
  assign N13538 = N13537 | data_masked[9067];
  assign N13537 = N13536 | data_masked[9195];
  assign N13536 = N13535 | data_masked[9323];
  assign N13535 = N13534 | data_masked[9451];
  assign N13534 = N13533 | data_masked[9579];
  assign N13533 = N13532 | data_masked[9707];
  assign N13532 = N13531 | data_masked[9835];
  assign N13531 = N13530 | data_masked[9963];
  assign N13530 = N13529 | data_masked[10091];
  assign N13529 = N13528 | data_masked[10219];
  assign N13528 = N13527 | data_masked[10347];
  assign N13527 = N13526 | data_masked[10475];
  assign N13526 = N13525 | data_masked[10603];
  assign N13525 = N13524 | data_masked[10731];
  assign N13524 = N13523 | data_masked[10859];
  assign N13523 = N13522 | data_masked[10987];
  assign N13522 = N13521 | data_masked[11115];
  assign N13521 = N13520 | data_masked[11243];
  assign N13520 = N13519 | data_masked[11371];
  assign N13519 = N13518 | data_masked[11499];
  assign N13518 = N13517 | data_masked[11627];
  assign N13517 = N13516 | data_masked[11755];
  assign N13516 = N13515 | data_masked[11883];
  assign N13515 = N13514 | data_masked[12011];
  assign N13514 = N13513 | data_masked[12139];
  assign N13513 = N13512 | data_masked[12267];
  assign N13512 = N13511 | data_masked[12395];
  assign N13511 = N13510 | data_masked[12523];
  assign N13510 = N13509 | data_masked[12651];
  assign N13509 = N13508 | data_masked[12779];
  assign N13508 = N13507 | data_masked[12907];
  assign N13507 = N13506 | data_masked[13035];
  assign N13506 = N13505 | data_masked[13163];
  assign N13505 = N13504 | data_masked[13291];
  assign N13504 = N13503 | data_masked[13419];
  assign N13503 = N13502 | data_masked[13547];
  assign N13502 = N13501 | data_masked[13675];
  assign N13501 = N13500 | data_masked[13803];
  assign N13500 = N13499 | data_masked[13931];
  assign N13499 = N13498 | data_masked[14059];
  assign N13498 = N13497 | data_masked[14187];
  assign N13497 = N13496 | data_masked[14315];
  assign N13496 = N13495 | data_masked[14443];
  assign N13495 = N13494 | data_masked[14571];
  assign N13494 = N13493 | data_masked[14699];
  assign N13493 = N13492 | data_masked[14827];
  assign N13492 = N13491 | data_masked[14955];
  assign N13491 = N13490 | data_masked[15083];
  assign N13490 = N13489 | data_masked[15211];
  assign N13489 = N13488 | data_masked[15339];
  assign N13488 = N13487 | data_masked[15467];
  assign N13487 = N13486 | data_masked[15595];
  assign N13486 = N13485 | data_masked[15723];
  assign N13485 = N13484 | data_masked[15851];
  assign N13484 = N13483 | data_masked[15979];
  assign N13483 = N13482 | data_masked[16107];
  assign N13482 = data_masked[16363] | data_masked[16235];
  assign data_o[108] = N13733 | data_masked[108];
  assign N13733 = N13732 | data_masked[236];
  assign N13732 = N13731 | data_masked[364];
  assign N13731 = N13730 | data_masked[492];
  assign N13730 = N13729 | data_masked[620];
  assign N13729 = N13728 | data_masked[748];
  assign N13728 = N13727 | data_masked[876];
  assign N13727 = N13726 | data_masked[1004];
  assign N13726 = N13725 | data_masked[1132];
  assign N13725 = N13724 | data_masked[1260];
  assign N13724 = N13723 | data_masked[1388];
  assign N13723 = N13722 | data_masked[1516];
  assign N13722 = N13721 | data_masked[1644];
  assign N13721 = N13720 | data_masked[1772];
  assign N13720 = N13719 | data_masked[1900];
  assign N13719 = N13718 | data_masked[2028];
  assign N13718 = N13717 | data_masked[2156];
  assign N13717 = N13716 | data_masked[2284];
  assign N13716 = N13715 | data_masked[2412];
  assign N13715 = N13714 | data_masked[2540];
  assign N13714 = N13713 | data_masked[2668];
  assign N13713 = N13712 | data_masked[2796];
  assign N13712 = N13711 | data_masked[2924];
  assign N13711 = N13710 | data_masked[3052];
  assign N13710 = N13709 | data_masked[3180];
  assign N13709 = N13708 | data_masked[3308];
  assign N13708 = N13707 | data_masked[3436];
  assign N13707 = N13706 | data_masked[3564];
  assign N13706 = N13705 | data_masked[3692];
  assign N13705 = N13704 | data_masked[3820];
  assign N13704 = N13703 | data_masked[3948];
  assign N13703 = N13702 | data_masked[4076];
  assign N13702 = N13701 | data_masked[4204];
  assign N13701 = N13700 | data_masked[4332];
  assign N13700 = N13699 | data_masked[4460];
  assign N13699 = N13698 | data_masked[4588];
  assign N13698 = N13697 | data_masked[4716];
  assign N13697 = N13696 | data_masked[4844];
  assign N13696 = N13695 | data_masked[4972];
  assign N13695 = N13694 | data_masked[5100];
  assign N13694 = N13693 | data_masked[5228];
  assign N13693 = N13692 | data_masked[5356];
  assign N13692 = N13691 | data_masked[5484];
  assign N13691 = N13690 | data_masked[5612];
  assign N13690 = N13689 | data_masked[5740];
  assign N13689 = N13688 | data_masked[5868];
  assign N13688 = N13687 | data_masked[5996];
  assign N13687 = N13686 | data_masked[6124];
  assign N13686 = N13685 | data_masked[6252];
  assign N13685 = N13684 | data_masked[6380];
  assign N13684 = N13683 | data_masked[6508];
  assign N13683 = N13682 | data_masked[6636];
  assign N13682 = N13681 | data_masked[6764];
  assign N13681 = N13680 | data_masked[6892];
  assign N13680 = N13679 | data_masked[7020];
  assign N13679 = N13678 | data_masked[7148];
  assign N13678 = N13677 | data_masked[7276];
  assign N13677 = N13676 | data_masked[7404];
  assign N13676 = N13675 | data_masked[7532];
  assign N13675 = N13674 | data_masked[7660];
  assign N13674 = N13673 | data_masked[7788];
  assign N13673 = N13672 | data_masked[7916];
  assign N13672 = N13671 | data_masked[8044];
  assign N13671 = N13670 | data_masked[8172];
  assign N13670 = N13669 | data_masked[8300];
  assign N13669 = N13668 | data_masked[8428];
  assign N13668 = N13667 | data_masked[8556];
  assign N13667 = N13666 | data_masked[8684];
  assign N13666 = N13665 | data_masked[8812];
  assign N13665 = N13664 | data_masked[8940];
  assign N13664 = N13663 | data_masked[9068];
  assign N13663 = N13662 | data_masked[9196];
  assign N13662 = N13661 | data_masked[9324];
  assign N13661 = N13660 | data_masked[9452];
  assign N13660 = N13659 | data_masked[9580];
  assign N13659 = N13658 | data_masked[9708];
  assign N13658 = N13657 | data_masked[9836];
  assign N13657 = N13656 | data_masked[9964];
  assign N13656 = N13655 | data_masked[10092];
  assign N13655 = N13654 | data_masked[10220];
  assign N13654 = N13653 | data_masked[10348];
  assign N13653 = N13652 | data_masked[10476];
  assign N13652 = N13651 | data_masked[10604];
  assign N13651 = N13650 | data_masked[10732];
  assign N13650 = N13649 | data_masked[10860];
  assign N13649 = N13648 | data_masked[10988];
  assign N13648 = N13647 | data_masked[11116];
  assign N13647 = N13646 | data_masked[11244];
  assign N13646 = N13645 | data_masked[11372];
  assign N13645 = N13644 | data_masked[11500];
  assign N13644 = N13643 | data_masked[11628];
  assign N13643 = N13642 | data_masked[11756];
  assign N13642 = N13641 | data_masked[11884];
  assign N13641 = N13640 | data_masked[12012];
  assign N13640 = N13639 | data_masked[12140];
  assign N13639 = N13638 | data_masked[12268];
  assign N13638 = N13637 | data_masked[12396];
  assign N13637 = N13636 | data_masked[12524];
  assign N13636 = N13635 | data_masked[12652];
  assign N13635 = N13634 | data_masked[12780];
  assign N13634 = N13633 | data_masked[12908];
  assign N13633 = N13632 | data_masked[13036];
  assign N13632 = N13631 | data_masked[13164];
  assign N13631 = N13630 | data_masked[13292];
  assign N13630 = N13629 | data_masked[13420];
  assign N13629 = N13628 | data_masked[13548];
  assign N13628 = N13627 | data_masked[13676];
  assign N13627 = N13626 | data_masked[13804];
  assign N13626 = N13625 | data_masked[13932];
  assign N13625 = N13624 | data_masked[14060];
  assign N13624 = N13623 | data_masked[14188];
  assign N13623 = N13622 | data_masked[14316];
  assign N13622 = N13621 | data_masked[14444];
  assign N13621 = N13620 | data_masked[14572];
  assign N13620 = N13619 | data_masked[14700];
  assign N13619 = N13618 | data_masked[14828];
  assign N13618 = N13617 | data_masked[14956];
  assign N13617 = N13616 | data_masked[15084];
  assign N13616 = N13615 | data_masked[15212];
  assign N13615 = N13614 | data_masked[15340];
  assign N13614 = N13613 | data_masked[15468];
  assign N13613 = N13612 | data_masked[15596];
  assign N13612 = N13611 | data_masked[15724];
  assign N13611 = N13610 | data_masked[15852];
  assign N13610 = N13609 | data_masked[15980];
  assign N13609 = N13608 | data_masked[16108];
  assign N13608 = data_masked[16364] | data_masked[16236];
  assign data_o[109] = N13859 | data_masked[109];
  assign N13859 = N13858 | data_masked[237];
  assign N13858 = N13857 | data_masked[365];
  assign N13857 = N13856 | data_masked[493];
  assign N13856 = N13855 | data_masked[621];
  assign N13855 = N13854 | data_masked[749];
  assign N13854 = N13853 | data_masked[877];
  assign N13853 = N13852 | data_masked[1005];
  assign N13852 = N13851 | data_masked[1133];
  assign N13851 = N13850 | data_masked[1261];
  assign N13850 = N13849 | data_masked[1389];
  assign N13849 = N13848 | data_masked[1517];
  assign N13848 = N13847 | data_masked[1645];
  assign N13847 = N13846 | data_masked[1773];
  assign N13846 = N13845 | data_masked[1901];
  assign N13845 = N13844 | data_masked[2029];
  assign N13844 = N13843 | data_masked[2157];
  assign N13843 = N13842 | data_masked[2285];
  assign N13842 = N13841 | data_masked[2413];
  assign N13841 = N13840 | data_masked[2541];
  assign N13840 = N13839 | data_masked[2669];
  assign N13839 = N13838 | data_masked[2797];
  assign N13838 = N13837 | data_masked[2925];
  assign N13837 = N13836 | data_masked[3053];
  assign N13836 = N13835 | data_masked[3181];
  assign N13835 = N13834 | data_masked[3309];
  assign N13834 = N13833 | data_masked[3437];
  assign N13833 = N13832 | data_masked[3565];
  assign N13832 = N13831 | data_masked[3693];
  assign N13831 = N13830 | data_masked[3821];
  assign N13830 = N13829 | data_masked[3949];
  assign N13829 = N13828 | data_masked[4077];
  assign N13828 = N13827 | data_masked[4205];
  assign N13827 = N13826 | data_masked[4333];
  assign N13826 = N13825 | data_masked[4461];
  assign N13825 = N13824 | data_masked[4589];
  assign N13824 = N13823 | data_masked[4717];
  assign N13823 = N13822 | data_masked[4845];
  assign N13822 = N13821 | data_masked[4973];
  assign N13821 = N13820 | data_masked[5101];
  assign N13820 = N13819 | data_masked[5229];
  assign N13819 = N13818 | data_masked[5357];
  assign N13818 = N13817 | data_masked[5485];
  assign N13817 = N13816 | data_masked[5613];
  assign N13816 = N13815 | data_masked[5741];
  assign N13815 = N13814 | data_masked[5869];
  assign N13814 = N13813 | data_masked[5997];
  assign N13813 = N13812 | data_masked[6125];
  assign N13812 = N13811 | data_masked[6253];
  assign N13811 = N13810 | data_masked[6381];
  assign N13810 = N13809 | data_masked[6509];
  assign N13809 = N13808 | data_masked[6637];
  assign N13808 = N13807 | data_masked[6765];
  assign N13807 = N13806 | data_masked[6893];
  assign N13806 = N13805 | data_masked[7021];
  assign N13805 = N13804 | data_masked[7149];
  assign N13804 = N13803 | data_masked[7277];
  assign N13803 = N13802 | data_masked[7405];
  assign N13802 = N13801 | data_masked[7533];
  assign N13801 = N13800 | data_masked[7661];
  assign N13800 = N13799 | data_masked[7789];
  assign N13799 = N13798 | data_masked[7917];
  assign N13798 = N13797 | data_masked[8045];
  assign N13797 = N13796 | data_masked[8173];
  assign N13796 = N13795 | data_masked[8301];
  assign N13795 = N13794 | data_masked[8429];
  assign N13794 = N13793 | data_masked[8557];
  assign N13793 = N13792 | data_masked[8685];
  assign N13792 = N13791 | data_masked[8813];
  assign N13791 = N13790 | data_masked[8941];
  assign N13790 = N13789 | data_masked[9069];
  assign N13789 = N13788 | data_masked[9197];
  assign N13788 = N13787 | data_masked[9325];
  assign N13787 = N13786 | data_masked[9453];
  assign N13786 = N13785 | data_masked[9581];
  assign N13785 = N13784 | data_masked[9709];
  assign N13784 = N13783 | data_masked[9837];
  assign N13783 = N13782 | data_masked[9965];
  assign N13782 = N13781 | data_masked[10093];
  assign N13781 = N13780 | data_masked[10221];
  assign N13780 = N13779 | data_masked[10349];
  assign N13779 = N13778 | data_masked[10477];
  assign N13778 = N13777 | data_masked[10605];
  assign N13777 = N13776 | data_masked[10733];
  assign N13776 = N13775 | data_masked[10861];
  assign N13775 = N13774 | data_masked[10989];
  assign N13774 = N13773 | data_masked[11117];
  assign N13773 = N13772 | data_masked[11245];
  assign N13772 = N13771 | data_masked[11373];
  assign N13771 = N13770 | data_masked[11501];
  assign N13770 = N13769 | data_masked[11629];
  assign N13769 = N13768 | data_masked[11757];
  assign N13768 = N13767 | data_masked[11885];
  assign N13767 = N13766 | data_masked[12013];
  assign N13766 = N13765 | data_masked[12141];
  assign N13765 = N13764 | data_masked[12269];
  assign N13764 = N13763 | data_masked[12397];
  assign N13763 = N13762 | data_masked[12525];
  assign N13762 = N13761 | data_masked[12653];
  assign N13761 = N13760 | data_masked[12781];
  assign N13760 = N13759 | data_masked[12909];
  assign N13759 = N13758 | data_masked[13037];
  assign N13758 = N13757 | data_masked[13165];
  assign N13757 = N13756 | data_masked[13293];
  assign N13756 = N13755 | data_masked[13421];
  assign N13755 = N13754 | data_masked[13549];
  assign N13754 = N13753 | data_masked[13677];
  assign N13753 = N13752 | data_masked[13805];
  assign N13752 = N13751 | data_masked[13933];
  assign N13751 = N13750 | data_masked[14061];
  assign N13750 = N13749 | data_masked[14189];
  assign N13749 = N13748 | data_masked[14317];
  assign N13748 = N13747 | data_masked[14445];
  assign N13747 = N13746 | data_masked[14573];
  assign N13746 = N13745 | data_masked[14701];
  assign N13745 = N13744 | data_masked[14829];
  assign N13744 = N13743 | data_masked[14957];
  assign N13743 = N13742 | data_masked[15085];
  assign N13742 = N13741 | data_masked[15213];
  assign N13741 = N13740 | data_masked[15341];
  assign N13740 = N13739 | data_masked[15469];
  assign N13739 = N13738 | data_masked[15597];
  assign N13738 = N13737 | data_masked[15725];
  assign N13737 = N13736 | data_masked[15853];
  assign N13736 = N13735 | data_masked[15981];
  assign N13735 = N13734 | data_masked[16109];
  assign N13734 = data_masked[16365] | data_masked[16237];
  assign data_o[110] = N13985 | data_masked[110];
  assign N13985 = N13984 | data_masked[238];
  assign N13984 = N13983 | data_masked[366];
  assign N13983 = N13982 | data_masked[494];
  assign N13982 = N13981 | data_masked[622];
  assign N13981 = N13980 | data_masked[750];
  assign N13980 = N13979 | data_masked[878];
  assign N13979 = N13978 | data_masked[1006];
  assign N13978 = N13977 | data_masked[1134];
  assign N13977 = N13976 | data_masked[1262];
  assign N13976 = N13975 | data_masked[1390];
  assign N13975 = N13974 | data_masked[1518];
  assign N13974 = N13973 | data_masked[1646];
  assign N13973 = N13972 | data_masked[1774];
  assign N13972 = N13971 | data_masked[1902];
  assign N13971 = N13970 | data_masked[2030];
  assign N13970 = N13969 | data_masked[2158];
  assign N13969 = N13968 | data_masked[2286];
  assign N13968 = N13967 | data_masked[2414];
  assign N13967 = N13966 | data_masked[2542];
  assign N13966 = N13965 | data_masked[2670];
  assign N13965 = N13964 | data_masked[2798];
  assign N13964 = N13963 | data_masked[2926];
  assign N13963 = N13962 | data_masked[3054];
  assign N13962 = N13961 | data_masked[3182];
  assign N13961 = N13960 | data_masked[3310];
  assign N13960 = N13959 | data_masked[3438];
  assign N13959 = N13958 | data_masked[3566];
  assign N13958 = N13957 | data_masked[3694];
  assign N13957 = N13956 | data_masked[3822];
  assign N13956 = N13955 | data_masked[3950];
  assign N13955 = N13954 | data_masked[4078];
  assign N13954 = N13953 | data_masked[4206];
  assign N13953 = N13952 | data_masked[4334];
  assign N13952 = N13951 | data_masked[4462];
  assign N13951 = N13950 | data_masked[4590];
  assign N13950 = N13949 | data_masked[4718];
  assign N13949 = N13948 | data_masked[4846];
  assign N13948 = N13947 | data_masked[4974];
  assign N13947 = N13946 | data_masked[5102];
  assign N13946 = N13945 | data_masked[5230];
  assign N13945 = N13944 | data_masked[5358];
  assign N13944 = N13943 | data_masked[5486];
  assign N13943 = N13942 | data_masked[5614];
  assign N13942 = N13941 | data_masked[5742];
  assign N13941 = N13940 | data_masked[5870];
  assign N13940 = N13939 | data_masked[5998];
  assign N13939 = N13938 | data_masked[6126];
  assign N13938 = N13937 | data_masked[6254];
  assign N13937 = N13936 | data_masked[6382];
  assign N13936 = N13935 | data_masked[6510];
  assign N13935 = N13934 | data_masked[6638];
  assign N13934 = N13933 | data_masked[6766];
  assign N13933 = N13932 | data_masked[6894];
  assign N13932 = N13931 | data_masked[7022];
  assign N13931 = N13930 | data_masked[7150];
  assign N13930 = N13929 | data_masked[7278];
  assign N13929 = N13928 | data_masked[7406];
  assign N13928 = N13927 | data_masked[7534];
  assign N13927 = N13926 | data_masked[7662];
  assign N13926 = N13925 | data_masked[7790];
  assign N13925 = N13924 | data_masked[7918];
  assign N13924 = N13923 | data_masked[8046];
  assign N13923 = N13922 | data_masked[8174];
  assign N13922 = N13921 | data_masked[8302];
  assign N13921 = N13920 | data_masked[8430];
  assign N13920 = N13919 | data_masked[8558];
  assign N13919 = N13918 | data_masked[8686];
  assign N13918 = N13917 | data_masked[8814];
  assign N13917 = N13916 | data_masked[8942];
  assign N13916 = N13915 | data_masked[9070];
  assign N13915 = N13914 | data_masked[9198];
  assign N13914 = N13913 | data_masked[9326];
  assign N13913 = N13912 | data_masked[9454];
  assign N13912 = N13911 | data_masked[9582];
  assign N13911 = N13910 | data_masked[9710];
  assign N13910 = N13909 | data_masked[9838];
  assign N13909 = N13908 | data_masked[9966];
  assign N13908 = N13907 | data_masked[10094];
  assign N13907 = N13906 | data_masked[10222];
  assign N13906 = N13905 | data_masked[10350];
  assign N13905 = N13904 | data_masked[10478];
  assign N13904 = N13903 | data_masked[10606];
  assign N13903 = N13902 | data_masked[10734];
  assign N13902 = N13901 | data_masked[10862];
  assign N13901 = N13900 | data_masked[10990];
  assign N13900 = N13899 | data_masked[11118];
  assign N13899 = N13898 | data_masked[11246];
  assign N13898 = N13897 | data_masked[11374];
  assign N13897 = N13896 | data_masked[11502];
  assign N13896 = N13895 | data_masked[11630];
  assign N13895 = N13894 | data_masked[11758];
  assign N13894 = N13893 | data_masked[11886];
  assign N13893 = N13892 | data_masked[12014];
  assign N13892 = N13891 | data_masked[12142];
  assign N13891 = N13890 | data_masked[12270];
  assign N13890 = N13889 | data_masked[12398];
  assign N13889 = N13888 | data_masked[12526];
  assign N13888 = N13887 | data_masked[12654];
  assign N13887 = N13886 | data_masked[12782];
  assign N13886 = N13885 | data_masked[12910];
  assign N13885 = N13884 | data_masked[13038];
  assign N13884 = N13883 | data_masked[13166];
  assign N13883 = N13882 | data_masked[13294];
  assign N13882 = N13881 | data_masked[13422];
  assign N13881 = N13880 | data_masked[13550];
  assign N13880 = N13879 | data_masked[13678];
  assign N13879 = N13878 | data_masked[13806];
  assign N13878 = N13877 | data_masked[13934];
  assign N13877 = N13876 | data_masked[14062];
  assign N13876 = N13875 | data_masked[14190];
  assign N13875 = N13874 | data_masked[14318];
  assign N13874 = N13873 | data_masked[14446];
  assign N13873 = N13872 | data_masked[14574];
  assign N13872 = N13871 | data_masked[14702];
  assign N13871 = N13870 | data_masked[14830];
  assign N13870 = N13869 | data_masked[14958];
  assign N13869 = N13868 | data_masked[15086];
  assign N13868 = N13867 | data_masked[15214];
  assign N13867 = N13866 | data_masked[15342];
  assign N13866 = N13865 | data_masked[15470];
  assign N13865 = N13864 | data_masked[15598];
  assign N13864 = N13863 | data_masked[15726];
  assign N13863 = N13862 | data_masked[15854];
  assign N13862 = N13861 | data_masked[15982];
  assign N13861 = N13860 | data_masked[16110];
  assign N13860 = data_masked[16366] | data_masked[16238];
  assign data_o[111] = N14111 | data_masked[111];
  assign N14111 = N14110 | data_masked[239];
  assign N14110 = N14109 | data_masked[367];
  assign N14109 = N14108 | data_masked[495];
  assign N14108 = N14107 | data_masked[623];
  assign N14107 = N14106 | data_masked[751];
  assign N14106 = N14105 | data_masked[879];
  assign N14105 = N14104 | data_masked[1007];
  assign N14104 = N14103 | data_masked[1135];
  assign N14103 = N14102 | data_masked[1263];
  assign N14102 = N14101 | data_masked[1391];
  assign N14101 = N14100 | data_masked[1519];
  assign N14100 = N14099 | data_masked[1647];
  assign N14099 = N14098 | data_masked[1775];
  assign N14098 = N14097 | data_masked[1903];
  assign N14097 = N14096 | data_masked[2031];
  assign N14096 = N14095 | data_masked[2159];
  assign N14095 = N14094 | data_masked[2287];
  assign N14094 = N14093 | data_masked[2415];
  assign N14093 = N14092 | data_masked[2543];
  assign N14092 = N14091 | data_masked[2671];
  assign N14091 = N14090 | data_masked[2799];
  assign N14090 = N14089 | data_masked[2927];
  assign N14089 = N14088 | data_masked[3055];
  assign N14088 = N14087 | data_masked[3183];
  assign N14087 = N14086 | data_masked[3311];
  assign N14086 = N14085 | data_masked[3439];
  assign N14085 = N14084 | data_masked[3567];
  assign N14084 = N14083 | data_masked[3695];
  assign N14083 = N14082 | data_masked[3823];
  assign N14082 = N14081 | data_masked[3951];
  assign N14081 = N14080 | data_masked[4079];
  assign N14080 = N14079 | data_masked[4207];
  assign N14079 = N14078 | data_masked[4335];
  assign N14078 = N14077 | data_masked[4463];
  assign N14077 = N14076 | data_masked[4591];
  assign N14076 = N14075 | data_masked[4719];
  assign N14075 = N14074 | data_masked[4847];
  assign N14074 = N14073 | data_masked[4975];
  assign N14073 = N14072 | data_masked[5103];
  assign N14072 = N14071 | data_masked[5231];
  assign N14071 = N14070 | data_masked[5359];
  assign N14070 = N14069 | data_masked[5487];
  assign N14069 = N14068 | data_masked[5615];
  assign N14068 = N14067 | data_masked[5743];
  assign N14067 = N14066 | data_masked[5871];
  assign N14066 = N14065 | data_masked[5999];
  assign N14065 = N14064 | data_masked[6127];
  assign N14064 = N14063 | data_masked[6255];
  assign N14063 = N14062 | data_masked[6383];
  assign N14062 = N14061 | data_masked[6511];
  assign N14061 = N14060 | data_masked[6639];
  assign N14060 = N14059 | data_masked[6767];
  assign N14059 = N14058 | data_masked[6895];
  assign N14058 = N14057 | data_masked[7023];
  assign N14057 = N14056 | data_masked[7151];
  assign N14056 = N14055 | data_masked[7279];
  assign N14055 = N14054 | data_masked[7407];
  assign N14054 = N14053 | data_masked[7535];
  assign N14053 = N14052 | data_masked[7663];
  assign N14052 = N14051 | data_masked[7791];
  assign N14051 = N14050 | data_masked[7919];
  assign N14050 = N14049 | data_masked[8047];
  assign N14049 = N14048 | data_masked[8175];
  assign N14048 = N14047 | data_masked[8303];
  assign N14047 = N14046 | data_masked[8431];
  assign N14046 = N14045 | data_masked[8559];
  assign N14045 = N14044 | data_masked[8687];
  assign N14044 = N14043 | data_masked[8815];
  assign N14043 = N14042 | data_masked[8943];
  assign N14042 = N14041 | data_masked[9071];
  assign N14041 = N14040 | data_masked[9199];
  assign N14040 = N14039 | data_masked[9327];
  assign N14039 = N14038 | data_masked[9455];
  assign N14038 = N14037 | data_masked[9583];
  assign N14037 = N14036 | data_masked[9711];
  assign N14036 = N14035 | data_masked[9839];
  assign N14035 = N14034 | data_masked[9967];
  assign N14034 = N14033 | data_masked[10095];
  assign N14033 = N14032 | data_masked[10223];
  assign N14032 = N14031 | data_masked[10351];
  assign N14031 = N14030 | data_masked[10479];
  assign N14030 = N14029 | data_masked[10607];
  assign N14029 = N14028 | data_masked[10735];
  assign N14028 = N14027 | data_masked[10863];
  assign N14027 = N14026 | data_masked[10991];
  assign N14026 = N14025 | data_masked[11119];
  assign N14025 = N14024 | data_masked[11247];
  assign N14024 = N14023 | data_masked[11375];
  assign N14023 = N14022 | data_masked[11503];
  assign N14022 = N14021 | data_masked[11631];
  assign N14021 = N14020 | data_masked[11759];
  assign N14020 = N14019 | data_masked[11887];
  assign N14019 = N14018 | data_masked[12015];
  assign N14018 = N14017 | data_masked[12143];
  assign N14017 = N14016 | data_masked[12271];
  assign N14016 = N14015 | data_masked[12399];
  assign N14015 = N14014 | data_masked[12527];
  assign N14014 = N14013 | data_masked[12655];
  assign N14013 = N14012 | data_masked[12783];
  assign N14012 = N14011 | data_masked[12911];
  assign N14011 = N14010 | data_masked[13039];
  assign N14010 = N14009 | data_masked[13167];
  assign N14009 = N14008 | data_masked[13295];
  assign N14008 = N14007 | data_masked[13423];
  assign N14007 = N14006 | data_masked[13551];
  assign N14006 = N14005 | data_masked[13679];
  assign N14005 = N14004 | data_masked[13807];
  assign N14004 = N14003 | data_masked[13935];
  assign N14003 = N14002 | data_masked[14063];
  assign N14002 = N14001 | data_masked[14191];
  assign N14001 = N14000 | data_masked[14319];
  assign N14000 = N13999 | data_masked[14447];
  assign N13999 = N13998 | data_masked[14575];
  assign N13998 = N13997 | data_masked[14703];
  assign N13997 = N13996 | data_masked[14831];
  assign N13996 = N13995 | data_masked[14959];
  assign N13995 = N13994 | data_masked[15087];
  assign N13994 = N13993 | data_masked[15215];
  assign N13993 = N13992 | data_masked[15343];
  assign N13992 = N13991 | data_masked[15471];
  assign N13991 = N13990 | data_masked[15599];
  assign N13990 = N13989 | data_masked[15727];
  assign N13989 = N13988 | data_masked[15855];
  assign N13988 = N13987 | data_masked[15983];
  assign N13987 = N13986 | data_masked[16111];
  assign N13986 = data_masked[16367] | data_masked[16239];
  assign data_o[112] = N14237 | data_masked[112];
  assign N14237 = N14236 | data_masked[240];
  assign N14236 = N14235 | data_masked[368];
  assign N14235 = N14234 | data_masked[496];
  assign N14234 = N14233 | data_masked[624];
  assign N14233 = N14232 | data_masked[752];
  assign N14232 = N14231 | data_masked[880];
  assign N14231 = N14230 | data_masked[1008];
  assign N14230 = N14229 | data_masked[1136];
  assign N14229 = N14228 | data_masked[1264];
  assign N14228 = N14227 | data_masked[1392];
  assign N14227 = N14226 | data_masked[1520];
  assign N14226 = N14225 | data_masked[1648];
  assign N14225 = N14224 | data_masked[1776];
  assign N14224 = N14223 | data_masked[1904];
  assign N14223 = N14222 | data_masked[2032];
  assign N14222 = N14221 | data_masked[2160];
  assign N14221 = N14220 | data_masked[2288];
  assign N14220 = N14219 | data_masked[2416];
  assign N14219 = N14218 | data_masked[2544];
  assign N14218 = N14217 | data_masked[2672];
  assign N14217 = N14216 | data_masked[2800];
  assign N14216 = N14215 | data_masked[2928];
  assign N14215 = N14214 | data_masked[3056];
  assign N14214 = N14213 | data_masked[3184];
  assign N14213 = N14212 | data_masked[3312];
  assign N14212 = N14211 | data_masked[3440];
  assign N14211 = N14210 | data_masked[3568];
  assign N14210 = N14209 | data_masked[3696];
  assign N14209 = N14208 | data_masked[3824];
  assign N14208 = N14207 | data_masked[3952];
  assign N14207 = N14206 | data_masked[4080];
  assign N14206 = N14205 | data_masked[4208];
  assign N14205 = N14204 | data_masked[4336];
  assign N14204 = N14203 | data_masked[4464];
  assign N14203 = N14202 | data_masked[4592];
  assign N14202 = N14201 | data_masked[4720];
  assign N14201 = N14200 | data_masked[4848];
  assign N14200 = N14199 | data_masked[4976];
  assign N14199 = N14198 | data_masked[5104];
  assign N14198 = N14197 | data_masked[5232];
  assign N14197 = N14196 | data_masked[5360];
  assign N14196 = N14195 | data_masked[5488];
  assign N14195 = N14194 | data_masked[5616];
  assign N14194 = N14193 | data_masked[5744];
  assign N14193 = N14192 | data_masked[5872];
  assign N14192 = N14191 | data_masked[6000];
  assign N14191 = N14190 | data_masked[6128];
  assign N14190 = N14189 | data_masked[6256];
  assign N14189 = N14188 | data_masked[6384];
  assign N14188 = N14187 | data_masked[6512];
  assign N14187 = N14186 | data_masked[6640];
  assign N14186 = N14185 | data_masked[6768];
  assign N14185 = N14184 | data_masked[6896];
  assign N14184 = N14183 | data_masked[7024];
  assign N14183 = N14182 | data_masked[7152];
  assign N14182 = N14181 | data_masked[7280];
  assign N14181 = N14180 | data_masked[7408];
  assign N14180 = N14179 | data_masked[7536];
  assign N14179 = N14178 | data_masked[7664];
  assign N14178 = N14177 | data_masked[7792];
  assign N14177 = N14176 | data_masked[7920];
  assign N14176 = N14175 | data_masked[8048];
  assign N14175 = N14174 | data_masked[8176];
  assign N14174 = N14173 | data_masked[8304];
  assign N14173 = N14172 | data_masked[8432];
  assign N14172 = N14171 | data_masked[8560];
  assign N14171 = N14170 | data_masked[8688];
  assign N14170 = N14169 | data_masked[8816];
  assign N14169 = N14168 | data_masked[8944];
  assign N14168 = N14167 | data_masked[9072];
  assign N14167 = N14166 | data_masked[9200];
  assign N14166 = N14165 | data_masked[9328];
  assign N14165 = N14164 | data_masked[9456];
  assign N14164 = N14163 | data_masked[9584];
  assign N14163 = N14162 | data_masked[9712];
  assign N14162 = N14161 | data_masked[9840];
  assign N14161 = N14160 | data_masked[9968];
  assign N14160 = N14159 | data_masked[10096];
  assign N14159 = N14158 | data_masked[10224];
  assign N14158 = N14157 | data_masked[10352];
  assign N14157 = N14156 | data_masked[10480];
  assign N14156 = N14155 | data_masked[10608];
  assign N14155 = N14154 | data_masked[10736];
  assign N14154 = N14153 | data_masked[10864];
  assign N14153 = N14152 | data_masked[10992];
  assign N14152 = N14151 | data_masked[11120];
  assign N14151 = N14150 | data_masked[11248];
  assign N14150 = N14149 | data_masked[11376];
  assign N14149 = N14148 | data_masked[11504];
  assign N14148 = N14147 | data_masked[11632];
  assign N14147 = N14146 | data_masked[11760];
  assign N14146 = N14145 | data_masked[11888];
  assign N14145 = N14144 | data_masked[12016];
  assign N14144 = N14143 | data_masked[12144];
  assign N14143 = N14142 | data_masked[12272];
  assign N14142 = N14141 | data_masked[12400];
  assign N14141 = N14140 | data_masked[12528];
  assign N14140 = N14139 | data_masked[12656];
  assign N14139 = N14138 | data_masked[12784];
  assign N14138 = N14137 | data_masked[12912];
  assign N14137 = N14136 | data_masked[13040];
  assign N14136 = N14135 | data_masked[13168];
  assign N14135 = N14134 | data_masked[13296];
  assign N14134 = N14133 | data_masked[13424];
  assign N14133 = N14132 | data_masked[13552];
  assign N14132 = N14131 | data_masked[13680];
  assign N14131 = N14130 | data_masked[13808];
  assign N14130 = N14129 | data_masked[13936];
  assign N14129 = N14128 | data_masked[14064];
  assign N14128 = N14127 | data_masked[14192];
  assign N14127 = N14126 | data_masked[14320];
  assign N14126 = N14125 | data_masked[14448];
  assign N14125 = N14124 | data_masked[14576];
  assign N14124 = N14123 | data_masked[14704];
  assign N14123 = N14122 | data_masked[14832];
  assign N14122 = N14121 | data_masked[14960];
  assign N14121 = N14120 | data_masked[15088];
  assign N14120 = N14119 | data_masked[15216];
  assign N14119 = N14118 | data_masked[15344];
  assign N14118 = N14117 | data_masked[15472];
  assign N14117 = N14116 | data_masked[15600];
  assign N14116 = N14115 | data_masked[15728];
  assign N14115 = N14114 | data_masked[15856];
  assign N14114 = N14113 | data_masked[15984];
  assign N14113 = N14112 | data_masked[16112];
  assign N14112 = data_masked[16368] | data_masked[16240];
  assign data_o[113] = N14363 | data_masked[113];
  assign N14363 = N14362 | data_masked[241];
  assign N14362 = N14361 | data_masked[369];
  assign N14361 = N14360 | data_masked[497];
  assign N14360 = N14359 | data_masked[625];
  assign N14359 = N14358 | data_masked[753];
  assign N14358 = N14357 | data_masked[881];
  assign N14357 = N14356 | data_masked[1009];
  assign N14356 = N14355 | data_masked[1137];
  assign N14355 = N14354 | data_masked[1265];
  assign N14354 = N14353 | data_masked[1393];
  assign N14353 = N14352 | data_masked[1521];
  assign N14352 = N14351 | data_masked[1649];
  assign N14351 = N14350 | data_masked[1777];
  assign N14350 = N14349 | data_masked[1905];
  assign N14349 = N14348 | data_masked[2033];
  assign N14348 = N14347 | data_masked[2161];
  assign N14347 = N14346 | data_masked[2289];
  assign N14346 = N14345 | data_masked[2417];
  assign N14345 = N14344 | data_masked[2545];
  assign N14344 = N14343 | data_masked[2673];
  assign N14343 = N14342 | data_masked[2801];
  assign N14342 = N14341 | data_masked[2929];
  assign N14341 = N14340 | data_masked[3057];
  assign N14340 = N14339 | data_masked[3185];
  assign N14339 = N14338 | data_masked[3313];
  assign N14338 = N14337 | data_masked[3441];
  assign N14337 = N14336 | data_masked[3569];
  assign N14336 = N14335 | data_masked[3697];
  assign N14335 = N14334 | data_masked[3825];
  assign N14334 = N14333 | data_masked[3953];
  assign N14333 = N14332 | data_masked[4081];
  assign N14332 = N14331 | data_masked[4209];
  assign N14331 = N14330 | data_masked[4337];
  assign N14330 = N14329 | data_masked[4465];
  assign N14329 = N14328 | data_masked[4593];
  assign N14328 = N14327 | data_masked[4721];
  assign N14327 = N14326 | data_masked[4849];
  assign N14326 = N14325 | data_masked[4977];
  assign N14325 = N14324 | data_masked[5105];
  assign N14324 = N14323 | data_masked[5233];
  assign N14323 = N14322 | data_masked[5361];
  assign N14322 = N14321 | data_masked[5489];
  assign N14321 = N14320 | data_masked[5617];
  assign N14320 = N14319 | data_masked[5745];
  assign N14319 = N14318 | data_masked[5873];
  assign N14318 = N14317 | data_masked[6001];
  assign N14317 = N14316 | data_masked[6129];
  assign N14316 = N14315 | data_masked[6257];
  assign N14315 = N14314 | data_masked[6385];
  assign N14314 = N14313 | data_masked[6513];
  assign N14313 = N14312 | data_masked[6641];
  assign N14312 = N14311 | data_masked[6769];
  assign N14311 = N14310 | data_masked[6897];
  assign N14310 = N14309 | data_masked[7025];
  assign N14309 = N14308 | data_masked[7153];
  assign N14308 = N14307 | data_masked[7281];
  assign N14307 = N14306 | data_masked[7409];
  assign N14306 = N14305 | data_masked[7537];
  assign N14305 = N14304 | data_masked[7665];
  assign N14304 = N14303 | data_masked[7793];
  assign N14303 = N14302 | data_masked[7921];
  assign N14302 = N14301 | data_masked[8049];
  assign N14301 = N14300 | data_masked[8177];
  assign N14300 = N14299 | data_masked[8305];
  assign N14299 = N14298 | data_masked[8433];
  assign N14298 = N14297 | data_masked[8561];
  assign N14297 = N14296 | data_masked[8689];
  assign N14296 = N14295 | data_masked[8817];
  assign N14295 = N14294 | data_masked[8945];
  assign N14294 = N14293 | data_masked[9073];
  assign N14293 = N14292 | data_masked[9201];
  assign N14292 = N14291 | data_masked[9329];
  assign N14291 = N14290 | data_masked[9457];
  assign N14290 = N14289 | data_masked[9585];
  assign N14289 = N14288 | data_masked[9713];
  assign N14288 = N14287 | data_masked[9841];
  assign N14287 = N14286 | data_masked[9969];
  assign N14286 = N14285 | data_masked[10097];
  assign N14285 = N14284 | data_masked[10225];
  assign N14284 = N14283 | data_masked[10353];
  assign N14283 = N14282 | data_masked[10481];
  assign N14282 = N14281 | data_masked[10609];
  assign N14281 = N14280 | data_masked[10737];
  assign N14280 = N14279 | data_masked[10865];
  assign N14279 = N14278 | data_masked[10993];
  assign N14278 = N14277 | data_masked[11121];
  assign N14277 = N14276 | data_masked[11249];
  assign N14276 = N14275 | data_masked[11377];
  assign N14275 = N14274 | data_masked[11505];
  assign N14274 = N14273 | data_masked[11633];
  assign N14273 = N14272 | data_masked[11761];
  assign N14272 = N14271 | data_masked[11889];
  assign N14271 = N14270 | data_masked[12017];
  assign N14270 = N14269 | data_masked[12145];
  assign N14269 = N14268 | data_masked[12273];
  assign N14268 = N14267 | data_masked[12401];
  assign N14267 = N14266 | data_masked[12529];
  assign N14266 = N14265 | data_masked[12657];
  assign N14265 = N14264 | data_masked[12785];
  assign N14264 = N14263 | data_masked[12913];
  assign N14263 = N14262 | data_masked[13041];
  assign N14262 = N14261 | data_masked[13169];
  assign N14261 = N14260 | data_masked[13297];
  assign N14260 = N14259 | data_masked[13425];
  assign N14259 = N14258 | data_masked[13553];
  assign N14258 = N14257 | data_masked[13681];
  assign N14257 = N14256 | data_masked[13809];
  assign N14256 = N14255 | data_masked[13937];
  assign N14255 = N14254 | data_masked[14065];
  assign N14254 = N14253 | data_masked[14193];
  assign N14253 = N14252 | data_masked[14321];
  assign N14252 = N14251 | data_masked[14449];
  assign N14251 = N14250 | data_masked[14577];
  assign N14250 = N14249 | data_masked[14705];
  assign N14249 = N14248 | data_masked[14833];
  assign N14248 = N14247 | data_masked[14961];
  assign N14247 = N14246 | data_masked[15089];
  assign N14246 = N14245 | data_masked[15217];
  assign N14245 = N14244 | data_masked[15345];
  assign N14244 = N14243 | data_masked[15473];
  assign N14243 = N14242 | data_masked[15601];
  assign N14242 = N14241 | data_masked[15729];
  assign N14241 = N14240 | data_masked[15857];
  assign N14240 = N14239 | data_masked[15985];
  assign N14239 = N14238 | data_masked[16113];
  assign N14238 = data_masked[16369] | data_masked[16241];
  assign data_o[114] = N14489 | data_masked[114];
  assign N14489 = N14488 | data_masked[242];
  assign N14488 = N14487 | data_masked[370];
  assign N14487 = N14486 | data_masked[498];
  assign N14486 = N14485 | data_masked[626];
  assign N14485 = N14484 | data_masked[754];
  assign N14484 = N14483 | data_masked[882];
  assign N14483 = N14482 | data_masked[1010];
  assign N14482 = N14481 | data_masked[1138];
  assign N14481 = N14480 | data_masked[1266];
  assign N14480 = N14479 | data_masked[1394];
  assign N14479 = N14478 | data_masked[1522];
  assign N14478 = N14477 | data_masked[1650];
  assign N14477 = N14476 | data_masked[1778];
  assign N14476 = N14475 | data_masked[1906];
  assign N14475 = N14474 | data_masked[2034];
  assign N14474 = N14473 | data_masked[2162];
  assign N14473 = N14472 | data_masked[2290];
  assign N14472 = N14471 | data_masked[2418];
  assign N14471 = N14470 | data_masked[2546];
  assign N14470 = N14469 | data_masked[2674];
  assign N14469 = N14468 | data_masked[2802];
  assign N14468 = N14467 | data_masked[2930];
  assign N14467 = N14466 | data_masked[3058];
  assign N14466 = N14465 | data_masked[3186];
  assign N14465 = N14464 | data_masked[3314];
  assign N14464 = N14463 | data_masked[3442];
  assign N14463 = N14462 | data_masked[3570];
  assign N14462 = N14461 | data_masked[3698];
  assign N14461 = N14460 | data_masked[3826];
  assign N14460 = N14459 | data_masked[3954];
  assign N14459 = N14458 | data_masked[4082];
  assign N14458 = N14457 | data_masked[4210];
  assign N14457 = N14456 | data_masked[4338];
  assign N14456 = N14455 | data_masked[4466];
  assign N14455 = N14454 | data_masked[4594];
  assign N14454 = N14453 | data_masked[4722];
  assign N14453 = N14452 | data_masked[4850];
  assign N14452 = N14451 | data_masked[4978];
  assign N14451 = N14450 | data_masked[5106];
  assign N14450 = N14449 | data_masked[5234];
  assign N14449 = N14448 | data_masked[5362];
  assign N14448 = N14447 | data_masked[5490];
  assign N14447 = N14446 | data_masked[5618];
  assign N14446 = N14445 | data_masked[5746];
  assign N14445 = N14444 | data_masked[5874];
  assign N14444 = N14443 | data_masked[6002];
  assign N14443 = N14442 | data_masked[6130];
  assign N14442 = N14441 | data_masked[6258];
  assign N14441 = N14440 | data_masked[6386];
  assign N14440 = N14439 | data_masked[6514];
  assign N14439 = N14438 | data_masked[6642];
  assign N14438 = N14437 | data_masked[6770];
  assign N14437 = N14436 | data_masked[6898];
  assign N14436 = N14435 | data_masked[7026];
  assign N14435 = N14434 | data_masked[7154];
  assign N14434 = N14433 | data_masked[7282];
  assign N14433 = N14432 | data_masked[7410];
  assign N14432 = N14431 | data_masked[7538];
  assign N14431 = N14430 | data_masked[7666];
  assign N14430 = N14429 | data_masked[7794];
  assign N14429 = N14428 | data_masked[7922];
  assign N14428 = N14427 | data_masked[8050];
  assign N14427 = N14426 | data_masked[8178];
  assign N14426 = N14425 | data_masked[8306];
  assign N14425 = N14424 | data_masked[8434];
  assign N14424 = N14423 | data_masked[8562];
  assign N14423 = N14422 | data_masked[8690];
  assign N14422 = N14421 | data_masked[8818];
  assign N14421 = N14420 | data_masked[8946];
  assign N14420 = N14419 | data_masked[9074];
  assign N14419 = N14418 | data_masked[9202];
  assign N14418 = N14417 | data_masked[9330];
  assign N14417 = N14416 | data_masked[9458];
  assign N14416 = N14415 | data_masked[9586];
  assign N14415 = N14414 | data_masked[9714];
  assign N14414 = N14413 | data_masked[9842];
  assign N14413 = N14412 | data_masked[9970];
  assign N14412 = N14411 | data_masked[10098];
  assign N14411 = N14410 | data_masked[10226];
  assign N14410 = N14409 | data_masked[10354];
  assign N14409 = N14408 | data_masked[10482];
  assign N14408 = N14407 | data_masked[10610];
  assign N14407 = N14406 | data_masked[10738];
  assign N14406 = N14405 | data_masked[10866];
  assign N14405 = N14404 | data_masked[10994];
  assign N14404 = N14403 | data_masked[11122];
  assign N14403 = N14402 | data_masked[11250];
  assign N14402 = N14401 | data_masked[11378];
  assign N14401 = N14400 | data_masked[11506];
  assign N14400 = N14399 | data_masked[11634];
  assign N14399 = N14398 | data_masked[11762];
  assign N14398 = N14397 | data_masked[11890];
  assign N14397 = N14396 | data_masked[12018];
  assign N14396 = N14395 | data_masked[12146];
  assign N14395 = N14394 | data_masked[12274];
  assign N14394 = N14393 | data_masked[12402];
  assign N14393 = N14392 | data_masked[12530];
  assign N14392 = N14391 | data_masked[12658];
  assign N14391 = N14390 | data_masked[12786];
  assign N14390 = N14389 | data_masked[12914];
  assign N14389 = N14388 | data_masked[13042];
  assign N14388 = N14387 | data_masked[13170];
  assign N14387 = N14386 | data_masked[13298];
  assign N14386 = N14385 | data_masked[13426];
  assign N14385 = N14384 | data_masked[13554];
  assign N14384 = N14383 | data_masked[13682];
  assign N14383 = N14382 | data_masked[13810];
  assign N14382 = N14381 | data_masked[13938];
  assign N14381 = N14380 | data_masked[14066];
  assign N14380 = N14379 | data_masked[14194];
  assign N14379 = N14378 | data_masked[14322];
  assign N14378 = N14377 | data_masked[14450];
  assign N14377 = N14376 | data_masked[14578];
  assign N14376 = N14375 | data_masked[14706];
  assign N14375 = N14374 | data_masked[14834];
  assign N14374 = N14373 | data_masked[14962];
  assign N14373 = N14372 | data_masked[15090];
  assign N14372 = N14371 | data_masked[15218];
  assign N14371 = N14370 | data_masked[15346];
  assign N14370 = N14369 | data_masked[15474];
  assign N14369 = N14368 | data_masked[15602];
  assign N14368 = N14367 | data_masked[15730];
  assign N14367 = N14366 | data_masked[15858];
  assign N14366 = N14365 | data_masked[15986];
  assign N14365 = N14364 | data_masked[16114];
  assign N14364 = data_masked[16370] | data_masked[16242];
  assign data_o[115] = N14615 | data_masked[115];
  assign N14615 = N14614 | data_masked[243];
  assign N14614 = N14613 | data_masked[371];
  assign N14613 = N14612 | data_masked[499];
  assign N14612 = N14611 | data_masked[627];
  assign N14611 = N14610 | data_masked[755];
  assign N14610 = N14609 | data_masked[883];
  assign N14609 = N14608 | data_masked[1011];
  assign N14608 = N14607 | data_masked[1139];
  assign N14607 = N14606 | data_masked[1267];
  assign N14606 = N14605 | data_masked[1395];
  assign N14605 = N14604 | data_masked[1523];
  assign N14604 = N14603 | data_masked[1651];
  assign N14603 = N14602 | data_masked[1779];
  assign N14602 = N14601 | data_masked[1907];
  assign N14601 = N14600 | data_masked[2035];
  assign N14600 = N14599 | data_masked[2163];
  assign N14599 = N14598 | data_masked[2291];
  assign N14598 = N14597 | data_masked[2419];
  assign N14597 = N14596 | data_masked[2547];
  assign N14596 = N14595 | data_masked[2675];
  assign N14595 = N14594 | data_masked[2803];
  assign N14594 = N14593 | data_masked[2931];
  assign N14593 = N14592 | data_masked[3059];
  assign N14592 = N14591 | data_masked[3187];
  assign N14591 = N14590 | data_masked[3315];
  assign N14590 = N14589 | data_masked[3443];
  assign N14589 = N14588 | data_masked[3571];
  assign N14588 = N14587 | data_masked[3699];
  assign N14587 = N14586 | data_masked[3827];
  assign N14586 = N14585 | data_masked[3955];
  assign N14585 = N14584 | data_masked[4083];
  assign N14584 = N14583 | data_masked[4211];
  assign N14583 = N14582 | data_masked[4339];
  assign N14582 = N14581 | data_masked[4467];
  assign N14581 = N14580 | data_masked[4595];
  assign N14580 = N14579 | data_masked[4723];
  assign N14579 = N14578 | data_masked[4851];
  assign N14578 = N14577 | data_masked[4979];
  assign N14577 = N14576 | data_masked[5107];
  assign N14576 = N14575 | data_masked[5235];
  assign N14575 = N14574 | data_masked[5363];
  assign N14574 = N14573 | data_masked[5491];
  assign N14573 = N14572 | data_masked[5619];
  assign N14572 = N14571 | data_masked[5747];
  assign N14571 = N14570 | data_masked[5875];
  assign N14570 = N14569 | data_masked[6003];
  assign N14569 = N14568 | data_masked[6131];
  assign N14568 = N14567 | data_masked[6259];
  assign N14567 = N14566 | data_masked[6387];
  assign N14566 = N14565 | data_masked[6515];
  assign N14565 = N14564 | data_masked[6643];
  assign N14564 = N14563 | data_masked[6771];
  assign N14563 = N14562 | data_masked[6899];
  assign N14562 = N14561 | data_masked[7027];
  assign N14561 = N14560 | data_masked[7155];
  assign N14560 = N14559 | data_masked[7283];
  assign N14559 = N14558 | data_masked[7411];
  assign N14558 = N14557 | data_masked[7539];
  assign N14557 = N14556 | data_masked[7667];
  assign N14556 = N14555 | data_masked[7795];
  assign N14555 = N14554 | data_masked[7923];
  assign N14554 = N14553 | data_masked[8051];
  assign N14553 = N14552 | data_masked[8179];
  assign N14552 = N14551 | data_masked[8307];
  assign N14551 = N14550 | data_masked[8435];
  assign N14550 = N14549 | data_masked[8563];
  assign N14549 = N14548 | data_masked[8691];
  assign N14548 = N14547 | data_masked[8819];
  assign N14547 = N14546 | data_masked[8947];
  assign N14546 = N14545 | data_masked[9075];
  assign N14545 = N14544 | data_masked[9203];
  assign N14544 = N14543 | data_masked[9331];
  assign N14543 = N14542 | data_masked[9459];
  assign N14542 = N14541 | data_masked[9587];
  assign N14541 = N14540 | data_masked[9715];
  assign N14540 = N14539 | data_masked[9843];
  assign N14539 = N14538 | data_masked[9971];
  assign N14538 = N14537 | data_masked[10099];
  assign N14537 = N14536 | data_masked[10227];
  assign N14536 = N14535 | data_masked[10355];
  assign N14535 = N14534 | data_masked[10483];
  assign N14534 = N14533 | data_masked[10611];
  assign N14533 = N14532 | data_masked[10739];
  assign N14532 = N14531 | data_masked[10867];
  assign N14531 = N14530 | data_masked[10995];
  assign N14530 = N14529 | data_masked[11123];
  assign N14529 = N14528 | data_masked[11251];
  assign N14528 = N14527 | data_masked[11379];
  assign N14527 = N14526 | data_masked[11507];
  assign N14526 = N14525 | data_masked[11635];
  assign N14525 = N14524 | data_masked[11763];
  assign N14524 = N14523 | data_masked[11891];
  assign N14523 = N14522 | data_masked[12019];
  assign N14522 = N14521 | data_masked[12147];
  assign N14521 = N14520 | data_masked[12275];
  assign N14520 = N14519 | data_masked[12403];
  assign N14519 = N14518 | data_masked[12531];
  assign N14518 = N14517 | data_masked[12659];
  assign N14517 = N14516 | data_masked[12787];
  assign N14516 = N14515 | data_masked[12915];
  assign N14515 = N14514 | data_masked[13043];
  assign N14514 = N14513 | data_masked[13171];
  assign N14513 = N14512 | data_masked[13299];
  assign N14512 = N14511 | data_masked[13427];
  assign N14511 = N14510 | data_masked[13555];
  assign N14510 = N14509 | data_masked[13683];
  assign N14509 = N14508 | data_masked[13811];
  assign N14508 = N14507 | data_masked[13939];
  assign N14507 = N14506 | data_masked[14067];
  assign N14506 = N14505 | data_masked[14195];
  assign N14505 = N14504 | data_masked[14323];
  assign N14504 = N14503 | data_masked[14451];
  assign N14503 = N14502 | data_masked[14579];
  assign N14502 = N14501 | data_masked[14707];
  assign N14501 = N14500 | data_masked[14835];
  assign N14500 = N14499 | data_masked[14963];
  assign N14499 = N14498 | data_masked[15091];
  assign N14498 = N14497 | data_masked[15219];
  assign N14497 = N14496 | data_masked[15347];
  assign N14496 = N14495 | data_masked[15475];
  assign N14495 = N14494 | data_masked[15603];
  assign N14494 = N14493 | data_masked[15731];
  assign N14493 = N14492 | data_masked[15859];
  assign N14492 = N14491 | data_masked[15987];
  assign N14491 = N14490 | data_masked[16115];
  assign N14490 = data_masked[16371] | data_masked[16243];
  assign data_o[116] = N14741 | data_masked[116];
  assign N14741 = N14740 | data_masked[244];
  assign N14740 = N14739 | data_masked[372];
  assign N14739 = N14738 | data_masked[500];
  assign N14738 = N14737 | data_masked[628];
  assign N14737 = N14736 | data_masked[756];
  assign N14736 = N14735 | data_masked[884];
  assign N14735 = N14734 | data_masked[1012];
  assign N14734 = N14733 | data_masked[1140];
  assign N14733 = N14732 | data_masked[1268];
  assign N14732 = N14731 | data_masked[1396];
  assign N14731 = N14730 | data_masked[1524];
  assign N14730 = N14729 | data_masked[1652];
  assign N14729 = N14728 | data_masked[1780];
  assign N14728 = N14727 | data_masked[1908];
  assign N14727 = N14726 | data_masked[2036];
  assign N14726 = N14725 | data_masked[2164];
  assign N14725 = N14724 | data_masked[2292];
  assign N14724 = N14723 | data_masked[2420];
  assign N14723 = N14722 | data_masked[2548];
  assign N14722 = N14721 | data_masked[2676];
  assign N14721 = N14720 | data_masked[2804];
  assign N14720 = N14719 | data_masked[2932];
  assign N14719 = N14718 | data_masked[3060];
  assign N14718 = N14717 | data_masked[3188];
  assign N14717 = N14716 | data_masked[3316];
  assign N14716 = N14715 | data_masked[3444];
  assign N14715 = N14714 | data_masked[3572];
  assign N14714 = N14713 | data_masked[3700];
  assign N14713 = N14712 | data_masked[3828];
  assign N14712 = N14711 | data_masked[3956];
  assign N14711 = N14710 | data_masked[4084];
  assign N14710 = N14709 | data_masked[4212];
  assign N14709 = N14708 | data_masked[4340];
  assign N14708 = N14707 | data_masked[4468];
  assign N14707 = N14706 | data_masked[4596];
  assign N14706 = N14705 | data_masked[4724];
  assign N14705 = N14704 | data_masked[4852];
  assign N14704 = N14703 | data_masked[4980];
  assign N14703 = N14702 | data_masked[5108];
  assign N14702 = N14701 | data_masked[5236];
  assign N14701 = N14700 | data_masked[5364];
  assign N14700 = N14699 | data_masked[5492];
  assign N14699 = N14698 | data_masked[5620];
  assign N14698 = N14697 | data_masked[5748];
  assign N14697 = N14696 | data_masked[5876];
  assign N14696 = N14695 | data_masked[6004];
  assign N14695 = N14694 | data_masked[6132];
  assign N14694 = N14693 | data_masked[6260];
  assign N14693 = N14692 | data_masked[6388];
  assign N14692 = N14691 | data_masked[6516];
  assign N14691 = N14690 | data_masked[6644];
  assign N14690 = N14689 | data_masked[6772];
  assign N14689 = N14688 | data_masked[6900];
  assign N14688 = N14687 | data_masked[7028];
  assign N14687 = N14686 | data_masked[7156];
  assign N14686 = N14685 | data_masked[7284];
  assign N14685 = N14684 | data_masked[7412];
  assign N14684 = N14683 | data_masked[7540];
  assign N14683 = N14682 | data_masked[7668];
  assign N14682 = N14681 | data_masked[7796];
  assign N14681 = N14680 | data_masked[7924];
  assign N14680 = N14679 | data_masked[8052];
  assign N14679 = N14678 | data_masked[8180];
  assign N14678 = N14677 | data_masked[8308];
  assign N14677 = N14676 | data_masked[8436];
  assign N14676 = N14675 | data_masked[8564];
  assign N14675 = N14674 | data_masked[8692];
  assign N14674 = N14673 | data_masked[8820];
  assign N14673 = N14672 | data_masked[8948];
  assign N14672 = N14671 | data_masked[9076];
  assign N14671 = N14670 | data_masked[9204];
  assign N14670 = N14669 | data_masked[9332];
  assign N14669 = N14668 | data_masked[9460];
  assign N14668 = N14667 | data_masked[9588];
  assign N14667 = N14666 | data_masked[9716];
  assign N14666 = N14665 | data_masked[9844];
  assign N14665 = N14664 | data_masked[9972];
  assign N14664 = N14663 | data_masked[10100];
  assign N14663 = N14662 | data_masked[10228];
  assign N14662 = N14661 | data_masked[10356];
  assign N14661 = N14660 | data_masked[10484];
  assign N14660 = N14659 | data_masked[10612];
  assign N14659 = N14658 | data_masked[10740];
  assign N14658 = N14657 | data_masked[10868];
  assign N14657 = N14656 | data_masked[10996];
  assign N14656 = N14655 | data_masked[11124];
  assign N14655 = N14654 | data_masked[11252];
  assign N14654 = N14653 | data_masked[11380];
  assign N14653 = N14652 | data_masked[11508];
  assign N14652 = N14651 | data_masked[11636];
  assign N14651 = N14650 | data_masked[11764];
  assign N14650 = N14649 | data_masked[11892];
  assign N14649 = N14648 | data_masked[12020];
  assign N14648 = N14647 | data_masked[12148];
  assign N14647 = N14646 | data_masked[12276];
  assign N14646 = N14645 | data_masked[12404];
  assign N14645 = N14644 | data_masked[12532];
  assign N14644 = N14643 | data_masked[12660];
  assign N14643 = N14642 | data_masked[12788];
  assign N14642 = N14641 | data_masked[12916];
  assign N14641 = N14640 | data_masked[13044];
  assign N14640 = N14639 | data_masked[13172];
  assign N14639 = N14638 | data_masked[13300];
  assign N14638 = N14637 | data_masked[13428];
  assign N14637 = N14636 | data_masked[13556];
  assign N14636 = N14635 | data_masked[13684];
  assign N14635 = N14634 | data_masked[13812];
  assign N14634 = N14633 | data_masked[13940];
  assign N14633 = N14632 | data_masked[14068];
  assign N14632 = N14631 | data_masked[14196];
  assign N14631 = N14630 | data_masked[14324];
  assign N14630 = N14629 | data_masked[14452];
  assign N14629 = N14628 | data_masked[14580];
  assign N14628 = N14627 | data_masked[14708];
  assign N14627 = N14626 | data_masked[14836];
  assign N14626 = N14625 | data_masked[14964];
  assign N14625 = N14624 | data_masked[15092];
  assign N14624 = N14623 | data_masked[15220];
  assign N14623 = N14622 | data_masked[15348];
  assign N14622 = N14621 | data_masked[15476];
  assign N14621 = N14620 | data_masked[15604];
  assign N14620 = N14619 | data_masked[15732];
  assign N14619 = N14618 | data_masked[15860];
  assign N14618 = N14617 | data_masked[15988];
  assign N14617 = N14616 | data_masked[16116];
  assign N14616 = data_masked[16372] | data_masked[16244];
  assign data_o[117] = N14867 | data_masked[117];
  assign N14867 = N14866 | data_masked[245];
  assign N14866 = N14865 | data_masked[373];
  assign N14865 = N14864 | data_masked[501];
  assign N14864 = N14863 | data_masked[629];
  assign N14863 = N14862 | data_masked[757];
  assign N14862 = N14861 | data_masked[885];
  assign N14861 = N14860 | data_masked[1013];
  assign N14860 = N14859 | data_masked[1141];
  assign N14859 = N14858 | data_masked[1269];
  assign N14858 = N14857 | data_masked[1397];
  assign N14857 = N14856 | data_masked[1525];
  assign N14856 = N14855 | data_masked[1653];
  assign N14855 = N14854 | data_masked[1781];
  assign N14854 = N14853 | data_masked[1909];
  assign N14853 = N14852 | data_masked[2037];
  assign N14852 = N14851 | data_masked[2165];
  assign N14851 = N14850 | data_masked[2293];
  assign N14850 = N14849 | data_masked[2421];
  assign N14849 = N14848 | data_masked[2549];
  assign N14848 = N14847 | data_masked[2677];
  assign N14847 = N14846 | data_masked[2805];
  assign N14846 = N14845 | data_masked[2933];
  assign N14845 = N14844 | data_masked[3061];
  assign N14844 = N14843 | data_masked[3189];
  assign N14843 = N14842 | data_masked[3317];
  assign N14842 = N14841 | data_masked[3445];
  assign N14841 = N14840 | data_masked[3573];
  assign N14840 = N14839 | data_masked[3701];
  assign N14839 = N14838 | data_masked[3829];
  assign N14838 = N14837 | data_masked[3957];
  assign N14837 = N14836 | data_masked[4085];
  assign N14836 = N14835 | data_masked[4213];
  assign N14835 = N14834 | data_masked[4341];
  assign N14834 = N14833 | data_masked[4469];
  assign N14833 = N14832 | data_masked[4597];
  assign N14832 = N14831 | data_masked[4725];
  assign N14831 = N14830 | data_masked[4853];
  assign N14830 = N14829 | data_masked[4981];
  assign N14829 = N14828 | data_masked[5109];
  assign N14828 = N14827 | data_masked[5237];
  assign N14827 = N14826 | data_masked[5365];
  assign N14826 = N14825 | data_masked[5493];
  assign N14825 = N14824 | data_masked[5621];
  assign N14824 = N14823 | data_masked[5749];
  assign N14823 = N14822 | data_masked[5877];
  assign N14822 = N14821 | data_masked[6005];
  assign N14821 = N14820 | data_masked[6133];
  assign N14820 = N14819 | data_masked[6261];
  assign N14819 = N14818 | data_masked[6389];
  assign N14818 = N14817 | data_masked[6517];
  assign N14817 = N14816 | data_masked[6645];
  assign N14816 = N14815 | data_masked[6773];
  assign N14815 = N14814 | data_masked[6901];
  assign N14814 = N14813 | data_masked[7029];
  assign N14813 = N14812 | data_masked[7157];
  assign N14812 = N14811 | data_masked[7285];
  assign N14811 = N14810 | data_masked[7413];
  assign N14810 = N14809 | data_masked[7541];
  assign N14809 = N14808 | data_masked[7669];
  assign N14808 = N14807 | data_masked[7797];
  assign N14807 = N14806 | data_masked[7925];
  assign N14806 = N14805 | data_masked[8053];
  assign N14805 = N14804 | data_masked[8181];
  assign N14804 = N14803 | data_masked[8309];
  assign N14803 = N14802 | data_masked[8437];
  assign N14802 = N14801 | data_masked[8565];
  assign N14801 = N14800 | data_masked[8693];
  assign N14800 = N14799 | data_masked[8821];
  assign N14799 = N14798 | data_masked[8949];
  assign N14798 = N14797 | data_masked[9077];
  assign N14797 = N14796 | data_masked[9205];
  assign N14796 = N14795 | data_masked[9333];
  assign N14795 = N14794 | data_masked[9461];
  assign N14794 = N14793 | data_masked[9589];
  assign N14793 = N14792 | data_masked[9717];
  assign N14792 = N14791 | data_masked[9845];
  assign N14791 = N14790 | data_masked[9973];
  assign N14790 = N14789 | data_masked[10101];
  assign N14789 = N14788 | data_masked[10229];
  assign N14788 = N14787 | data_masked[10357];
  assign N14787 = N14786 | data_masked[10485];
  assign N14786 = N14785 | data_masked[10613];
  assign N14785 = N14784 | data_masked[10741];
  assign N14784 = N14783 | data_masked[10869];
  assign N14783 = N14782 | data_masked[10997];
  assign N14782 = N14781 | data_masked[11125];
  assign N14781 = N14780 | data_masked[11253];
  assign N14780 = N14779 | data_masked[11381];
  assign N14779 = N14778 | data_masked[11509];
  assign N14778 = N14777 | data_masked[11637];
  assign N14777 = N14776 | data_masked[11765];
  assign N14776 = N14775 | data_masked[11893];
  assign N14775 = N14774 | data_masked[12021];
  assign N14774 = N14773 | data_masked[12149];
  assign N14773 = N14772 | data_masked[12277];
  assign N14772 = N14771 | data_masked[12405];
  assign N14771 = N14770 | data_masked[12533];
  assign N14770 = N14769 | data_masked[12661];
  assign N14769 = N14768 | data_masked[12789];
  assign N14768 = N14767 | data_masked[12917];
  assign N14767 = N14766 | data_masked[13045];
  assign N14766 = N14765 | data_masked[13173];
  assign N14765 = N14764 | data_masked[13301];
  assign N14764 = N14763 | data_masked[13429];
  assign N14763 = N14762 | data_masked[13557];
  assign N14762 = N14761 | data_masked[13685];
  assign N14761 = N14760 | data_masked[13813];
  assign N14760 = N14759 | data_masked[13941];
  assign N14759 = N14758 | data_masked[14069];
  assign N14758 = N14757 | data_masked[14197];
  assign N14757 = N14756 | data_masked[14325];
  assign N14756 = N14755 | data_masked[14453];
  assign N14755 = N14754 | data_masked[14581];
  assign N14754 = N14753 | data_masked[14709];
  assign N14753 = N14752 | data_masked[14837];
  assign N14752 = N14751 | data_masked[14965];
  assign N14751 = N14750 | data_masked[15093];
  assign N14750 = N14749 | data_masked[15221];
  assign N14749 = N14748 | data_masked[15349];
  assign N14748 = N14747 | data_masked[15477];
  assign N14747 = N14746 | data_masked[15605];
  assign N14746 = N14745 | data_masked[15733];
  assign N14745 = N14744 | data_masked[15861];
  assign N14744 = N14743 | data_masked[15989];
  assign N14743 = N14742 | data_masked[16117];
  assign N14742 = data_masked[16373] | data_masked[16245];
  assign data_o[118] = N14993 | data_masked[118];
  assign N14993 = N14992 | data_masked[246];
  assign N14992 = N14991 | data_masked[374];
  assign N14991 = N14990 | data_masked[502];
  assign N14990 = N14989 | data_masked[630];
  assign N14989 = N14988 | data_masked[758];
  assign N14988 = N14987 | data_masked[886];
  assign N14987 = N14986 | data_masked[1014];
  assign N14986 = N14985 | data_masked[1142];
  assign N14985 = N14984 | data_masked[1270];
  assign N14984 = N14983 | data_masked[1398];
  assign N14983 = N14982 | data_masked[1526];
  assign N14982 = N14981 | data_masked[1654];
  assign N14981 = N14980 | data_masked[1782];
  assign N14980 = N14979 | data_masked[1910];
  assign N14979 = N14978 | data_masked[2038];
  assign N14978 = N14977 | data_masked[2166];
  assign N14977 = N14976 | data_masked[2294];
  assign N14976 = N14975 | data_masked[2422];
  assign N14975 = N14974 | data_masked[2550];
  assign N14974 = N14973 | data_masked[2678];
  assign N14973 = N14972 | data_masked[2806];
  assign N14972 = N14971 | data_masked[2934];
  assign N14971 = N14970 | data_masked[3062];
  assign N14970 = N14969 | data_masked[3190];
  assign N14969 = N14968 | data_masked[3318];
  assign N14968 = N14967 | data_masked[3446];
  assign N14967 = N14966 | data_masked[3574];
  assign N14966 = N14965 | data_masked[3702];
  assign N14965 = N14964 | data_masked[3830];
  assign N14964 = N14963 | data_masked[3958];
  assign N14963 = N14962 | data_masked[4086];
  assign N14962 = N14961 | data_masked[4214];
  assign N14961 = N14960 | data_masked[4342];
  assign N14960 = N14959 | data_masked[4470];
  assign N14959 = N14958 | data_masked[4598];
  assign N14958 = N14957 | data_masked[4726];
  assign N14957 = N14956 | data_masked[4854];
  assign N14956 = N14955 | data_masked[4982];
  assign N14955 = N14954 | data_masked[5110];
  assign N14954 = N14953 | data_masked[5238];
  assign N14953 = N14952 | data_masked[5366];
  assign N14952 = N14951 | data_masked[5494];
  assign N14951 = N14950 | data_masked[5622];
  assign N14950 = N14949 | data_masked[5750];
  assign N14949 = N14948 | data_masked[5878];
  assign N14948 = N14947 | data_masked[6006];
  assign N14947 = N14946 | data_masked[6134];
  assign N14946 = N14945 | data_masked[6262];
  assign N14945 = N14944 | data_masked[6390];
  assign N14944 = N14943 | data_masked[6518];
  assign N14943 = N14942 | data_masked[6646];
  assign N14942 = N14941 | data_masked[6774];
  assign N14941 = N14940 | data_masked[6902];
  assign N14940 = N14939 | data_masked[7030];
  assign N14939 = N14938 | data_masked[7158];
  assign N14938 = N14937 | data_masked[7286];
  assign N14937 = N14936 | data_masked[7414];
  assign N14936 = N14935 | data_masked[7542];
  assign N14935 = N14934 | data_masked[7670];
  assign N14934 = N14933 | data_masked[7798];
  assign N14933 = N14932 | data_masked[7926];
  assign N14932 = N14931 | data_masked[8054];
  assign N14931 = N14930 | data_masked[8182];
  assign N14930 = N14929 | data_masked[8310];
  assign N14929 = N14928 | data_masked[8438];
  assign N14928 = N14927 | data_masked[8566];
  assign N14927 = N14926 | data_masked[8694];
  assign N14926 = N14925 | data_masked[8822];
  assign N14925 = N14924 | data_masked[8950];
  assign N14924 = N14923 | data_masked[9078];
  assign N14923 = N14922 | data_masked[9206];
  assign N14922 = N14921 | data_masked[9334];
  assign N14921 = N14920 | data_masked[9462];
  assign N14920 = N14919 | data_masked[9590];
  assign N14919 = N14918 | data_masked[9718];
  assign N14918 = N14917 | data_masked[9846];
  assign N14917 = N14916 | data_masked[9974];
  assign N14916 = N14915 | data_masked[10102];
  assign N14915 = N14914 | data_masked[10230];
  assign N14914 = N14913 | data_masked[10358];
  assign N14913 = N14912 | data_masked[10486];
  assign N14912 = N14911 | data_masked[10614];
  assign N14911 = N14910 | data_masked[10742];
  assign N14910 = N14909 | data_masked[10870];
  assign N14909 = N14908 | data_masked[10998];
  assign N14908 = N14907 | data_masked[11126];
  assign N14907 = N14906 | data_masked[11254];
  assign N14906 = N14905 | data_masked[11382];
  assign N14905 = N14904 | data_masked[11510];
  assign N14904 = N14903 | data_masked[11638];
  assign N14903 = N14902 | data_masked[11766];
  assign N14902 = N14901 | data_masked[11894];
  assign N14901 = N14900 | data_masked[12022];
  assign N14900 = N14899 | data_masked[12150];
  assign N14899 = N14898 | data_masked[12278];
  assign N14898 = N14897 | data_masked[12406];
  assign N14897 = N14896 | data_masked[12534];
  assign N14896 = N14895 | data_masked[12662];
  assign N14895 = N14894 | data_masked[12790];
  assign N14894 = N14893 | data_masked[12918];
  assign N14893 = N14892 | data_masked[13046];
  assign N14892 = N14891 | data_masked[13174];
  assign N14891 = N14890 | data_masked[13302];
  assign N14890 = N14889 | data_masked[13430];
  assign N14889 = N14888 | data_masked[13558];
  assign N14888 = N14887 | data_masked[13686];
  assign N14887 = N14886 | data_masked[13814];
  assign N14886 = N14885 | data_masked[13942];
  assign N14885 = N14884 | data_masked[14070];
  assign N14884 = N14883 | data_masked[14198];
  assign N14883 = N14882 | data_masked[14326];
  assign N14882 = N14881 | data_masked[14454];
  assign N14881 = N14880 | data_masked[14582];
  assign N14880 = N14879 | data_masked[14710];
  assign N14879 = N14878 | data_masked[14838];
  assign N14878 = N14877 | data_masked[14966];
  assign N14877 = N14876 | data_masked[15094];
  assign N14876 = N14875 | data_masked[15222];
  assign N14875 = N14874 | data_masked[15350];
  assign N14874 = N14873 | data_masked[15478];
  assign N14873 = N14872 | data_masked[15606];
  assign N14872 = N14871 | data_masked[15734];
  assign N14871 = N14870 | data_masked[15862];
  assign N14870 = N14869 | data_masked[15990];
  assign N14869 = N14868 | data_masked[16118];
  assign N14868 = data_masked[16374] | data_masked[16246];
  assign data_o[119] = N15119 | data_masked[119];
  assign N15119 = N15118 | data_masked[247];
  assign N15118 = N15117 | data_masked[375];
  assign N15117 = N15116 | data_masked[503];
  assign N15116 = N15115 | data_masked[631];
  assign N15115 = N15114 | data_masked[759];
  assign N15114 = N15113 | data_masked[887];
  assign N15113 = N15112 | data_masked[1015];
  assign N15112 = N15111 | data_masked[1143];
  assign N15111 = N15110 | data_masked[1271];
  assign N15110 = N15109 | data_masked[1399];
  assign N15109 = N15108 | data_masked[1527];
  assign N15108 = N15107 | data_masked[1655];
  assign N15107 = N15106 | data_masked[1783];
  assign N15106 = N15105 | data_masked[1911];
  assign N15105 = N15104 | data_masked[2039];
  assign N15104 = N15103 | data_masked[2167];
  assign N15103 = N15102 | data_masked[2295];
  assign N15102 = N15101 | data_masked[2423];
  assign N15101 = N15100 | data_masked[2551];
  assign N15100 = N15099 | data_masked[2679];
  assign N15099 = N15098 | data_masked[2807];
  assign N15098 = N15097 | data_masked[2935];
  assign N15097 = N15096 | data_masked[3063];
  assign N15096 = N15095 | data_masked[3191];
  assign N15095 = N15094 | data_masked[3319];
  assign N15094 = N15093 | data_masked[3447];
  assign N15093 = N15092 | data_masked[3575];
  assign N15092 = N15091 | data_masked[3703];
  assign N15091 = N15090 | data_masked[3831];
  assign N15090 = N15089 | data_masked[3959];
  assign N15089 = N15088 | data_masked[4087];
  assign N15088 = N15087 | data_masked[4215];
  assign N15087 = N15086 | data_masked[4343];
  assign N15086 = N15085 | data_masked[4471];
  assign N15085 = N15084 | data_masked[4599];
  assign N15084 = N15083 | data_masked[4727];
  assign N15083 = N15082 | data_masked[4855];
  assign N15082 = N15081 | data_masked[4983];
  assign N15081 = N15080 | data_masked[5111];
  assign N15080 = N15079 | data_masked[5239];
  assign N15079 = N15078 | data_masked[5367];
  assign N15078 = N15077 | data_masked[5495];
  assign N15077 = N15076 | data_masked[5623];
  assign N15076 = N15075 | data_masked[5751];
  assign N15075 = N15074 | data_masked[5879];
  assign N15074 = N15073 | data_masked[6007];
  assign N15073 = N15072 | data_masked[6135];
  assign N15072 = N15071 | data_masked[6263];
  assign N15071 = N15070 | data_masked[6391];
  assign N15070 = N15069 | data_masked[6519];
  assign N15069 = N15068 | data_masked[6647];
  assign N15068 = N15067 | data_masked[6775];
  assign N15067 = N15066 | data_masked[6903];
  assign N15066 = N15065 | data_masked[7031];
  assign N15065 = N15064 | data_masked[7159];
  assign N15064 = N15063 | data_masked[7287];
  assign N15063 = N15062 | data_masked[7415];
  assign N15062 = N15061 | data_masked[7543];
  assign N15061 = N15060 | data_masked[7671];
  assign N15060 = N15059 | data_masked[7799];
  assign N15059 = N15058 | data_masked[7927];
  assign N15058 = N15057 | data_masked[8055];
  assign N15057 = N15056 | data_masked[8183];
  assign N15056 = N15055 | data_masked[8311];
  assign N15055 = N15054 | data_masked[8439];
  assign N15054 = N15053 | data_masked[8567];
  assign N15053 = N15052 | data_masked[8695];
  assign N15052 = N15051 | data_masked[8823];
  assign N15051 = N15050 | data_masked[8951];
  assign N15050 = N15049 | data_masked[9079];
  assign N15049 = N15048 | data_masked[9207];
  assign N15048 = N15047 | data_masked[9335];
  assign N15047 = N15046 | data_masked[9463];
  assign N15046 = N15045 | data_masked[9591];
  assign N15045 = N15044 | data_masked[9719];
  assign N15044 = N15043 | data_masked[9847];
  assign N15043 = N15042 | data_masked[9975];
  assign N15042 = N15041 | data_masked[10103];
  assign N15041 = N15040 | data_masked[10231];
  assign N15040 = N15039 | data_masked[10359];
  assign N15039 = N15038 | data_masked[10487];
  assign N15038 = N15037 | data_masked[10615];
  assign N15037 = N15036 | data_masked[10743];
  assign N15036 = N15035 | data_masked[10871];
  assign N15035 = N15034 | data_masked[10999];
  assign N15034 = N15033 | data_masked[11127];
  assign N15033 = N15032 | data_masked[11255];
  assign N15032 = N15031 | data_masked[11383];
  assign N15031 = N15030 | data_masked[11511];
  assign N15030 = N15029 | data_masked[11639];
  assign N15029 = N15028 | data_masked[11767];
  assign N15028 = N15027 | data_masked[11895];
  assign N15027 = N15026 | data_masked[12023];
  assign N15026 = N15025 | data_masked[12151];
  assign N15025 = N15024 | data_masked[12279];
  assign N15024 = N15023 | data_masked[12407];
  assign N15023 = N15022 | data_masked[12535];
  assign N15022 = N15021 | data_masked[12663];
  assign N15021 = N15020 | data_masked[12791];
  assign N15020 = N15019 | data_masked[12919];
  assign N15019 = N15018 | data_masked[13047];
  assign N15018 = N15017 | data_masked[13175];
  assign N15017 = N15016 | data_masked[13303];
  assign N15016 = N15015 | data_masked[13431];
  assign N15015 = N15014 | data_masked[13559];
  assign N15014 = N15013 | data_masked[13687];
  assign N15013 = N15012 | data_masked[13815];
  assign N15012 = N15011 | data_masked[13943];
  assign N15011 = N15010 | data_masked[14071];
  assign N15010 = N15009 | data_masked[14199];
  assign N15009 = N15008 | data_masked[14327];
  assign N15008 = N15007 | data_masked[14455];
  assign N15007 = N15006 | data_masked[14583];
  assign N15006 = N15005 | data_masked[14711];
  assign N15005 = N15004 | data_masked[14839];
  assign N15004 = N15003 | data_masked[14967];
  assign N15003 = N15002 | data_masked[15095];
  assign N15002 = N15001 | data_masked[15223];
  assign N15001 = N15000 | data_masked[15351];
  assign N15000 = N14999 | data_masked[15479];
  assign N14999 = N14998 | data_masked[15607];
  assign N14998 = N14997 | data_masked[15735];
  assign N14997 = N14996 | data_masked[15863];
  assign N14996 = N14995 | data_masked[15991];
  assign N14995 = N14994 | data_masked[16119];
  assign N14994 = data_masked[16375] | data_masked[16247];
  assign data_o[120] = N15245 | data_masked[120];
  assign N15245 = N15244 | data_masked[248];
  assign N15244 = N15243 | data_masked[376];
  assign N15243 = N15242 | data_masked[504];
  assign N15242 = N15241 | data_masked[632];
  assign N15241 = N15240 | data_masked[760];
  assign N15240 = N15239 | data_masked[888];
  assign N15239 = N15238 | data_masked[1016];
  assign N15238 = N15237 | data_masked[1144];
  assign N15237 = N15236 | data_masked[1272];
  assign N15236 = N15235 | data_masked[1400];
  assign N15235 = N15234 | data_masked[1528];
  assign N15234 = N15233 | data_masked[1656];
  assign N15233 = N15232 | data_masked[1784];
  assign N15232 = N15231 | data_masked[1912];
  assign N15231 = N15230 | data_masked[2040];
  assign N15230 = N15229 | data_masked[2168];
  assign N15229 = N15228 | data_masked[2296];
  assign N15228 = N15227 | data_masked[2424];
  assign N15227 = N15226 | data_masked[2552];
  assign N15226 = N15225 | data_masked[2680];
  assign N15225 = N15224 | data_masked[2808];
  assign N15224 = N15223 | data_masked[2936];
  assign N15223 = N15222 | data_masked[3064];
  assign N15222 = N15221 | data_masked[3192];
  assign N15221 = N15220 | data_masked[3320];
  assign N15220 = N15219 | data_masked[3448];
  assign N15219 = N15218 | data_masked[3576];
  assign N15218 = N15217 | data_masked[3704];
  assign N15217 = N15216 | data_masked[3832];
  assign N15216 = N15215 | data_masked[3960];
  assign N15215 = N15214 | data_masked[4088];
  assign N15214 = N15213 | data_masked[4216];
  assign N15213 = N15212 | data_masked[4344];
  assign N15212 = N15211 | data_masked[4472];
  assign N15211 = N15210 | data_masked[4600];
  assign N15210 = N15209 | data_masked[4728];
  assign N15209 = N15208 | data_masked[4856];
  assign N15208 = N15207 | data_masked[4984];
  assign N15207 = N15206 | data_masked[5112];
  assign N15206 = N15205 | data_masked[5240];
  assign N15205 = N15204 | data_masked[5368];
  assign N15204 = N15203 | data_masked[5496];
  assign N15203 = N15202 | data_masked[5624];
  assign N15202 = N15201 | data_masked[5752];
  assign N15201 = N15200 | data_masked[5880];
  assign N15200 = N15199 | data_masked[6008];
  assign N15199 = N15198 | data_masked[6136];
  assign N15198 = N15197 | data_masked[6264];
  assign N15197 = N15196 | data_masked[6392];
  assign N15196 = N15195 | data_masked[6520];
  assign N15195 = N15194 | data_masked[6648];
  assign N15194 = N15193 | data_masked[6776];
  assign N15193 = N15192 | data_masked[6904];
  assign N15192 = N15191 | data_masked[7032];
  assign N15191 = N15190 | data_masked[7160];
  assign N15190 = N15189 | data_masked[7288];
  assign N15189 = N15188 | data_masked[7416];
  assign N15188 = N15187 | data_masked[7544];
  assign N15187 = N15186 | data_masked[7672];
  assign N15186 = N15185 | data_masked[7800];
  assign N15185 = N15184 | data_masked[7928];
  assign N15184 = N15183 | data_masked[8056];
  assign N15183 = N15182 | data_masked[8184];
  assign N15182 = N15181 | data_masked[8312];
  assign N15181 = N15180 | data_masked[8440];
  assign N15180 = N15179 | data_masked[8568];
  assign N15179 = N15178 | data_masked[8696];
  assign N15178 = N15177 | data_masked[8824];
  assign N15177 = N15176 | data_masked[8952];
  assign N15176 = N15175 | data_masked[9080];
  assign N15175 = N15174 | data_masked[9208];
  assign N15174 = N15173 | data_masked[9336];
  assign N15173 = N15172 | data_masked[9464];
  assign N15172 = N15171 | data_masked[9592];
  assign N15171 = N15170 | data_masked[9720];
  assign N15170 = N15169 | data_masked[9848];
  assign N15169 = N15168 | data_masked[9976];
  assign N15168 = N15167 | data_masked[10104];
  assign N15167 = N15166 | data_masked[10232];
  assign N15166 = N15165 | data_masked[10360];
  assign N15165 = N15164 | data_masked[10488];
  assign N15164 = N15163 | data_masked[10616];
  assign N15163 = N15162 | data_masked[10744];
  assign N15162 = N15161 | data_masked[10872];
  assign N15161 = N15160 | data_masked[11000];
  assign N15160 = N15159 | data_masked[11128];
  assign N15159 = N15158 | data_masked[11256];
  assign N15158 = N15157 | data_masked[11384];
  assign N15157 = N15156 | data_masked[11512];
  assign N15156 = N15155 | data_masked[11640];
  assign N15155 = N15154 | data_masked[11768];
  assign N15154 = N15153 | data_masked[11896];
  assign N15153 = N15152 | data_masked[12024];
  assign N15152 = N15151 | data_masked[12152];
  assign N15151 = N15150 | data_masked[12280];
  assign N15150 = N15149 | data_masked[12408];
  assign N15149 = N15148 | data_masked[12536];
  assign N15148 = N15147 | data_masked[12664];
  assign N15147 = N15146 | data_masked[12792];
  assign N15146 = N15145 | data_masked[12920];
  assign N15145 = N15144 | data_masked[13048];
  assign N15144 = N15143 | data_masked[13176];
  assign N15143 = N15142 | data_masked[13304];
  assign N15142 = N15141 | data_masked[13432];
  assign N15141 = N15140 | data_masked[13560];
  assign N15140 = N15139 | data_masked[13688];
  assign N15139 = N15138 | data_masked[13816];
  assign N15138 = N15137 | data_masked[13944];
  assign N15137 = N15136 | data_masked[14072];
  assign N15136 = N15135 | data_masked[14200];
  assign N15135 = N15134 | data_masked[14328];
  assign N15134 = N15133 | data_masked[14456];
  assign N15133 = N15132 | data_masked[14584];
  assign N15132 = N15131 | data_masked[14712];
  assign N15131 = N15130 | data_masked[14840];
  assign N15130 = N15129 | data_masked[14968];
  assign N15129 = N15128 | data_masked[15096];
  assign N15128 = N15127 | data_masked[15224];
  assign N15127 = N15126 | data_masked[15352];
  assign N15126 = N15125 | data_masked[15480];
  assign N15125 = N15124 | data_masked[15608];
  assign N15124 = N15123 | data_masked[15736];
  assign N15123 = N15122 | data_masked[15864];
  assign N15122 = N15121 | data_masked[15992];
  assign N15121 = N15120 | data_masked[16120];
  assign N15120 = data_masked[16376] | data_masked[16248];
  assign data_o[121] = N15371 | data_masked[121];
  assign N15371 = N15370 | data_masked[249];
  assign N15370 = N15369 | data_masked[377];
  assign N15369 = N15368 | data_masked[505];
  assign N15368 = N15367 | data_masked[633];
  assign N15367 = N15366 | data_masked[761];
  assign N15366 = N15365 | data_masked[889];
  assign N15365 = N15364 | data_masked[1017];
  assign N15364 = N15363 | data_masked[1145];
  assign N15363 = N15362 | data_masked[1273];
  assign N15362 = N15361 | data_masked[1401];
  assign N15361 = N15360 | data_masked[1529];
  assign N15360 = N15359 | data_masked[1657];
  assign N15359 = N15358 | data_masked[1785];
  assign N15358 = N15357 | data_masked[1913];
  assign N15357 = N15356 | data_masked[2041];
  assign N15356 = N15355 | data_masked[2169];
  assign N15355 = N15354 | data_masked[2297];
  assign N15354 = N15353 | data_masked[2425];
  assign N15353 = N15352 | data_masked[2553];
  assign N15352 = N15351 | data_masked[2681];
  assign N15351 = N15350 | data_masked[2809];
  assign N15350 = N15349 | data_masked[2937];
  assign N15349 = N15348 | data_masked[3065];
  assign N15348 = N15347 | data_masked[3193];
  assign N15347 = N15346 | data_masked[3321];
  assign N15346 = N15345 | data_masked[3449];
  assign N15345 = N15344 | data_masked[3577];
  assign N15344 = N15343 | data_masked[3705];
  assign N15343 = N15342 | data_masked[3833];
  assign N15342 = N15341 | data_masked[3961];
  assign N15341 = N15340 | data_masked[4089];
  assign N15340 = N15339 | data_masked[4217];
  assign N15339 = N15338 | data_masked[4345];
  assign N15338 = N15337 | data_masked[4473];
  assign N15337 = N15336 | data_masked[4601];
  assign N15336 = N15335 | data_masked[4729];
  assign N15335 = N15334 | data_masked[4857];
  assign N15334 = N15333 | data_masked[4985];
  assign N15333 = N15332 | data_masked[5113];
  assign N15332 = N15331 | data_masked[5241];
  assign N15331 = N15330 | data_masked[5369];
  assign N15330 = N15329 | data_masked[5497];
  assign N15329 = N15328 | data_masked[5625];
  assign N15328 = N15327 | data_masked[5753];
  assign N15327 = N15326 | data_masked[5881];
  assign N15326 = N15325 | data_masked[6009];
  assign N15325 = N15324 | data_masked[6137];
  assign N15324 = N15323 | data_masked[6265];
  assign N15323 = N15322 | data_masked[6393];
  assign N15322 = N15321 | data_masked[6521];
  assign N15321 = N15320 | data_masked[6649];
  assign N15320 = N15319 | data_masked[6777];
  assign N15319 = N15318 | data_masked[6905];
  assign N15318 = N15317 | data_masked[7033];
  assign N15317 = N15316 | data_masked[7161];
  assign N15316 = N15315 | data_masked[7289];
  assign N15315 = N15314 | data_masked[7417];
  assign N15314 = N15313 | data_masked[7545];
  assign N15313 = N15312 | data_masked[7673];
  assign N15312 = N15311 | data_masked[7801];
  assign N15311 = N15310 | data_masked[7929];
  assign N15310 = N15309 | data_masked[8057];
  assign N15309 = N15308 | data_masked[8185];
  assign N15308 = N15307 | data_masked[8313];
  assign N15307 = N15306 | data_masked[8441];
  assign N15306 = N15305 | data_masked[8569];
  assign N15305 = N15304 | data_masked[8697];
  assign N15304 = N15303 | data_masked[8825];
  assign N15303 = N15302 | data_masked[8953];
  assign N15302 = N15301 | data_masked[9081];
  assign N15301 = N15300 | data_masked[9209];
  assign N15300 = N15299 | data_masked[9337];
  assign N15299 = N15298 | data_masked[9465];
  assign N15298 = N15297 | data_masked[9593];
  assign N15297 = N15296 | data_masked[9721];
  assign N15296 = N15295 | data_masked[9849];
  assign N15295 = N15294 | data_masked[9977];
  assign N15294 = N15293 | data_masked[10105];
  assign N15293 = N15292 | data_masked[10233];
  assign N15292 = N15291 | data_masked[10361];
  assign N15291 = N15290 | data_masked[10489];
  assign N15290 = N15289 | data_masked[10617];
  assign N15289 = N15288 | data_masked[10745];
  assign N15288 = N15287 | data_masked[10873];
  assign N15287 = N15286 | data_masked[11001];
  assign N15286 = N15285 | data_masked[11129];
  assign N15285 = N15284 | data_masked[11257];
  assign N15284 = N15283 | data_masked[11385];
  assign N15283 = N15282 | data_masked[11513];
  assign N15282 = N15281 | data_masked[11641];
  assign N15281 = N15280 | data_masked[11769];
  assign N15280 = N15279 | data_masked[11897];
  assign N15279 = N15278 | data_masked[12025];
  assign N15278 = N15277 | data_masked[12153];
  assign N15277 = N15276 | data_masked[12281];
  assign N15276 = N15275 | data_masked[12409];
  assign N15275 = N15274 | data_masked[12537];
  assign N15274 = N15273 | data_masked[12665];
  assign N15273 = N15272 | data_masked[12793];
  assign N15272 = N15271 | data_masked[12921];
  assign N15271 = N15270 | data_masked[13049];
  assign N15270 = N15269 | data_masked[13177];
  assign N15269 = N15268 | data_masked[13305];
  assign N15268 = N15267 | data_masked[13433];
  assign N15267 = N15266 | data_masked[13561];
  assign N15266 = N15265 | data_masked[13689];
  assign N15265 = N15264 | data_masked[13817];
  assign N15264 = N15263 | data_masked[13945];
  assign N15263 = N15262 | data_masked[14073];
  assign N15262 = N15261 | data_masked[14201];
  assign N15261 = N15260 | data_masked[14329];
  assign N15260 = N15259 | data_masked[14457];
  assign N15259 = N15258 | data_masked[14585];
  assign N15258 = N15257 | data_masked[14713];
  assign N15257 = N15256 | data_masked[14841];
  assign N15256 = N15255 | data_masked[14969];
  assign N15255 = N15254 | data_masked[15097];
  assign N15254 = N15253 | data_masked[15225];
  assign N15253 = N15252 | data_masked[15353];
  assign N15252 = N15251 | data_masked[15481];
  assign N15251 = N15250 | data_masked[15609];
  assign N15250 = N15249 | data_masked[15737];
  assign N15249 = N15248 | data_masked[15865];
  assign N15248 = N15247 | data_masked[15993];
  assign N15247 = N15246 | data_masked[16121];
  assign N15246 = data_masked[16377] | data_masked[16249];
  assign data_o[122] = N15497 | data_masked[122];
  assign N15497 = N15496 | data_masked[250];
  assign N15496 = N15495 | data_masked[378];
  assign N15495 = N15494 | data_masked[506];
  assign N15494 = N15493 | data_masked[634];
  assign N15493 = N15492 | data_masked[762];
  assign N15492 = N15491 | data_masked[890];
  assign N15491 = N15490 | data_masked[1018];
  assign N15490 = N15489 | data_masked[1146];
  assign N15489 = N15488 | data_masked[1274];
  assign N15488 = N15487 | data_masked[1402];
  assign N15487 = N15486 | data_masked[1530];
  assign N15486 = N15485 | data_masked[1658];
  assign N15485 = N15484 | data_masked[1786];
  assign N15484 = N15483 | data_masked[1914];
  assign N15483 = N15482 | data_masked[2042];
  assign N15482 = N15481 | data_masked[2170];
  assign N15481 = N15480 | data_masked[2298];
  assign N15480 = N15479 | data_masked[2426];
  assign N15479 = N15478 | data_masked[2554];
  assign N15478 = N15477 | data_masked[2682];
  assign N15477 = N15476 | data_masked[2810];
  assign N15476 = N15475 | data_masked[2938];
  assign N15475 = N15474 | data_masked[3066];
  assign N15474 = N15473 | data_masked[3194];
  assign N15473 = N15472 | data_masked[3322];
  assign N15472 = N15471 | data_masked[3450];
  assign N15471 = N15470 | data_masked[3578];
  assign N15470 = N15469 | data_masked[3706];
  assign N15469 = N15468 | data_masked[3834];
  assign N15468 = N15467 | data_masked[3962];
  assign N15467 = N15466 | data_masked[4090];
  assign N15466 = N15465 | data_masked[4218];
  assign N15465 = N15464 | data_masked[4346];
  assign N15464 = N15463 | data_masked[4474];
  assign N15463 = N15462 | data_masked[4602];
  assign N15462 = N15461 | data_masked[4730];
  assign N15461 = N15460 | data_masked[4858];
  assign N15460 = N15459 | data_masked[4986];
  assign N15459 = N15458 | data_masked[5114];
  assign N15458 = N15457 | data_masked[5242];
  assign N15457 = N15456 | data_masked[5370];
  assign N15456 = N15455 | data_masked[5498];
  assign N15455 = N15454 | data_masked[5626];
  assign N15454 = N15453 | data_masked[5754];
  assign N15453 = N15452 | data_masked[5882];
  assign N15452 = N15451 | data_masked[6010];
  assign N15451 = N15450 | data_masked[6138];
  assign N15450 = N15449 | data_masked[6266];
  assign N15449 = N15448 | data_masked[6394];
  assign N15448 = N15447 | data_masked[6522];
  assign N15447 = N15446 | data_masked[6650];
  assign N15446 = N15445 | data_masked[6778];
  assign N15445 = N15444 | data_masked[6906];
  assign N15444 = N15443 | data_masked[7034];
  assign N15443 = N15442 | data_masked[7162];
  assign N15442 = N15441 | data_masked[7290];
  assign N15441 = N15440 | data_masked[7418];
  assign N15440 = N15439 | data_masked[7546];
  assign N15439 = N15438 | data_masked[7674];
  assign N15438 = N15437 | data_masked[7802];
  assign N15437 = N15436 | data_masked[7930];
  assign N15436 = N15435 | data_masked[8058];
  assign N15435 = N15434 | data_masked[8186];
  assign N15434 = N15433 | data_masked[8314];
  assign N15433 = N15432 | data_masked[8442];
  assign N15432 = N15431 | data_masked[8570];
  assign N15431 = N15430 | data_masked[8698];
  assign N15430 = N15429 | data_masked[8826];
  assign N15429 = N15428 | data_masked[8954];
  assign N15428 = N15427 | data_masked[9082];
  assign N15427 = N15426 | data_masked[9210];
  assign N15426 = N15425 | data_masked[9338];
  assign N15425 = N15424 | data_masked[9466];
  assign N15424 = N15423 | data_masked[9594];
  assign N15423 = N15422 | data_masked[9722];
  assign N15422 = N15421 | data_masked[9850];
  assign N15421 = N15420 | data_masked[9978];
  assign N15420 = N15419 | data_masked[10106];
  assign N15419 = N15418 | data_masked[10234];
  assign N15418 = N15417 | data_masked[10362];
  assign N15417 = N15416 | data_masked[10490];
  assign N15416 = N15415 | data_masked[10618];
  assign N15415 = N15414 | data_masked[10746];
  assign N15414 = N15413 | data_masked[10874];
  assign N15413 = N15412 | data_masked[11002];
  assign N15412 = N15411 | data_masked[11130];
  assign N15411 = N15410 | data_masked[11258];
  assign N15410 = N15409 | data_masked[11386];
  assign N15409 = N15408 | data_masked[11514];
  assign N15408 = N15407 | data_masked[11642];
  assign N15407 = N15406 | data_masked[11770];
  assign N15406 = N15405 | data_masked[11898];
  assign N15405 = N15404 | data_masked[12026];
  assign N15404 = N15403 | data_masked[12154];
  assign N15403 = N15402 | data_masked[12282];
  assign N15402 = N15401 | data_masked[12410];
  assign N15401 = N15400 | data_masked[12538];
  assign N15400 = N15399 | data_masked[12666];
  assign N15399 = N15398 | data_masked[12794];
  assign N15398 = N15397 | data_masked[12922];
  assign N15397 = N15396 | data_masked[13050];
  assign N15396 = N15395 | data_masked[13178];
  assign N15395 = N15394 | data_masked[13306];
  assign N15394 = N15393 | data_masked[13434];
  assign N15393 = N15392 | data_masked[13562];
  assign N15392 = N15391 | data_masked[13690];
  assign N15391 = N15390 | data_masked[13818];
  assign N15390 = N15389 | data_masked[13946];
  assign N15389 = N15388 | data_masked[14074];
  assign N15388 = N15387 | data_masked[14202];
  assign N15387 = N15386 | data_masked[14330];
  assign N15386 = N15385 | data_masked[14458];
  assign N15385 = N15384 | data_masked[14586];
  assign N15384 = N15383 | data_masked[14714];
  assign N15383 = N15382 | data_masked[14842];
  assign N15382 = N15381 | data_masked[14970];
  assign N15381 = N15380 | data_masked[15098];
  assign N15380 = N15379 | data_masked[15226];
  assign N15379 = N15378 | data_masked[15354];
  assign N15378 = N15377 | data_masked[15482];
  assign N15377 = N15376 | data_masked[15610];
  assign N15376 = N15375 | data_masked[15738];
  assign N15375 = N15374 | data_masked[15866];
  assign N15374 = N15373 | data_masked[15994];
  assign N15373 = N15372 | data_masked[16122];
  assign N15372 = data_masked[16378] | data_masked[16250];
  assign data_o[123] = N15623 | data_masked[123];
  assign N15623 = N15622 | data_masked[251];
  assign N15622 = N15621 | data_masked[379];
  assign N15621 = N15620 | data_masked[507];
  assign N15620 = N15619 | data_masked[635];
  assign N15619 = N15618 | data_masked[763];
  assign N15618 = N15617 | data_masked[891];
  assign N15617 = N15616 | data_masked[1019];
  assign N15616 = N15615 | data_masked[1147];
  assign N15615 = N15614 | data_masked[1275];
  assign N15614 = N15613 | data_masked[1403];
  assign N15613 = N15612 | data_masked[1531];
  assign N15612 = N15611 | data_masked[1659];
  assign N15611 = N15610 | data_masked[1787];
  assign N15610 = N15609 | data_masked[1915];
  assign N15609 = N15608 | data_masked[2043];
  assign N15608 = N15607 | data_masked[2171];
  assign N15607 = N15606 | data_masked[2299];
  assign N15606 = N15605 | data_masked[2427];
  assign N15605 = N15604 | data_masked[2555];
  assign N15604 = N15603 | data_masked[2683];
  assign N15603 = N15602 | data_masked[2811];
  assign N15602 = N15601 | data_masked[2939];
  assign N15601 = N15600 | data_masked[3067];
  assign N15600 = N15599 | data_masked[3195];
  assign N15599 = N15598 | data_masked[3323];
  assign N15598 = N15597 | data_masked[3451];
  assign N15597 = N15596 | data_masked[3579];
  assign N15596 = N15595 | data_masked[3707];
  assign N15595 = N15594 | data_masked[3835];
  assign N15594 = N15593 | data_masked[3963];
  assign N15593 = N15592 | data_masked[4091];
  assign N15592 = N15591 | data_masked[4219];
  assign N15591 = N15590 | data_masked[4347];
  assign N15590 = N15589 | data_masked[4475];
  assign N15589 = N15588 | data_masked[4603];
  assign N15588 = N15587 | data_masked[4731];
  assign N15587 = N15586 | data_masked[4859];
  assign N15586 = N15585 | data_masked[4987];
  assign N15585 = N15584 | data_masked[5115];
  assign N15584 = N15583 | data_masked[5243];
  assign N15583 = N15582 | data_masked[5371];
  assign N15582 = N15581 | data_masked[5499];
  assign N15581 = N15580 | data_masked[5627];
  assign N15580 = N15579 | data_masked[5755];
  assign N15579 = N15578 | data_masked[5883];
  assign N15578 = N15577 | data_masked[6011];
  assign N15577 = N15576 | data_masked[6139];
  assign N15576 = N15575 | data_masked[6267];
  assign N15575 = N15574 | data_masked[6395];
  assign N15574 = N15573 | data_masked[6523];
  assign N15573 = N15572 | data_masked[6651];
  assign N15572 = N15571 | data_masked[6779];
  assign N15571 = N15570 | data_masked[6907];
  assign N15570 = N15569 | data_masked[7035];
  assign N15569 = N15568 | data_masked[7163];
  assign N15568 = N15567 | data_masked[7291];
  assign N15567 = N15566 | data_masked[7419];
  assign N15566 = N15565 | data_masked[7547];
  assign N15565 = N15564 | data_masked[7675];
  assign N15564 = N15563 | data_masked[7803];
  assign N15563 = N15562 | data_masked[7931];
  assign N15562 = N15561 | data_masked[8059];
  assign N15561 = N15560 | data_masked[8187];
  assign N15560 = N15559 | data_masked[8315];
  assign N15559 = N15558 | data_masked[8443];
  assign N15558 = N15557 | data_masked[8571];
  assign N15557 = N15556 | data_masked[8699];
  assign N15556 = N15555 | data_masked[8827];
  assign N15555 = N15554 | data_masked[8955];
  assign N15554 = N15553 | data_masked[9083];
  assign N15553 = N15552 | data_masked[9211];
  assign N15552 = N15551 | data_masked[9339];
  assign N15551 = N15550 | data_masked[9467];
  assign N15550 = N15549 | data_masked[9595];
  assign N15549 = N15548 | data_masked[9723];
  assign N15548 = N15547 | data_masked[9851];
  assign N15547 = N15546 | data_masked[9979];
  assign N15546 = N15545 | data_masked[10107];
  assign N15545 = N15544 | data_masked[10235];
  assign N15544 = N15543 | data_masked[10363];
  assign N15543 = N15542 | data_masked[10491];
  assign N15542 = N15541 | data_masked[10619];
  assign N15541 = N15540 | data_masked[10747];
  assign N15540 = N15539 | data_masked[10875];
  assign N15539 = N15538 | data_masked[11003];
  assign N15538 = N15537 | data_masked[11131];
  assign N15537 = N15536 | data_masked[11259];
  assign N15536 = N15535 | data_masked[11387];
  assign N15535 = N15534 | data_masked[11515];
  assign N15534 = N15533 | data_masked[11643];
  assign N15533 = N15532 | data_masked[11771];
  assign N15532 = N15531 | data_masked[11899];
  assign N15531 = N15530 | data_masked[12027];
  assign N15530 = N15529 | data_masked[12155];
  assign N15529 = N15528 | data_masked[12283];
  assign N15528 = N15527 | data_masked[12411];
  assign N15527 = N15526 | data_masked[12539];
  assign N15526 = N15525 | data_masked[12667];
  assign N15525 = N15524 | data_masked[12795];
  assign N15524 = N15523 | data_masked[12923];
  assign N15523 = N15522 | data_masked[13051];
  assign N15522 = N15521 | data_masked[13179];
  assign N15521 = N15520 | data_masked[13307];
  assign N15520 = N15519 | data_masked[13435];
  assign N15519 = N15518 | data_masked[13563];
  assign N15518 = N15517 | data_masked[13691];
  assign N15517 = N15516 | data_masked[13819];
  assign N15516 = N15515 | data_masked[13947];
  assign N15515 = N15514 | data_masked[14075];
  assign N15514 = N15513 | data_masked[14203];
  assign N15513 = N15512 | data_masked[14331];
  assign N15512 = N15511 | data_masked[14459];
  assign N15511 = N15510 | data_masked[14587];
  assign N15510 = N15509 | data_masked[14715];
  assign N15509 = N15508 | data_masked[14843];
  assign N15508 = N15507 | data_masked[14971];
  assign N15507 = N15506 | data_masked[15099];
  assign N15506 = N15505 | data_masked[15227];
  assign N15505 = N15504 | data_masked[15355];
  assign N15504 = N15503 | data_masked[15483];
  assign N15503 = N15502 | data_masked[15611];
  assign N15502 = N15501 | data_masked[15739];
  assign N15501 = N15500 | data_masked[15867];
  assign N15500 = N15499 | data_masked[15995];
  assign N15499 = N15498 | data_masked[16123];
  assign N15498 = data_masked[16379] | data_masked[16251];
  assign data_o[124] = N15749 | data_masked[124];
  assign N15749 = N15748 | data_masked[252];
  assign N15748 = N15747 | data_masked[380];
  assign N15747 = N15746 | data_masked[508];
  assign N15746 = N15745 | data_masked[636];
  assign N15745 = N15744 | data_masked[764];
  assign N15744 = N15743 | data_masked[892];
  assign N15743 = N15742 | data_masked[1020];
  assign N15742 = N15741 | data_masked[1148];
  assign N15741 = N15740 | data_masked[1276];
  assign N15740 = N15739 | data_masked[1404];
  assign N15739 = N15738 | data_masked[1532];
  assign N15738 = N15737 | data_masked[1660];
  assign N15737 = N15736 | data_masked[1788];
  assign N15736 = N15735 | data_masked[1916];
  assign N15735 = N15734 | data_masked[2044];
  assign N15734 = N15733 | data_masked[2172];
  assign N15733 = N15732 | data_masked[2300];
  assign N15732 = N15731 | data_masked[2428];
  assign N15731 = N15730 | data_masked[2556];
  assign N15730 = N15729 | data_masked[2684];
  assign N15729 = N15728 | data_masked[2812];
  assign N15728 = N15727 | data_masked[2940];
  assign N15727 = N15726 | data_masked[3068];
  assign N15726 = N15725 | data_masked[3196];
  assign N15725 = N15724 | data_masked[3324];
  assign N15724 = N15723 | data_masked[3452];
  assign N15723 = N15722 | data_masked[3580];
  assign N15722 = N15721 | data_masked[3708];
  assign N15721 = N15720 | data_masked[3836];
  assign N15720 = N15719 | data_masked[3964];
  assign N15719 = N15718 | data_masked[4092];
  assign N15718 = N15717 | data_masked[4220];
  assign N15717 = N15716 | data_masked[4348];
  assign N15716 = N15715 | data_masked[4476];
  assign N15715 = N15714 | data_masked[4604];
  assign N15714 = N15713 | data_masked[4732];
  assign N15713 = N15712 | data_masked[4860];
  assign N15712 = N15711 | data_masked[4988];
  assign N15711 = N15710 | data_masked[5116];
  assign N15710 = N15709 | data_masked[5244];
  assign N15709 = N15708 | data_masked[5372];
  assign N15708 = N15707 | data_masked[5500];
  assign N15707 = N15706 | data_masked[5628];
  assign N15706 = N15705 | data_masked[5756];
  assign N15705 = N15704 | data_masked[5884];
  assign N15704 = N15703 | data_masked[6012];
  assign N15703 = N15702 | data_masked[6140];
  assign N15702 = N15701 | data_masked[6268];
  assign N15701 = N15700 | data_masked[6396];
  assign N15700 = N15699 | data_masked[6524];
  assign N15699 = N15698 | data_masked[6652];
  assign N15698 = N15697 | data_masked[6780];
  assign N15697 = N15696 | data_masked[6908];
  assign N15696 = N15695 | data_masked[7036];
  assign N15695 = N15694 | data_masked[7164];
  assign N15694 = N15693 | data_masked[7292];
  assign N15693 = N15692 | data_masked[7420];
  assign N15692 = N15691 | data_masked[7548];
  assign N15691 = N15690 | data_masked[7676];
  assign N15690 = N15689 | data_masked[7804];
  assign N15689 = N15688 | data_masked[7932];
  assign N15688 = N15687 | data_masked[8060];
  assign N15687 = N15686 | data_masked[8188];
  assign N15686 = N15685 | data_masked[8316];
  assign N15685 = N15684 | data_masked[8444];
  assign N15684 = N15683 | data_masked[8572];
  assign N15683 = N15682 | data_masked[8700];
  assign N15682 = N15681 | data_masked[8828];
  assign N15681 = N15680 | data_masked[8956];
  assign N15680 = N15679 | data_masked[9084];
  assign N15679 = N15678 | data_masked[9212];
  assign N15678 = N15677 | data_masked[9340];
  assign N15677 = N15676 | data_masked[9468];
  assign N15676 = N15675 | data_masked[9596];
  assign N15675 = N15674 | data_masked[9724];
  assign N15674 = N15673 | data_masked[9852];
  assign N15673 = N15672 | data_masked[9980];
  assign N15672 = N15671 | data_masked[10108];
  assign N15671 = N15670 | data_masked[10236];
  assign N15670 = N15669 | data_masked[10364];
  assign N15669 = N15668 | data_masked[10492];
  assign N15668 = N15667 | data_masked[10620];
  assign N15667 = N15666 | data_masked[10748];
  assign N15666 = N15665 | data_masked[10876];
  assign N15665 = N15664 | data_masked[11004];
  assign N15664 = N15663 | data_masked[11132];
  assign N15663 = N15662 | data_masked[11260];
  assign N15662 = N15661 | data_masked[11388];
  assign N15661 = N15660 | data_masked[11516];
  assign N15660 = N15659 | data_masked[11644];
  assign N15659 = N15658 | data_masked[11772];
  assign N15658 = N15657 | data_masked[11900];
  assign N15657 = N15656 | data_masked[12028];
  assign N15656 = N15655 | data_masked[12156];
  assign N15655 = N15654 | data_masked[12284];
  assign N15654 = N15653 | data_masked[12412];
  assign N15653 = N15652 | data_masked[12540];
  assign N15652 = N15651 | data_masked[12668];
  assign N15651 = N15650 | data_masked[12796];
  assign N15650 = N15649 | data_masked[12924];
  assign N15649 = N15648 | data_masked[13052];
  assign N15648 = N15647 | data_masked[13180];
  assign N15647 = N15646 | data_masked[13308];
  assign N15646 = N15645 | data_masked[13436];
  assign N15645 = N15644 | data_masked[13564];
  assign N15644 = N15643 | data_masked[13692];
  assign N15643 = N15642 | data_masked[13820];
  assign N15642 = N15641 | data_masked[13948];
  assign N15641 = N15640 | data_masked[14076];
  assign N15640 = N15639 | data_masked[14204];
  assign N15639 = N15638 | data_masked[14332];
  assign N15638 = N15637 | data_masked[14460];
  assign N15637 = N15636 | data_masked[14588];
  assign N15636 = N15635 | data_masked[14716];
  assign N15635 = N15634 | data_masked[14844];
  assign N15634 = N15633 | data_masked[14972];
  assign N15633 = N15632 | data_masked[15100];
  assign N15632 = N15631 | data_masked[15228];
  assign N15631 = N15630 | data_masked[15356];
  assign N15630 = N15629 | data_masked[15484];
  assign N15629 = N15628 | data_masked[15612];
  assign N15628 = N15627 | data_masked[15740];
  assign N15627 = N15626 | data_masked[15868];
  assign N15626 = N15625 | data_masked[15996];
  assign N15625 = N15624 | data_masked[16124];
  assign N15624 = data_masked[16380] | data_masked[16252];
  assign data_o[125] = N15875 | data_masked[125];
  assign N15875 = N15874 | data_masked[253];
  assign N15874 = N15873 | data_masked[381];
  assign N15873 = N15872 | data_masked[509];
  assign N15872 = N15871 | data_masked[637];
  assign N15871 = N15870 | data_masked[765];
  assign N15870 = N15869 | data_masked[893];
  assign N15869 = N15868 | data_masked[1021];
  assign N15868 = N15867 | data_masked[1149];
  assign N15867 = N15866 | data_masked[1277];
  assign N15866 = N15865 | data_masked[1405];
  assign N15865 = N15864 | data_masked[1533];
  assign N15864 = N15863 | data_masked[1661];
  assign N15863 = N15862 | data_masked[1789];
  assign N15862 = N15861 | data_masked[1917];
  assign N15861 = N15860 | data_masked[2045];
  assign N15860 = N15859 | data_masked[2173];
  assign N15859 = N15858 | data_masked[2301];
  assign N15858 = N15857 | data_masked[2429];
  assign N15857 = N15856 | data_masked[2557];
  assign N15856 = N15855 | data_masked[2685];
  assign N15855 = N15854 | data_masked[2813];
  assign N15854 = N15853 | data_masked[2941];
  assign N15853 = N15852 | data_masked[3069];
  assign N15852 = N15851 | data_masked[3197];
  assign N15851 = N15850 | data_masked[3325];
  assign N15850 = N15849 | data_masked[3453];
  assign N15849 = N15848 | data_masked[3581];
  assign N15848 = N15847 | data_masked[3709];
  assign N15847 = N15846 | data_masked[3837];
  assign N15846 = N15845 | data_masked[3965];
  assign N15845 = N15844 | data_masked[4093];
  assign N15844 = N15843 | data_masked[4221];
  assign N15843 = N15842 | data_masked[4349];
  assign N15842 = N15841 | data_masked[4477];
  assign N15841 = N15840 | data_masked[4605];
  assign N15840 = N15839 | data_masked[4733];
  assign N15839 = N15838 | data_masked[4861];
  assign N15838 = N15837 | data_masked[4989];
  assign N15837 = N15836 | data_masked[5117];
  assign N15836 = N15835 | data_masked[5245];
  assign N15835 = N15834 | data_masked[5373];
  assign N15834 = N15833 | data_masked[5501];
  assign N15833 = N15832 | data_masked[5629];
  assign N15832 = N15831 | data_masked[5757];
  assign N15831 = N15830 | data_masked[5885];
  assign N15830 = N15829 | data_masked[6013];
  assign N15829 = N15828 | data_masked[6141];
  assign N15828 = N15827 | data_masked[6269];
  assign N15827 = N15826 | data_masked[6397];
  assign N15826 = N15825 | data_masked[6525];
  assign N15825 = N15824 | data_masked[6653];
  assign N15824 = N15823 | data_masked[6781];
  assign N15823 = N15822 | data_masked[6909];
  assign N15822 = N15821 | data_masked[7037];
  assign N15821 = N15820 | data_masked[7165];
  assign N15820 = N15819 | data_masked[7293];
  assign N15819 = N15818 | data_masked[7421];
  assign N15818 = N15817 | data_masked[7549];
  assign N15817 = N15816 | data_masked[7677];
  assign N15816 = N15815 | data_masked[7805];
  assign N15815 = N15814 | data_masked[7933];
  assign N15814 = N15813 | data_masked[8061];
  assign N15813 = N15812 | data_masked[8189];
  assign N15812 = N15811 | data_masked[8317];
  assign N15811 = N15810 | data_masked[8445];
  assign N15810 = N15809 | data_masked[8573];
  assign N15809 = N15808 | data_masked[8701];
  assign N15808 = N15807 | data_masked[8829];
  assign N15807 = N15806 | data_masked[8957];
  assign N15806 = N15805 | data_masked[9085];
  assign N15805 = N15804 | data_masked[9213];
  assign N15804 = N15803 | data_masked[9341];
  assign N15803 = N15802 | data_masked[9469];
  assign N15802 = N15801 | data_masked[9597];
  assign N15801 = N15800 | data_masked[9725];
  assign N15800 = N15799 | data_masked[9853];
  assign N15799 = N15798 | data_masked[9981];
  assign N15798 = N15797 | data_masked[10109];
  assign N15797 = N15796 | data_masked[10237];
  assign N15796 = N15795 | data_masked[10365];
  assign N15795 = N15794 | data_masked[10493];
  assign N15794 = N15793 | data_masked[10621];
  assign N15793 = N15792 | data_masked[10749];
  assign N15792 = N15791 | data_masked[10877];
  assign N15791 = N15790 | data_masked[11005];
  assign N15790 = N15789 | data_masked[11133];
  assign N15789 = N15788 | data_masked[11261];
  assign N15788 = N15787 | data_masked[11389];
  assign N15787 = N15786 | data_masked[11517];
  assign N15786 = N15785 | data_masked[11645];
  assign N15785 = N15784 | data_masked[11773];
  assign N15784 = N15783 | data_masked[11901];
  assign N15783 = N15782 | data_masked[12029];
  assign N15782 = N15781 | data_masked[12157];
  assign N15781 = N15780 | data_masked[12285];
  assign N15780 = N15779 | data_masked[12413];
  assign N15779 = N15778 | data_masked[12541];
  assign N15778 = N15777 | data_masked[12669];
  assign N15777 = N15776 | data_masked[12797];
  assign N15776 = N15775 | data_masked[12925];
  assign N15775 = N15774 | data_masked[13053];
  assign N15774 = N15773 | data_masked[13181];
  assign N15773 = N15772 | data_masked[13309];
  assign N15772 = N15771 | data_masked[13437];
  assign N15771 = N15770 | data_masked[13565];
  assign N15770 = N15769 | data_masked[13693];
  assign N15769 = N15768 | data_masked[13821];
  assign N15768 = N15767 | data_masked[13949];
  assign N15767 = N15766 | data_masked[14077];
  assign N15766 = N15765 | data_masked[14205];
  assign N15765 = N15764 | data_masked[14333];
  assign N15764 = N15763 | data_masked[14461];
  assign N15763 = N15762 | data_masked[14589];
  assign N15762 = N15761 | data_masked[14717];
  assign N15761 = N15760 | data_masked[14845];
  assign N15760 = N15759 | data_masked[14973];
  assign N15759 = N15758 | data_masked[15101];
  assign N15758 = N15757 | data_masked[15229];
  assign N15757 = N15756 | data_masked[15357];
  assign N15756 = N15755 | data_masked[15485];
  assign N15755 = N15754 | data_masked[15613];
  assign N15754 = N15753 | data_masked[15741];
  assign N15753 = N15752 | data_masked[15869];
  assign N15752 = N15751 | data_masked[15997];
  assign N15751 = N15750 | data_masked[16125];
  assign N15750 = data_masked[16381] | data_masked[16253];
  assign data_o[126] = N16001 | data_masked[126];
  assign N16001 = N16000 | data_masked[254];
  assign N16000 = N15999 | data_masked[382];
  assign N15999 = N15998 | data_masked[510];
  assign N15998 = N15997 | data_masked[638];
  assign N15997 = N15996 | data_masked[766];
  assign N15996 = N15995 | data_masked[894];
  assign N15995 = N15994 | data_masked[1022];
  assign N15994 = N15993 | data_masked[1150];
  assign N15993 = N15992 | data_masked[1278];
  assign N15992 = N15991 | data_masked[1406];
  assign N15991 = N15990 | data_masked[1534];
  assign N15990 = N15989 | data_masked[1662];
  assign N15989 = N15988 | data_masked[1790];
  assign N15988 = N15987 | data_masked[1918];
  assign N15987 = N15986 | data_masked[2046];
  assign N15986 = N15985 | data_masked[2174];
  assign N15985 = N15984 | data_masked[2302];
  assign N15984 = N15983 | data_masked[2430];
  assign N15983 = N15982 | data_masked[2558];
  assign N15982 = N15981 | data_masked[2686];
  assign N15981 = N15980 | data_masked[2814];
  assign N15980 = N15979 | data_masked[2942];
  assign N15979 = N15978 | data_masked[3070];
  assign N15978 = N15977 | data_masked[3198];
  assign N15977 = N15976 | data_masked[3326];
  assign N15976 = N15975 | data_masked[3454];
  assign N15975 = N15974 | data_masked[3582];
  assign N15974 = N15973 | data_masked[3710];
  assign N15973 = N15972 | data_masked[3838];
  assign N15972 = N15971 | data_masked[3966];
  assign N15971 = N15970 | data_masked[4094];
  assign N15970 = N15969 | data_masked[4222];
  assign N15969 = N15968 | data_masked[4350];
  assign N15968 = N15967 | data_masked[4478];
  assign N15967 = N15966 | data_masked[4606];
  assign N15966 = N15965 | data_masked[4734];
  assign N15965 = N15964 | data_masked[4862];
  assign N15964 = N15963 | data_masked[4990];
  assign N15963 = N15962 | data_masked[5118];
  assign N15962 = N15961 | data_masked[5246];
  assign N15961 = N15960 | data_masked[5374];
  assign N15960 = N15959 | data_masked[5502];
  assign N15959 = N15958 | data_masked[5630];
  assign N15958 = N15957 | data_masked[5758];
  assign N15957 = N15956 | data_masked[5886];
  assign N15956 = N15955 | data_masked[6014];
  assign N15955 = N15954 | data_masked[6142];
  assign N15954 = N15953 | data_masked[6270];
  assign N15953 = N15952 | data_masked[6398];
  assign N15952 = N15951 | data_masked[6526];
  assign N15951 = N15950 | data_masked[6654];
  assign N15950 = N15949 | data_masked[6782];
  assign N15949 = N15948 | data_masked[6910];
  assign N15948 = N15947 | data_masked[7038];
  assign N15947 = N15946 | data_masked[7166];
  assign N15946 = N15945 | data_masked[7294];
  assign N15945 = N15944 | data_masked[7422];
  assign N15944 = N15943 | data_masked[7550];
  assign N15943 = N15942 | data_masked[7678];
  assign N15942 = N15941 | data_masked[7806];
  assign N15941 = N15940 | data_masked[7934];
  assign N15940 = N15939 | data_masked[8062];
  assign N15939 = N15938 | data_masked[8190];
  assign N15938 = N15937 | data_masked[8318];
  assign N15937 = N15936 | data_masked[8446];
  assign N15936 = N15935 | data_masked[8574];
  assign N15935 = N15934 | data_masked[8702];
  assign N15934 = N15933 | data_masked[8830];
  assign N15933 = N15932 | data_masked[8958];
  assign N15932 = N15931 | data_masked[9086];
  assign N15931 = N15930 | data_masked[9214];
  assign N15930 = N15929 | data_masked[9342];
  assign N15929 = N15928 | data_masked[9470];
  assign N15928 = N15927 | data_masked[9598];
  assign N15927 = N15926 | data_masked[9726];
  assign N15926 = N15925 | data_masked[9854];
  assign N15925 = N15924 | data_masked[9982];
  assign N15924 = N15923 | data_masked[10110];
  assign N15923 = N15922 | data_masked[10238];
  assign N15922 = N15921 | data_masked[10366];
  assign N15921 = N15920 | data_masked[10494];
  assign N15920 = N15919 | data_masked[10622];
  assign N15919 = N15918 | data_masked[10750];
  assign N15918 = N15917 | data_masked[10878];
  assign N15917 = N15916 | data_masked[11006];
  assign N15916 = N15915 | data_masked[11134];
  assign N15915 = N15914 | data_masked[11262];
  assign N15914 = N15913 | data_masked[11390];
  assign N15913 = N15912 | data_masked[11518];
  assign N15912 = N15911 | data_masked[11646];
  assign N15911 = N15910 | data_masked[11774];
  assign N15910 = N15909 | data_masked[11902];
  assign N15909 = N15908 | data_masked[12030];
  assign N15908 = N15907 | data_masked[12158];
  assign N15907 = N15906 | data_masked[12286];
  assign N15906 = N15905 | data_masked[12414];
  assign N15905 = N15904 | data_masked[12542];
  assign N15904 = N15903 | data_masked[12670];
  assign N15903 = N15902 | data_masked[12798];
  assign N15902 = N15901 | data_masked[12926];
  assign N15901 = N15900 | data_masked[13054];
  assign N15900 = N15899 | data_masked[13182];
  assign N15899 = N15898 | data_masked[13310];
  assign N15898 = N15897 | data_masked[13438];
  assign N15897 = N15896 | data_masked[13566];
  assign N15896 = N15895 | data_masked[13694];
  assign N15895 = N15894 | data_masked[13822];
  assign N15894 = N15893 | data_masked[13950];
  assign N15893 = N15892 | data_masked[14078];
  assign N15892 = N15891 | data_masked[14206];
  assign N15891 = N15890 | data_masked[14334];
  assign N15890 = N15889 | data_masked[14462];
  assign N15889 = N15888 | data_masked[14590];
  assign N15888 = N15887 | data_masked[14718];
  assign N15887 = N15886 | data_masked[14846];
  assign N15886 = N15885 | data_masked[14974];
  assign N15885 = N15884 | data_masked[15102];
  assign N15884 = N15883 | data_masked[15230];
  assign N15883 = N15882 | data_masked[15358];
  assign N15882 = N15881 | data_masked[15486];
  assign N15881 = N15880 | data_masked[15614];
  assign N15880 = N15879 | data_masked[15742];
  assign N15879 = N15878 | data_masked[15870];
  assign N15878 = N15877 | data_masked[15998];
  assign N15877 = N15876 | data_masked[16126];
  assign N15876 = data_masked[16382] | data_masked[16254];
  assign data_o[127] = N16127 | data_masked[127];
  assign N16127 = N16126 | data_masked[255];
  assign N16126 = N16125 | data_masked[383];
  assign N16125 = N16124 | data_masked[511];
  assign N16124 = N16123 | data_masked[639];
  assign N16123 = N16122 | data_masked[767];
  assign N16122 = N16121 | data_masked[895];
  assign N16121 = N16120 | data_masked[1023];
  assign N16120 = N16119 | data_masked[1151];
  assign N16119 = N16118 | data_masked[1279];
  assign N16118 = N16117 | data_masked[1407];
  assign N16117 = N16116 | data_masked[1535];
  assign N16116 = N16115 | data_masked[1663];
  assign N16115 = N16114 | data_masked[1791];
  assign N16114 = N16113 | data_masked[1919];
  assign N16113 = N16112 | data_masked[2047];
  assign N16112 = N16111 | data_masked[2175];
  assign N16111 = N16110 | data_masked[2303];
  assign N16110 = N16109 | data_masked[2431];
  assign N16109 = N16108 | data_masked[2559];
  assign N16108 = N16107 | data_masked[2687];
  assign N16107 = N16106 | data_masked[2815];
  assign N16106 = N16105 | data_masked[2943];
  assign N16105 = N16104 | data_masked[3071];
  assign N16104 = N16103 | data_masked[3199];
  assign N16103 = N16102 | data_masked[3327];
  assign N16102 = N16101 | data_masked[3455];
  assign N16101 = N16100 | data_masked[3583];
  assign N16100 = N16099 | data_masked[3711];
  assign N16099 = N16098 | data_masked[3839];
  assign N16098 = N16097 | data_masked[3967];
  assign N16097 = N16096 | data_masked[4095];
  assign N16096 = N16095 | data_masked[4223];
  assign N16095 = N16094 | data_masked[4351];
  assign N16094 = N16093 | data_masked[4479];
  assign N16093 = N16092 | data_masked[4607];
  assign N16092 = N16091 | data_masked[4735];
  assign N16091 = N16090 | data_masked[4863];
  assign N16090 = N16089 | data_masked[4991];
  assign N16089 = N16088 | data_masked[5119];
  assign N16088 = N16087 | data_masked[5247];
  assign N16087 = N16086 | data_masked[5375];
  assign N16086 = N16085 | data_masked[5503];
  assign N16085 = N16084 | data_masked[5631];
  assign N16084 = N16083 | data_masked[5759];
  assign N16083 = N16082 | data_masked[5887];
  assign N16082 = N16081 | data_masked[6015];
  assign N16081 = N16080 | data_masked[6143];
  assign N16080 = N16079 | data_masked[6271];
  assign N16079 = N16078 | data_masked[6399];
  assign N16078 = N16077 | data_masked[6527];
  assign N16077 = N16076 | data_masked[6655];
  assign N16076 = N16075 | data_masked[6783];
  assign N16075 = N16074 | data_masked[6911];
  assign N16074 = N16073 | data_masked[7039];
  assign N16073 = N16072 | data_masked[7167];
  assign N16072 = N16071 | data_masked[7295];
  assign N16071 = N16070 | data_masked[7423];
  assign N16070 = N16069 | data_masked[7551];
  assign N16069 = N16068 | data_masked[7679];
  assign N16068 = N16067 | data_masked[7807];
  assign N16067 = N16066 | data_masked[7935];
  assign N16066 = N16065 | data_masked[8063];
  assign N16065 = N16064 | data_masked[8191];
  assign N16064 = N16063 | data_masked[8319];
  assign N16063 = N16062 | data_masked[8447];
  assign N16062 = N16061 | data_masked[8575];
  assign N16061 = N16060 | data_masked[8703];
  assign N16060 = N16059 | data_masked[8831];
  assign N16059 = N16058 | data_masked[8959];
  assign N16058 = N16057 | data_masked[9087];
  assign N16057 = N16056 | data_masked[9215];
  assign N16056 = N16055 | data_masked[9343];
  assign N16055 = N16054 | data_masked[9471];
  assign N16054 = N16053 | data_masked[9599];
  assign N16053 = N16052 | data_masked[9727];
  assign N16052 = N16051 | data_masked[9855];
  assign N16051 = N16050 | data_masked[9983];
  assign N16050 = N16049 | data_masked[10111];
  assign N16049 = N16048 | data_masked[10239];
  assign N16048 = N16047 | data_masked[10367];
  assign N16047 = N16046 | data_masked[10495];
  assign N16046 = N16045 | data_masked[10623];
  assign N16045 = N16044 | data_masked[10751];
  assign N16044 = N16043 | data_masked[10879];
  assign N16043 = N16042 | data_masked[11007];
  assign N16042 = N16041 | data_masked[11135];
  assign N16041 = N16040 | data_masked[11263];
  assign N16040 = N16039 | data_masked[11391];
  assign N16039 = N16038 | data_masked[11519];
  assign N16038 = N16037 | data_masked[11647];
  assign N16037 = N16036 | data_masked[11775];
  assign N16036 = N16035 | data_masked[11903];
  assign N16035 = N16034 | data_masked[12031];
  assign N16034 = N16033 | data_masked[12159];
  assign N16033 = N16032 | data_masked[12287];
  assign N16032 = N16031 | data_masked[12415];
  assign N16031 = N16030 | data_masked[12543];
  assign N16030 = N16029 | data_masked[12671];
  assign N16029 = N16028 | data_masked[12799];
  assign N16028 = N16027 | data_masked[12927];
  assign N16027 = N16026 | data_masked[13055];
  assign N16026 = N16025 | data_masked[13183];
  assign N16025 = N16024 | data_masked[13311];
  assign N16024 = N16023 | data_masked[13439];
  assign N16023 = N16022 | data_masked[13567];
  assign N16022 = N16021 | data_masked[13695];
  assign N16021 = N16020 | data_masked[13823];
  assign N16020 = N16019 | data_masked[13951];
  assign N16019 = N16018 | data_masked[14079];
  assign N16018 = N16017 | data_masked[14207];
  assign N16017 = N16016 | data_masked[14335];
  assign N16016 = N16015 | data_masked[14463];
  assign N16015 = N16014 | data_masked[14591];
  assign N16014 = N16013 | data_masked[14719];
  assign N16013 = N16012 | data_masked[14847];
  assign N16012 = N16011 | data_masked[14975];
  assign N16011 = N16010 | data_masked[15103];
  assign N16010 = N16009 | data_masked[15231];
  assign N16009 = N16008 | data_masked[15359];
  assign N16008 = N16007 | data_masked[15487];
  assign N16007 = N16006 | data_masked[15615];
  assign N16006 = N16005 | data_masked[15743];
  assign N16005 = N16004 | data_masked[15871];
  assign N16004 = N16003 | data_masked[15999];
  assign N16003 = N16002 | data_masked[16127];
  assign N16002 = data_masked[16383] | data_masked[16255];

endmodule



module bsg_crossbar_o_by_i
(
  i,
  sel_oi_one_hot_i,
  o
);

  input [16383:0] i;
  input [16383:0] sel_oi_one_hot_i;
  output [16383:0] o;
  wire [16383:0] o;

  bsg_mux_one_hot_width_p128_els_p128
  genblk1_0__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[127:0]),
    .data_o(o[127:0])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_1__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[255:128]),
    .data_o(o[255:128])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_2__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[383:256]),
    .data_o(o[383:256])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_3__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[511:384]),
    .data_o(o[511:384])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_4__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[639:512]),
    .data_o(o[639:512])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_5__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[767:640]),
    .data_o(o[767:640])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_6__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[895:768]),
    .data_o(o[895:768])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_7__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1023:896]),
    .data_o(o[1023:896])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_8__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1151:1024]),
    .data_o(o[1151:1024])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_9__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1279:1152]),
    .data_o(o[1279:1152])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_10__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1407:1280]),
    .data_o(o[1407:1280])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_11__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1535:1408]),
    .data_o(o[1535:1408])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_12__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1663:1536]),
    .data_o(o[1663:1536])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_13__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1791:1664]),
    .data_o(o[1791:1664])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_14__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1919:1792]),
    .data_o(o[1919:1792])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_15__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2047:1920]),
    .data_o(o[2047:1920])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_16__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2175:2048]),
    .data_o(o[2175:2048])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_17__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2303:2176]),
    .data_o(o[2303:2176])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_18__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2431:2304]),
    .data_o(o[2431:2304])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_19__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2559:2432]),
    .data_o(o[2559:2432])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_20__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2687:2560]),
    .data_o(o[2687:2560])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_21__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2815:2688]),
    .data_o(o[2815:2688])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_22__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2943:2816]),
    .data_o(o[2943:2816])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_23__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3071:2944]),
    .data_o(o[3071:2944])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_24__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3199:3072]),
    .data_o(o[3199:3072])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_25__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3327:3200]),
    .data_o(o[3327:3200])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_26__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3455:3328]),
    .data_o(o[3455:3328])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_27__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3583:3456]),
    .data_o(o[3583:3456])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_28__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3711:3584]),
    .data_o(o[3711:3584])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_29__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3839:3712]),
    .data_o(o[3839:3712])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_30__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3967:3840]),
    .data_o(o[3967:3840])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_31__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[4095:3968]),
    .data_o(o[4095:3968])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_32__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[4223:4096]),
    .data_o(o[4223:4096])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_33__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[4351:4224]),
    .data_o(o[4351:4224])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_34__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[4479:4352]),
    .data_o(o[4479:4352])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_35__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[4607:4480]),
    .data_o(o[4607:4480])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_36__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[4735:4608]),
    .data_o(o[4735:4608])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_37__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[4863:4736]),
    .data_o(o[4863:4736])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_38__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[4991:4864]),
    .data_o(o[4991:4864])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_39__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[5119:4992]),
    .data_o(o[5119:4992])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_40__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[5247:5120]),
    .data_o(o[5247:5120])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_41__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[5375:5248]),
    .data_o(o[5375:5248])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_42__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[5503:5376]),
    .data_o(o[5503:5376])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_43__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[5631:5504]),
    .data_o(o[5631:5504])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_44__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[5759:5632]),
    .data_o(o[5759:5632])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_45__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[5887:5760]),
    .data_o(o[5887:5760])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_46__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[6015:5888]),
    .data_o(o[6015:5888])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_47__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[6143:6016]),
    .data_o(o[6143:6016])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_48__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[6271:6144]),
    .data_o(o[6271:6144])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_49__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[6399:6272]),
    .data_o(o[6399:6272])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_50__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[6527:6400]),
    .data_o(o[6527:6400])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_51__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[6655:6528]),
    .data_o(o[6655:6528])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_52__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[6783:6656]),
    .data_o(o[6783:6656])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_53__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[6911:6784]),
    .data_o(o[6911:6784])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_54__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[7039:6912]),
    .data_o(o[7039:6912])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_55__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[7167:7040]),
    .data_o(o[7167:7040])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_56__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[7295:7168]),
    .data_o(o[7295:7168])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_57__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[7423:7296]),
    .data_o(o[7423:7296])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_58__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[7551:7424]),
    .data_o(o[7551:7424])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_59__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[7679:7552]),
    .data_o(o[7679:7552])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_60__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[7807:7680]),
    .data_o(o[7807:7680])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_61__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[7935:7808]),
    .data_o(o[7935:7808])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_62__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[8063:7936]),
    .data_o(o[8063:7936])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_63__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[8191:8064]),
    .data_o(o[8191:8064])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_64__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[8319:8192]),
    .data_o(o[8319:8192])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_65__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[8447:8320]),
    .data_o(o[8447:8320])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_66__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[8575:8448]),
    .data_o(o[8575:8448])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_67__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[8703:8576]),
    .data_o(o[8703:8576])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_68__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[8831:8704]),
    .data_o(o[8831:8704])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_69__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[8959:8832]),
    .data_o(o[8959:8832])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_70__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[9087:8960]),
    .data_o(o[9087:8960])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_71__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[9215:9088]),
    .data_o(o[9215:9088])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_72__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[9343:9216]),
    .data_o(o[9343:9216])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_73__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[9471:9344]),
    .data_o(o[9471:9344])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_74__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[9599:9472]),
    .data_o(o[9599:9472])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_75__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[9727:9600]),
    .data_o(o[9727:9600])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_76__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[9855:9728]),
    .data_o(o[9855:9728])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_77__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[9983:9856]),
    .data_o(o[9983:9856])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_78__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[10111:9984]),
    .data_o(o[10111:9984])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_79__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[10239:10112]),
    .data_o(o[10239:10112])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_80__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[10367:10240]),
    .data_o(o[10367:10240])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_81__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[10495:10368]),
    .data_o(o[10495:10368])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_82__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[10623:10496]),
    .data_o(o[10623:10496])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_83__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[10751:10624]),
    .data_o(o[10751:10624])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_84__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[10879:10752]),
    .data_o(o[10879:10752])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_85__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[11007:10880]),
    .data_o(o[11007:10880])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_86__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[11135:11008]),
    .data_o(o[11135:11008])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_87__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[11263:11136]),
    .data_o(o[11263:11136])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_88__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[11391:11264]),
    .data_o(o[11391:11264])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_89__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[11519:11392]),
    .data_o(o[11519:11392])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_90__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[11647:11520]),
    .data_o(o[11647:11520])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_91__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[11775:11648]),
    .data_o(o[11775:11648])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_92__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[11903:11776]),
    .data_o(o[11903:11776])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_93__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[12031:11904]),
    .data_o(o[12031:11904])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_94__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[12159:12032]),
    .data_o(o[12159:12032])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_95__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[12287:12160]),
    .data_o(o[12287:12160])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_96__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[12415:12288]),
    .data_o(o[12415:12288])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_97__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[12543:12416]),
    .data_o(o[12543:12416])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_98__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[12671:12544]),
    .data_o(o[12671:12544])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_99__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[12799:12672]),
    .data_o(o[12799:12672])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_100__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[12927:12800]),
    .data_o(o[12927:12800])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_101__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[13055:12928]),
    .data_o(o[13055:12928])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_102__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[13183:13056]),
    .data_o(o[13183:13056])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_103__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[13311:13184]),
    .data_o(o[13311:13184])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_104__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[13439:13312]),
    .data_o(o[13439:13312])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_105__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[13567:13440]),
    .data_o(o[13567:13440])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_106__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[13695:13568]),
    .data_o(o[13695:13568])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_107__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[13823:13696]),
    .data_o(o[13823:13696])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_108__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[13951:13824]),
    .data_o(o[13951:13824])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_109__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[14079:13952]),
    .data_o(o[14079:13952])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_110__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[14207:14080]),
    .data_o(o[14207:14080])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_111__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[14335:14208]),
    .data_o(o[14335:14208])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_112__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[14463:14336]),
    .data_o(o[14463:14336])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_113__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[14591:14464]),
    .data_o(o[14591:14464])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_114__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[14719:14592]),
    .data_o(o[14719:14592])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_115__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[14847:14720]),
    .data_o(o[14847:14720])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_116__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[14975:14848]),
    .data_o(o[14975:14848])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_117__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[15103:14976]),
    .data_o(o[15103:14976])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_118__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[15231:15104]),
    .data_o(o[15231:15104])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_119__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[15359:15232]),
    .data_o(o[15359:15232])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_120__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[15487:15360]),
    .data_o(o[15487:15360])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_121__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[15615:15488]),
    .data_o(o[15615:15488])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_122__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[15743:15616]),
    .data_o(o[15743:15616])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_123__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[15871:15744]),
    .data_o(o[15871:15744])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_124__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[15999:15872]),
    .data_o(o[15999:15872])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_125__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[16127:16000]),
    .data_o(o[16127:16000])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_126__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[16255:16128]),
    .data_o(o[16255:16128])
  );


  bsg_mux_one_hot_width_p128_els_p128
  genblk1_127__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[16383:16256]),
    .data_o(o[16383:16256])
  );


endmodule

