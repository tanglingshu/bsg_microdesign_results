

module top
(
  clk_i,
  reset_i,
  v_i,
  tag_i,
  yumi_o,
  v_o,
  ready_i
);

  input [6:0] tag_i;
  output [127:0] v_o;
  input [127:0] ready_i;
  input clk_i;
  input reset_i;
  input v_i;
  output yumi_o;

  bsg_1_to_n_tagged
  wrapper
  (
    .tag_i(tag_i),
    .v_o(v_o),
    .ready_i(ready_i),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .yumi_o(yumi_o)
  );


endmodule



module bsg_decode_num_out_p128
(
  i,
  o
);

  input [6:0] i;
  output [127:0] o;
  wire [127:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_decode_with_v_num_out_p128
(
  i,
  v_i,
  o
);

  input [6:0] i;
  output [127:0] o;
  input v_i;
  wire [127:0] o,lo;

  bsg_decode_num_out_p128
  bd
  (
    .i(i),
    .o(lo)
  );

  assign o[127] = v_i & lo[127];
  assign o[126] = v_i & lo[126];
  assign o[125] = v_i & lo[125];
  assign o[124] = v_i & lo[124];
  assign o[123] = v_i & lo[123];
  assign o[122] = v_i & lo[122];
  assign o[121] = v_i & lo[121];
  assign o[120] = v_i & lo[120];
  assign o[119] = v_i & lo[119];
  assign o[118] = v_i & lo[118];
  assign o[117] = v_i & lo[117];
  assign o[116] = v_i & lo[116];
  assign o[115] = v_i & lo[115];
  assign o[114] = v_i & lo[114];
  assign o[113] = v_i & lo[113];
  assign o[112] = v_i & lo[112];
  assign o[111] = v_i & lo[111];
  assign o[110] = v_i & lo[110];
  assign o[109] = v_i & lo[109];
  assign o[108] = v_i & lo[108];
  assign o[107] = v_i & lo[107];
  assign o[106] = v_i & lo[106];
  assign o[105] = v_i & lo[105];
  assign o[104] = v_i & lo[104];
  assign o[103] = v_i & lo[103];
  assign o[102] = v_i & lo[102];
  assign o[101] = v_i & lo[101];
  assign o[100] = v_i & lo[100];
  assign o[99] = v_i & lo[99];
  assign o[98] = v_i & lo[98];
  assign o[97] = v_i & lo[97];
  assign o[96] = v_i & lo[96];
  assign o[95] = v_i & lo[95];
  assign o[94] = v_i & lo[94];
  assign o[93] = v_i & lo[93];
  assign o[92] = v_i & lo[92];
  assign o[91] = v_i & lo[91];
  assign o[90] = v_i & lo[90];
  assign o[89] = v_i & lo[89];
  assign o[88] = v_i & lo[88];
  assign o[87] = v_i & lo[87];
  assign o[86] = v_i & lo[86];
  assign o[85] = v_i & lo[85];
  assign o[84] = v_i & lo[84];
  assign o[83] = v_i & lo[83];
  assign o[82] = v_i & lo[82];
  assign o[81] = v_i & lo[81];
  assign o[80] = v_i & lo[80];
  assign o[79] = v_i & lo[79];
  assign o[78] = v_i & lo[78];
  assign o[77] = v_i & lo[77];
  assign o[76] = v_i & lo[76];
  assign o[75] = v_i & lo[75];
  assign o[74] = v_i & lo[74];
  assign o[73] = v_i & lo[73];
  assign o[72] = v_i & lo[72];
  assign o[71] = v_i & lo[71];
  assign o[70] = v_i & lo[70];
  assign o[69] = v_i & lo[69];
  assign o[68] = v_i & lo[68];
  assign o[67] = v_i & lo[67];
  assign o[66] = v_i & lo[66];
  assign o[65] = v_i & lo[65];
  assign o[64] = v_i & lo[64];
  assign o[63] = v_i & lo[63];
  assign o[62] = v_i & lo[62];
  assign o[61] = v_i & lo[61];
  assign o[60] = v_i & lo[60];
  assign o[59] = v_i & lo[59];
  assign o[58] = v_i & lo[58];
  assign o[57] = v_i & lo[57];
  assign o[56] = v_i & lo[56];
  assign o[55] = v_i & lo[55];
  assign o[54] = v_i & lo[54];
  assign o[53] = v_i & lo[53];
  assign o[52] = v_i & lo[52];
  assign o[51] = v_i & lo[51];
  assign o[50] = v_i & lo[50];
  assign o[49] = v_i & lo[49];
  assign o[48] = v_i & lo[48];
  assign o[47] = v_i & lo[47];
  assign o[46] = v_i & lo[46];
  assign o[45] = v_i & lo[45];
  assign o[44] = v_i & lo[44];
  assign o[43] = v_i & lo[43];
  assign o[42] = v_i & lo[42];
  assign o[41] = v_i & lo[41];
  assign o[40] = v_i & lo[40];
  assign o[39] = v_i & lo[39];
  assign o[38] = v_i & lo[38];
  assign o[37] = v_i & lo[37];
  assign o[36] = v_i & lo[36];
  assign o[35] = v_i & lo[35];
  assign o[34] = v_i & lo[34];
  assign o[33] = v_i & lo[33];
  assign o[32] = v_i & lo[32];
  assign o[31] = v_i & lo[31];
  assign o[30] = v_i & lo[30];
  assign o[29] = v_i & lo[29];
  assign o[28] = v_i & lo[28];
  assign o[27] = v_i & lo[27];
  assign o[26] = v_i & lo[26];
  assign o[25] = v_i & lo[25];
  assign o[24] = v_i & lo[24];
  assign o[23] = v_i & lo[23];
  assign o[22] = v_i & lo[22];
  assign o[21] = v_i & lo[21];
  assign o[20] = v_i & lo[20];
  assign o[19] = v_i & lo[19];
  assign o[18] = v_i & lo[18];
  assign o[17] = v_i & lo[17];
  assign o[16] = v_i & lo[16];
  assign o[15] = v_i & lo[15];
  assign o[14] = v_i & lo[14];
  assign o[13] = v_i & lo[13];
  assign o[12] = v_i & lo[12];
  assign o[11] = v_i & lo[11];
  assign o[10] = v_i & lo[10];
  assign o[9] = v_i & lo[9];
  assign o[8] = v_i & lo[8];
  assign o[7] = v_i & lo[7];
  assign o[6] = v_i & lo[6];
  assign o[5] = v_i & lo[5];
  assign o[4] = v_i & lo[4];
  assign o[3] = v_i & lo[3];
  assign o[2] = v_i & lo[2];
  assign o[1] = v_i & lo[1];
  assign o[0] = v_i & lo[0];

endmodule



module bsg_1_to_n_tagged
(
  clk_i,
  reset_i,
  v_i,
  tag_i,
  yumi_o,
  v_o,
  ready_i
);

  input [6:0] tag_i;
  output [127:0] v_o;
  input [127:0] ready_i;
  input clk_i;
  input reset_i;
  input v_i;
  output yumi_o;
  wire [127:0] v_o;
  wire yumi_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259;

  bsg_decode_with_v_num_out_p128
  many_bdv
  (
    .i(tag_i),
    .v_i(v_i),
    .o(v_o)
  );

  assign N259 = (N131)? ready_i[0] : 
                (N133)? ready_i[1] : 
                (N135)? ready_i[2] : 
                (N137)? ready_i[3] : 
                (N139)? ready_i[4] : 
                (N141)? ready_i[5] : 
                (N143)? ready_i[6] : 
                (N145)? ready_i[7] : 
                (N147)? ready_i[8] : 
                (N149)? ready_i[9] : 
                (N151)? ready_i[10] : 
                (N153)? ready_i[11] : 
                (N155)? ready_i[12] : 
                (N157)? ready_i[13] : 
                (N159)? ready_i[14] : 
                (N161)? ready_i[15] : 
                (N163)? ready_i[16] : 
                (N165)? ready_i[17] : 
                (N167)? ready_i[18] : 
                (N169)? ready_i[19] : 
                (N171)? ready_i[20] : 
                (N173)? ready_i[21] : 
                (N175)? ready_i[22] : 
                (N177)? ready_i[23] : 
                (N179)? ready_i[24] : 
                (N181)? ready_i[25] : 
                (N183)? ready_i[26] : 
                (N185)? ready_i[27] : 
                (N187)? ready_i[28] : 
                (N189)? ready_i[29] : 
                (N191)? ready_i[30] : 
                (N193)? ready_i[31] : 
                (N195)? ready_i[32] : 
                (N197)? ready_i[33] : 
                (N199)? ready_i[34] : 
                (N201)? ready_i[35] : 
                (N203)? ready_i[36] : 
                (N205)? ready_i[37] : 
                (N207)? ready_i[38] : 
                (N209)? ready_i[39] : 
                (N211)? ready_i[40] : 
                (N213)? ready_i[41] : 
                (N215)? ready_i[42] : 
                (N217)? ready_i[43] : 
                (N219)? ready_i[44] : 
                (N221)? ready_i[45] : 
                (N223)? ready_i[46] : 
                (N225)? ready_i[47] : 
                (N227)? ready_i[48] : 
                (N229)? ready_i[49] : 
                (N231)? ready_i[50] : 
                (N233)? ready_i[51] : 
                (N235)? ready_i[52] : 
                (N237)? ready_i[53] : 
                (N239)? ready_i[54] : 
                (N241)? ready_i[55] : 
                (N243)? ready_i[56] : 
                (N245)? ready_i[57] : 
                (N247)? ready_i[58] : 
                (N249)? ready_i[59] : 
                (N251)? ready_i[60] : 
                (N253)? ready_i[61] : 
                (N255)? ready_i[62] : 
                (N257)? ready_i[63] : 
                (N132)? ready_i[64] : 
                (N134)? ready_i[65] : 
                (N136)? ready_i[66] : 
                (N138)? ready_i[67] : 
                (N140)? ready_i[68] : 
                (N142)? ready_i[69] : 
                (N144)? ready_i[70] : 
                (N146)? ready_i[71] : 
                (N148)? ready_i[72] : 
                (N150)? ready_i[73] : 
                (N152)? ready_i[74] : 
                (N154)? ready_i[75] : 
                (N156)? ready_i[76] : 
                (N158)? ready_i[77] : 
                (N160)? ready_i[78] : 
                (N162)? ready_i[79] : 
                (N164)? ready_i[80] : 
                (N166)? ready_i[81] : 
                (N168)? ready_i[82] : 
                (N170)? ready_i[83] : 
                (N172)? ready_i[84] : 
                (N174)? ready_i[85] : 
                (N176)? ready_i[86] : 
                (N178)? ready_i[87] : 
                (N180)? ready_i[88] : 
                (N182)? ready_i[89] : 
                (N184)? ready_i[90] : 
                (N186)? ready_i[91] : 
                (N188)? ready_i[92] : 
                (N190)? ready_i[93] : 
                (N192)? ready_i[94] : 
                (N194)? ready_i[95] : 
                (N196)? ready_i[96] : 
                (N198)? ready_i[97] : 
                (N200)? ready_i[98] : 
                (N202)? ready_i[99] : 
                (N204)? ready_i[100] : 
                (N206)? ready_i[101] : 
                (N208)? ready_i[102] : 
                (N210)? ready_i[103] : 
                (N212)? ready_i[104] : 
                (N214)? ready_i[105] : 
                (N216)? ready_i[106] : 
                (N218)? ready_i[107] : 
                (N220)? ready_i[108] : 
                (N222)? ready_i[109] : 
                (N224)? ready_i[110] : 
                (N226)? ready_i[111] : 
                (N228)? ready_i[112] : 
                (N230)? ready_i[113] : 
                (N232)? ready_i[114] : 
                (N234)? ready_i[115] : 
                (N236)? ready_i[116] : 
                (N238)? ready_i[117] : 
                (N240)? ready_i[118] : 
                (N242)? ready_i[119] : 
                (N244)? ready_i[120] : 
                (N246)? ready_i[121] : 
                (N248)? ready_i[122] : 
                (N250)? ready_i[123] : 
                (N252)? ready_i[124] : 
                (N254)? ready_i[125] : 
                (N256)? ready_i[126] : 
                (N258)? ready_i[127] : 1'b0;
  assign N0 = ~tag_i[0];
  assign N1 = ~tag_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & tag_i[1];
  assign N4 = tag_i[0] & N1;
  assign N5 = tag_i[0] & tag_i[1];
  assign N6 = ~tag_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & tag_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & tag_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & tag_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & tag_i[2];
  assign N15 = ~tag_i[3];
  assign N16 = N7 & N15;
  assign N17 = N7 & tag_i[3];
  assign N18 = N9 & N15;
  assign N19 = N9 & tag_i[3];
  assign N20 = N11 & N15;
  assign N21 = N11 & tag_i[3];
  assign N22 = N13 & N15;
  assign N23 = N13 & tag_i[3];
  assign N24 = N8 & N15;
  assign N25 = N8 & tag_i[3];
  assign N26 = N10 & N15;
  assign N27 = N10 & tag_i[3];
  assign N28 = N12 & N15;
  assign N29 = N12 & tag_i[3];
  assign N30 = N14 & N15;
  assign N31 = N14 & tag_i[3];
  assign N32 = ~tag_i[4];
  assign N33 = N16 & N32;
  assign N34 = N16 & tag_i[4];
  assign N35 = N18 & N32;
  assign N36 = N18 & tag_i[4];
  assign N37 = N20 & N32;
  assign N38 = N20 & tag_i[4];
  assign N39 = N22 & N32;
  assign N40 = N22 & tag_i[4];
  assign N41 = N24 & N32;
  assign N42 = N24 & tag_i[4];
  assign N43 = N26 & N32;
  assign N44 = N26 & tag_i[4];
  assign N45 = N28 & N32;
  assign N46 = N28 & tag_i[4];
  assign N47 = N30 & N32;
  assign N48 = N30 & tag_i[4];
  assign N49 = N17 & N32;
  assign N50 = N17 & tag_i[4];
  assign N51 = N19 & N32;
  assign N52 = N19 & tag_i[4];
  assign N53 = N21 & N32;
  assign N54 = N21 & tag_i[4];
  assign N55 = N23 & N32;
  assign N56 = N23 & tag_i[4];
  assign N57 = N25 & N32;
  assign N58 = N25 & tag_i[4];
  assign N59 = N27 & N32;
  assign N60 = N27 & tag_i[4];
  assign N61 = N29 & N32;
  assign N62 = N29 & tag_i[4];
  assign N63 = N31 & N32;
  assign N64 = N31 & tag_i[4];
  assign N65 = ~tag_i[5];
  assign N66 = N33 & N65;
  assign N67 = N33 & tag_i[5];
  assign N68 = N35 & N65;
  assign N69 = N35 & tag_i[5];
  assign N70 = N37 & N65;
  assign N71 = N37 & tag_i[5];
  assign N72 = N39 & N65;
  assign N73 = N39 & tag_i[5];
  assign N74 = N41 & N65;
  assign N75 = N41 & tag_i[5];
  assign N76 = N43 & N65;
  assign N77 = N43 & tag_i[5];
  assign N78 = N45 & N65;
  assign N79 = N45 & tag_i[5];
  assign N80 = N47 & N65;
  assign N81 = N47 & tag_i[5];
  assign N82 = N49 & N65;
  assign N83 = N49 & tag_i[5];
  assign N84 = N51 & N65;
  assign N85 = N51 & tag_i[5];
  assign N86 = N53 & N65;
  assign N87 = N53 & tag_i[5];
  assign N88 = N55 & N65;
  assign N89 = N55 & tag_i[5];
  assign N90 = N57 & N65;
  assign N91 = N57 & tag_i[5];
  assign N92 = N59 & N65;
  assign N93 = N59 & tag_i[5];
  assign N94 = N61 & N65;
  assign N95 = N61 & tag_i[5];
  assign N96 = N63 & N65;
  assign N97 = N63 & tag_i[5];
  assign N98 = N34 & N65;
  assign N99 = N34 & tag_i[5];
  assign N100 = N36 & N65;
  assign N101 = N36 & tag_i[5];
  assign N102 = N38 & N65;
  assign N103 = N38 & tag_i[5];
  assign N104 = N40 & N65;
  assign N105 = N40 & tag_i[5];
  assign N106 = N42 & N65;
  assign N107 = N42 & tag_i[5];
  assign N108 = N44 & N65;
  assign N109 = N44 & tag_i[5];
  assign N110 = N46 & N65;
  assign N111 = N46 & tag_i[5];
  assign N112 = N48 & N65;
  assign N113 = N48 & tag_i[5];
  assign N114 = N50 & N65;
  assign N115 = N50 & tag_i[5];
  assign N116 = N52 & N65;
  assign N117 = N52 & tag_i[5];
  assign N118 = N54 & N65;
  assign N119 = N54 & tag_i[5];
  assign N120 = N56 & N65;
  assign N121 = N56 & tag_i[5];
  assign N122 = N58 & N65;
  assign N123 = N58 & tag_i[5];
  assign N124 = N60 & N65;
  assign N125 = N60 & tag_i[5];
  assign N126 = N62 & N65;
  assign N127 = N62 & tag_i[5];
  assign N128 = N64 & N65;
  assign N129 = N64 & tag_i[5];
  assign N130 = ~tag_i[6];
  assign N131 = N66 & N130;
  assign N132 = N66 & tag_i[6];
  assign N133 = N68 & N130;
  assign N134 = N68 & tag_i[6];
  assign N135 = N70 & N130;
  assign N136 = N70 & tag_i[6];
  assign N137 = N72 & N130;
  assign N138 = N72 & tag_i[6];
  assign N139 = N74 & N130;
  assign N140 = N74 & tag_i[6];
  assign N141 = N76 & N130;
  assign N142 = N76 & tag_i[6];
  assign N143 = N78 & N130;
  assign N144 = N78 & tag_i[6];
  assign N145 = N80 & N130;
  assign N146 = N80 & tag_i[6];
  assign N147 = N82 & N130;
  assign N148 = N82 & tag_i[6];
  assign N149 = N84 & N130;
  assign N150 = N84 & tag_i[6];
  assign N151 = N86 & N130;
  assign N152 = N86 & tag_i[6];
  assign N153 = N88 & N130;
  assign N154 = N88 & tag_i[6];
  assign N155 = N90 & N130;
  assign N156 = N90 & tag_i[6];
  assign N157 = N92 & N130;
  assign N158 = N92 & tag_i[6];
  assign N159 = N94 & N130;
  assign N160 = N94 & tag_i[6];
  assign N161 = N96 & N130;
  assign N162 = N96 & tag_i[6];
  assign N163 = N98 & N130;
  assign N164 = N98 & tag_i[6];
  assign N165 = N100 & N130;
  assign N166 = N100 & tag_i[6];
  assign N167 = N102 & N130;
  assign N168 = N102 & tag_i[6];
  assign N169 = N104 & N130;
  assign N170 = N104 & tag_i[6];
  assign N171 = N106 & N130;
  assign N172 = N106 & tag_i[6];
  assign N173 = N108 & N130;
  assign N174 = N108 & tag_i[6];
  assign N175 = N110 & N130;
  assign N176 = N110 & tag_i[6];
  assign N177 = N112 & N130;
  assign N178 = N112 & tag_i[6];
  assign N179 = N114 & N130;
  assign N180 = N114 & tag_i[6];
  assign N181 = N116 & N130;
  assign N182 = N116 & tag_i[6];
  assign N183 = N118 & N130;
  assign N184 = N118 & tag_i[6];
  assign N185 = N120 & N130;
  assign N186 = N120 & tag_i[6];
  assign N187 = N122 & N130;
  assign N188 = N122 & tag_i[6];
  assign N189 = N124 & N130;
  assign N190 = N124 & tag_i[6];
  assign N191 = N126 & N130;
  assign N192 = N126 & tag_i[6];
  assign N193 = N128 & N130;
  assign N194 = N128 & tag_i[6];
  assign N195 = N67 & N130;
  assign N196 = N67 & tag_i[6];
  assign N197 = N69 & N130;
  assign N198 = N69 & tag_i[6];
  assign N199 = N71 & N130;
  assign N200 = N71 & tag_i[6];
  assign N201 = N73 & N130;
  assign N202 = N73 & tag_i[6];
  assign N203 = N75 & N130;
  assign N204 = N75 & tag_i[6];
  assign N205 = N77 & N130;
  assign N206 = N77 & tag_i[6];
  assign N207 = N79 & N130;
  assign N208 = N79 & tag_i[6];
  assign N209 = N81 & N130;
  assign N210 = N81 & tag_i[6];
  assign N211 = N83 & N130;
  assign N212 = N83 & tag_i[6];
  assign N213 = N85 & N130;
  assign N214 = N85 & tag_i[6];
  assign N215 = N87 & N130;
  assign N216 = N87 & tag_i[6];
  assign N217 = N89 & N130;
  assign N218 = N89 & tag_i[6];
  assign N219 = N91 & N130;
  assign N220 = N91 & tag_i[6];
  assign N221 = N93 & N130;
  assign N222 = N93 & tag_i[6];
  assign N223 = N95 & N130;
  assign N224 = N95 & tag_i[6];
  assign N225 = N97 & N130;
  assign N226 = N97 & tag_i[6];
  assign N227 = N99 & N130;
  assign N228 = N99 & tag_i[6];
  assign N229 = N101 & N130;
  assign N230 = N101 & tag_i[6];
  assign N231 = N103 & N130;
  assign N232 = N103 & tag_i[6];
  assign N233 = N105 & N130;
  assign N234 = N105 & tag_i[6];
  assign N235 = N107 & N130;
  assign N236 = N107 & tag_i[6];
  assign N237 = N109 & N130;
  assign N238 = N109 & tag_i[6];
  assign N239 = N111 & N130;
  assign N240 = N111 & tag_i[6];
  assign N241 = N113 & N130;
  assign N242 = N113 & tag_i[6];
  assign N243 = N115 & N130;
  assign N244 = N115 & tag_i[6];
  assign N245 = N117 & N130;
  assign N246 = N117 & tag_i[6];
  assign N247 = N119 & N130;
  assign N248 = N119 & tag_i[6];
  assign N249 = N121 & N130;
  assign N250 = N121 & tag_i[6];
  assign N251 = N123 & N130;
  assign N252 = N123 & tag_i[6];
  assign N253 = N125 & N130;
  assign N254 = N125 & tag_i[6];
  assign N255 = N127 & N130;
  assign N256 = N127 & tag_i[6];
  assign N257 = N129 & N130;
  assign N258 = N129 & tag_i[6];
  assign yumi_o = N259 & v_i;

endmodule

