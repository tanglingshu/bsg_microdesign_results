

module top
(
  lru_i,
  way_id_o
);

  input [62:0] lru_i;
  output [5:0] way_id_o;

  bsg_lru_pseudo_tree_encode
  wrapper
  (
    .lru_i(lru_i),
    .way_id_o(way_id_o)
  );


endmodule



module bsg_lru_pseudo_tree_encode
(
  lru_i,
  way_id_o
);

  input [62:0] lru_i;
  output [5:0] way_id_o;
  wire [5:0] way_id_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
  N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,
  N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,
  N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,
  N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,
  N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,
  N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,
  N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,
  N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,
  N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,
  N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,
  N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,
  N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,
  N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,
  N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,
  N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,
  N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,
  N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
  N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,
  N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,
  N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,
  N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,
  N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,
  N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,
  N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,
  N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,
  N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,
  N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,
  N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,
  N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,
  N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,
  N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,
  N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,
  N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,
  N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,
  N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,
  N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,
  N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,
  N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,
  N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,
  N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,
  N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,
  N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,
  N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,
  N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,
  N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,
  N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,
  N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,
  N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,
  N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,
  N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,
  N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,
  N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,
  N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,
  N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,
  N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,
  N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,
  N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,
  N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,
  N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,
  N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,
  N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,
  N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,
  N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,
  N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,
  N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,
  N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,
  N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,
  N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,
  N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,
  N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,
  N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,
  N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,
  N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,
  N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,
  N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,
  N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,
  N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,
  N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,
  N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,
  N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,
  N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,
  N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,
  N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144,
  N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,
  N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,N2170,
  N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,N2184,
  N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197,
  N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,N2210,
  N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,N2224,
  N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,
  N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,
  N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,N2264,
  N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,
  N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290,
  N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302,N2303,N2304,
  N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,
  N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,
  N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,
  N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,
  N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2369,N2370,
  N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382,N2383,N2384,
  pe_o_5__5_,pe_o_5__4_,pe_o_5__3_,pe_o_5__2_,pe_o_5__1_,pe_o_5__0_,pe_o_4__5_,
  pe_o_4__4_,pe_o_4__3_,pe_o_4__2_,pe_o_4__1_,pe_o_4__0_,pe_o_3__5_,pe_o_3__4_,
  pe_o_3__3_,pe_o_3__2_,pe_o_3__1_,pe_o_3__0_,pe_o_2__5_,pe_o_2__4_,pe_o_2__3_,
  pe_o_2__2_,pe_o_2__1_,pe_o_2__0_,pe_o_1__5_,pe_o_1__4_,pe_o_1__3_,pe_o_1__2_,pe_o_1__1_,
  pe_o_1__0_,N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,N2394,N2395,
  N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407,N2408,N2409,
  N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422,
  N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2435,
  N2436,N2437,N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447,N2448,N2449,
  N2450,N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,N2460,N2461,N2462,
  N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,N2474,N2475,
  N2476,N2477,N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,N2488,N2489,
  N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,N2500,N2501,N2502,
  N2503,N2504,N2505,N2506,N2507,N2508,pe_i_5__62_,pe_i_5__61_,pe_i_5__60_,
  pe_i_5__59_,pe_i_5__58_,pe_i_5__57_,pe_i_5__56_,pe_i_5__55_,pe_i_5__54_,pe_i_5__53_,
  pe_i_5__52_,pe_i_5__51_,pe_i_5__50_,pe_i_5__49_,pe_i_5__48_,pe_i_5__47_,pe_i_5__46_,
  pe_i_5__45_,pe_i_5__44_,pe_i_5__43_,pe_i_5__42_,pe_i_5__41_,pe_i_5__40_,
  pe_i_5__39_,pe_i_5__38_,pe_i_5__37_,pe_i_5__36_,pe_i_5__35_,pe_i_5__34_,pe_i_5__33_,
  pe_i_5__32_,pe_i_5__31_,pe_i_5__30_,pe_i_5__29_,pe_i_5__28_,pe_i_5__27_,pe_i_5__26_,
  pe_i_5__25_,pe_i_5__24_,pe_i_5__23_,pe_i_5__22_,pe_i_5__21_,pe_i_5__20_,
  pe_i_5__19_,pe_i_5__18_,pe_i_5__17_,pe_i_5__16_,pe_i_5__15_,pe_i_5__14_,pe_i_5__13_,
  pe_i_5__12_,pe_i_5__11_,pe_i_5__10_,pe_i_5__9_,pe_i_5__8_,pe_i_5__7_,pe_i_5__6_,
  pe_i_5__5_,pe_i_5__4_,pe_i_5__3_,pe_i_5__2_,pe_i_5__1_,pe_i_5__0_,pe_i_4__62_,
  pe_i_4__61_,pe_i_4__60_,pe_i_4__59_,pe_i_4__58_,pe_i_4__57_,pe_i_4__56_,pe_i_4__55_,
  pe_i_4__54_,pe_i_4__53_,pe_i_4__52_,pe_i_4__51_,pe_i_4__50_,pe_i_4__49_,pe_i_4__48_,
  pe_i_4__47_,pe_i_4__46_,pe_i_4__45_,pe_i_4__44_,pe_i_4__43_,pe_i_4__42_,
  pe_i_4__41_,pe_i_4__40_,pe_i_4__39_,pe_i_4__38_,pe_i_4__37_,pe_i_4__36_,pe_i_4__35_,
  pe_i_4__34_,pe_i_4__33_,pe_i_4__32_,pe_i_4__31_,pe_i_4__30_,pe_i_4__29_,pe_i_4__28_,
  pe_i_4__27_,pe_i_4__26_,pe_i_4__25_,pe_i_4__24_,pe_i_4__23_,pe_i_4__22_,
  pe_i_4__21_,pe_i_4__20_,pe_i_4__19_,pe_i_4__18_,pe_i_4__17_,pe_i_4__16_,pe_i_4__15_,
  pe_i_4__14_,pe_i_4__13_,pe_i_4__12_,pe_i_4__11_,pe_i_4__10_,pe_i_4__9_,pe_i_4__8_,
  pe_i_4__7_,pe_i_4__6_,pe_i_4__5_,pe_i_4__4_,pe_i_4__3_,pe_i_4__2_,pe_i_4__1_,
  pe_i_4__0_,pe_i_3__62_,pe_i_3__61_,pe_i_3__60_,pe_i_3__59_,pe_i_3__58_,pe_i_3__57_,
  pe_i_3__56_,pe_i_3__55_,pe_i_3__54_,pe_i_3__53_,pe_i_3__52_,pe_i_3__51_,
  pe_i_3__50_,pe_i_3__49_,pe_i_3__48_,pe_i_3__47_,pe_i_3__46_,pe_i_3__45_,pe_i_3__44_,
  pe_i_3__43_,pe_i_3__42_,pe_i_3__41_,pe_i_3__40_,pe_i_3__39_,pe_i_3__38_,pe_i_3__37_,
  pe_i_3__36_,pe_i_3__35_,pe_i_3__34_,pe_i_3__33_,pe_i_3__32_,pe_i_3__31_,
  pe_i_3__30_,pe_i_3__29_,pe_i_3__28_,pe_i_3__27_,pe_i_3__26_,pe_i_3__25_,pe_i_3__24_,
  pe_i_3__23_,pe_i_3__22_,pe_i_3__21_,pe_i_3__20_,pe_i_3__19_,pe_i_3__18_,pe_i_3__17_,
  pe_i_3__16_,pe_i_3__15_,pe_i_3__14_,pe_i_3__13_,pe_i_3__12_,pe_i_3__11_,
  pe_i_3__10_,pe_i_3__9_,pe_i_3__8_,pe_i_3__7_,pe_i_3__6_,pe_i_3__5_,pe_i_3__4_,pe_i_3__3_,
  pe_i_3__2_,pe_i_3__1_,pe_i_3__0_,pe_i_2__62_,pe_i_2__61_,pe_i_2__60_,pe_i_2__59_,
  pe_i_2__58_,pe_i_2__57_,pe_i_2__56_,pe_i_2__55_,pe_i_2__54_,pe_i_2__53_,
  pe_i_2__52_,pe_i_2__51_,pe_i_2__50_,pe_i_2__49_,pe_i_2__48_,pe_i_2__47_,pe_i_2__46_,
  pe_i_2__45_,pe_i_2__44_,pe_i_2__43_,pe_i_2__42_,pe_i_2__41_,pe_i_2__40_,pe_i_2__39_,
  pe_i_2__38_,pe_i_2__37_,pe_i_2__36_,pe_i_2__35_,pe_i_2__34_,pe_i_2__33_,
  pe_i_2__32_,pe_i_2__31_,pe_i_2__30_,pe_i_2__29_,pe_i_2__28_,pe_i_2__27_,pe_i_2__26_,
  pe_i_2__25_,pe_i_2__24_,pe_i_2__23_,pe_i_2__22_,pe_i_2__21_,pe_i_2__20_,pe_i_2__19_,
  pe_i_2__18_,pe_i_2__17_,pe_i_2__16_,pe_i_2__15_,pe_i_2__14_,pe_i_2__13_,
  pe_i_2__12_,pe_i_2__11_,pe_i_2__10_,pe_i_2__9_,pe_i_2__8_,pe_i_2__7_,pe_i_2__6_,
  pe_i_2__5_,pe_i_2__4_,pe_i_2__3_,pe_i_2__2_,pe_i_2__1_,pe_i_2__0_,pe_i_1__62_,
  pe_i_1__61_,pe_i_1__60_,pe_i_1__59_,pe_i_1__58_,pe_i_1__57_,pe_i_1__56_,pe_i_1__55_,
  pe_i_1__54_,pe_i_1__53_,pe_i_1__52_,pe_i_1__51_,pe_i_1__50_,pe_i_1__49_,pe_i_1__48_,
  pe_i_1__47_,pe_i_1__46_,pe_i_1__45_,pe_i_1__44_,pe_i_1__43_,pe_i_1__42_,
  pe_i_1__41_,pe_i_1__40_,pe_i_1__39_,pe_i_1__38_,pe_i_1__37_,pe_i_1__36_,pe_i_1__35_,
  pe_i_1__34_,pe_i_1__33_,pe_i_1__32_,pe_i_1__31_,pe_i_1__30_,pe_i_1__29_,pe_i_1__28_,
  pe_i_1__27_,pe_i_1__26_,pe_i_1__25_,pe_i_1__24_,pe_i_1__23_,pe_i_1__22_,
  pe_i_1__21_,pe_i_1__20_,pe_i_1__19_,pe_i_1__18_,pe_i_1__17_,pe_i_1__16_,pe_i_1__15_,
  pe_i_1__14_,pe_i_1__13_,pe_i_1__12_,pe_i_1__11_,pe_i_1__10_,pe_i_1__9_,pe_i_1__8_,
  pe_i_1__7_,pe_i_1__6_,pe_i_1__5_,pe_i_1__4_,pe_i_1__3_,pe_i_1__2_,pe_i_1__1_,
  pe_i_1__0_,N2509,N2510,N2511,N2512,N2513,N2514,N2515,N2516,N2517,N2518,N2519,N2520,
  N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528,N2529,N2530,N2531,N2532,N2533,N2534,
  N2535,N2536,N2537,N2538,N2539,N2540,N2541,N2542,N2543,N2544,N2545,N2546,N2547,
  N2548,N2549,N2550,N2551,N2552,N2553,N2554,N2555,N2556,N2557,N2558,N2559,N2560,
  N2561,N2562,N2563,N2564,N2565,N2566,N2567,N2568,N2569,N2570,N2571,N2572,N2573,N2574,
  N2575,N2576,N2577,N2578,N2579,N2580,N2581,N2582,N2583,N2584,N2585,N2586,N2587,
  N2588,N2589,N2590,N2591,N2592,N2593,N2594,N2595,N2596,N2597,N2598,N2599,N2600,
  N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2614,
  N2615,N2616,N2617,N2618,N2619,N2620,N2621,N2622,N2623,N2624,N2625,N2626,N2627,
  N2628,N2629,N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2637,N2638,N2639,N2640,
  N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,N2649,N2650,N2651,N2652,N2653,N2654,
  N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662,N2663,N2664,N2665,N2666,N2667,
  N2668,N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,N2678,N2679,N2680,
  N2681,N2682,N2683,N2684,N2685,N2686,N2687,N2688,N2689,N2690,N2691,N2692,N2693,N2694,
  N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2704,N2705,N2706,N2707,
  N2708,N2709,N2710,N2711,N2712,N2713,N2714,N2715,N2716,N2717,N2718,N2719,N2720,
  N2721,N2722,N2723,N2724,N2725,N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,
  N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2747,
  N2748,N2749,N2750,N2751,N2752,N2753,N2754,N2755,N2756,N2757,N2758,N2759,N2760,
  N2761,N2762,N2763,N2764,N2765,N2766,N2767,N2768,N2769,N2770,N2771,N2772,N2773,N2774,
  N2775,N2776,N2777,N2778,N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,
  N2788,N2789,N2790,N2791,N2792,N2793,N2794,N2795,N2796,N2797,N2798,N2799,N2800,
  N2801,N2802,N2803,N2804,N2805,N2806,N2807,N2808,N2809,N2810,N2811,N2812,N2813,N2814,
  N2815,N2816,N2817,N2818,N2819,N2820,N2821,N2822,N2823,N2824,N2825,N2826,N2827,
  N2828,N2829,N2830,N2831,N2832,N2833,N2834,N2835,N2836,N2837,N2838,N2839,N2840,
  N2841,N2842,N2843,N2844,N2845,N2846,N2847,N2848,N2849,N2850,N2851,N2852,N2853,N2854,
  N2855,N2856,N2857,N2858,N2859,N2860,N2861,N2862,N2863,N2864,N2865,N2866,N2867,
  N2868,N2869,N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,
  N2881,N2882,N2883,N2884,N2885,N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2893,N2894,
  N2895,N2896,N2897,N2898,N2899,N2900,N2901,N2902,N2903,N2904,N2905,N2906,N2907,
  N2908,N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,N2917,N2918,N2919,N2920,
  N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,
  N2935,N2936,N2937,N2938,N2939,N2940,N2941,N2942,N2943,N2944,N2945,N2946,N2947,
  N2948,N2949,N2950,N2951,N2952,N2953,N2954,N2955,N2956,N2957,N2958,N2959,N2960,
  N2961,N2962,N2963,N2964,N2965,N2966,N2967,N2968,N2969,N2970,N2971,N2972,N2973,N2974,
  N2975,N2976,N2977,N2978,N2979,N2980,N2981,N2982,N2983,N2984,N2985,N2986,N2987,
  N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,
  N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,N3010,N3011,N3012,N3013,N3014,
  N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,
  N3028,N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,
  N3041,N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,N3050,N3051,N3052,N3053,N3054,
  N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3062,N3063,N3064,N3065,N3066,N3067,
  N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,N3076,N3077,N3078,N3079,N3080,
  N3081,N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,N3090,N3091,N3092,N3093,N3094,
  N3095,N3096,N3097,N3098,N3099,N3100,N3101,N3102,N3103,N3104,N3105,N3106;
  wire [62:1] mask;

  bsg_priority_encode
  rof2_1__fi3_pe
  (
    .i({ pe_i_1__62_, pe_i_1__61_, pe_i_1__60_, pe_i_1__59_, pe_i_1__58_, pe_i_1__57_, pe_i_1__56_, pe_i_1__55_, pe_i_1__54_, pe_i_1__53_, pe_i_1__52_, pe_i_1__51_, pe_i_1__50_, pe_i_1__49_, pe_i_1__48_, pe_i_1__47_, pe_i_1__46_, pe_i_1__45_, pe_i_1__44_, pe_i_1__43_, pe_i_1__42_, pe_i_1__41_, pe_i_1__40_, pe_i_1__39_, pe_i_1__38_, pe_i_1__37_, pe_i_1__36_, pe_i_1__35_, pe_i_1__34_, pe_i_1__33_, pe_i_1__32_, pe_i_1__31_, pe_i_1__30_, pe_i_1__29_, pe_i_1__28_, pe_i_1__27_, pe_i_1__26_, pe_i_1__25_, pe_i_1__24_, pe_i_1__23_, pe_i_1__22_, pe_i_1__21_, pe_i_1__20_, pe_i_1__19_, pe_i_1__18_, pe_i_1__17_, pe_i_1__16_, pe_i_1__15_, pe_i_1__14_, pe_i_1__13_, pe_i_1__12_, pe_i_1__11_, pe_i_1__10_, pe_i_1__9_, pe_i_1__8_, pe_i_1__7_, pe_i_1__6_, pe_i_1__5_, pe_i_1__4_, pe_i_1__3_, pe_i_1__2_, pe_i_1__1_, pe_i_1__0_ }),
    .addr_o({ pe_o_1__5_, pe_o_1__4_, pe_o_1__3_, pe_o_1__2_, pe_o_1__1_, pe_o_1__0_ })
  );

  assign { N2697, N2696, N2695, N2694, N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, N2668, N2667, N2666, N2665, N2664, N2663, N2662, N2661, N2660, N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << { pe_o_1__5_, pe_o_1__4_, pe_o_1__3_, pe_o_1__2_, pe_o_1__1_, pe_o_1__0_ };

  bsg_priority_encode
  rof2_2__fi3_pe
  (
    .i({ pe_i_2__62_, pe_i_2__61_, pe_i_2__60_, pe_i_2__59_, pe_i_2__58_, pe_i_2__57_, pe_i_2__56_, pe_i_2__55_, pe_i_2__54_, pe_i_2__53_, pe_i_2__52_, pe_i_2__51_, pe_i_2__50_, pe_i_2__49_, pe_i_2__48_, pe_i_2__47_, pe_i_2__46_, pe_i_2__45_, pe_i_2__44_, pe_i_2__43_, pe_i_2__42_, pe_i_2__41_, pe_i_2__40_, pe_i_2__39_, pe_i_2__38_, pe_i_2__37_, pe_i_2__36_, pe_i_2__35_, pe_i_2__34_, pe_i_2__33_, pe_i_2__32_, pe_i_2__31_, pe_i_2__30_, pe_i_2__29_, pe_i_2__28_, pe_i_2__27_, pe_i_2__26_, pe_i_2__25_, pe_i_2__24_, pe_i_2__23_, pe_i_2__22_, pe_i_2__21_, pe_i_2__20_, pe_i_2__19_, pe_i_2__18_, pe_i_2__17_, pe_i_2__16_, pe_i_2__15_, pe_i_2__14_, pe_i_2__13_, pe_i_2__12_, pe_i_2__11_, pe_i_2__10_, pe_i_2__9_, pe_i_2__8_, pe_i_2__7_, pe_i_2__6_, pe_i_2__5_, pe_i_2__4_, pe_i_2__3_, pe_i_2__2_, pe_i_2__1_, pe_i_2__0_ }),
    .addr_o({ pe_o_2__5_, pe_o_2__4_, pe_o_2__3_, pe_o_2__2_, pe_o_2__1_, pe_o_2__0_ })
  );

  assign { N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N2806, N2805, N2804, N2803, N2802, N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, N2778, N2777, N2776, N2775, N2774, N2773, N2772, N2771, N2770, N2769, N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << { pe_o_2__5_, pe_o_2__4_, pe_o_2__3_, pe_o_2__2_, pe_o_2__1_, pe_o_2__0_ };

  bsg_priority_encode
  rof2_3__fi3_pe
  (
    .i({ pe_i_3__62_, pe_i_3__61_, pe_i_3__60_, pe_i_3__59_, pe_i_3__58_, pe_i_3__57_, pe_i_3__56_, pe_i_3__55_, pe_i_3__54_, pe_i_3__53_, pe_i_3__52_, pe_i_3__51_, pe_i_3__50_, pe_i_3__49_, pe_i_3__48_, pe_i_3__47_, pe_i_3__46_, pe_i_3__45_, pe_i_3__44_, pe_i_3__43_, pe_i_3__42_, pe_i_3__41_, pe_i_3__40_, pe_i_3__39_, pe_i_3__38_, pe_i_3__37_, pe_i_3__36_, pe_i_3__35_, pe_i_3__34_, pe_i_3__33_, pe_i_3__32_, pe_i_3__31_, pe_i_3__30_, pe_i_3__29_, pe_i_3__28_, pe_i_3__27_, pe_i_3__26_, pe_i_3__25_, pe_i_3__24_, pe_i_3__23_, pe_i_3__22_, pe_i_3__21_, pe_i_3__20_, pe_i_3__19_, pe_i_3__18_, pe_i_3__17_, pe_i_3__16_, pe_i_3__15_, pe_i_3__14_, pe_i_3__13_, pe_i_3__12_, pe_i_3__11_, pe_i_3__10_, pe_i_3__9_, pe_i_3__8_, pe_i_3__7_, pe_i_3__6_, pe_i_3__5_, pe_i_3__4_, pe_i_3__3_, pe_i_3__2_, pe_i_3__1_, pe_i_3__0_ }),
    .addr_o({ pe_o_3__5_, pe_o_3__4_, pe_o_3__3_, pe_o_3__2_, pe_o_3__1_, pe_o_3__0_ })
  );

  assign { N2949, N2948, N2947, N2946, N2945, N2944, N2943, N2942, N2941, N2940, N2939, N2938, N2937, N2936, N2935, N2934, N2933, N2932, N2931, N2930, N2929, N2928, N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908, N2907, N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << { pe_o_3__5_, pe_o_3__4_, pe_o_3__3_, pe_o_3__2_, pe_o_3__1_, pe_o_3__0_ };

  bsg_priority_encode
  rof2_4__fi3_pe
  (
    .i({ pe_i_4__62_, pe_i_4__61_, pe_i_4__60_, pe_i_4__59_, pe_i_4__58_, pe_i_4__57_, pe_i_4__56_, pe_i_4__55_, pe_i_4__54_, pe_i_4__53_, pe_i_4__52_, pe_i_4__51_, pe_i_4__50_, pe_i_4__49_, pe_i_4__48_, pe_i_4__47_, pe_i_4__46_, pe_i_4__45_, pe_i_4__44_, pe_i_4__43_, pe_i_4__42_, pe_i_4__41_, pe_i_4__40_, pe_i_4__39_, pe_i_4__38_, pe_i_4__37_, pe_i_4__36_, pe_i_4__35_, pe_i_4__34_, pe_i_4__33_, pe_i_4__32_, pe_i_4__31_, pe_i_4__30_, pe_i_4__29_, pe_i_4__28_, pe_i_4__27_, pe_i_4__26_, pe_i_4__25_, pe_i_4__24_, pe_i_4__23_, pe_i_4__22_, pe_i_4__21_, pe_i_4__20_, pe_i_4__19_, pe_i_4__18_, pe_i_4__17_, pe_i_4__16_, pe_i_4__15_, pe_i_4__14_, pe_i_4__13_, pe_i_4__12_, pe_i_4__11_, pe_i_4__10_, pe_i_4__9_, pe_i_4__8_, pe_i_4__7_, pe_i_4__6_, pe_i_4__5_, pe_i_4__4_, pe_i_4__3_, pe_i_4__2_, pe_i_4__1_, pe_i_4__0_ }),
    .addr_o({ pe_o_4__5_, pe_o_4__4_, pe_o_4__3_, pe_o_4__2_, pe_o_4__1_, pe_o_4__0_ })
  );

  assign { N3075, N3074, N3073, N3072, N3071, N3070, N3069, N3068, N3067, N3066, N3065, N3064, N3063, N3062, N3061, N3060, N3059, N3058, N3057, N3056, N3055, N3054, N3053, N3052, N3051, N3050, N3049, N3048, N3047, N3046, N3045, N3044, N3043, N3042, N3041, N3040, N3039, N3038, N3037, N3036, N3035, N3034, N3033, N3032, N3031, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N3023, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N3015, N3014, N3013 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << { pe_o_4__5_, pe_o_4__4_, pe_o_4__3_, pe_o_4__2_, pe_o_4__1_, pe_o_4__0_ };

  bsg_priority_encode
  rof2_5__fi3_pe
  (
    .i({ pe_i_5__62_, pe_i_5__61_, pe_i_5__60_, pe_i_5__59_, pe_i_5__58_, pe_i_5__57_, pe_i_5__56_, pe_i_5__55_, pe_i_5__54_, pe_i_5__53_, pe_i_5__52_, pe_i_5__51_, pe_i_5__50_, pe_i_5__49_, pe_i_5__48_, pe_i_5__47_, pe_i_5__46_, pe_i_5__45_, pe_i_5__44_, pe_i_5__43_, pe_i_5__42_, pe_i_5__41_, pe_i_5__40_, pe_i_5__39_, pe_i_5__38_, pe_i_5__37_, pe_i_5__36_, pe_i_5__35_, pe_i_5__34_, pe_i_5__33_, pe_i_5__32_, pe_i_5__31_, pe_i_5__30_, pe_i_5__29_, pe_i_5__28_, pe_i_5__27_, pe_i_5__26_, pe_i_5__25_, pe_i_5__24_, pe_i_5__23_, pe_i_5__22_, pe_i_5__21_, pe_i_5__20_, pe_i_5__19_, pe_i_5__18_, pe_i_5__17_, pe_i_5__16_, pe_i_5__15_, pe_i_5__14_, pe_i_5__13_, pe_i_5__12_, pe_i_5__11_, pe_i_5__10_, pe_i_5__9_, pe_i_5__8_, pe_i_5__7_, pe_i_5__6_, pe_i_5__5_, pe_i_5__4_, pe_i_5__3_, pe_i_5__2_, pe_i_5__1_, pe_i_5__0_ }),
    .addr_o({ pe_o_5__5_, pe_o_5__4_, pe_o_5__3_, pe_o_5__2_, pe_o_5__1_, pe_o_5__0_ })
  );

  assign N0 = N4 & N5;
  assign N1 = N0 & N6;
  assign N2 = N1 & N7;
  assign N3 = N2 & N8;
  assign N2509 = N3 & N9;
  assign N4 = ~pe_o_1__5_;
  assign N5 = ~pe_o_1__4_;
  assign N6 = ~pe_o_1__3_;
  assign N7 = ~pe_o_1__2_;
  assign N8 = ~pe_o_1__0_;
  assign N9 = ~pe_o_1__1_;
  assign N10 = pe_o_1__5_ & N14;
  assign N11 = N10 & N15;
  assign N12 = N11 & N16;
  assign N13 = N12 & N17;
  assign N2510 = N13 & N18;
  assign N14 = ~pe_o_1__4_;
  assign N15 = ~pe_o_1__3_;
  assign N16 = ~pe_o_1__2_;
  assign N17 = ~pe_o_1__0_;
  assign N18 = ~pe_o_1__1_;
  assign N19 = N23 & N24;
  assign N20 = N19 & N25;
  assign N21 = N20 & N26;
  assign N22 = N21 & pe_o_1__0_;
  assign N2511 = N22 & N27;
  assign N23 = ~pe_o_1__5_;
  assign N24 = ~pe_o_1__4_;
  assign N25 = ~pe_o_1__3_;
  assign N26 = ~pe_o_1__2_;
  assign N27 = ~pe_o_1__1_;
  assign N28 = N32 & N33;
  assign N29 = N28 & N34;
  assign N30 = N29 & N35;
  assign N31 = N30 & N36;
  assign N2513 = N31 & pe_o_1__1_;
  assign N32 = ~pe_o_1__5_;
  assign N33 = ~pe_o_1__4_;
  assign N34 = ~pe_o_1__3_;
  assign N35 = ~pe_o_1__2_;
  assign N36 = ~pe_o_1__0_;
  assign N37 = N41 & N42;
  assign N38 = N37 & N43;
  assign N39 = N38 & N44;
  assign N40 = N39 & pe_o_1__0_;
  assign N2515 = N40 & pe_o_1__1_;
  assign N41 = ~pe_o_1__5_;
  assign N42 = ~pe_o_1__4_;
  assign N43 = ~pe_o_1__3_;
  assign N44 = ~pe_o_1__2_;
  assign N45 = N49 & N50;
  assign N46 = N45 & N51;
  assign N47 = N46 & pe_o_1__2_;
  assign N48 = N47 & N52;
  assign N2517 = N48 & N53;
  assign N49 = ~pe_o_1__5_;
  assign N50 = ~pe_o_1__4_;
  assign N51 = ~pe_o_1__3_;
  assign N52 = ~pe_o_1__0_;
  assign N53 = ~pe_o_1__1_;
  assign N54 = N58 & N59;
  assign N55 = N54 & N60;
  assign N56 = N55 & pe_o_1__2_;
  assign N57 = N56 & pe_o_1__0_;
  assign N2519 = N57 & N61;
  assign N58 = ~pe_o_1__5_;
  assign N59 = ~pe_o_1__4_;
  assign N60 = ~pe_o_1__3_;
  assign N61 = ~pe_o_1__1_;
  assign N62 = N66 & N67;
  assign N63 = N62 & N68;
  assign N64 = N63 & pe_o_1__2_;
  assign N65 = N64 & N69;
  assign N2521 = N65 & pe_o_1__1_;
  assign N66 = ~pe_o_1__5_;
  assign N67 = ~pe_o_1__4_;
  assign N68 = ~pe_o_1__3_;
  assign N69 = ~pe_o_1__0_;
  assign N70 = N74 & N75;
  assign N71 = N70 & N76;
  assign N72 = N71 & pe_o_1__2_;
  assign N73 = N72 & pe_o_1__0_;
  assign N2523 = N73 & pe_o_1__1_;
  assign N74 = ~pe_o_1__5_;
  assign N75 = ~pe_o_1__4_;
  assign N76 = ~pe_o_1__3_;
  assign N77 = N81 & N82;
  assign N78 = N77 & pe_o_1__3_;
  assign N79 = N78 & N83;
  assign N80 = N79 & N84;
  assign N2525 = N80 & N85;
  assign N81 = ~pe_o_1__5_;
  assign N82 = ~pe_o_1__4_;
  assign N83 = ~pe_o_1__2_;
  assign N84 = ~pe_o_1__0_;
  assign N85 = ~pe_o_1__1_;
  assign N86 = N90 & N91;
  assign N87 = N86 & pe_o_1__3_;
  assign N88 = N87 & N92;
  assign N89 = N88 & pe_o_1__0_;
  assign N2527 = N89 & N93;
  assign N90 = ~pe_o_1__5_;
  assign N91 = ~pe_o_1__4_;
  assign N92 = ~pe_o_1__2_;
  assign N93 = ~pe_o_1__1_;
  assign N94 = N98 & N99;
  assign N95 = N94 & pe_o_1__3_;
  assign N96 = N95 & N100;
  assign N97 = N96 & N101;
  assign N2529 = N97 & pe_o_1__1_;
  assign N98 = ~pe_o_1__5_;
  assign N99 = ~pe_o_1__4_;
  assign N100 = ~pe_o_1__2_;
  assign N101 = ~pe_o_1__0_;
  assign N102 = N106 & N107;
  assign N103 = N102 & pe_o_1__3_;
  assign N104 = N103 & N108;
  assign N105 = N104 & pe_o_1__0_;
  assign N2531 = N105 & pe_o_1__1_;
  assign N106 = ~pe_o_1__5_;
  assign N107 = ~pe_o_1__4_;
  assign N108 = ~pe_o_1__2_;
  assign N109 = N113 & N114;
  assign N110 = N109 & pe_o_1__3_;
  assign N111 = N110 & pe_o_1__2_;
  assign N112 = N111 & N115;
  assign N2533 = N112 & N116;
  assign N113 = ~pe_o_1__5_;
  assign N114 = ~pe_o_1__4_;
  assign N115 = ~pe_o_1__0_;
  assign N116 = ~pe_o_1__1_;
  assign N117 = N121 & N122;
  assign N118 = N117 & pe_o_1__3_;
  assign N119 = N118 & pe_o_1__2_;
  assign N120 = N119 & pe_o_1__0_;
  assign N2535 = N120 & N123;
  assign N121 = ~pe_o_1__5_;
  assign N122 = ~pe_o_1__4_;
  assign N123 = ~pe_o_1__1_;
  assign N124 = N128 & N129;
  assign N125 = N124 & pe_o_1__3_;
  assign N126 = N125 & pe_o_1__2_;
  assign N127 = N126 & N130;
  assign N2537 = N127 & pe_o_1__1_;
  assign N128 = ~pe_o_1__5_;
  assign N129 = ~pe_o_1__4_;
  assign N130 = ~pe_o_1__0_;
  assign N131 = N135 & N136;
  assign N132 = N131 & pe_o_1__3_;
  assign N133 = N132 & pe_o_1__2_;
  assign N134 = N133 & pe_o_1__0_;
  assign N2539 = N134 & pe_o_1__1_;
  assign N135 = ~pe_o_1__5_;
  assign N136 = ~pe_o_1__4_;
  assign N137 = N141 & pe_o_1__4_;
  assign N138 = N137 & N142;
  assign N139 = N138 & N143;
  assign N140 = N139 & N144;
  assign N2541 = N140 & N145;
  assign N141 = ~pe_o_1__5_;
  assign N142 = ~pe_o_1__3_;
  assign N143 = ~pe_o_1__2_;
  assign N144 = ~pe_o_1__0_;
  assign N145 = ~pe_o_1__1_;
  assign N146 = N150 & pe_o_1__4_;
  assign N147 = N146 & N151;
  assign N148 = N147 & N152;
  assign N149 = N148 & pe_o_1__0_;
  assign N2543 = N149 & N153;
  assign N150 = ~pe_o_1__5_;
  assign N151 = ~pe_o_1__3_;
  assign N152 = ~pe_o_1__2_;
  assign N153 = ~pe_o_1__1_;
  assign N154 = N158 & pe_o_1__4_;
  assign N155 = N154 & N159;
  assign N156 = N155 & N160;
  assign N157 = N156 & N161;
  assign N2545 = N157 & pe_o_1__1_;
  assign N158 = ~pe_o_1__5_;
  assign N159 = ~pe_o_1__3_;
  assign N160 = ~pe_o_1__2_;
  assign N161 = ~pe_o_1__0_;
  assign N162 = N166 & pe_o_1__4_;
  assign N163 = N162 & N167;
  assign N164 = N163 & N168;
  assign N165 = N164 & pe_o_1__0_;
  assign N2547 = N165 & pe_o_1__1_;
  assign N166 = ~pe_o_1__5_;
  assign N167 = ~pe_o_1__3_;
  assign N168 = ~pe_o_1__2_;
  assign N169 = N173 & pe_o_1__4_;
  assign N170 = N169 & N174;
  assign N171 = N170 & pe_o_1__2_;
  assign N172 = N171 & N175;
  assign N2549 = N172 & N176;
  assign N173 = ~pe_o_1__5_;
  assign N174 = ~pe_o_1__3_;
  assign N175 = ~pe_o_1__0_;
  assign N176 = ~pe_o_1__1_;
  assign N177 = N181 & pe_o_1__4_;
  assign N178 = N177 & N182;
  assign N179 = N178 & pe_o_1__2_;
  assign N180 = N179 & pe_o_1__0_;
  assign N2551 = N180 & N183;
  assign N181 = ~pe_o_1__5_;
  assign N182 = ~pe_o_1__3_;
  assign N183 = ~pe_o_1__1_;
  assign N184 = N188 & pe_o_1__4_;
  assign N185 = N184 & N189;
  assign N186 = N185 & pe_o_1__2_;
  assign N187 = N186 & N190;
  assign N2553 = N187 & pe_o_1__1_;
  assign N188 = ~pe_o_1__5_;
  assign N189 = ~pe_o_1__3_;
  assign N190 = ~pe_o_1__0_;
  assign N191 = N195 & pe_o_1__4_;
  assign N192 = N191 & N196;
  assign N193 = N192 & pe_o_1__2_;
  assign N194 = N193 & pe_o_1__0_;
  assign N2555 = N194 & pe_o_1__1_;
  assign N195 = ~pe_o_1__5_;
  assign N196 = ~pe_o_1__3_;
  assign N197 = N201 & pe_o_1__4_;
  assign N198 = N197 & pe_o_1__3_;
  assign N199 = N198 & N202;
  assign N200 = N199 & N203;
  assign N2557 = N200 & N204;
  assign N201 = ~pe_o_1__5_;
  assign N202 = ~pe_o_1__2_;
  assign N203 = ~pe_o_1__0_;
  assign N204 = ~pe_o_1__1_;
  assign N205 = N209 & pe_o_1__4_;
  assign N206 = N205 & pe_o_1__3_;
  assign N207 = N206 & N210;
  assign N208 = N207 & pe_o_1__0_;
  assign N2559 = N208 & N211;
  assign N209 = ~pe_o_1__5_;
  assign N210 = ~pe_o_1__2_;
  assign N211 = ~pe_o_1__1_;
  assign N212 = N216 & pe_o_1__4_;
  assign N213 = N212 & pe_o_1__3_;
  assign N214 = N213 & N217;
  assign N215 = N214 & N218;
  assign N2561 = N215 & pe_o_1__1_;
  assign N216 = ~pe_o_1__5_;
  assign N217 = ~pe_o_1__2_;
  assign N218 = ~pe_o_1__0_;
  assign N219 = N223 & pe_o_1__4_;
  assign N220 = N219 & pe_o_1__3_;
  assign N221 = N220 & N224;
  assign N222 = N221 & pe_o_1__0_;
  assign N2563 = N222 & pe_o_1__1_;
  assign N223 = ~pe_o_1__5_;
  assign N224 = ~pe_o_1__2_;
  assign N225 = N229 & pe_o_1__4_;
  assign N226 = N225 & pe_o_1__3_;
  assign N227 = N226 & pe_o_1__2_;
  assign N228 = N227 & N230;
  assign N2565 = N228 & N231;
  assign N229 = ~pe_o_1__5_;
  assign N230 = ~pe_o_1__0_;
  assign N231 = ~pe_o_1__1_;
  assign N232 = N236 & pe_o_1__4_;
  assign N233 = N232 & pe_o_1__3_;
  assign N234 = N233 & pe_o_1__2_;
  assign N235 = N234 & pe_o_1__0_;
  assign N2567 = N235 & N237;
  assign N236 = ~pe_o_1__5_;
  assign N237 = ~pe_o_1__1_;
  assign N238 = N242 & pe_o_1__4_;
  assign N239 = N238 & pe_o_1__3_;
  assign N240 = N239 & pe_o_1__2_;
  assign N241 = N240 & N243;
  assign N2569 = N241 & pe_o_1__1_;
  assign N242 = ~pe_o_1__5_;
  assign N243 = ~pe_o_1__0_;
  assign N2571 = pe_o_1__4_ & pe_o_1__3_ & (pe_o_1__2_ & pe_o_1__0_) & pe_o_1__1_;
  assign N244 = pe_o_1__5_ & N248;
  assign N245 = N244 & N249;
  assign N246 = N245 & N250;
  assign N247 = N246 & pe_o_1__0_;
  assign N2512 = N247 & N251;
  assign N248 = ~pe_o_1__4_;
  assign N249 = ~pe_o_1__3_;
  assign N250 = ~pe_o_1__2_;
  assign N251 = ~pe_o_1__1_;
  assign N252 = pe_o_1__5_ & N256;
  assign N253 = N252 & N257;
  assign N254 = N253 & N258;
  assign N255 = N254 & N259;
  assign N2514 = N255 & pe_o_1__1_;
  assign N256 = ~pe_o_1__4_;
  assign N257 = ~pe_o_1__3_;
  assign N258 = ~pe_o_1__2_;
  assign N259 = ~pe_o_1__0_;
  assign N260 = pe_o_1__5_ & N264;
  assign N261 = N260 & N265;
  assign N262 = N261 & N266;
  assign N263 = N262 & pe_o_1__0_;
  assign N2516 = N263 & pe_o_1__1_;
  assign N264 = ~pe_o_1__4_;
  assign N265 = ~pe_o_1__3_;
  assign N266 = ~pe_o_1__2_;
  assign N267 = pe_o_1__5_ & N271;
  assign N268 = N267 & N272;
  assign N269 = N268 & pe_o_1__2_;
  assign N270 = N269 & N273;
  assign N2518 = N270 & N274;
  assign N271 = ~pe_o_1__4_;
  assign N272 = ~pe_o_1__3_;
  assign N273 = ~pe_o_1__0_;
  assign N274 = ~pe_o_1__1_;
  assign N275 = pe_o_1__5_ & N279;
  assign N276 = N275 & N280;
  assign N277 = N276 & pe_o_1__2_;
  assign N278 = N277 & pe_o_1__0_;
  assign N2520 = N278 & N281;
  assign N279 = ~pe_o_1__4_;
  assign N280 = ~pe_o_1__3_;
  assign N281 = ~pe_o_1__1_;
  assign N282 = pe_o_1__5_ & N286;
  assign N283 = N282 & N287;
  assign N284 = N283 & pe_o_1__2_;
  assign N285 = N284 & N288;
  assign N2522 = N285 & pe_o_1__1_;
  assign N286 = ~pe_o_1__4_;
  assign N287 = ~pe_o_1__3_;
  assign N288 = ~pe_o_1__0_;
  assign N289 = pe_o_1__5_ & N293;
  assign N290 = N289 & N294;
  assign N291 = N290 & pe_o_1__2_;
  assign N292 = N291 & pe_o_1__0_;
  assign N2524 = N292 & pe_o_1__1_;
  assign N293 = ~pe_o_1__4_;
  assign N294 = ~pe_o_1__3_;
  assign N295 = pe_o_1__5_ & N299;
  assign N296 = N295 & pe_o_1__3_;
  assign N297 = N296 & N300;
  assign N298 = N297 & N301;
  assign N2526 = N298 & N302;
  assign N299 = ~pe_o_1__4_;
  assign N300 = ~pe_o_1__2_;
  assign N301 = ~pe_o_1__0_;
  assign N302 = ~pe_o_1__1_;
  assign N303 = pe_o_1__5_ & N307;
  assign N304 = N303 & pe_o_1__3_;
  assign N305 = N304 & N308;
  assign N306 = N305 & pe_o_1__0_;
  assign N2528 = N306 & N309;
  assign N307 = ~pe_o_1__4_;
  assign N308 = ~pe_o_1__2_;
  assign N309 = ~pe_o_1__1_;
  assign N310 = pe_o_1__5_ & N314;
  assign N311 = N310 & pe_o_1__3_;
  assign N312 = N311 & N315;
  assign N313 = N312 & N316;
  assign N2530 = N313 & pe_o_1__1_;
  assign N314 = ~pe_o_1__4_;
  assign N315 = ~pe_o_1__2_;
  assign N316 = ~pe_o_1__0_;
  assign N317 = pe_o_1__5_ & N321;
  assign N318 = N317 & pe_o_1__3_;
  assign N319 = N318 & N322;
  assign N320 = N319 & pe_o_1__0_;
  assign N2532 = N320 & pe_o_1__1_;
  assign N321 = ~pe_o_1__4_;
  assign N322 = ~pe_o_1__2_;
  assign N323 = pe_o_1__5_ & N327;
  assign N324 = N323 & pe_o_1__3_;
  assign N325 = N324 & pe_o_1__2_;
  assign N326 = N325 & N328;
  assign N2534 = N326 & N329;
  assign N327 = ~pe_o_1__4_;
  assign N328 = ~pe_o_1__0_;
  assign N329 = ~pe_o_1__1_;
  assign N330 = pe_o_1__5_ & N334;
  assign N331 = N330 & pe_o_1__3_;
  assign N332 = N331 & pe_o_1__2_;
  assign N333 = N332 & pe_o_1__0_;
  assign N2536 = N333 & N335;
  assign N334 = ~pe_o_1__4_;
  assign N335 = ~pe_o_1__1_;
  assign N336 = pe_o_1__5_ & N340;
  assign N337 = N336 & pe_o_1__3_;
  assign N338 = N337 & pe_o_1__2_;
  assign N339 = N338 & N341;
  assign N2538 = N339 & pe_o_1__1_;
  assign N340 = ~pe_o_1__4_;
  assign N341 = ~pe_o_1__0_;
  assign N2540 = pe_o_1__5_ & pe_o_1__3_ & (pe_o_1__2_ & pe_o_1__0_) & pe_o_1__1_;
  assign N342 = pe_o_1__5_ & pe_o_1__4_;
  assign N343 = N342 & N346;
  assign N344 = N343 & N347;
  assign N345 = N344 & N348;
  assign N2542 = N345 & N349;
  assign N346 = ~pe_o_1__3_;
  assign N347 = ~pe_o_1__2_;
  assign N348 = ~pe_o_1__0_;
  assign N349 = ~pe_o_1__1_;
  assign N350 = pe_o_1__5_ & pe_o_1__4_;
  assign N351 = N350 & N354;
  assign N352 = N351 & N355;
  assign N353 = N352 & pe_o_1__0_;
  assign N2544 = N353 & N356;
  assign N354 = ~pe_o_1__3_;
  assign N355 = ~pe_o_1__2_;
  assign N356 = ~pe_o_1__1_;
  assign N357 = pe_o_1__5_ & pe_o_1__4_;
  assign N358 = N357 & N361;
  assign N359 = N358 & N362;
  assign N360 = N359 & N363;
  assign N2546 = N360 & pe_o_1__1_;
  assign N361 = ~pe_o_1__3_;
  assign N362 = ~pe_o_1__2_;
  assign N363 = ~pe_o_1__0_;
  assign N364 = pe_o_1__5_ & pe_o_1__4_;
  assign N365 = N364 & N368;
  assign N366 = N365 & N369;
  assign N367 = N366 & pe_o_1__0_;
  assign N2548 = N367 & pe_o_1__1_;
  assign N368 = ~pe_o_1__3_;
  assign N369 = ~pe_o_1__2_;
  assign N370 = pe_o_1__5_ & pe_o_1__4_;
  assign N371 = N370 & N374;
  assign N372 = N371 & pe_o_1__2_;
  assign N373 = N372 & N375;
  assign N2550 = N373 & N376;
  assign N374 = ~pe_o_1__3_;
  assign N375 = ~pe_o_1__0_;
  assign N376 = ~pe_o_1__1_;
  assign N377 = pe_o_1__5_ & pe_o_1__4_;
  assign N378 = N377 & N381;
  assign N379 = N378 & pe_o_1__2_;
  assign N380 = N379 & pe_o_1__0_;
  assign N2552 = N380 & N382;
  assign N381 = ~pe_o_1__3_;
  assign N382 = ~pe_o_1__1_;
  assign N383 = pe_o_1__5_ & pe_o_1__4_;
  assign N384 = N383 & N387;
  assign N385 = N384 & pe_o_1__2_;
  assign N386 = N385 & N388;
  assign N2554 = N386 & pe_o_1__1_;
  assign N387 = ~pe_o_1__3_;
  assign N388 = ~pe_o_1__0_;
  assign N2556 = pe_o_1__5_ & pe_o_1__4_ & (pe_o_1__2_ & pe_o_1__0_) & pe_o_1__1_;
  assign N389 = pe_o_1__5_ & pe_o_1__4_;
  assign N390 = N389 & pe_o_1__3_;
  assign N391 = N390 & N393;
  assign N392 = N391 & N394;
  assign N2558 = N392 & N395;
  assign N393 = ~pe_o_1__2_;
  assign N394 = ~pe_o_1__0_;
  assign N395 = ~pe_o_1__1_;
  assign N396 = pe_o_1__5_ & pe_o_1__4_;
  assign N397 = N396 & pe_o_1__3_;
  assign N398 = N397 & N400;
  assign N399 = N398 & pe_o_1__0_;
  assign N2560 = N399 & N401;
  assign N400 = ~pe_o_1__2_;
  assign N401 = ~pe_o_1__1_;
  assign N402 = pe_o_1__5_ & pe_o_1__4_;
  assign N403 = N402 & pe_o_1__3_;
  assign N404 = N403 & N406;
  assign N405 = N404 & N407;
  assign N2562 = N405 & pe_o_1__1_;
  assign N406 = ~pe_o_1__2_;
  assign N407 = ~pe_o_1__0_;
  assign N2564 = pe_o_1__5_ & pe_o_1__4_ & (pe_o_1__3_ & pe_o_1__0_) & pe_o_1__1_;
  assign N408 = pe_o_1__5_ & pe_o_1__4_;
  assign N409 = N408 & pe_o_1__3_;
  assign N410 = N409 & pe_o_1__2_;
  assign N411 = N410 & N412;
  assign N2566 = N411 & N413;
  assign N412 = ~pe_o_1__0_;
  assign N413 = ~pe_o_1__1_;
  assign N2568 = pe_o_1__5_ & pe_o_1__4_ & (pe_o_1__3_ & pe_o_1__2_) & pe_o_1__0_;
  assign N2570 = pe_o_1__5_ & pe_o_1__4_ & (pe_o_1__3_ & pe_o_1__2_) & pe_o_1__1_;
  assign N414 = N418 & N419;
  assign N415 = N414 & N420;
  assign N416 = N415 & N421;
  assign N417 = N416 & N422;
  assign N2572 = N417 & N423;
  assign N418 = ~pe_o_2__5_;
  assign N419 = ~pe_o_2__4_;
  assign N420 = ~pe_o_2__3_;
  assign N421 = ~pe_o_2__2_;
  assign N422 = ~pe_o_2__0_;
  assign N423 = ~pe_o_2__1_;
  assign N424 = pe_o_2__5_ & N428;
  assign N425 = N424 & N429;
  assign N426 = N425 & N430;
  assign N427 = N426 & N431;
  assign N2573 = N427 & N432;
  assign N428 = ~pe_o_2__4_;
  assign N429 = ~pe_o_2__3_;
  assign N430 = ~pe_o_2__2_;
  assign N431 = ~pe_o_2__0_;
  assign N432 = ~pe_o_2__1_;
  assign N433 = N437 & N438;
  assign N434 = N433 & N439;
  assign N435 = N434 & N440;
  assign N436 = N435 & pe_o_2__0_;
  assign N2574 = N436 & N441;
  assign N437 = ~pe_o_2__5_;
  assign N438 = ~pe_o_2__4_;
  assign N439 = ~pe_o_2__3_;
  assign N440 = ~pe_o_2__2_;
  assign N441 = ~pe_o_2__1_;
  assign N442 = N446 & N447;
  assign N443 = N442 & N448;
  assign N444 = N443 & N449;
  assign N445 = N444 & N450;
  assign N2576 = N445 & pe_o_2__1_;
  assign N446 = ~pe_o_2__5_;
  assign N447 = ~pe_o_2__4_;
  assign N448 = ~pe_o_2__3_;
  assign N449 = ~pe_o_2__2_;
  assign N450 = ~pe_o_2__0_;
  assign N451 = N455 & N456;
  assign N452 = N451 & N457;
  assign N453 = N452 & N458;
  assign N454 = N453 & pe_o_2__0_;
  assign N2578 = N454 & pe_o_2__1_;
  assign N455 = ~pe_o_2__5_;
  assign N456 = ~pe_o_2__4_;
  assign N457 = ~pe_o_2__3_;
  assign N458 = ~pe_o_2__2_;
  assign N459 = N463 & N464;
  assign N460 = N459 & N465;
  assign N461 = N460 & pe_o_2__2_;
  assign N462 = N461 & N466;
  assign N2580 = N462 & N467;
  assign N463 = ~pe_o_2__5_;
  assign N464 = ~pe_o_2__4_;
  assign N465 = ~pe_o_2__3_;
  assign N466 = ~pe_o_2__0_;
  assign N467 = ~pe_o_2__1_;
  assign N468 = N472 & N473;
  assign N469 = N468 & N474;
  assign N470 = N469 & pe_o_2__2_;
  assign N471 = N470 & pe_o_2__0_;
  assign N2582 = N471 & N475;
  assign N472 = ~pe_o_2__5_;
  assign N473 = ~pe_o_2__4_;
  assign N474 = ~pe_o_2__3_;
  assign N475 = ~pe_o_2__1_;
  assign N476 = N480 & N481;
  assign N477 = N476 & N482;
  assign N478 = N477 & pe_o_2__2_;
  assign N479 = N478 & N483;
  assign N2584 = N479 & pe_o_2__1_;
  assign N480 = ~pe_o_2__5_;
  assign N481 = ~pe_o_2__4_;
  assign N482 = ~pe_o_2__3_;
  assign N483 = ~pe_o_2__0_;
  assign N484 = N488 & N489;
  assign N485 = N484 & N490;
  assign N486 = N485 & pe_o_2__2_;
  assign N487 = N486 & pe_o_2__0_;
  assign N2586 = N487 & pe_o_2__1_;
  assign N488 = ~pe_o_2__5_;
  assign N489 = ~pe_o_2__4_;
  assign N490 = ~pe_o_2__3_;
  assign N491 = N495 & N496;
  assign N492 = N491 & pe_o_2__3_;
  assign N493 = N492 & N497;
  assign N494 = N493 & N498;
  assign N2588 = N494 & N499;
  assign N495 = ~pe_o_2__5_;
  assign N496 = ~pe_o_2__4_;
  assign N497 = ~pe_o_2__2_;
  assign N498 = ~pe_o_2__0_;
  assign N499 = ~pe_o_2__1_;
  assign N500 = N504 & N505;
  assign N501 = N500 & pe_o_2__3_;
  assign N502 = N501 & N506;
  assign N503 = N502 & pe_o_2__0_;
  assign N2590 = N503 & N507;
  assign N504 = ~pe_o_2__5_;
  assign N505 = ~pe_o_2__4_;
  assign N506 = ~pe_o_2__2_;
  assign N507 = ~pe_o_2__1_;
  assign N508 = N512 & N513;
  assign N509 = N508 & pe_o_2__3_;
  assign N510 = N509 & N514;
  assign N511 = N510 & N515;
  assign N2592 = N511 & pe_o_2__1_;
  assign N512 = ~pe_o_2__5_;
  assign N513 = ~pe_o_2__4_;
  assign N514 = ~pe_o_2__2_;
  assign N515 = ~pe_o_2__0_;
  assign N516 = N520 & N521;
  assign N517 = N516 & pe_o_2__3_;
  assign N518 = N517 & N522;
  assign N519 = N518 & pe_o_2__0_;
  assign N2594 = N519 & pe_o_2__1_;
  assign N520 = ~pe_o_2__5_;
  assign N521 = ~pe_o_2__4_;
  assign N522 = ~pe_o_2__2_;
  assign N523 = N527 & N528;
  assign N524 = N523 & pe_o_2__3_;
  assign N525 = N524 & pe_o_2__2_;
  assign N526 = N525 & N529;
  assign N2596 = N526 & N530;
  assign N527 = ~pe_o_2__5_;
  assign N528 = ~pe_o_2__4_;
  assign N529 = ~pe_o_2__0_;
  assign N530 = ~pe_o_2__1_;
  assign N531 = N535 & N536;
  assign N532 = N531 & pe_o_2__3_;
  assign N533 = N532 & pe_o_2__2_;
  assign N534 = N533 & pe_o_2__0_;
  assign N2598 = N534 & N537;
  assign N535 = ~pe_o_2__5_;
  assign N536 = ~pe_o_2__4_;
  assign N537 = ~pe_o_2__1_;
  assign N538 = N542 & N543;
  assign N539 = N538 & pe_o_2__3_;
  assign N540 = N539 & pe_o_2__2_;
  assign N541 = N540 & N544;
  assign N2600 = N541 & pe_o_2__1_;
  assign N542 = ~pe_o_2__5_;
  assign N543 = ~pe_o_2__4_;
  assign N544 = ~pe_o_2__0_;
  assign N545 = N549 & N550;
  assign N546 = N545 & pe_o_2__3_;
  assign N547 = N546 & pe_o_2__2_;
  assign N548 = N547 & pe_o_2__0_;
  assign N2602 = N548 & pe_o_2__1_;
  assign N549 = ~pe_o_2__5_;
  assign N550 = ~pe_o_2__4_;
  assign N551 = N555 & pe_o_2__4_;
  assign N552 = N551 & N556;
  assign N553 = N552 & N557;
  assign N554 = N553 & N558;
  assign N2604 = N554 & N559;
  assign N555 = ~pe_o_2__5_;
  assign N556 = ~pe_o_2__3_;
  assign N557 = ~pe_o_2__2_;
  assign N558 = ~pe_o_2__0_;
  assign N559 = ~pe_o_2__1_;
  assign N560 = N564 & pe_o_2__4_;
  assign N561 = N560 & N565;
  assign N562 = N561 & N566;
  assign N563 = N562 & pe_o_2__0_;
  assign N2606 = N563 & N567;
  assign N564 = ~pe_o_2__5_;
  assign N565 = ~pe_o_2__3_;
  assign N566 = ~pe_o_2__2_;
  assign N567 = ~pe_o_2__1_;
  assign N568 = N572 & pe_o_2__4_;
  assign N569 = N568 & N573;
  assign N570 = N569 & N574;
  assign N571 = N570 & N575;
  assign N2608 = N571 & pe_o_2__1_;
  assign N572 = ~pe_o_2__5_;
  assign N573 = ~pe_o_2__3_;
  assign N574 = ~pe_o_2__2_;
  assign N575 = ~pe_o_2__0_;
  assign N576 = N580 & pe_o_2__4_;
  assign N577 = N576 & N581;
  assign N578 = N577 & N582;
  assign N579 = N578 & pe_o_2__0_;
  assign N2610 = N579 & pe_o_2__1_;
  assign N580 = ~pe_o_2__5_;
  assign N581 = ~pe_o_2__3_;
  assign N582 = ~pe_o_2__2_;
  assign N583 = N587 & pe_o_2__4_;
  assign N584 = N583 & N588;
  assign N585 = N584 & pe_o_2__2_;
  assign N586 = N585 & N589;
  assign N2612 = N586 & N590;
  assign N587 = ~pe_o_2__5_;
  assign N588 = ~pe_o_2__3_;
  assign N589 = ~pe_o_2__0_;
  assign N590 = ~pe_o_2__1_;
  assign N591 = N595 & pe_o_2__4_;
  assign N592 = N591 & N596;
  assign N593 = N592 & pe_o_2__2_;
  assign N594 = N593 & pe_o_2__0_;
  assign N2614 = N594 & N597;
  assign N595 = ~pe_o_2__5_;
  assign N596 = ~pe_o_2__3_;
  assign N597 = ~pe_o_2__1_;
  assign N598 = N602 & pe_o_2__4_;
  assign N599 = N598 & N603;
  assign N600 = N599 & pe_o_2__2_;
  assign N601 = N600 & N604;
  assign N2616 = N601 & pe_o_2__1_;
  assign N602 = ~pe_o_2__5_;
  assign N603 = ~pe_o_2__3_;
  assign N604 = ~pe_o_2__0_;
  assign N605 = N609 & pe_o_2__4_;
  assign N606 = N605 & N610;
  assign N607 = N606 & pe_o_2__2_;
  assign N608 = N607 & pe_o_2__0_;
  assign N2618 = N608 & pe_o_2__1_;
  assign N609 = ~pe_o_2__5_;
  assign N610 = ~pe_o_2__3_;
  assign N611 = N615 & pe_o_2__4_;
  assign N612 = N611 & pe_o_2__3_;
  assign N613 = N612 & N616;
  assign N614 = N613 & N617;
  assign N2620 = N614 & N618;
  assign N615 = ~pe_o_2__5_;
  assign N616 = ~pe_o_2__2_;
  assign N617 = ~pe_o_2__0_;
  assign N618 = ~pe_o_2__1_;
  assign N619 = N623 & pe_o_2__4_;
  assign N620 = N619 & pe_o_2__3_;
  assign N621 = N620 & N624;
  assign N622 = N621 & pe_o_2__0_;
  assign N2622 = N622 & N625;
  assign N623 = ~pe_o_2__5_;
  assign N624 = ~pe_o_2__2_;
  assign N625 = ~pe_o_2__1_;
  assign N626 = N630 & pe_o_2__4_;
  assign N627 = N626 & pe_o_2__3_;
  assign N628 = N627 & N631;
  assign N629 = N628 & N632;
  assign N2624 = N629 & pe_o_2__1_;
  assign N630 = ~pe_o_2__5_;
  assign N631 = ~pe_o_2__2_;
  assign N632 = ~pe_o_2__0_;
  assign N633 = N637 & pe_o_2__4_;
  assign N634 = N633 & pe_o_2__3_;
  assign N635 = N634 & N638;
  assign N636 = N635 & pe_o_2__0_;
  assign N2626 = N636 & pe_o_2__1_;
  assign N637 = ~pe_o_2__5_;
  assign N638 = ~pe_o_2__2_;
  assign N639 = N643 & pe_o_2__4_;
  assign N640 = N639 & pe_o_2__3_;
  assign N641 = N640 & pe_o_2__2_;
  assign N642 = N641 & N644;
  assign N2628 = N642 & N645;
  assign N643 = ~pe_o_2__5_;
  assign N644 = ~pe_o_2__0_;
  assign N645 = ~pe_o_2__1_;
  assign N646 = N650 & pe_o_2__4_;
  assign N647 = N646 & pe_o_2__3_;
  assign N648 = N647 & pe_o_2__2_;
  assign N649 = N648 & pe_o_2__0_;
  assign N2630 = N649 & N651;
  assign N650 = ~pe_o_2__5_;
  assign N651 = ~pe_o_2__1_;
  assign N652 = N656 & pe_o_2__4_;
  assign N653 = N652 & pe_o_2__3_;
  assign N654 = N653 & pe_o_2__2_;
  assign N655 = N654 & N657;
  assign N2632 = N655 & pe_o_2__1_;
  assign N656 = ~pe_o_2__5_;
  assign N657 = ~pe_o_2__0_;
  assign N2634 = pe_o_2__4_ & pe_o_2__3_ & (pe_o_2__2_ & pe_o_2__0_) & pe_o_2__1_;
  assign N658 = pe_o_2__5_ & N662;
  assign N659 = N658 & N663;
  assign N660 = N659 & N664;
  assign N661 = N660 & pe_o_2__0_;
  assign N2575 = N661 & N665;
  assign N662 = ~pe_o_2__4_;
  assign N663 = ~pe_o_2__3_;
  assign N664 = ~pe_o_2__2_;
  assign N665 = ~pe_o_2__1_;
  assign N666 = pe_o_2__5_ & N670;
  assign N667 = N666 & N671;
  assign N668 = N667 & N672;
  assign N669 = N668 & N673;
  assign N2577 = N669 & pe_o_2__1_;
  assign N670 = ~pe_o_2__4_;
  assign N671 = ~pe_o_2__3_;
  assign N672 = ~pe_o_2__2_;
  assign N673 = ~pe_o_2__0_;
  assign N674 = pe_o_2__5_ & N678;
  assign N675 = N674 & N679;
  assign N676 = N675 & N680;
  assign N677 = N676 & pe_o_2__0_;
  assign N2579 = N677 & pe_o_2__1_;
  assign N678 = ~pe_o_2__4_;
  assign N679 = ~pe_o_2__3_;
  assign N680 = ~pe_o_2__2_;
  assign N681 = pe_o_2__5_ & N685;
  assign N682 = N681 & N686;
  assign N683 = N682 & pe_o_2__2_;
  assign N684 = N683 & N687;
  assign N2581 = N684 & N688;
  assign N685 = ~pe_o_2__4_;
  assign N686 = ~pe_o_2__3_;
  assign N687 = ~pe_o_2__0_;
  assign N688 = ~pe_o_2__1_;
  assign N689 = pe_o_2__5_ & N693;
  assign N690 = N689 & N694;
  assign N691 = N690 & pe_o_2__2_;
  assign N692 = N691 & pe_o_2__0_;
  assign N2583 = N692 & N695;
  assign N693 = ~pe_o_2__4_;
  assign N694 = ~pe_o_2__3_;
  assign N695 = ~pe_o_2__1_;
  assign N696 = pe_o_2__5_ & N700;
  assign N697 = N696 & N701;
  assign N698 = N697 & pe_o_2__2_;
  assign N699 = N698 & N702;
  assign N2585 = N699 & pe_o_2__1_;
  assign N700 = ~pe_o_2__4_;
  assign N701 = ~pe_o_2__3_;
  assign N702 = ~pe_o_2__0_;
  assign N703 = pe_o_2__5_ & N707;
  assign N704 = N703 & N708;
  assign N705 = N704 & pe_o_2__2_;
  assign N706 = N705 & pe_o_2__0_;
  assign N2587 = N706 & pe_o_2__1_;
  assign N707 = ~pe_o_2__4_;
  assign N708 = ~pe_o_2__3_;
  assign N709 = pe_o_2__5_ & N713;
  assign N710 = N709 & pe_o_2__3_;
  assign N711 = N710 & N714;
  assign N712 = N711 & N715;
  assign N2589 = N712 & N716;
  assign N713 = ~pe_o_2__4_;
  assign N714 = ~pe_o_2__2_;
  assign N715 = ~pe_o_2__0_;
  assign N716 = ~pe_o_2__1_;
  assign N717 = pe_o_2__5_ & N721;
  assign N718 = N717 & pe_o_2__3_;
  assign N719 = N718 & N722;
  assign N720 = N719 & pe_o_2__0_;
  assign N2591 = N720 & N723;
  assign N721 = ~pe_o_2__4_;
  assign N722 = ~pe_o_2__2_;
  assign N723 = ~pe_o_2__1_;
  assign N724 = pe_o_2__5_ & N728;
  assign N725 = N724 & pe_o_2__3_;
  assign N726 = N725 & N729;
  assign N727 = N726 & N730;
  assign N2593 = N727 & pe_o_2__1_;
  assign N728 = ~pe_o_2__4_;
  assign N729 = ~pe_o_2__2_;
  assign N730 = ~pe_o_2__0_;
  assign N731 = pe_o_2__5_ & N735;
  assign N732 = N731 & pe_o_2__3_;
  assign N733 = N732 & N736;
  assign N734 = N733 & pe_o_2__0_;
  assign N2595 = N734 & pe_o_2__1_;
  assign N735 = ~pe_o_2__4_;
  assign N736 = ~pe_o_2__2_;
  assign N737 = pe_o_2__5_ & N741;
  assign N738 = N737 & pe_o_2__3_;
  assign N739 = N738 & pe_o_2__2_;
  assign N740 = N739 & N742;
  assign N2597 = N740 & N743;
  assign N741 = ~pe_o_2__4_;
  assign N742 = ~pe_o_2__0_;
  assign N743 = ~pe_o_2__1_;
  assign N744 = pe_o_2__5_ & N748;
  assign N745 = N744 & pe_o_2__3_;
  assign N746 = N745 & pe_o_2__2_;
  assign N747 = N746 & pe_o_2__0_;
  assign N2599 = N747 & N749;
  assign N748 = ~pe_o_2__4_;
  assign N749 = ~pe_o_2__1_;
  assign N750 = pe_o_2__5_ & N754;
  assign N751 = N750 & pe_o_2__3_;
  assign N752 = N751 & pe_o_2__2_;
  assign N753 = N752 & N755;
  assign N2601 = N753 & pe_o_2__1_;
  assign N754 = ~pe_o_2__4_;
  assign N755 = ~pe_o_2__0_;
  assign N2603 = pe_o_2__5_ & pe_o_2__3_ & (pe_o_2__2_ & pe_o_2__0_) & pe_o_2__1_;
  assign N756 = pe_o_2__5_ & pe_o_2__4_;
  assign N757 = N756 & N760;
  assign N758 = N757 & N761;
  assign N759 = N758 & N762;
  assign N2605 = N759 & N763;
  assign N760 = ~pe_o_2__3_;
  assign N761 = ~pe_o_2__2_;
  assign N762 = ~pe_o_2__0_;
  assign N763 = ~pe_o_2__1_;
  assign N764 = pe_o_2__5_ & pe_o_2__4_;
  assign N765 = N764 & N768;
  assign N766 = N765 & N769;
  assign N767 = N766 & pe_o_2__0_;
  assign N2607 = N767 & N770;
  assign N768 = ~pe_o_2__3_;
  assign N769 = ~pe_o_2__2_;
  assign N770 = ~pe_o_2__1_;
  assign N771 = pe_o_2__5_ & pe_o_2__4_;
  assign N772 = N771 & N775;
  assign N773 = N772 & N776;
  assign N774 = N773 & N777;
  assign N2609 = N774 & pe_o_2__1_;
  assign N775 = ~pe_o_2__3_;
  assign N776 = ~pe_o_2__2_;
  assign N777 = ~pe_o_2__0_;
  assign N778 = pe_o_2__5_ & pe_o_2__4_;
  assign N779 = N778 & N782;
  assign N780 = N779 & N783;
  assign N781 = N780 & pe_o_2__0_;
  assign N2611 = N781 & pe_o_2__1_;
  assign N782 = ~pe_o_2__3_;
  assign N783 = ~pe_o_2__2_;
  assign N784 = pe_o_2__5_ & pe_o_2__4_;
  assign N785 = N784 & N788;
  assign N786 = N785 & pe_o_2__2_;
  assign N787 = N786 & N789;
  assign N2613 = N787 & N790;
  assign N788 = ~pe_o_2__3_;
  assign N789 = ~pe_o_2__0_;
  assign N790 = ~pe_o_2__1_;
  assign N791 = pe_o_2__5_ & pe_o_2__4_;
  assign N792 = N791 & N795;
  assign N793 = N792 & pe_o_2__2_;
  assign N794 = N793 & pe_o_2__0_;
  assign N2615 = N794 & N796;
  assign N795 = ~pe_o_2__3_;
  assign N796 = ~pe_o_2__1_;
  assign N797 = pe_o_2__5_ & pe_o_2__4_;
  assign N798 = N797 & N801;
  assign N799 = N798 & pe_o_2__2_;
  assign N800 = N799 & N802;
  assign N2617 = N800 & pe_o_2__1_;
  assign N801 = ~pe_o_2__3_;
  assign N802 = ~pe_o_2__0_;
  assign N2619 = pe_o_2__5_ & pe_o_2__4_ & (pe_o_2__2_ & pe_o_2__0_) & pe_o_2__1_;
  assign N803 = pe_o_2__5_ & pe_o_2__4_;
  assign N804 = N803 & pe_o_2__3_;
  assign N805 = N804 & N807;
  assign N806 = N805 & N808;
  assign N2621 = N806 & N809;
  assign N807 = ~pe_o_2__2_;
  assign N808 = ~pe_o_2__0_;
  assign N809 = ~pe_o_2__1_;
  assign N810 = pe_o_2__5_ & pe_o_2__4_;
  assign N811 = N810 & pe_o_2__3_;
  assign N812 = N811 & N814;
  assign N813 = N812 & pe_o_2__0_;
  assign N2623 = N813 & N815;
  assign N814 = ~pe_o_2__2_;
  assign N815 = ~pe_o_2__1_;
  assign N816 = pe_o_2__5_ & pe_o_2__4_;
  assign N817 = N816 & pe_o_2__3_;
  assign N818 = N817 & N820;
  assign N819 = N818 & N821;
  assign N2625 = N819 & pe_o_2__1_;
  assign N820 = ~pe_o_2__2_;
  assign N821 = ~pe_o_2__0_;
  assign N2627 = pe_o_2__5_ & pe_o_2__4_ & (pe_o_2__3_ & pe_o_2__0_) & pe_o_2__1_;
  assign N822 = pe_o_2__5_ & pe_o_2__4_;
  assign N823 = N822 & pe_o_2__3_;
  assign N824 = N823 & pe_o_2__2_;
  assign N825 = N824 & N826;
  assign N2629 = N825 & N827;
  assign N826 = ~pe_o_2__0_;
  assign N827 = ~pe_o_2__1_;
  assign N2631 = pe_o_2__5_ & pe_o_2__4_ & (pe_o_2__3_ & pe_o_2__2_) & pe_o_2__0_;
  assign N2633 = pe_o_2__5_ & pe_o_2__4_ & (pe_o_2__3_ & pe_o_2__2_) & pe_o_2__1_;
  assign N828 = N832 & N833;
  assign N829 = N828 & N834;
  assign N830 = N829 & N835;
  assign N831 = N830 & N836;
  assign N2698 = N831 & N837;
  assign N832 = ~pe_o_3__5_;
  assign N833 = ~pe_o_3__4_;
  assign N834 = ~pe_o_3__3_;
  assign N835 = ~pe_o_3__2_;
  assign N836 = ~pe_o_3__0_;
  assign N837 = ~pe_o_3__1_;
  assign N838 = pe_o_3__5_ & N842;
  assign N839 = N838 & N843;
  assign N840 = N839 & N844;
  assign N841 = N840 & N845;
  assign N2699 = N841 & N846;
  assign N842 = ~pe_o_3__4_;
  assign N843 = ~pe_o_3__3_;
  assign N844 = ~pe_o_3__2_;
  assign N845 = ~pe_o_3__0_;
  assign N846 = ~pe_o_3__1_;
  assign N847 = N851 & N852;
  assign N848 = N847 & N853;
  assign N849 = N848 & N854;
  assign N850 = N849 & pe_o_3__0_;
  assign N2700 = N850 & N855;
  assign N851 = ~pe_o_3__5_;
  assign N852 = ~pe_o_3__4_;
  assign N853 = ~pe_o_3__3_;
  assign N854 = ~pe_o_3__2_;
  assign N855 = ~pe_o_3__1_;
  assign N856 = N860 & N861;
  assign N857 = N856 & N862;
  assign N858 = N857 & N863;
  assign N859 = N858 & N864;
  assign N2702 = N859 & pe_o_3__1_;
  assign N860 = ~pe_o_3__5_;
  assign N861 = ~pe_o_3__4_;
  assign N862 = ~pe_o_3__3_;
  assign N863 = ~pe_o_3__2_;
  assign N864 = ~pe_o_3__0_;
  assign N865 = N869 & N870;
  assign N866 = N865 & N871;
  assign N867 = N866 & N872;
  assign N868 = N867 & pe_o_3__0_;
  assign N2704 = N868 & pe_o_3__1_;
  assign N869 = ~pe_o_3__5_;
  assign N870 = ~pe_o_3__4_;
  assign N871 = ~pe_o_3__3_;
  assign N872 = ~pe_o_3__2_;
  assign N873 = N877 & N878;
  assign N874 = N873 & N879;
  assign N875 = N874 & pe_o_3__2_;
  assign N876 = N875 & N880;
  assign N2706 = N876 & N881;
  assign N877 = ~pe_o_3__5_;
  assign N878 = ~pe_o_3__4_;
  assign N879 = ~pe_o_3__3_;
  assign N880 = ~pe_o_3__0_;
  assign N881 = ~pe_o_3__1_;
  assign N882 = N886 & N887;
  assign N883 = N882 & N888;
  assign N884 = N883 & pe_o_3__2_;
  assign N885 = N884 & pe_o_3__0_;
  assign N2708 = N885 & N889;
  assign N886 = ~pe_o_3__5_;
  assign N887 = ~pe_o_3__4_;
  assign N888 = ~pe_o_3__3_;
  assign N889 = ~pe_o_3__1_;
  assign N890 = N894 & N895;
  assign N891 = N890 & N896;
  assign N892 = N891 & pe_o_3__2_;
  assign N893 = N892 & N897;
  assign N2710 = N893 & pe_o_3__1_;
  assign N894 = ~pe_o_3__5_;
  assign N895 = ~pe_o_3__4_;
  assign N896 = ~pe_o_3__3_;
  assign N897 = ~pe_o_3__0_;
  assign N898 = N902 & N903;
  assign N899 = N898 & N904;
  assign N900 = N899 & pe_o_3__2_;
  assign N901 = N900 & pe_o_3__0_;
  assign N2712 = N901 & pe_o_3__1_;
  assign N902 = ~pe_o_3__5_;
  assign N903 = ~pe_o_3__4_;
  assign N904 = ~pe_o_3__3_;
  assign N905 = N909 & N910;
  assign N906 = N905 & pe_o_3__3_;
  assign N907 = N906 & N911;
  assign N908 = N907 & N912;
  assign N2714 = N908 & N913;
  assign N909 = ~pe_o_3__5_;
  assign N910 = ~pe_o_3__4_;
  assign N911 = ~pe_o_3__2_;
  assign N912 = ~pe_o_3__0_;
  assign N913 = ~pe_o_3__1_;
  assign N914 = N918 & N919;
  assign N915 = N914 & pe_o_3__3_;
  assign N916 = N915 & N920;
  assign N917 = N916 & pe_o_3__0_;
  assign N2716 = N917 & N921;
  assign N918 = ~pe_o_3__5_;
  assign N919 = ~pe_o_3__4_;
  assign N920 = ~pe_o_3__2_;
  assign N921 = ~pe_o_3__1_;
  assign N922 = N926 & N927;
  assign N923 = N922 & pe_o_3__3_;
  assign N924 = N923 & N928;
  assign N925 = N924 & N929;
  assign N2718 = N925 & pe_o_3__1_;
  assign N926 = ~pe_o_3__5_;
  assign N927 = ~pe_o_3__4_;
  assign N928 = ~pe_o_3__2_;
  assign N929 = ~pe_o_3__0_;
  assign N930 = N934 & N935;
  assign N931 = N930 & pe_o_3__3_;
  assign N932 = N931 & N936;
  assign N933 = N932 & pe_o_3__0_;
  assign N2720 = N933 & pe_o_3__1_;
  assign N934 = ~pe_o_3__5_;
  assign N935 = ~pe_o_3__4_;
  assign N936 = ~pe_o_3__2_;
  assign N937 = N941 & N942;
  assign N938 = N937 & pe_o_3__3_;
  assign N939 = N938 & pe_o_3__2_;
  assign N940 = N939 & N943;
  assign N2722 = N940 & N944;
  assign N941 = ~pe_o_3__5_;
  assign N942 = ~pe_o_3__4_;
  assign N943 = ~pe_o_3__0_;
  assign N944 = ~pe_o_3__1_;
  assign N945 = N949 & N950;
  assign N946 = N945 & pe_o_3__3_;
  assign N947 = N946 & pe_o_3__2_;
  assign N948 = N947 & pe_o_3__0_;
  assign N2724 = N948 & N951;
  assign N949 = ~pe_o_3__5_;
  assign N950 = ~pe_o_3__4_;
  assign N951 = ~pe_o_3__1_;
  assign N952 = N956 & N957;
  assign N953 = N952 & pe_o_3__3_;
  assign N954 = N953 & pe_o_3__2_;
  assign N955 = N954 & N958;
  assign N2726 = N955 & pe_o_3__1_;
  assign N956 = ~pe_o_3__5_;
  assign N957 = ~pe_o_3__4_;
  assign N958 = ~pe_o_3__0_;
  assign N959 = N963 & N964;
  assign N960 = N959 & pe_o_3__3_;
  assign N961 = N960 & pe_o_3__2_;
  assign N962 = N961 & pe_o_3__0_;
  assign N2728 = N962 & pe_o_3__1_;
  assign N963 = ~pe_o_3__5_;
  assign N964 = ~pe_o_3__4_;
  assign N965 = N969 & pe_o_3__4_;
  assign N966 = N965 & N970;
  assign N967 = N966 & N971;
  assign N968 = N967 & N972;
  assign N2730 = N968 & N973;
  assign N969 = ~pe_o_3__5_;
  assign N970 = ~pe_o_3__3_;
  assign N971 = ~pe_o_3__2_;
  assign N972 = ~pe_o_3__0_;
  assign N973 = ~pe_o_3__1_;
  assign N974 = N978 & pe_o_3__4_;
  assign N975 = N974 & N979;
  assign N976 = N975 & N980;
  assign N977 = N976 & pe_o_3__0_;
  assign N2732 = N977 & N981;
  assign N978 = ~pe_o_3__5_;
  assign N979 = ~pe_o_3__3_;
  assign N980 = ~pe_o_3__2_;
  assign N981 = ~pe_o_3__1_;
  assign N982 = N986 & pe_o_3__4_;
  assign N983 = N982 & N987;
  assign N984 = N983 & N988;
  assign N985 = N984 & N989;
  assign N2734 = N985 & pe_o_3__1_;
  assign N986 = ~pe_o_3__5_;
  assign N987 = ~pe_o_3__3_;
  assign N988 = ~pe_o_3__2_;
  assign N989 = ~pe_o_3__0_;
  assign N990 = N994 & pe_o_3__4_;
  assign N991 = N990 & N995;
  assign N992 = N991 & N996;
  assign N993 = N992 & pe_o_3__0_;
  assign N2736 = N993 & pe_o_3__1_;
  assign N994 = ~pe_o_3__5_;
  assign N995 = ~pe_o_3__3_;
  assign N996 = ~pe_o_3__2_;
  assign N997 = N1001 & pe_o_3__4_;
  assign N998 = N997 & N1002;
  assign N999 = N998 & pe_o_3__2_;
  assign N1000 = N999 & N1003;
  assign N2738 = N1000 & N1004;
  assign N1001 = ~pe_o_3__5_;
  assign N1002 = ~pe_o_3__3_;
  assign N1003 = ~pe_o_3__0_;
  assign N1004 = ~pe_o_3__1_;
  assign N1005 = N1009 & pe_o_3__4_;
  assign N1006 = N1005 & N1010;
  assign N1007 = N1006 & pe_o_3__2_;
  assign N1008 = N1007 & pe_o_3__0_;
  assign N2740 = N1008 & N1011;
  assign N1009 = ~pe_o_3__5_;
  assign N1010 = ~pe_o_3__3_;
  assign N1011 = ~pe_o_3__1_;
  assign N1012 = N1016 & pe_o_3__4_;
  assign N1013 = N1012 & N1017;
  assign N1014 = N1013 & pe_o_3__2_;
  assign N1015 = N1014 & N1018;
  assign N2742 = N1015 & pe_o_3__1_;
  assign N1016 = ~pe_o_3__5_;
  assign N1017 = ~pe_o_3__3_;
  assign N1018 = ~pe_o_3__0_;
  assign N1019 = N1023 & pe_o_3__4_;
  assign N1020 = N1019 & N1024;
  assign N1021 = N1020 & pe_o_3__2_;
  assign N1022 = N1021 & pe_o_3__0_;
  assign N2744 = N1022 & pe_o_3__1_;
  assign N1023 = ~pe_o_3__5_;
  assign N1024 = ~pe_o_3__3_;
  assign N1025 = N1029 & pe_o_3__4_;
  assign N1026 = N1025 & pe_o_3__3_;
  assign N1027 = N1026 & N1030;
  assign N1028 = N1027 & N1031;
  assign N2746 = N1028 & N1032;
  assign N1029 = ~pe_o_3__5_;
  assign N1030 = ~pe_o_3__2_;
  assign N1031 = ~pe_o_3__0_;
  assign N1032 = ~pe_o_3__1_;
  assign N1033 = N1037 & pe_o_3__4_;
  assign N1034 = N1033 & pe_o_3__3_;
  assign N1035 = N1034 & N1038;
  assign N1036 = N1035 & pe_o_3__0_;
  assign N2748 = N1036 & N1039;
  assign N1037 = ~pe_o_3__5_;
  assign N1038 = ~pe_o_3__2_;
  assign N1039 = ~pe_o_3__1_;
  assign N1040 = N1044 & pe_o_3__4_;
  assign N1041 = N1040 & pe_o_3__3_;
  assign N1042 = N1041 & N1045;
  assign N1043 = N1042 & N1046;
  assign N2750 = N1043 & pe_o_3__1_;
  assign N1044 = ~pe_o_3__5_;
  assign N1045 = ~pe_o_3__2_;
  assign N1046 = ~pe_o_3__0_;
  assign N1047 = N1051 & pe_o_3__4_;
  assign N1048 = N1047 & pe_o_3__3_;
  assign N1049 = N1048 & N1052;
  assign N1050 = N1049 & pe_o_3__0_;
  assign N2752 = N1050 & pe_o_3__1_;
  assign N1051 = ~pe_o_3__5_;
  assign N1052 = ~pe_o_3__2_;
  assign N1053 = N1057 & pe_o_3__4_;
  assign N1054 = N1053 & pe_o_3__3_;
  assign N1055 = N1054 & pe_o_3__2_;
  assign N1056 = N1055 & N1058;
  assign N2754 = N1056 & N1059;
  assign N1057 = ~pe_o_3__5_;
  assign N1058 = ~pe_o_3__0_;
  assign N1059 = ~pe_o_3__1_;
  assign N1060 = N1064 & pe_o_3__4_;
  assign N1061 = N1060 & pe_o_3__3_;
  assign N1062 = N1061 & pe_o_3__2_;
  assign N1063 = N1062 & pe_o_3__0_;
  assign N2756 = N1063 & N1065;
  assign N1064 = ~pe_o_3__5_;
  assign N1065 = ~pe_o_3__1_;
  assign N1066 = N1070 & pe_o_3__4_;
  assign N1067 = N1066 & pe_o_3__3_;
  assign N1068 = N1067 & pe_o_3__2_;
  assign N1069 = N1068 & N1071;
  assign N2758 = N1069 & pe_o_3__1_;
  assign N1070 = ~pe_o_3__5_;
  assign N1071 = ~pe_o_3__0_;
  assign N2760 = pe_o_3__4_ & pe_o_3__3_ & (pe_o_3__2_ & pe_o_3__0_) & pe_o_3__1_;
  assign N1072 = pe_o_3__5_ & N1076;
  assign N1073 = N1072 & N1077;
  assign N1074 = N1073 & N1078;
  assign N1075 = N1074 & pe_o_3__0_;
  assign N2701 = N1075 & N1079;
  assign N1076 = ~pe_o_3__4_;
  assign N1077 = ~pe_o_3__3_;
  assign N1078 = ~pe_o_3__2_;
  assign N1079 = ~pe_o_3__1_;
  assign N1080 = pe_o_3__5_ & N1084;
  assign N1081 = N1080 & N1085;
  assign N1082 = N1081 & N1086;
  assign N1083 = N1082 & N1087;
  assign N2703 = N1083 & pe_o_3__1_;
  assign N1084 = ~pe_o_3__4_;
  assign N1085 = ~pe_o_3__3_;
  assign N1086 = ~pe_o_3__2_;
  assign N1087 = ~pe_o_3__0_;
  assign N1088 = pe_o_3__5_ & N1092;
  assign N1089 = N1088 & N1093;
  assign N1090 = N1089 & N1094;
  assign N1091 = N1090 & pe_o_3__0_;
  assign N2705 = N1091 & pe_o_3__1_;
  assign N1092 = ~pe_o_3__4_;
  assign N1093 = ~pe_o_3__3_;
  assign N1094 = ~pe_o_3__2_;
  assign N1095 = pe_o_3__5_ & N1099;
  assign N1096 = N1095 & N1100;
  assign N1097 = N1096 & pe_o_3__2_;
  assign N1098 = N1097 & N1101;
  assign N2707 = N1098 & N1102;
  assign N1099 = ~pe_o_3__4_;
  assign N1100 = ~pe_o_3__3_;
  assign N1101 = ~pe_o_3__0_;
  assign N1102 = ~pe_o_3__1_;
  assign N1103 = pe_o_3__5_ & N1107;
  assign N1104 = N1103 & N1108;
  assign N1105 = N1104 & pe_o_3__2_;
  assign N1106 = N1105 & pe_o_3__0_;
  assign N2709 = N1106 & N1109;
  assign N1107 = ~pe_o_3__4_;
  assign N1108 = ~pe_o_3__3_;
  assign N1109 = ~pe_o_3__1_;
  assign N1110 = pe_o_3__5_ & N1114;
  assign N1111 = N1110 & N1115;
  assign N1112 = N1111 & pe_o_3__2_;
  assign N1113 = N1112 & N1116;
  assign N2711 = N1113 & pe_o_3__1_;
  assign N1114 = ~pe_o_3__4_;
  assign N1115 = ~pe_o_3__3_;
  assign N1116 = ~pe_o_3__0_;
  assign N1117 = pe_o_3__5_ & N1121;
  assign N1118 = N1117 & N1122;
  assign N1119 = N1118 & pe_o_3__2_;
  assign N1120 = N1119 & pe_o_3__0_;
  assign N2713 = N1120 & pe_o_3__1_;
  assign N1121 = ~pe_o_3__4_;
  assign N1122 = ~pe_o_3__3_;
  assign N1123 = pe_o_3__5_ & N1127;
  assign N1124 = N1123 & pe_o_3__3_;
  assign N1125 = N1124 & N1128;
  assign N1126 = N1125 & N1129;
  assign N2715 = N1126 & N1130;
  assign N1127 = ~pe_o_3__4_;
  assign N1128 = ~pe_o_3__2_;
  assign N1129 = ~pe_o_3__0_;
  assign N1130 = ~pe_o_3__1_;
  assign N1131 = pe_o_3__5_ & N1135;
  assign N1132 = N1131 & pe_o_3__3_;
  assign N1133 = N1132 & N1136;
  assign N1134 = N1133 & pe_o_3__0_;
  assign N2717 = N1134 & N1137;
  assign N1135 = ~pe_o_3__4_;
  assign N1136 = ~pe_o_3__2_;
  assign N1137 = ~pe_o_3__1_;
  assign N1138 = pe_o_3__5_ & N1142;
  assign N1139 = N1138 & pe_o_3__3_;
  assign N1140 = N1139 & N1143;
  assign N1141 = N1140 & N1144;
  assign N2719 = N1141 & pe_o_3__1_;
  assign N1142 = ~pe_o_3__4_;
  assign N1143 = ~pe_o_3__2_;
  assign N1144 = ~pe_o_3__0_;
  assign N1145 = pe_o_3__5_ & N1149;
  assign N1146 = N1145 & pe_o_3__3_;
  assign N1147 = N1146 & N1150;
  assign N1148 = N1147 & pe_o_3__0_;
  assign N2721 = N1148 & pe_o_3__1_;
  assign N1149 = ~pe_o_3__4_;
  assign N1150 = ~pe_o_3__2_;
  assign N1151 = pe_o_3__5_ & N1155;
  assign N1152 = N1151 & pe_o_3__3_;
  assign N1153 = N1152 & pe_o_3__2_;
  assign N1154 = N1153 & N1156;
  assign N2723 = N1154 & N1157;
  assign N1155 = ~pe_o_3__4_;
  assign N1156 = ~pe_o_3__0_;
  assign N1157 = ~pe_o_3__1_;
  assign N1158 = pe_o_3__5_ & N1162;
  assign N1159 = N1158 & pe_o_3__3_;
  assign N1160 = N1159 & pe_o_3__2_;
  assign N1161 = N1160 & pe_o_3__0_;
  assign N2725 = N1161 & N1163;
  assign N1162 = ~pe_o_3__4_;
  assign N1163 = ~pe_o_3__1_;
  assign N1164 = pe_o_3__5_ & N1168;
  assign N1165 = N1164 & pe_o_3__3_;
  assign N1166 = N1165 & pe_o_3__2_;
  assign N1167 = N1166 & N1169;
  assign N2727 = N1167 & pe_o_3__1_;
  assign N1168 = ~pe_o_3__4_;
  assign N1169 = ~pe_o_3__0_;
  assign N2729 = pe_o_3__5_ & pe_o_3__3_ & (pe_o_3__2_ & pe_o_3__0_) & pe_o_3__1_;
  assign N1170 = pe_o_3__5_ & pe_o_3__4_;
  assign N1171 = N1170 & N1174;
  assign N1172 = N1171 & N1175;
  assign N1173 = N1172 & N1176;
  assign N2731 = N1173 & N1177;
  assign N1174 = ~pe_o_3__3_;
  assign N1175 = ~pe_o_3__2_;
  assign N1176 = ~pe_o_3__0_;
  assign N1177 = ~pe_o_3__1_;
  assign N1178 = pe_o_3__5_ & pe_o_3__4_;
  assign N1179 = N1178 & N1182;
  assign N1180 = N1179 & N1183;
  assign N1181 = N1180 & pe_o_3__0_;
  assign N2733 = N1181 & N1184;
  assign N1182 = ~pe_o_3__3_;
  assign N1183 = ~pe_o_3__2_;
  assign N1184 = ~pe_o_3__1_;
  assign N1185 = pe_o_3__5_ & pe_o_3__4_;
  assign N1186 = N1185 & N1189;
  assign N1187 = N1186 & N1190;
  assign N1188 = N1187 & N1191;
  assign N2735 = N1188 & pe_o_3__1_;
  assign N1189 = ~pe_o_3__3_;
  assign N1190 = ~pe_o_3__2_;
  assign N1191 = ~pe_o_3__0_;
  assign N1192 = pe_o_3__5_ & pe_o_3__4_;
  assign N1193 = N1192 & N1196;
  assign N1194 = N1193 & N1197;
  assign N1195 = N1194 & pe_o_3__0_;
  assign N2737 = N1195 & pe_o_3__1_;
  assign N1196 = ~pe_o_3__3_;
  assign N1197 = ~pe_o_3__2_;
  assign N1198 = pe_o_3__5_ & pe_o_3__4_;
  assign N1199 = N1198 & N1202;
  assign N1200 = N1199 & pe_o_3__2_;
  assign N1201 = N1200 & N1203;
  assign N2739 = N1201 & N1204;
  assign N1202 = ~pe_o_3__3_;
  assign N1203 = ~pe_o_3__0_;
  assign N1204 = ~pe_o_3__1_;
  assign N1205 = pe_o_3__5_ & pe_o_3__4_;
  assign N1206 = N1205 & N1209;
  assign N1207 = N1206 & pe_o_3__2_;
  assign N1208 = N1207 & pe_o_3__0_;
  assign N2741 = N1208 & N1210;
  assign N1209 = ~pe_o_3__3_;
  assign N1210 = ~pe_o_3__1_;
  assign N1211 = pe_o_3__5_ & pe_o_3__4_;
  assign N1212 = N1211 & N1215;
  assign N1213 = N1212 & pe_o_3__2_;
  assign N1214 = N1213 & N1216;
  assign N2743 = N1214 & pe_o_3__1_;
  assign N1215 = ~pe_o_3__3_;
  assign N1216 = ~pe_o_3__0_;
  assign N2745 = pe_o_3__5_ & pe_o_3__4_ & (pe_o_3__2_ & pe_o_3__0_) & pe_o_3__1_;
  assign N1217 = pe_o_3__5_ & pe_o_3__4_;
  assign N1218 = N1217 & pe_o_3__3_;
  assign N1219 = N1218 & N1221;
  assign N1220 = N1219 & N1222;
  assign N2747 = N1220 & N1223;
  assign N1221 = ~pe_o_3__2_;
  assign N1222 = ~pe_o_3__0_;
  assign N1223 = ~pe_o_3__1_;
  assign N1224 = pe_o_3__5_ & pe_o_3__4_;
  assign N1225 = N1224 & pe_o_3__3_;
  assign N1226 = N1225 & N1228;
  assign N1227 = N1226 & pe_o_3__0_;
  assign N2749 = N1227 & N1229;
  assign N1228 = ~pe_o_3__2_;
  assign N1229 = ~pe_o_3__1_;
  assign N1230 = pe_o_3__5_ & pe_o_3__4_;
  assign N1231 = N1230 & pe_o_3__3_;
  assign N1232 = N1231 & N1234;
  assign N1233 = N1232 & N1235;
  assign N2751 = N1233 & pe_o_3__1_;
  assign N1234 = ~pe_o_3__2_;
  assign N1235 = ~pe_o_3__0_;
  assign N2753 = pe_o_3__5_ & pe_o_3__4_ & (pe_o_3__3_ & pe_o_3__0_) & pe_o_3__1_;
  assign N1236 = pe_o_3__5_ & pe_o_3__4_;
  assign N1237 = N1236 & pe_o_3__3_;
  assign N1238 = N1237 & pe_o_3__2_;
  assign N1239 = N1238 & N1240;
  assign N2755 = N1239 & N1241;
  assign N1240 = ~pe_o_3__0_;
  assign N1241 = ~pe_o_3__1_;
  assign N2757 = pe_o_3__5_ & pe_o_3__4_ & (pe_o_3__3_ & pe_o_3__2_) & pe_o_3__0_;
  assign N2759 = pe_o_3__5_ & pe_o_3__4_ & (pe_o_3__3_ & pe_o_3__2_) & pe_o_3__1_;
  assign N1242 = N1246 & N1247;
  assign N1243 = N1242 & N1248;
  assign N1244 = N1243 & N1249;
  assign N1245 = N1244 & N1250;
  assign N2824 = N1245 & N1251;
  assign N1246 = ~pe_o_4__5_;
  assign N1247 = ~pe_o_4__4_;
  assign N1248 = ~pe_o_4__3_;
  assign N1249 = ~pe_o_4__2_;
  assign N1250 = ~pe_o_4__0_;
  assign N1251 = ~pe_o_4__1_;
  assign N1252 = pe_o_4__5_ & N1256;
  assign N1253 = N1252 & N1257;
  assign N1254 = N1253 & N1258;
  assign N1255 = N1254 & N1259;
  assign N2825 = N1255 & N1260;
  assign N1256 = ~pe_o_4__4_;
  assign N1257 = ~pe_o_4__3_;
  assign N1258 = ~pe_o_4__2_;
  assign N1259 = ~pe_o_4__0_;
  assign N1260 = ~pe_o_4__1_;
  assign N1261 = N1265 & N1266;
  assign N1262 = N1261 & N1267;
  assign N1263 = N1262 & N1268;
  assign N1264 = N1263 & pe_o_4__0_;
  assign N2826 = N1264 & N1269;
  assign N1265 = ~pe_o_4__5_;
  assign N1266 = ~pe_o_4__4_;
  assign N1267 = ~pe_o_4__3_;
  assign N1268 = ~pe_o_4__2_;
  assign N1269 = ~pe_o_4__1_;
  assign N1270 = N1274 & N1275;
  assign N1271 = N1270 & N1276;
  assign N1272 = N1271 & N1277;
  assign N1273 = N1272 & N1278;
  assign N2828 = N1273 & pe_o_4__1_;
  assign N1274 = ~pe_o_4__5_;
  assign N1275 = ~pe_o_4__4_;
  assign N1276 = ~pe_o_4__3_;
  assign N1277 = ~pe_o_4__2_;
  assign N1278 = ~pe_o_4__0_;
  assign N1279 = N1283 & N1284;
  assign N1280 = N1279 & N1285;
  assign N1281 = N1280 & N1286;
  assign N1282 = N1281 & pe_o_4__0_;
  assign N2830 = N1282 & pe_o_4__1_;
  assign N1283 = ~pe_o_4__5_;
  assign N1284 = ~pe_o_4__4_;
  assign N1285 = ~pe_o_4__3_;
  assign N1286 = ~pe_o_4__2_;
  assign N1287 = N1291 & N1292;
  assign N1288 = N1287 & N1293;
  assign N1289 = N1288 & pe_o_4__2_;
  assign N1290 = N1289 & N1294;
  assign N2832 = N1290 & N1295;
  assign N1291 = ~pe_o_4__5_;
  assign N1292 = ~pe_o_4__4_;
  assign N1293 = ~pe_o_4__3_;
  assign N1294 = ~pe_o_4__0_;
  assign N1295 = ~pe_o_4__1_;
  assign N1296 = N1300 & N1301;
  assign N1297 = N1296 & N1302;
  assign N1298 = N1297 & pe_o_4__2_;
  assign N1299 = N1298 & pe_o_4__0_;
  assign N2834 = N1299 & N1303;
  assign N1300 = ~pe_o_4__5_;
  assign N1301 = ~pe_o_4__4_;
  assign N1302 = ~pe_o_4__3_;
  assign N1303 = ~pe_o_4__1_;
  assign N1304 = N1308 & N1309;
  assign N1305 = N1304 & N1310;
  assign N1306 = N1305 & pe_o_4__2_;
  assign N1307 = N1306 & N1311;
  assign N2836 = N1307 & pe_o_4__1_;
  assign N1308 = ~pe_o_4__5_;
  assign N1309 = ~pe_o_4__4_;
  assign N1310 = ~pe_o_4__3_;
  assign N1311 = ~pe_o_4__0_;
  assign N1312 = N1316 & N1317;
  assign N1313 = N1312 & N1318;
  assign N1314 = N1313 & pe_o_4__2_;
  assign N1315 = N1314 & pe_o_4__0_;
  assign N2838 = N1315 & pe_o_4__1_;
  assign N1316 = ~pe_o_4__5_;
  assign N1317 = ~pe_o_4__4_;
  assign N1318 = ~pe_o_4__3_;
  assign N1319 = N1323 & N1324;
  assign N1320 = N1319 & pe_o_4__3_;
  assign N1321 = N1320 & N1325;
  assign N1322 = N1321 & N1326;
  assign N2840 = N1322 & N1327;
  assign N1323 = ~pe_o_4__5_;
  assign N1324 = ~pe_o_4__4_;
  assign N1325 = ~pe_o_4__2_;
  assign N1326 = ~pe_o_4__0_;
  assign N1327 = ~pe_o_4__1_;
  assign N1328 = N1332 & N1333;
  assign N1329 = N1328 & pe_o_4__3_;
  assign N1330 = N1329 & N1334;
  assign N1331 = N1330 & pe_o_4__0_;
  assign N2842 = N1331 & N1335;
  assign N1332 = ~pe_o_4__5_;
  assign N1333 = ~pe_o_4__4_;
  assign N1334 = ~pe_o_4__2_;
  assign N1335 = ~pe_o_4__1_;
  assign N1336 = N1340 & N1341;
  assign N1337 = N1336 & pe_o_4__3_;
  assign N1338 = N1337 & N1342;
  assign N1339 = N1338 & N1343;
  assign N2844 = N1339 & pe_o_4__1_;
  assign N1340 = ~pe_o_4__5_;
  assign N1341 = ~pe_o_4__4_;
  assign N1342 = ~pe_o_4__2_;
  assign N1343 = ~pe_o_4__0_;
  assign N1344 = N1348 & N1349;
  assign N1345 = N1344 & pe_o_4__3_;
  assign N1346 = N1345 & N1350;
  assign N1347 = N1346 & pe_o_4__0_;
  assign N2846 = N1347 & pe_o_4__1_;
  assign N1348 = ~pe_o_4__5_;
  assign N1349 = ~pe_o_4__4_;
  assign N1350 = ~pe_o_4__2_;
  assign N1351 = N1355 & N1356;
  assign N1352 = N1351 & pe_o_4__3_;
  assign N1353 = N1352 & pe_o_4__2_;
  assign N1354 = N1353 & N1357;
  assign N2848 = N1354 & N1358;
  assign N1355 = ~pe_o_4__5_;
  assign N1356 = ~pe_o_4__4_;
  assign N1357 = ~pe_o_4__0_;
  assign N1358 = ~pe_o_4__1_;
  assign N1359 = N1363 & N1364;
  assign N1360 = N1359 & pe_o_4__3_;
  assign N1361 = N1360 & pe_o_4__2_;
  assign N1362 = N1361 & pe_o_4__0_;
  assign N2850 = N1362 & N1365;
  assign N1363 = ~pe_o_4__5_;
  assign N1364 = ~pe_o_4__4_;
  assign N1365 = ~pe_o_4__1_;
  assign N1366 = N1370 & N1371;
  assign N1367 = N1366 & pe_o_4__3_;
  assign N1368 = N1367 & pe_o_4__2_;
  assign N1369 = N1368 & N1372;
  assign N2852 = N1369 & pe_o_4__1_;
  assign N1370 = ~pe_o_4__5_;
  assign N1371 = ~pe_o_4__4_;
  assign N1372 = ~pe_o_4__0_;
  assign N1373 = N1377 & N1378;
  assign N1374 = N1373 & pe_o_4__3_;
  assign N1375 = N1374 & pe_o_4__2_;
  assign N1376 = N1375 & pe_o_4__0_;
  assign N2854 = N1376 & pe_o_4__1_;
  assign N1377 = ~pe_o_4__5_;
  assign N1378 = ~pe_o_4__4_;
  assign N1379 = N1383 & pe_o_4__4_;
  assign N1380 = N1379 & N1384;
  assign N1381 = N1380 & N1385;
  assign N1382 = N1381 & N1386;
  assign N2856 = N1382 & N1387;
  assign N1383 = ~pe_o_4__5_;
  assign N1384 = ~pe_o_4__3_;
  assign N1385 = ~pe_o_4__2_;
  assign N1386 = ~pe_o_4__0_;
  assign N1387 = ~pe_o_4__1_;
  assign N1388 = N1392 & pe_o_4__4_;
  assign N1389 = N1388 & N1393;
  assign N1390 = N1389 & N1394;
  assign N1391 = N1390 & pe_o_4__0_;
  assign N2858 = N1391 & N1395;
  assign N1392 = ~pe_o_4__5_;
  assign N1393 = ~pe_o_4__3_;
  assign N1394 = ~pe_o_4__2_;
  assign N1395 = ~pe_o_4__1_;
  assign N1396 = N1400 & pe_o_4__4_;
  assign N1397 = N1396 & N1401;
  assign N1398 = N1397 & N1402;
  assign N1399 = N1398 & N1403;
  assign N2860 = N1399 & pe_o_4__1_;
  assign N1400 = ~pe_o_4__5_;
  assign N1401 = ~pe_o_4__3_;
  assign N1402 = ~pe_o_4__2_;
  assign N1403 = ~pe_o_4__0_;
  assign N1404 = N1408 & pe_o_4__4_;
  assign N1405 = N1404 & N1409;
  assign N1406 = N1405 & N1410;
  assign N1407 = N1406 & pe_o_4__0_;
  assign N2862 = N1407 & pe_o_4__1_;
  assign N1408 = ~pe_o_4__5_;
  assign N1409 = ~pe_o_4__3_;
  assign N1410 = ~pe_o_4__2_;
  assign N1411 = N1415 & pe_o_4__4_;
  assign N1412 = N1411 & N1416;
  assign N1413 = N1412 & pe_o_4__2_;
  assign N1414 = N1413 & N1417;
  assign N2864 = N1414 & N1418;
  assign N1415 = ~pe_o_4__5_;
  assign N1416 = ~pe_o_4__3_;
  assign N1417 = ~pe_o_4__0_;
  assign N1418 = ~pe_o_4__1_;
  assign N1419 = N1423 & pe_o_4__4_;
  assign N1420 = N1419 & N1424;
  assign N1421 = N1420 & pe_o_4__2_;
  assign N1422 = N1421 & pe_o_4__0_;
  assign N2866 = N1422 & N1425;
  assign N1423 = ~pe_o_4__5_;
  assign N1424 = ~pe_o_4__3_;
  assign N1425 = ~pe_o_4__1_;
  assign N1426 = N1430 & pe_o_4__4_;
  assign N1427 = N1426 & N1431;
  assign N1428 = N1427 & pe_o_4__2_;
  assign N1429 = N1428 & N1432;
  assign N2868 = N1429 & pe_o_4__1_;
  assign N1430 = ~pe_o_4__5_;
  assign N1431 = ~pe_o_4__3_;
  assign N1432 = ~pe_o_4__0_;
  assign N1433 = N1437 & pe_o_4__4_;
  assign N1434 = N1433 & N1438;
  assign N1435 = N1434 & pe_o_4__2_;
  assign N1436 = N1435 & pe_o_4__0_;
  assign N2870 = N1436 & pe_o_4__1_;
  assign N1437 = ~pe_o_4__5_;
  assign N1438 = ~pe_o_4__3_;
  assign N1439 = N1443 & pe_o_4__4_;
  assign N1440 = N1439 & pe_o_4__3_;
  assign N1441 = N1440 & N1444;
  assign N1442 = N1441 & N1445;
  assign N2872 = N1442 & N1446;
  assign N1443 = ~pe_o_4__5_;
  assign N1444 = ~pe_o_4__2_;
  assign N1445 = ~pe_o_4__0_;
  assign N1446 = ~pe_o_4__1_;
  assign N1447 = N1451 & pe_o_4__4_;
  assign N1448 = N1447 & pe_o_4__3_;
  assign N1449 = N1448 & N1452;
  assign N1450 = N1449 & pe_o_4__0_;
  assign N2874 = N1450 & N1453;
  assign N1451 = ~pe_o_4__5_;
  assign N1452 = ~pe_o_4__2_;
  assign N1453 = ~pe_o_4__1_;
  assign N1454 = N1458 & pe_o_4__4_;
  assign N1455 = N1454 & pe_o_4__3_;
  assign N1456 = N1455 & N1459;
  assign N1457 = N1456 & N1460;
  assign N2876 = N1457 & pe_o_4__1_;
  assign N1458 = ~pe_o_4__5_;
  assign N1459 = ~pe_o_4__2_;
  assign N1460 = ~pe_o_4__0_;
  assign N1461 = N1465 & pe_o_4__4_;
  assign N1462 = N1461 & pe_o_4__3_;
  assign N1463 = N1462 & N1466;
  assign N1464 = N1463 & pe_o_4__0_;
  assign N2878 = N1464 & pe_o_4__1_;
  assign N1465 = ~pe_o_4__5_;
  assign N1466 = ~pe_o_4__2_;
  assign N1467 = N1471 & pe_o_4__4_;
  assign N1468 = N1467 & pe_o_4__3_;
  assign N1469 = N1468 & pe_o_4__2_;
  assign N1470 = N1469 & N1472;
  assign N2880 = N1470 & N1473;
  assign N1471 = ~pe_o_4__5_;
  assign N1472 = ~pe_o_4__0_;
  assign N1473 = ~pe_o_4__1_;
  assign N1474 = N1478 & pe_o_4__4_;
  assign N1475 = N1474 & pe_o_4__3_;
  assign N1476 = N1475 & pe_o_4__2_;
  assign N1477 = N1476 & pe_o_4__0_;
  assign N2882 = N1477 & N1479;
  assign N1478 = ~pe_o_4__5_;
  assign N1479 = ~pe_o_4__1_;
  assign N1480 = N1484 & pe_o_4__4_;
  assign N1481 = N1480 & pe_o_4__3_;
  assign N1482 = N1481 & pe_o_4__2_;
  assign N1483 = N1482 & N1485;
  assign N2884 = N1483 & pe_o_4__1_;
  assign N1484 = ~pe_o_4__5_;
  assign N1485 = ~pe_o_4__0_;
  assign N2886 = pe_o_4__4_ & pe_o_4__3_ & (pe_o_4__2_ & pe_o_4__0_) & pe_o_4__1_;
  assign N1486 = pe_o_4__5_ & N1490;
  assign N1487 = N1486 & N1491;
  assign N1488 = N1487 & N1492;
  assign N1489 = N1488 & pe_o_4__0_;
  assign N2827 = N1489 & N1493;
  assign N1490 = ~pe_o_4__4_;
  assign N1491 = ~pe_o_4__3_;
  assign N1492 = ~pe_o_4__2_;
  assign N1493 = ~pe_o_4__1_;
  assign N1494 = pe_o_4__5_ & N1498;
  assign N1495 = N1494 & N1499;
  assign N1496 = N1495 & N1500;
  assign N1497 = N1496 & N1501;
  assign N2829 = N1497 & pe_o_4__1_;
  assign N1498 = ~pe_o_4__4_;
  assign N1499 = ~pe_o_4__3_;
  assign N1500 = ~pe_o_4__2_;
  assign N1501 = ~pe_o_4__0_;
  assign N1502 = pe_o_4__5_ & N1506;
  assign N1503 = N1502 & N1507;
  assign N1504 = N1503 & N1508;
  assign N1505 = N1504 & pe_o_4__0_;
  assign N2831 = N1505 & pe_o_4__1_;
  assign N1506 = ~pe_o_4__4_;
  assign N1507 = ~pe_o_4__3_;
  assign N1508 = ~pe_o_4__2_;
  assign N1509 = pe_o_4__5_ & N1513;
  assign N1510 = N1509 & N1514;
  assign N1511 = N1510 & pe_o_4__2_;
  assign N1512 = N1511 & N1515;
  assign N2833 = N1512 & N1516;
  assign N1513 = ~pe_o_4__4_;
  assign N1514 = ~pe_o_4__3_;
  assign N1515 = ~pe_o_4__0_;
  assign N1516 = ~pe_o_4__1_;
  assign N1517 = pe_o_4__5_ & N1521;
  assign N1518 = N1517 & N1522;
  assign N1519 = N1518 & pe_o_4__2_;
  assign N1520 = N1519 & pe_o_4__0_;
  assign N2835 = N1520 & N1523;
  assign N1521 = ~pe_o_4__4_;
  assign N1522 = ~pe_o_4__3_;
  assign N1523 = ~pe_o_4__1_;
  assign N1524 = pe_o_4__5_ & N1528;
  assign N1525 = N1524 & N1529;
  assign N1526 = N1525 & pe_o_4__2_;
  assign N1527 = N1526 & N1530;
  assign N2837 = N1527 & pe_o_4__1_;
  assign N1528 = ~pe_o_4__4_;
  assign N1529 = ~pe_o_4__3_;
  assign N1530 = ~pe_o_4__0_;
  assign N1531 = pe_o_4__5_ & N1535;
  assign N1532 = N1531 & N1536;
  assign N1533 = N1532 & pe_o_4__2_;
  assign N1534 = N1533 & pe_o_4__0_;
  assign N2839 = N1534 & pe_o_4__1_;
  assign N1535 = ~pe_o_4__4_;
  assign N1536 = ~pe_o_4__3_;
  assign N1537 = pe_o_4__5_ & N1541;
  assign N1538 = N1537 & pe_o_4__3_;
  assign N1539 = N1538 & N1542;
  assign N1540 = N1539 & N1543;
  assign N2841 = N1540 & N1544;
  assign N1541 = ~pe_o_4__4_;
  assign N1542 = ~pe_o_4__2_;
  assign N1543 = ~pe_o_4__0_;
  assign N1544 = ~pe_o_4__1_;
  assign N1545 = pe_o_4__5_ & N1549;
  assign N1546 = N1545 & pe_o_4__3_;
  assign N1547 = N1546 & N1550;
  assign N1548 = N1547 & pe_o_4__0_;
  assign N2843 = N1548 & N1551;
  assign N1549 = ~pe_o_4__4_;
  assign N1550 = ~pe_o_4__2_;
  assign N1551 = ~pe_o_4__1_;
  assign N1552 = pe_o_4__5_ & N1556;
  assign N1553 = N1552 & pe_o_4__3_;
  assign N1554 = N1553 & N1557;
  assign N1555 = N1554 & N1558;
  assign N2845 = N1555 & pe_o_4__1_;
  assign N1556 = ~pe_o_4__4_;
  assign N1557 = ~pe_o_4__2_;
  assign N1558 = ~pe_o_4__0_;
  assign N1559 = pe_o_4__5_ & N1563;
  assign N1560 = N1559 & pe_o_4__3_;
  assign N1561 = N1560 & N1564;
  assign N1562 = N1561 & pe_o_4__0_;
  assign N2847 = N1562 & pe_o_4__1_;
  assign N1563 = ~pe_o_4__4_;
  assign N1564 = ~pe_o_4__2_;
  assign N1565 = pe_o_4__5_ & N1569;
  assign N1566 = N1565 & pe_o_4__3_;
  assign N1567 = N1566 & pe_o_4__2_;
  assign N1568 = N1567 & N1570;
  assign N2849 = N1568 & N1571;
  assign N1569 = ~pe_o_4__4_;
  assign N1570 = ~pe_o_4__0_;
  assign N1571 = ~pe_o_4__1_;
  assign N1572 = pe_o_4__5_ & N1576;
  assign N1573 = N1572 & pe_o_4__3_;
  assign N1574 = N1573 & pe_o_4__2_;
  assign N1575 = N1574 & pe_o_4__0_;
  assign N2851 = N1575 & N1577;
  assign N1576 = ~pe_o_4__4_;
  assign N1577 = ~pe_o_4__1_;
  assign N1578 = pe_o_4__5_ & N1582;
  assign N1579 = N1578 & pe_o_4__3_;
  assign N1580 = N1579 & pe_o_4__2_;
  assign N1581 = N1580 & N1583;
  assign N2853 = N1581 & pe_o_4__1_;
  assign N1582 = ~pe_o_4__4_;
  assign N1583 = ~pe_o_4__0_;
  assign N2855 = pe_o_4__5_ & pe_o_4__3_ & (pe_o_4__2_ & pe_o_4__0_) & pe_o_4__1_;
  assign N1584 = pe_o_4__5_ & pe_o_4__4_;
  assign N1585 = N1584 & N1588;
  assign N1586 = N1585 & N1589;
  assign N1587 = N1586 & N1590;
  assign N2857 = N1587 & N1591;
  assign N1588 = ~pe_o_4__3_;
  assign N1589 = ~pe_o_4__2_;
  assign N1590 = ~pe_o_4__0_;
  assign N1591 = ~pe_o_4__1_;
  assign N1592 = pe_o_4__5_ & pe_o_4__4_;
  assign N1593 = N1592 & N1596;
  assign N1594 = N1593 & N1597;
  assign N1595 = N1594 & pe_o_4__0_;
  assign N2859 = N1595 & N1598;
  assign N1596 = ~pe_o_4__3_;
  assign N1597 = ~pe_o_4__2_;
  assign N1598 = ~pe_o_4__1_;
  assign N1599 = pe_o_4__5_ & pe_o_4__4_;
  assign N1600 = N1599 & N1603;
  assign N1601 = N1600 & N1604;
  assign N1602 = N1601 & N1605;
  assign N2861 = N1602 & pe_o_4__1_;
  assign N1603 = ~pe_o_4__3_;
  assign N1604 = ~pe_o_4__2_;
  assign N1605 = ~pe_o_4__0_;
  assign N1606 = pe_o_4__5_ & pe_o_4__4_;
  assign N1607 = N1606 & N1610;
  assign N1608 = N1607 & N1611;
  assign N1609 = N1608 & pe_o_4__0_;
  assign N2863 = N1609 & pe_o_4__1_;
  assign N1610 = ~pe_o_4__3_;
  assign N1611 = ~pe_o_4__2_;
  assign N1612 = pe_o_4__5_ & pe_o_4__4_;
  assign N1613 = N1612 & N1616;
  assign N1614 = N1613 & pe_o_4__2_;
  assign N1615 = N1614 & N1617;
  assign N2865 = N1615 & N1618;
  assign N1616 = ~pe_o_4__3_;
  assign N1617 = ~pe_o_4__0_;
  assign N1618 = ~pe_o_4__1_;
  assign N1619 = pe_o_4__5_ & pe_o_4__4_;
  assign N1620 = N1619 & N1623;
  assign N1621 = N1620 & pe_o_4__2_;
  assign N1622 = N1621 & pe_o_4__0_;
  assign N2867 = N1622 & N1624;
  assign N1623 = ~pe_o_4__3_;
  assign N1624 = ~pe_o_4__1_;
  assign N1625 = pe_o_4__5_ & pe_o_4__4_;
  assign N1626 = N1625 & N1629;
  assign N1627 = N1626 & pe_o_4__2_;
  assign N1628 = N1627 & N1630;
  assign N2869 = N1628 & pe_o_4__1_;
  assign N1629 = ~pe_o_4__3_;
  assign N1630 = ~pe_o_4__0_;
  assign N2871 = pe_o_4__5_ & pe_o_4__4_ & (pe_o_4__2_ & pe_o_4__0_) & pe_o_4__1_;
  assign N1631 = pe_o_4__5_ & pe_o_4__4_;
  assign N1632 = N1631 & pe_o_4__3_;
  assign N1633 = N1632 & N1635;
  assign N1634 = N1633 & N1636;
  assign N2873 = N1634 & N1637;
  assign N1635 = ~pe_o_4__2_;
  assign N1636 = ~pe_o_4__0_;
  assign N1637 = ~pe_o_4__1_;
  assign N1638 = pe_o_4__5_ & pe_o_4__4_;
  assign N1639 = N1638 & pe_o_4__3_;
  assign N1640 = N1639 & N1642;
  assign N1641 = N1640 & pe_o_4__0_;
  assign N2875 = N1641 & N1643;
  assign N1642 = ~pe_o_4__2_;
  assign N1643 = ~pe_o_4__1_;
  assign N1644 = pe_o_4__5_ & pe_o_4__4_;
  assign N1645 = N1644 & pe_o_4__3_;
  assign N1646 = N1645 & N1648;
  assign N1647 = N1646 & N1649;
  assign N2877 = N1647 & pe_o_4__1_;
  assign N1648 = ~pe_o_4__2_;
  assign N1649 = ~pe_o_4__0_;
  assign N2879 = pe_o_4__5_ & pe_o_4__4_ & (pe_o_4__3_ & pe_o_4__0_) & pe_o_4__1_;
  assign N1650 = pe_o_4__5_ & pe_o_4__4_;
  assign N1651 = N1650 & pe_o_4__3_;
  assign N1652 = N1651 & pe_o_4__2_;
  assign N1653 = N1652 & N1654;
  assign N2881 = N1653 & N1655;
  assign N1654 = ~pe_o_4__0_;
  assign N1655 = ~pe_o_4__1_;
  assign N2883 = pe_o_4__5_ & pe_o_4__4_ & (pe_o_4__3_ & pe_o_4__2_) & pe_o_4__0_;
  assign N2885 = pe_o_4__5_ & pe_o_4__4_ & (pe_o_4__3_ & pe_o_4__2_) & pe_o_4__1_;
  assign N1656 = N1660 & N1661;
  assign N1657 = N1656 & N1662;
  assign N1658 = N1657 & N1663;
  assign N1659 = N1658 & N1664;
  assign N2950 = N1659 & N1665;
  assign N1660 = ~pe_o_5__5_;
  assign N1661 = ~pe_o_5__4_;
  assign N1662 = ~pe_o_5__3_;
  assign N1663 = ~pe_o_5__2_;
  assign N1664 = ~pe_o_5__0_;
  assign N1665 = ~pe_o_5__1_;
  assign N1666 = pe_o_5__5_ & N1670;
  assign N1667 = N1666 & N1671;
  assign N1668 = N1667 & N1672;
  assign N1669 = N1668 & N1673;
  assign N2951 = N1669 & N1674;
  assign N1670 = ~pe_o_5__4_;
  assign N1671 = ~pe_o_5__3_;
  assign N1672 = ~pe_o_5__2_;
  assign N1673 = ~pe_o_5__0_;
  assign N1674 = ~pe_o_5__1_;
  assign N1675 = N1679 & N1680;
  assign N1676 = N1675 & N1681;
  assign N1677 = N1676 & N1682;
  assign N1678 = N1677 & pe_o_5__0_;
  assign N2952 = N1678 & N1683;
  assign N1679 = ~pe_o_5__5_;
  assign N1680 = ~pe_o_5__4_;
  assign N1681 = ~pe_o_5__3_;
  assign N1682 = ~pe_o_5__2_;
  assign N1683 = ~pe_o_5__1_;
  assign N1684 = N1688 & N1689;
  assign N1685 = N1684 & N1690;
  assign N1686 = N1685 & N1691;
  assign N1687 = N1686 & N1692;
  assign N2954 = N1687 & pe_o_5__1_;
  assign N1688 = ~pe_o_5__5_;
  assign N1689 = ~pe_o_5__4_;
  assign N1690 = ~pe_o_5__3_;
  assign N1691 = ~pe_o_5__2_;
  assign N1692 = ~pe_o_5__0_;
  assign N1693 = N1697 & N1698;
  assign N1694 = N1693 & N1699;
  assign N1695 = N1694 & N1700;
  assign N1696 = N1695 & pe_o_5__0_;
  assign N2956 = N1696 & pe_o_5__1_;
  assign N1697 = ~pe_o_5__5_;
  assign N1698 = ~pe_o_5__4_;
  assign N1699 = ~pe_o_5__3_;
  assign N1700 = ~pe_o_5__2_;
  assign N1701 = N1705 & N1706;
  assign N1702 = N1701 & N1707;
  assign N1703 = N1702 & pe_o_5__2_;
  assign N1704 = N1703 & N1708;
  assign N2958 = N1704 & N1709;
  assign N1705 = ~pe_o_5__5_;
  assign N1706 = ~pe_o_5__4_;
  assign N1707 = ~pe_o_5__3_;
  assign N1708 = ~pe_o_5__0_;
  assign N1709 = ~pe_o_5__1_;
  assign N1710 = N1714 & N1715;
  assign N1711 = N1710 & N1716;
  assign N1712 = N1711 & pe_o_5__2_;
  assign N1713 = N1712 & pe_o_5__0_;
  assign N2960 = N1713 & N1717;
  assign N1714 = ~pe_o_5__5_;
  assign N1715 = ~pe_o_5__4_;
  assign N1716 = ~pe_o_5__3_;
  assign N1717 = ~pe_o_5__1_;
  assign N1718 = N1722 & N1723;
  assign N1719 = N1718 & N1724;
  assign N1720 = N1719 & pe_o_5__2_;
  assign N1721 = N1720 & N1725;
  assign N2962 = N1721 & pe_o_5__1_;
  assign N1722 = ~pe_o_5__5_;
  assign N1723 = ~pe_o_5__4_;
  assign N1724 = ~pe_o_5__3_;
  assign N1725 = ~pe_o_5__0_;
  assign N1726 = N1730 & N1731;
  assign N1727 = N1726 & N1732;
  assign N1728 = N1727 & pe_o_5__2_;
  assign N1729 = N1728 & pe_o_5__0_;
  assign N2964 = N1729 & pe_o_5__1_;
  assign N1730 = ~pe_o_5__5_;
  assign N1731 = ~pe_o_5__4_;
  assign N1732 = ~pe_o_5__3_;
  assign N1733 = N1737 & N1738;
  assign N1734 = N1733 & pe_o_5__3_;
  assign N1735 = N1734 & N1739;
  assign N1736 = N1735 & N1740;
  assign N2966 = N1736 & N1741;
  assign N1737 = ~pe_o_5__5_;
  assign N1738 = ~pe_o_5__4_;
  assign N1739 = ~pe_o_5__2_;
  assign N1740 = ~pe_o_5__0_;
  assign N1741 = ~pe_o_5__1_;
  assign N1742 = N1746 & N1747;
  assign N1743 = N1742 & pe_o_5__3_;
  assign N1744 = N1743 & N1748;
  assign N1745 = N1744 & pe_o_5__0_;
  assign N2968 = N1745 & N1749;
  assign N1746 = ~pe_o_5__5_;
  assign N1747 = ~pe_o_5__4_;
  assign N1748 = ~pe_o_5__2_;
  assign N1749 = ~pe_o_5__1_;
  assign N1750 = N1754 & N1755;
  assign N1751 = N1750 & pe_o_5__3_;
  assign N1752 = N1751 & N1756;
  assign N1753 = N1752 & N1757;
  assign N2970 = N1753 & pe_o_5__1_;
  assign N1754 = ~pe_o_5__5_;
  assign N1755 = ~pe_o_5__4_;
  assign N1756 = ~pe_o_5__2_;
  assign N1757 = ~pe_o_5__0_;
  assign N1758 = N1762 & N1763;
  assign N1759 = N1758 & pe_o_5__3_;
  assign N1760 = N1759 & N1764;
  assign N1761 = N1760 & pe_o_5__0_;
  assign N2972 = N1761 & pe_o_5__1_;
  assign N1762 = ~pe_o_5__5_;
  assign N1763 = ~pe_o_5__4_;
  assign N1764 = ~pe_o_5__2_;
  assign N1765 = N1769 & N1770;
  assign N1766 = N1765 & pe_o_5__3_;
  assign N1767 = N1766 & pe_o_5__2_;
  assign N1768 = N1767 & N1771;
  assign N2974 = N1768 & N1772;
  assign N1769 = ~pe_o_5__5_;
  assign N1770 = ~pe_o_5__4_;
  assign N1771 = ~pe_o_5__0_;
  assign N1772 = ~pe_o_5__1_;
  assign N1773 = N1777 & N1778;
  assign N1774 = N1773 & pe_o_5__3_;
  assign N1775 = N1774 & pe_o_5__2_;
  assign N1776 = N1775 & pe_o_5__0_;
  assign N2976 = N1776 & N1779;
  assign N1777 = ~pe_o_5__5_;
  assign N1778 = ~pe_o_5__4_;
  assign N1779 = ~pe_o_5__1_;
  assign N1780 = N1784 & N1785;
  assign N1781 = N1780 & pe_o_5__3_;
  assign N1782 = N1781 & pe_o_5__2_;
  assign N1783 = N1782 & N1786;
  assign N2978 = N1783 & pe_o_5__1_;
  assign N1784 = ~pe_o_5__5_;
  assign N1785 = ~pe_o_5__4_;
  assign N1786 = ~pe_o_5__0_;
  assign N1787 = N1791 & N1792;
  assign N1788 = N1787 & pe_o_5__3_;
  assign N1789 = N1788 & pe_o_5__2_;
  assign N1790 = N1789 & pe_o_5__0_;
  assign N2980 = N1790 & pe_o_5__1_;
  assign N1791 = ~pe_o_5__5_;
  assign N1792 = ~pe_o_5__4_;
  assign N1793 = N1797 & pe_o_5__4_;
  assign N1794 = N1793 & N1798;
  assign N1795 = N1794 & N1799;
  assign N1796 = N1795 & N1800;
  assign N2982 = N1796 & N1801;
  assign N1797 = ~pe_o_5__5_;
  assign N1798 = ~pe_o_5__3_;
  assign N1799 = ~pe_o_5__2_;
  assign N1800 = ~pe_o_5__0_;
  assign N1801 = ~pe_o_5__1_;
  assign N1802 = N1806 & pe_o_5__4_;
  assign N1803 = N1802 & N1807;
  assign N1804 = N1803 & N1808;
  assign N1805 = N1804 & pe_o_5__0_;
  assign N2984 = N1805 & N1809;
  assign N1806 = ~pe_o_5__5_;
  assign N1807 = ~pe_o_5__3_;
  assign N1808 = ~pe_o_5__2_;
  assign N1809 = ~pe_o_5__1_;
  assign N1810 = N1814 & pe_o_5__4_;
  assign N1811 = N1810 & N1815;
  assign N1812 = N1811 & N1816;
  assign N1813 = N1812 & N1817;
  assign N2986 = N1813 & pe_o_5__1_;
  assign N1814 = ~pe_o_5__5_;
  assign N1815 = ~pe_o_5__3_;
  assign N1816 = ~pe_o_5__2_;
  assign N1817 = ~pe_o_5__0_;
  assign N1818 = N1822 & pe_o_5__4_;
  assign N1819 = N1818 & N1823;
  assign N1820 = N1819 & N1824;
  assign N1821 = N1820 & pe_o_5__0_;
  assign N2988 = N1821 & pe_o_5__1_;
  assign N1822 = ~pe_o_5__5_;
  assign N1823 = ~pe_o_5__3_;
  assign N1824 = ~pe_o_5__2_;
  assign N1825 = N1829 & pe_o_5__4_;
  assign N1826 = N1825 & N1830;
  assign N1827 = N1826 & pe_o_5__2_;
  assign N1828 = N1827 & N1831;
  assign N2990 = N1828 & N1832;
  assign N1829 = ~pe_o_5__5_;
  assign N1830 = ~pe_o_5__3_;
  assign N1831 = ~pe_o_5__0_;
  assign N1832 = ~pe_o_5__1_;
  assign N1833 = N1837 & pe_o_5__4_;
  assign N1834 = N1833 & N1838;
  assign N1835 = N1834 & pe_o_5__2_;
  assign N1836 = N1835 & pe_o_5__0_;
  assign N2992 = N1836 & N1839;
  assign N1837 = ~pe_o_5__5_;
  assign N1838 = ~pe_o_5__3_;
  assign N1839 = ~pe_o_5__1_;
  assign N1840 = N1844 & pe_o_5__4_;
  assign N1841 = N1840 & N1845;
  assign N1842 = N1841 & pe_o_5__2_;
  assign N1843 = N1842 & N1846;
  assign N2994 = N1843 & pe_o_5__1_;
  assign N1844 = ~pe_o_5__5_;
  assign N1845 = ~pe_o_5__3_;
  assign N1846 = ~pe_o_5__0_;
  assign N1847 = N1851 & pe_o_5__4_;
  assign N1848 = N1847 & N1852;
  assign N1849 = N1848 & pe_o_5__2_;
  assign N1850 = N1849 & pe_o_5__0_;
  assign N2996 = N1850 & pe_o_5__1_;
  assign N1851 = ~pe_o_5__5_;
  assign N1852 = ~pe_o_5__3_;
  assign N1853 = N1857 & pe_o_5__4_;
  assign N1854 = N1853 & pe_o_5__3_;
  assign N1855 = N1854 & N1858;
  assign N1856 = N1855 & N1859;
  assign N2998 = N1856 & N1860;
  assign N1857 = ~pe_o_5__5_;
  assign N1858 = ~pe_o_5__2_;
  assign N1859 = ~pe_o_5__0_;
  assign N1860 = ~pe_o_5__1_;
  assign N1861 = N1865 & pe_o_5__4_;
  assign N1862 = N1861 & pe_o_5__3_;
  assign N1863 = N1862 & N1866;
  assign N1864 = N1863 & pe_o_5__0_;
  assign N3000 = N1864 & N1867;
  assign N1865 = ~pe_o_5__5_;
  assign N1866 = ~pe_o_5__2_;
  assign N1867 = ~pe_o_5__1_;
  assign N1868 = N1872 & pe_o_5__4_;
  assign N1869 = N1868 & pe_o_5__3_;
  assign N1870 = N1869 & N1873;
  assign N1871 = N1870 & N1874;
  assign N3002 = N1871 & pe_o_5__1_;
  assign N1872 = ~pe_o_5__5_;
  assign N1873 = ~pe_o_5__2_;
  assign N1874 = ~pe_o_5__0_;
  assign N1875 = N1879 & pe_o_5__4_;
  assign N1876 = N1875 & pe_o_5__3_;
  assign N1877 = N1876 & N1880;
  assign N1878 = N1877 & pe_o_5__0_;
  assign N3004 = N1878 & pe_o_5__1_;
  assign N1879 = ~pe_o_5__5_;
  assign N1880 = ~pe_o_5__2_;
  assign N1881 = N1885 & pe_o_5__4_;
  assign N1882 = N1881 & pe_o_5__3_;
  assign N1883 = N1882 & pe_o_5__2_;
  assign N1884 = N1883 & N1886;
  assign N3006 = N1884 & N1887;
  assign N1885 = ~pe_o_5__5_;
  assign N1886 = ~pe_o_5__0_;
  assign N1887 = ~pe_o_5__1_;
  assign N1888 = N1892 & pe_o_5__4_;
  assign N1889 = N1888 & pe_o_5__3_;
  assign N1890 = N1889 & pe_o_5__2_;
  assign N1891 = N1890 & pe_o_5__0_;
  assign N3008 = N1891 & N1893;
  assign N1892 = ~pe_o_5__5_;
  assign N1893 = ~pe_o_5__1_;
  assign N1894 = N1898 & pe_o_5__4_;
  assign N1895 = N1894 & pe_o_5__3_;
  assign N1896 = N1895 & pe_o_5__2_;
  assign N1897 = N1896 & N1899;
  assign N3010 = N1897 & pe_o_5__1_;
  assign N1898 = ~pe_o_5__5_;
  assign N1899 = ~pe_o_5__0_;
  assign N3012 = pe_o_5__4_ & pe_o_5__3_ & (pe_o_5__2_ & pe_o_5__0_) & pe_o_5__1_;
  assign N1900 = pe_o_5__5_ & N1904;
  assign N1901 = N1900 & N1905;
  assign N1902 = N1901 & N1906;
  assign N1903 = N1902 & pe_o_5__0_;
  assign N2953 = N1903 & N1907;
  assign N1904 = ~pe_o_5__4_;
  assign N1905 = ~pe_o_5__3_;
  assign N1906 = ~pe_o_5__2_;
  assign N1907 = ~pe_o_5__1_;
  assign N1908 = pe_o_5__5_ & N1912;
  assign N1909 = N1908 & N1913;
  assign N1910 = N1909 & N1914;
  assign N1911 = N1910 & N1915;
  assign N2955 = N1911 & pe_o_5__1_;
  assign N1912 = ~pe_o_5__4_;
  assign N1913 = ~pe_o_5__3_;
  assign N1914 = ~pe_o_5__2_;
  assign N1915 = ~pe_o_5__0_;
  assign N1916 = pe_o_5__5_ & N1920;
  assign N1917 = N1916 & N1921;
  assign N1918 = N1917 & N1922;
  assign N1919 = N1918 & pe_o_5__0_;
  assign N2957 = N1919 & pe_o_5__1_;
  assign N1920 = ~pe_o_5__4_;
  assign N1921 = ~pe_o_5__3_;
  assign N1922 = ~pe_o_5__2_;
  assign N1923 = pe_o_5__5_ & N1927;
  assign N1924 = N1923 & N1928;
  assign N1925 = N1924 & pe_o_5__2_;
  assign N1926 = N1925 & N1929;
  assign N2959 = N1926 & N1930;
  assign N1927 = ~pe_o_5__4_;
  assign N1928 = ~pe_o_5__3_;
  assign N1929 = ~pe_o_5__0_;
  assign N1930 = ~pe_o_5__1_;
  assign N1931 = pe_o_5__5_ & N1935;
  assign N1932 = N1931 & N1936;
  assign N1933 = N1932 & pe_o_5__2_;
  assign N1934 = N1933 & pe_o_5__0_;
  assign N2961 = N1934 & N1937;
  assign N1935 = ~pe_o_5__4_;
  assign N1936 = ~pe_o_5__3_;
  assign N1937 = ~pe_o_5__1_;
  assign N1938 = pe_o_5__5_ & N1942;
  assign N1939 = N1938 & N1943;
  assign N1940 = N1939 & pe_o_5__2_;
  assign N1941 = N1940 & N1944;
  assign N2963 = N1941 & pe_o_5__1_;
  assign N1942 = ~pe_o_5__4_;
  assign N1943 = ~pe_o_5__3_;
  assign N1944 = ~pe_o_5__0_;
  assign N1945 = pe_o_5__5_ & N1949;
  assign N1946 = N1945 & N1950;
  assign N1947 = N1946 & pe_o_5__2_;
  assign N1948 = N1947 & pe_o_5__0_;
  assign N2965 = N1948 & pe_o_5__1_;
  assign N1949 = ~pe_o_5__4_;
  assign N1950 = ~pe_o_5__3_;
  assign N1951 = pe_o_5__5_ & N1955;
  assign N1952 = N1951 & pe_o_5__3_;
  assign N1953 = N1952 & N1956;
  assign N1954 = N1953 & N1957;
  assign N2967 = N1954 & N1958;
  assign N1955 = ~pe_o_5__4_;
  assign N1956 = ~pe_o_5__2_;
  assign N1957 = ~pe_o_5__0_;
  assign N1958 = ~pe_o_5__1_;
  assign N1959 = pe_o_5__5_ & N1963;
  assign N1960 = N1959 & pe_o_5__3_;
  assign N1961 = N1960 & N1964;
  assign N1962 = N1961 & pe_o_5__0_;
  assign N2969 = N1962 & N1965;
  assign N1963 = ~pe_o_5__4_;
  assign N1964 = ~pe_o_5__2_;
  assign N1965 = ~pe_o_5__1_;
  assign N1966 = pe_o_5__5_ & N1970;
  assign N1967 = N1966 & pe_o_5__3_;
  assign N1968 = N1967 & N1971;
  assign N1969 = N1968 & N1972;
  assign N2971 = N1969 & pe_o_5__1_;
  assign N1970 = ~pe_o_5__4_;
  assign N1971 = ~pe_o_5__2_;
  assign N1972 = ~pe_o_5__0_;
  assign N1973 = pe_o_5__5_ & N1977;
  assign N1974 = N1973 & pe_o_5__3_;
  assign N1975 = N1974 & N1978;
  assign N1976 = N1975 & pe_o_5__0_;
  assign N2973 = N1976 & pe_o_5__1_;
  assign N1977 = ~pe_o_5__4_;
  assign N1978 = ~pe_o_5__2_;
  assign N1979 = pe_o_5__5_ & N1983;
  assign N1980 = N1979 & pe_o_5__3_;
  assign N1981 = N1980 & pe_o_5__2_;
  assign N1982 = N1981 & N1984;
  assign N2975 = N1982 & N1985;
  assign N1983 = ~pe_o_5__4_;
  assign N1984 = ~pe_o_5__0_;
  assign N1985 = ~pe_o_5__1_;
  assign N1986 = pe_o_5__5_ & N1990;
  assign N1987 = N1986 & pe_o_5__3_;
  assign N1988 = N1987 & pe_o_5__2_;
  assign N1989 = N1988 & pe_o_5__0_;
  assign N2977 = N1989 & N1991;
  assign N1990 = ~pe_o_5__4_;
  assign N1991 = ~pe_o_5__1_;
  assign N1992 = pe_o_5__5_ & N1996;
  assign N1993 = N1992 & pe_o_5__3_;
  assign N1994 = N1993 & pe_o_5__2_;
  assign N1995 = N1994 & N1997;
  assign N2979 = N1995 & pe_o_5__1_;
  assign N1996 = ~pe_o_5__4_;
  assign N1997 = ~pe_o_5__0_;
  assign N2981 = pe_o_5__5_ & pe_o_5__3_ & (pe_o_5__2_ & pe_o_5__0_) & pe_o_5__1_;
  assign N1998 = pe_o_5__5_ & pe_o_5__4_;
  assign N1999 = N1998 & N2002;
  assign N2000 = N1999 & N2003;
  assign N2001 = N2000 & N2004;
  assign N2983 = N2001 & N2005;
  assign N2002 = ~pe_o_5__3_;
  assign N2003 = ~pe_o_5__2_;
  assign N2004 = ~pe_o_5__0_;
  assign N2005 = ~pe_o_5__1_;
  assign N2006 = pe_o_5__5_ & pe_o_5__4_;
  assign N2007 = N2006 & N2010;
  assign N2008 = N2007 & N2011;
  assign N2009 = N2008 & pe_o_5__0_;
  assign N2985 = N2009 & N2012;
  assign N2010 = ~pe_o_5__3_;
  assign N2011 = ~pe_o_5__2_;
  assign N2012 = ~pe_o_5__1_;
  assign N2013 = pe_o_5__5_ & pe_o_5__4_;
  assign N2014 = N2013 & N2017;
  assign N2015 = N2014 & N2018;
  assign N2016 = N2015 & N2019;
  assign N2987 = N2016 & pe_o_5__1_;
  assign N2017 = ~pe_o_5__3_;
  assign N2018 = ~pe_o_5__2_;
  assign N2019 = ~pe_o_5__0_;
  assign N2020 = pe_o_5__5_ & pe_o_5__4_;
  assign N2021 = N2020 & N2024;
  assign N2022 = N2021 & N2025;
  assign N2023 = N2022 & pe_o_5__0_;
  assign N2989 = N2023 & pe_o_5__1_;
  assign N2024 = ~pe_o_5__3_;
  assign N2025 = ~pe_o_5__2_;
  assign N2026 = pe_o_5__5_ & pe_o_5__4_;
  assign N2027 = N2026 & N2030;
  assign N2028 = N2027 & pe_o_5__2_;
  assign N2029 = N2028 & N2031;
  assign N2991 = N2029 & N2032;
  assign N2030 = ~pe_o_5__3_;
  assign N2031 = ~pe_o_5__0_;
  assign N2032 = ~pe_o_5__1_;
  assign N2033 = pe_o_5__5_ & pe_o_5__4_;
  assign N2034 = N2033 & N2037;
  assign N2035 = N2034 & pe_o_5__2_;
  assign N2036 = N2035 & pe_o_5__0_;
  assign N2993 = N2036 & N2038;
  assign N2037 = ~pe_o_5__3_;
  assign N2038 = ~pe_o_5__1_;
  assign N2039 = pe_o_5__5_ & pe_o_5__4_;
  assign N2040 = N2039 & N2043;
  assign N2041 = N2040 & pe_o_5__2_;
  assign N2042 = N2041 & N2044;
  assign N2995 = N2042 & pe_o_5__1_;
  assign N2043 = ~pe_o_5__3_;
  assign N2044 = ~pe_o_5__0_;
  assign N2997 = pe_o_5__5_ & pe_o_5__4_ & (pe_o_5__2_ & pe_o_5__0_) & pe_o_5__1_;
  assign N2045 = pe_o_5__5_ & pe_o_5__4_;
  assign N2046 = N2045 & pe_o_5__3_;
  assign N2047 = N2046 & N2049;
  assign N2048 = N2047 & N2050;
  assign N2999 = N2048 & N2051;
  assign N2049 = ~pe_o_5__2_;
  assign N2050 = ~pe_o_5__0_;
  assign N2051 = ~pe_o_5__1_;
  assign N2052 = pe_o_5__5_ & pe_o_5__4_;
  assign N2053 = N2052 & pe_o_5__3_;
  assign N2054 = N2053 & N2056;
  assign N2055 = N2054 & pe_o_5__0_;
  assign N3001 = N2055 & N2057;
  assign N2056 = ~pe_o_5__2_;
  assign N2057 = ~pe_o_5__1_;
  assign N2058 = pe_o_5__5_ & pe_o_5__4_;
  assign N2059 = N2058 & pe_o_5__3_;
  assign N2060 = N2059 & N2062;
  assign N2061 = N2060 & N2063;
  assign N3003 = N2061 & pe_o_5__1_;
  assign N2062 = ~pe_o_5__2_;
  assign N2063 = ~pe_o_5__0_;
  assign N3005 = pe_o_5__5_ & pe_o_5__4_ & (pe_o_5__3_ & pe_o_5__0_) & pe_o_5__1_;
  assign N2064 = pe_o_5__5_ & pe_o_5__4_;
  assign N2065 = N2064 & pe_o_5__3_;
  assign N2066 = N2065 & pe_o_5__2_;
  assign N2067 = N2066 & N2068;
  assign N3007 = N2067 & N2069;
  assign N2068 = ~pe_o_5__0_;
  assign N2069 = ~pe_o_5__1_;
  assign N3009 = pe_o_5__5_ & pe_o_5__4_ & (pe_o_5__3_ & pe_o_5__2_) & pe_o_5__0_;
  assign N3011 = pe_o_5__5_ & pe_o_5__4_ & (pe_o_5__3_ & pe_o_5__2_) & pe_o_5__1_;
  assign way_id_o[4] = (N2070)? lru_i[0] : 
                       (N2071)? lru_i[1] : 
                       (N2072)? lru_i[2] : 
                       (N2073)? lru_i[3] : 
                       (N2074)? lru_i[4] : 
                       (N2075)? lru_i[5] : 
                       (N2076)? lru_i[6] : 
                       (N2077)? lru_i[7] : 
                       (N2078)? lru_i[8] : 
                       (N2079)? lru_i[9] : 
                       (N2080)? lru_i[10] : 
                       (N2081)? lru_i[11] : 
                       (N2082)? lru_i[12] : 
                       (N2083)? lru_i[13] : 
                       (N2084)? lru_i[14] : 
                       (N2085)? lru_i[15] : 
                       (N2086)? lru_i[16] : 
                       (N2087)? lru_i[17] : 
                       (N2088)? lru_i[18] : 
                       (N2089)? lru_i[19] : 
                       (N2090)? lru_i[20] : 
                       (N2091)? lru_i[21] : 
                       (N2092)? lru_i[22] : 
                       (N2093)? lru_i[23] : 
                       (N2094)? lru_i[24] : 
                       (N2095)? lru_i[25] : 
                       (N2096)? lru_i[26] : 
                       (N2097)? lru_i[27] : 
                       (N2098)? lru_i[28] : 
                       (N2099)? lru_i[29] : 
                       (N2100)? lru_i[30] : 
                       (N2101)? lru_i[31] : 
                       (N2102)? lru_i[32] : 
                       (N2103)? lru_i[33] : 
                       (N2104)? lru_i[34] : 
                       (N2105)? lru_i[35] : 
                       (N2106)? lru_i[36] : 
                       (N2107)? lru_i[37] : 
                       (N2108)? lru_i[38] : 
                       (N2109)? lru_i[39] : 
                       (N2110)? lru_i[40] : 
                       (N2111)? lru_i[41] : 
                       (N2112)? lru_i[42] : 
                       (N2113)? lru_i[43] : 
                       (N2114)? lru_i[44] : 
                       (N2115)? lru_i[45] : 
                       (N2116)? lru_i[46] : 
                       (N2117)? lru_i[47] : 
                       (N2118)? lru_i[48] : 
                       (N2119)? lru_i[49] : 
                       (N2120)? lru_i[50] : 
                       (N2121)? lru_i[51] : 
                       (N2122)? lru_i[52] : 
                       (N2123)? lru_i[53] : 
                       (N2124)? lru_i[54] : 
                       (N2125)? lru_i[55] : 
                       (N2126)? lru_i[56] : 
                       (N2127)? lru_i[57] : 
                       (N2128)? lru_i[58] : 
                       (N2129)? lru_i[59] : 
                       (N2130)? lru_i[60] : 
                       (N2131)? lru_i[61] : 
                       (N2132)? lru_i[62] : 1'b0;
  assign N2070 = N2509;
  assign N2071 = N2511;
  assign N2072 = N2513;
  assign N2073 = N2515;
  assign N2074 = N2517;
  assign N2075 = N2519;
  assign N2076 = N2521;
  assign N2077 = N2523;
  assign N2078 = N2525;
  assign N2079 = N2527;
  assign N2080 = N2529;
  assign N2081 = N2531;
  assign N2082 = N2533;
  assign N2083 = N2535;
  assign N2084 = N2537;
  assign N2085 = N2539;
  assign N2086 = N2541;
  assign N2087 = N2543;
  assign N2088 = N2545;
  assign N2089 = N2547;
  assign N2090 = N2549;
  assign N2091 = N2551;
  assign N2092 = N2553;
  assign N2093 = N2555;
  assign N2094 = N2557;
  assign N2095 = N2559;
  assign N2096 = N2561;
  assign N2097 = N2563;
  assign N2098 = N2565;
  assign N2099 = N2567;
  assign N2100 = N2569;
  assign N2101 = N2571;
  assign N2102 = N2510;
  assign N2103 = N2512;
  assign N2104 = N2514;
  assign N2105 = N2516;
  assign N2106 = N2518;
  assign N2107 = N2520;
  assign N2108 = N2522;
  assign N2109 = N2524;
  assign N2110 = N2526;
  assign N2111 = N2528;
  assign N2112 = N2530;
  assign N2113 = N2532;
  assign N2114 = N2534;
  assign N2115 = N2536;
  assign N2116 = N2538;
  assign N2117 = N2540;
  assign N2118 = N2542;
  assign N2119 = N2544;
  assign N2120 = N2546;
  assign N2121 = N2548;
  assign N2122 = N2550;
  assign N2123 = N2552;
  assign N2124 = N2554;
  assign N2125 = N2556;
  assign N2126 = N2558;
  assign N2127 = N2560;
  assign N2128 = N2562;
  assign N2129 = N2564;
  assign N2130 = N2566;
  assign N2131 = N2568;
  assign N2132 = N2570;
  assign way_id_o[3] = (N2133)? lru_i[0] : 
                       (N2134)? lru_i[1] : 
                       (N2135)? lru_i[2] : 
                       (N2136)? lru_i[3] : 
                       (N2137)? lru_i[4] : 
                       (N2138)? lru_i[5] : 
                       (N2139)? lru_i[6] : 
                       (N2140)? lru_i[7] : 
                       (N2141)? lru_i[8] : 
                       (N2142)? lru_i[9] : 
                       (N2143)? lru_i[10] : 
                       (N2144)? lru_i[11] : 
                       (N2145)? lru_i[12] : 
                       (N2146)? lru_i[13] : 
                       (N2147)? lru_i[14] : 
                       (N2148)? lru_i[15] : 
                       (N2149)? lru_i[16] : 
                       (N2150)? lru_i[17] : 
                       (N2151)? lru_i[18] : 
                       (N2152)? lru_i[19] : 
                       (N2153)? lru_i[20] : 
                       (N2154)? lru_i[21] : 
                       (N2155)? lru_i[22] : 
                       (N2156)? lru_i[23] : 
                       (N2157)? lru_i[24] : 
                       (N2158)? lru_i[25] : 
                       (N2159)? lru_i[26] : 
                       (N2160)? lru_i[27] : 
                       (N2161)? lru_i[28] : 
                       (N2162)? lru_i[29] : 
                       (N2163)? lru_i[30] : 
                       (N2164)? lru_i[31] : 
                       (N2165)? lru_i[32] : 
                       (N2166)? lru_i[33] : 
                       (N2167)? lru_i[34] : 
                       (N2168)? lru_i[35] : 
                       (N2169)? lru_i[36] : 
                       (N2170)? lru_i[37] : 
                       (N2171)? lru_i[38] : 
                       (N2172)? lru_i[39] : 
                       (N2173)? lru_i[40] : 
                       (N2174)? lru_i[41] : 
                       (N2175)? lru_i[42] : 
                       (N2176)? lru_i[43] : 
                       (N2177)? lru_i[44] : 
                       (N2178)? lru_i[45] : 
                       (N2179)? lru_i[46] : 
                       (N2180)? lru_i[47] : 
                       (N2181)? lru_i[48] : 
                       (N2182)? lru_i[49] : 
                       (N2183)? lru_i[50] : 
                       (N2184)? lru_i[51] : 
                       (N2185)? lru_i[52] : 
                       (N2186)? lru_i[53] : 
                       (N2187)? lru_i[54] : 
                       (N2188)? lru_i[55] : 
                       (N2189)? lru_i[56] : 
                       (N2190)? lru_i[57] : 
                       (N2191)? lru_i[58] : 
                       (N2192)? lru_i[59] : 
                       (N2193)? lru_i[60] : 
                       (N2194)? lru_i[61] : 
                       (N2195)? lru_i[62] : 1'b0;
  assign N2133 = N2572;
  assign N2134 = N2574;
  assign N2135 = N2576;
  assign N2136 = N2578;
  assign N2137 = N2580;
  assign N2138 = N2582;
  assign N2139 = N2584;
  assign N2140 = N2586;
  assign N2141 = N2588;
  assign N2142 = N2590;
  assign N2143 = N2592;
  assign N2144 = N2594;
  assign N2145 = N2596;
  assign N2146 = N2598;
  assign N2147 = N2600;
  assign N2148 = N2602;
  assign N2149 = N2604;
  assign N2150 = N2606;
  assign N2151 = N2608;
  assign N2152 = N2610;
  assign N2153 = N2612;
  assign N2154 = N2614;
  assign N2155 = N2616;
  assign N2156 = N2618;
  assign N2157 = N2620;
  assign N2158 = N2622;
  assign N2159 = N2624;
  assign N2160 = N2626;
  assign N2161 = N2628;
  assign N2162 = N2630;
  assign N2163 = N2632;
  assign N2164 = N2634;
  assign N2165 = N2573;
  assign N2166 = N2575;
  assign N2167 = N2577;
  assign N2168 = N2579;
  assign N2169 = N2581;
  assign N2170 = N2583;
  assign N2171 = N2585;
  assign N2172 = N2587;
  assign N2173 = N2589;
  assign N2174 = N2591;
  assign N2175 = N2593;
  assign N2176 = N2595;
  assign N2177 = N2597;
  assign N2178 = N2599;
  assign N2179 = N2601;
  assign N2180 = N2603;
  assign N2181 = N2605;
  assign N2182 = N2607;
  assign N2183 = N2609;
  assign N2184 = N2611;
  assign N2185 = N2613;
  assign N2186 = N2615;
  assign N2187 = N2617;
  assign N2188 = N2619;
  assign N2189 = N2621;
  assign N2190 = N2623;
  assign N2191 = N2625;
  assign N2192 = N2627;
  assign N2193 = N2629;
  assign N2194 = N2631;
  assign N2195 = N2633;
  assign way_id_o[2] = (N2196)? lru_i[0] : 
                       (N2197)? lru_i[1] : 
                       (N2198)? lru_i[2] : 
                       (N2199)? lru_i[3] : 
                       (N2200)? lru_i[4] : 
                       (N2201)? lru_i[5] : 
                       (N2202)? lru_i[6] : 
                       (N2203)? lru_i[7] : 
                       (N2204)? lru_i[8] : 
                       (N2205)? lru_i[9] : 
                       (N2206)? lru_i[10] : 
                       (N2207)? lru_i[11] : 
                       (N2208)? lru_i[12] : 
                       (N2209)? lru_i[13] : 
                       (N2210)? lru_i[14] : 
                       (N2211)? lru_i[15] : 
                       (N2212)? lru_i[16] : 
                       (N2213)? lru_i[17] : 
                       (N2214)? lru_i[18] : 
                       (N2215)? lru_i[19] : 
                       (N2216)? lru_i[20] : 
                       (N2217)? lru_i[21] : 
                       (N2218)? lru_i[22] : 
                       (N2219)? lru_i[23] : 
                       (N2220)? lru_i[24] : 
                       (N2221)? lru_i[25] : 
                       (N2222)? lru_i[26] : 
                       (N2223)? lru_i[27] : 
                       (N2224)? lru_i[28] : 
                       (N2225)? lru_i[29] : 
                       (N2226)? lru_i[30] : 
                       (N2227)? lru_i[31] : 
                       (N2228)? lru_i[32] : 
                       (N2229)? lru_i[33] : 
                       (N2230)? lru_i[34] : 
                       (N2231)? lru_i[35] : 
                       (N2232)? lru_i[36] : 
                       (N2233)? lru_i[37] : 
                       (N2234)? lru_i[38] : 
                       (N2235)? lru_i[39] : 
                       (N2236)? lru_i[40] : 
                       (N2237)? lru_i[41] : 
                       (N2238)? lru_i[42] : 
                       (N2239)? lru_i[43] : 
                       (N2240)? lru_i[44] : 
                       (N2241)? lru_i[45] : 
                       (N2242)? lru_i[46] : 
                       (N2243)? lru_i[47] : 
                       (N2244)? lru_i[48] : 
                       (N2245)? lru_i[49] : 
                       (N2246)? lru_i[50] : 
                       (N2247)? lru_i[51] : 
                       (N2248)? lru_i[52] : 
                       (N2249)? lru_i[53] : 
                       (N2250)? lru_i[54] : 
                       (N2251)? lru_i[55] : 
                       (N2252)? lru_i[56] : 
                       (N2253)? lru_i[57] : 
                       (N2254)? lru_i[58] : 
                       (N2255)? lru_i[59] : 
                       (N2256)? lru_i[60] : 
                       (N2257)? lru_i[61] : 
                       (N2258)? lru_i[62] : 1'b0;
  assign N2196 = N2698;
  assign N2197 = N2700;
  assign N2198 = N2702;
  assign N2199 = N2704;
  assign N2200 = N2706;
  assign N2201 = N2708;
  assign N2202 = N2710;
  assign N2203 = N2712;
  assign N2204 = N2714;
  assign N2205 = N2716;
  assign N2206 = N2718;
  assign N2207 = N2720;
  assign N2208 = N2722;
  assign N2209 = N2724;
  assign N2210 = N2726;
  assign N2211 = N2728;
  assign N2212 = N2730;
  assign N2213 = N2732;
  assign N2214 = N2734;
  assign N2215 = N2736;
  assign N2216 = N2738;
  assign N2217 = N2740;
  assign N2218 = N2742;
  assign N2219 = N2744;
  assign N2220 = N2746;
  assign N2221 = N2748;
  assign N2222 = N2750;
  assign N2223 = N2752;
  assign N2224 = N2754;
  assign N2225 = N2756;
  assign N2226 = N2758;
  assign N2227 = N2760;
  assign N2228 = N2699;
  assign N2229 = N2701;
  assign N2230 = N2703;
  assign N2231 = N2705;
  assign N2232 = N2707;
  assign N2233 = N2709;
  assign N2234 = N2711;
  assign N2235 = N2713;
  assign N2236 = N2715;
  assign N2237 = N2717;
  assign N2238 = N2719;
  assign N2239 = N2721;
  assign N2240 = N2723;
  assign N2241 = N2725;
  assign N2242 = N2727;
  assign N2243 = N2729;
  assign N2244 = N2731;
  assign N2245 = N2733;
  assign N2246 = N2735;
  assign N2247 = N2737;
  assign N2248 = N2739;
  assign N2249 = N2741;
  assign N2250 = N2743;
  assign N2251 = N2745;
  assign N2252 = N2747;
  assign N2253 = N2749;
  assign N2254 = N2751;
  assign N2255 = N2753;
  assign N2256 = N2755;
  assign N2257 = N2757;
  assign N2258 = N2759;
  assign way_id_o[1] = (N2259)? lru_i[0] : 
                       (N2260)? lru_i[1] : 
                       (N2261)? lru_i[2] : 
                       (N2262)? lru_i[3] : 
                       (N2263)? lru_i[4] : 
                       (N2264)? lru_i[5] : 
                       (N2265)? lru_i[6] : 
                       (N2266)? lru_i[7] : 
                       (N2267)? lru_i[8] : 
                       (N2268)? lru_i[9] : 
                       (N2269)? lru_i[10] : 
                       (N2270)? lru_i[11] : 
                       (N2271)? lru_i[12] : 
                       (N2272)? lru_i[13] : 
                       (N2273)? lru_i[14] : 
                       (N2274)? lru_i[15] : 
                       (N2275)? lru_i[16] : 
                       (N2276)? lru_i[17] : 
                       (N2277)? lru_i[18] : 
                       (N2278)? lru_i[19] : 
                       (N2279)? lru_i[20] : 
                       (N2280)? lru_i[21] : 
                       (N2281)? lru_i[22] : 
                       (N2282)? lru_i[23] : 
                       (N2283)? lru_i[24] : 
                       (N2284)? lru_i[25] : 
                       (N2285)? lru_i[26] : 
                       (N2286)? lru_i[27] : 
                       (N2287)? lru_i[28] : 
                       (N2288)? lru_i[29] : 
                       (N2289)? lru_i[30] : 
                       (N2290)? lru_i[31] : 
                       (N2291)? lru_i[32] : 
                       (N2292)? lru_i[33] : 
                       (N2293)? lru_i[34] : 
                       (N2294)? lru_i[35] : 
                       (N2295)? lru_i[36] : 
                       (N2296)? lru_i[37] : 
                       (N2297)? lru_i[38] : 
                       (N2298)? lru_i[39] : 
                       (N2299)? lru_i[40] : 
                       (N2300)? lru_i[41] : 
                       (N2301)? lru_i[42] : 
                       (N2302)? lru_i[43] : 
                       (N2303)? lru_i[44] : 
                       (N2304)? lru_i[45] : 
                       (N2305)? lru_i[46] : 
                       (N2306)? lru_i[47] : 
                       (N2307)? lru_i[48] : 
                       (N2308)? lru_i[49] : 
                       (N2309)? lru_i[50] : 
                       (N2310)? lru_i[51] : 
                       (N2311)? lru_i[52] : 
                       (N2312)? lru_i[53] : 
                       (N2313)? lru_i[54] : 
                       (N2314)? lru_i[55] : 
                       (N2315)? lru_i[56] : 
                       (N2316)? lru_i[57] : 
                       (N2317)? lru_i[58] : 
                       (N2318)? lru_i[59] : 
                       (N2319)? lru_i[60] : 
                       (N2320)? lru_i[61] : 
                       (N2321)? lru_i[62] : 1'b0;
  assign N2259 = N2824;
  assign N2260 = N2826;
  assign N2261 = N2828;
  assign N2262 = N2830;
  assign N2263 = N2832;
  assign N2264 = N2834;
  assign N2265 = N2836;
  assign N2266 = N2838;
  assign N2267 = N2840;
  assign N2268 = N2842;
  assign N2269 = N2844;
  assign N2270 = N2846;
  assign N2271 = N2848;
  assign N2272 = N2850;
  assign N2273 = N2852;
  assign N2274 = N2854;
  assign N2275 = N2856;
  assign N2276 = N2858;
  assign N2277 = N2860;
  assign N2278 = N2862;
  assign N2279 = N2864;
  assign N2280 = N2866;
  assign N2281 = N2868;
  assign N2282 = N2870;
  assign N2283 = N2872;
  assign N2284 = N2874;
  assign N2285 = N2876;
  assign N2286 = N2878;
  assign N2287 = N2880;
  assign N2288 = N2882;
  assign N2289 = N2884;
  assign N2290 = N2886;
  assign N2291 = N2825;
  assign N2292 = N2827;
  assign N2293 = N2829;
  assign N2294 = N2831;
  assign N2295 = N2833;
  assign N2296 = N2835;
  assign N2297 = N2837;
  assign N2298 = N2839;
  assign N2299 = N2841;
  assign N2300 = N2843;
  assign N2301 = N2845;
  assign N2302 = N2847;
  assign N2303 = N2849;
  assign N2304 = N2851;
  assign N2305 = N2853;
  assign N2306 = N2855;
  assign N2307 = N2857;
  assign N2308 = N2859;
  assign N2309 = N2861;
  assign N2310 = N2863;
  assign N2311 = N2865;
  assign N2312 = N2867;
  assign N2313 = N2869;
  assign N2314 = N2871;
  assign N2315 = N2873;
  assign N2316 = N2875;
  assign N2317 = N2877;
  assign N2318 = N2879;
  assign N2319 = N2881;
  assign N2320 = N2883;
  assign N2321 = N2885;
  assign way_id_o[0] = (N2322)? lru_i[0] : 
                       (N2323)? lru_i[1] : 
                       (N2324)? lru_i[2] : 
                       (N2325)? lru_i[3] : 
                       (N2326)? lru_i[4] : 
                       (N2327)? lru_i[5] : 
                       (N2328)? lru_i[6] : 
                       (N2329)? lru_i[7] : 
                       (N2330)? lru_i[8] : 
                       (N2331)? lru_i[9] : 
                       (N2332)? lru_i[10] : 
                       (N2333)? lru_i[11] : 
                       (N2334)? lru_i[12] : 
                       (N2335)? lru_i[13] : 
                       (N2336)? lru_i[14] : 
                       (N2337)? lru_i[15] : 
                       (N2338)? lru_i[16] : 
                       (N2339)? lru_i[17] : 
                       (N2340)? lru_i[18] : 
                       (N2341)? lru_i[19] : 
                       (N2342)? lru_i[20] : 
                       (N2343)? lru_i[21] : 
                       (N2344)? lru_i[22] : 
                       (N2345)? lru_i[23] : 
                       (N2346)? lru_i[24] : 
                       (N2347)? lru_i[25] : 
                       (N2348)? lru_i[26] : 
                       (N2349)? lru_i[27] : 
                       (N2350)? lru_i[28] : 
                       (N2351)? lru_i[29] : 
                       (N2352)? lru_i[30] : 
                       (N2353)? lru_i[31] : 
                       (N2354)? lru_i[32] : 
                       (N2355)? lru_i[33] : 
                       (N2356)? lru_i[34] : 
                       (N2357)? lru_i[35] : 
                       (N2358)? lru_i[36] : 
                       (N2359)? lru_i[37] : 
                       (N2360)? lru_i[38] : 
                       (N2361)? lru_i[39] : 
                       (N2362)? lru_i[40] : 
                       (N2363)? lru_i[41] : 
                       (N2364)? lru_i[42] : 
                       (N2365)? lru_i[43] : 
                       (N2366)? lru_i[44] : 
                       (N2367)? lru_i[45] : 
                       (N2368)? lru_i[46] : 
                       (N2369)? lru_i[47] : 
                       (N2370)? lru_i[48] : 
                       (N2371)? lru_i[49] : 
                       (N2372)? lru_i[50] : 
                       (N2373)? lru_i[51] : 
                       (N2374)? lru_i[52] : 
                       (N2375)? lru_i[53] : 
                       (N2376)? lru_i[54] : 
                       (N2377)? lru_i[55] : 
                       (N2378)? lru_i[56] : 
                       (N2379)? lru_i[57] : 
                       (N2380)? lru_i[58] : 
                       (N2381)? lru_i[59] : 
                       (N2382)? lru_i[60] : 
                       (N2383)? lru_i[61] : 
                       (N2384)? lru_i[62] : 1'b0;
  assign N2322 = N2950;
  assign N2323 = N2952;
  assign N2324 = N2954;
  assign N2325 = N2956;
  assign N2326 = N2958;
  assign N2327 = N2960;
  assign N2328 = N2962;
  assign N2329 = N2964;
  assign N2330 = N2966;
  assign N2331 = N2968;
  assign N2332 = N2970;
  assign N2333 = N2972;
  assign N2334 = N2974;
  assign N2335 = N2976;
  assign N2336 = N2978;
  assign N2337 = N2980;
  assign N2338 = N2982;
  assign N2339 = N2984;
  assign N2340 = N2986;
  assign N2341 = N2988;
  assign N2342 = N2990;
  assign N2343 = N2992;
  assign N2344 = N2994;
  assign N2345 = N2996;
  assign N2346 = N2998;
  assign N2347 = N3000;
  assign N2348 = N3002;
  assign N2349 = N3004;
  assign N2350 = N3006;
  assign N2351 = N3008;
  assign N2352 = N3010;
  assign N2353 = N3012;
  assign N2354 = N2951;
  assign N2355 = N2953;
  assign N2356 = N2955;
  assign N2357 = N2957;
  assign N2358 = N2959;
  assign N2359 = N2961;
  assign N2360 = N2963;
  assign N2361 = N2965;
  assign N2362 = N2967;
  assign N2363 = N2969;
  assign N2364 = N2971;
  assign N2365 = N2973;
  assign N2366 = N2975;
  assign N2367 = N2977;
  assign N2368 = N2979;
  assign N2369 = N2981;
  assign N2370 = N2983;
  assign N2371 = N2985;
  assign N2372 = N2987;
  assign N2373 = N2989;
  assign N2374 = N2991;
  assign N2375 = N2993;
  assign N2376 = N2995;
  assign N2377 = N2997;
  assign N2378 = N2999;
  assign N2379 = N3001;
  assign N2380 = N3003;
  assign N2381 = N3005;
  assign N2382 = N3007;
  assign N2383 = N3009;
  assign N2384 = N3011;
  assign way_id_o[5] = (N2446)? lru_i[0] : 
                       (N2448)? lru_i[1] : 
                       (N2450)? lru_i[2] : 
                       (N2452)? lru_i[3] : 
                       (N2454)? lru_i[4] : 
                       (N2456)? lru_i[5] : 
                       (N2458)? lru_i[6] : 
                       (N2460)? lru_i[7] : 
                       (N2462)? lru_i[8] : 
                       (N2464)? lru_i[9] : 
                       (N2466)? lru_i[10] : 
                       (N2468)? lru_i[11] : 
                       (N2470)? lru_i[12] : 
                       (N2472)? lru_i[13] : 
                       (N2474)? lru_i[14] : 
                       (N2476)? lru_i[15] : 
                       (N2478)? lru_i[16] : 
                       (N2480)? lru_i[17] : 
                       (N2482)? lru_i[18] : 
                       (N2484)? lru_i[19] : 
                       (N2486)? lru_i[20] : 
                       (N2488)? lru_i[21] : 
                       (N2490)? lru_i[22] : 
                       (N2492)? lru_i[23] : 
                       (N2494)? lru_i[24] : 
                       (N2496)? lru_i[25] : 
                       (N2498)? lru_i[26] : 
                       (N2500)? lru_i[27] : 
                       (N2502)? lru_i[28] : 
                       (N2504)? lru_i[29] : 
                       (N2506)? lru_i[30] : 
                       (N2508)? lru_i[31] : 
                       (N2447)? lru_i[32] : 
                       (N2449)? lru_i[33] : 
                       (N2451)? lru_i[34] : 
                       (N2453)? lru_i[35] : 
                       (N2455)? lru_i[36] : 
                       (N2457)? lru_i[37] : 
                       (N2459)? lru_i[38] : 
                       (N2461)? lru_i[39] : 
                       (N2463)? lru_i[40] : 
                       (N2465)? lru_i[41] : 
                       (N2467)? lru_i[42] : 
                       (N2469)? lru_i[43] : 
                       (N2471)? lru_i[44] : 
                       (N2473)? lru_i[45] : 
                       (N2475)? lru_i[46] : 
                       (N2477)? lru_i[47] : 
                       (N2479)? lru_i[48] : 
                       (N2481)? lru_i[49] : 
                       (N2483)? lru_i[50] : 
                       (N2485)? lru_i[51] : 
                       (N2487)? lru_i[52] : 
                       (N2489)? lru_i[53] : 
                       (N2491)? lru_i[54] : 
                       (N2493)? lru_i[55] : 
                       (N2495)? lru_i[56] : 
                       (N2497)? lru_i[57] : 
                       (N2499)? lru_i[58] : 
                       (N2501)? lru_i[59] : 
                       (N2503)? lru_i[60] : 
                       (N2505)? lru_i[61] : 
                       (N2507)? lru_i[62] : 1'b0;
  assign mask[1] = 1'b1 & N3076;
  assign N3076 = ~lru_i[0];
  assign mask[2] = 1'b1 & lru_i[0];
  assign mask[3] = mask[1] & N3077;
  assign N3077 = ~lru_i[1];
  assign mask[4] = mask[1] & lru_i[1];
  assign mask[5] = mask[2] & N3078;
  assign N3078 = ~lru_i[2];
  assign mask[6] = mask[2] & lru_i[2];
  assign mask[7] = mask[3] & N3079;
  assign N3079 = ~lru_i[3];
  assign mask[8] = mask[3] & lru_i[3];
  assign mask[9] = mask[4] & N3080;
  assign N3080 = ~lru_i[4];
  assign mask[10] = mask[4] & lru_i[4];
  assign mask[11] = mask[5] & N3081;
  assign N3081 = ~lru_i[5];
  assign mask[12] = mask[5] & lru_i[5];
  assign mask[13] = mask[6] & N3082;
  assign N3082 = ~lru_i[6];
  assign mask[14] = mask[6] & lru_i[6];
  assign mask[15] = mask[7] & N3083;
  assign N3083 = ~lru_i[7];
  assign mask[16] = mask[7] & lru_i[7];
  assign mask[17] = mask[8] & N3084;
  assign N3084 = ~lru_i[8];
  assign mask[18] = mask[8] & lru_i[8];
  assign mask[19] = mask[9] & N3085;
  assign N3085 = ~lru_i[9];
  assign mask[20] = mask[9] & lru_i[9];
  assign mask[21] = mask[10] & N3086;
  assign N3086 = ~lru_i[10];
  assign mask[22] = mask[10] & lru_i[10];
  assign mask[23] = mask[11] & N3087;
  assign N3087 = ~lru_i[11];
  assign mask[24] = mask[11] & lru_i[11];
  assign mask[25] = mask[12] & N3088;
  assign N3088 = ~lru_i[12];
  assign mask[26] = mask[12] & lru_i[12];
  assign mask[27] = mask[13] & N3089;
  assign N3089 = ~lru_i[13];
  assign mask[28] = mask[13] & lru_i[13];
  assign mask[29] = mask[14] & N3090;
  assign N3090 = ~lru_i[14];
  assign mask[30] = mask[14] & lru_i[14];
  assign mask[31] = mask[15] & N3091;
  assign N3091 = ~lru_i[15];
  assign mask[32] = mask[15] & lru_i[15];
  assign mask[33] = mask[16] & N3092;
  assign N3092 = ~lru_i[16];
  assign mask[34] = mask[16] & lru_i[16];
  assign mask[35] = mask[17] & N3093;
  assign N3093 = ~lru_i[17];
  assign mask[36] = mask[17] & lru_i[17];
  assign mask[37] = mask[18] & N3094;
  assign N3094 = ~lru_i[18];
  assign mask[38] = mask[18] & lru_i[18];
  assign mask[39] = mask[19] & N3095;
  assign N3095 = ~lru_i[19];
  assign mask[40] = mask[19] & lru_i[19];
  assign mask[41] = mask[20] & N3096;
  assign N3096 = ~lru_i[20];
  assign mask[42] = mask[20] & lru_i[20];
  assign mask[43] = mask[21] & N3097;
  assign N3097 = ~lru_i[21];
  assign mask[44] = mask[21] & lru_i[21];
  assign mask[45] = mask[22] & N3098;
  assign N3098 = ~lru_i[22];
  assign mask[46] = mask[22] & lru_i[22];
  assign mask[47] = mask[23] & N3099;
  assign N3099 = ~lru_i[23];
  assign mask[48] = mask[23] & lru_i[23];
  assign mask[49] = mask[24] & N3100;
  assign N3100 = ~lru_i[24];
  assign mask[50] = mask[24] & lru_i[24];
  assign mask[51] = mask[25] & N3101;
  assign N3101 = ~lru_i[25];
  assign mask[52] = mask[25] & lru_i[25];
  assign mask[53] = mask[26] & N3102;
  assign N3102 = ~lru_i[26];
  assign mask[54] = mask[26] & lru_i[26];
  assign mask[55] = mask[27] & N3103;
  assign N3103 = ~lru_i[27];
  assign mask[56] = mask[27] & lru_i[27];
  assign mask[57] = mask[28] & N3104;
  assign N3104 = ~lru_i[28];
  assign mask[58] = mask[28] & lru_i[28];
  assign mask[59] = mask[29] & N3105;
  assign N3105 = ~lru_i[29];
  assign mask[60] = mask[29] & lru_i[29];
  assign mask[61] = mask[30] & N3106;
  assign N3106 = ~lru_i[30];
  assign mask[62] = mask[30] & lru_i[30];
  assign N2385 = N2445 & N2445;
  assign N2386 = N2445 & 1'b0;
  assign N2387 = 1'b0 & N2445;
  assign N2388 = 1'b0 & 1'b0;
  assign N2389 = N2385 & N2445;
  assign N2390 = N2385 & 1'b0;
  assign N2391 = N2387 & N2445;
  assign N2392 = N2387 & 1'b0;
  assign N2393 = N2386 & N2445;
  assign N2394 = N2386 & 1'b0;
  assign N2395 = N2388 & N2445;
  assign N2396 = N2388 & 1'b0;
  assign N2397 = N2389 & N2445;
  assign N2398 = N2389 & 1'b0;
  assign N2399 = N2391 & N2445;
  assign N2400 = N2391 & 1'b0;
  assign N2401 = N2393 & N2445;
  assign N2402 = N2393 & 1'b0;
  assign N2403 = N2395 & N2445;
  assign N2404 = N2395 & 1'b0;
  assign N2405 = N2390 & N2445;
  assign N2406 = N2390 & 1'b0;
  assign N2407 = N2392 & N2445;
  assign N2408 = N2392 & 1'b0;
  assign N2409 = N2394 & N2445;
  assign N2410 = N2394 & 1'b0;
  assign N2411 = N2396 & N2445;
  assign N2412 = N2396 & 1'b0;
  assign N2413 = N2397 & N2445;
  assign N2414 = N2397 & 1'b0;
  assign N2415 = N2399 & N2445;
  assign N2416 = N2399 & 1'b0;
  assign N2417 = N2401 & N2445;
  assign N2418 = N2401 & 1'b0;
  assign N2419 = N2403 & N2445;
  assign N2420 = N2403 & 1'b0;
  assign N2421 = N2405 & N2445;
  assign N2422 = N2405 & 1'b0;
  assign N2423 = N2407 & N2445;
  assign N2424 = N2407 & 1'b0;
  assign N2425 = N2409 & N2445;
  assign N2426 = N2409 & 1'b0;
  assign N2427 = N2411 & N2445;
  assign N2428 = N2411 & 1'b0;
  assign N2429 = N2398 & N2445;
  assign N2430 = N2398 & 1'b0;
  assign N2431 = N2400 & N2445;
  assign N2432 = N2400 & 1'b0;
  assign N2433 = N2402 & N2445;
  assign N2434 = N2402 & 1'b0;
  assign N2435 = N2404 & N2445;
  assign N2436 = N2404 & 1'b0;
  assign N2437 = N2406 & N2445;
  assign N2438 = N2406 & 1'b0;
  assign N2439 = N2408 & N2445;
  assign N2440 = N2408 & 1'b0;
  assign N2441 = N2410 & N2445;
  assign N2442 = N2410 & 1'b0;
  assign N2443 = N2412 & N2445;
  assign N2444 = N2412 & 1'b0;
  assign N2445 = ~1'b0;
  assign N2446 = N2413 & N2445;
  assign N2447 = N2413 & 1'b0;
  assign N2448 = N2415 & N2445;
  assign N2449 = N2415 & 1'b0;
  assign N2450 = N2417 & N2445;
  assign N2451 = N2417 & 1'b0;
  assign N2452 = N2419 & N2445;
  assign N2453 = N2419 & 1'b0;
  assign N2454 = N2421 & N2445;
  assign N2455 = N2421 & 1'b0;
  assign N2456 = N2423 & N2445;
  assign N2457 = N2423 & 1'b0;
  assign N2458 = N2425 & N2445;
  assign N2459 = N2425 & 1'b0;
  assign N2460 = N2427 & N2445;
  assign N2461 = N2427 & 1'b0;
  assign N2462 = N2429 & N2445;
  assign N2463 = N2429 & 1'b0;
  assign N2464 = N2431 & N2445;
  assign N2465 = N2431 & 1'b0;
  assign N2466 = N2433 & N2445;
  assign N2467 = N2433 & 1'b0;
  assign N2468 = N2435 & N2445;
  assign N2469 = N2435 & 1'b0;
  assign N2470 = N2437 & N2445;
  assign N2471 = N2437 & 1'b0;
  assign N2472 = N2439 & N2445;
  assign N2473 = N2439 & 1'b0;
  assign N2474 = N2441 & N2445;
  assign N2475 = N2441 & 1'b0;
  assign N2476 = N2443 & N2445;
  assign N2477 = N2443 & 1'b0;
  assign N2478 = N2414 & N2445;
  assign N2479 = N2414 & 1'b0;
  assign N2480 = N2416 & N2445;
  assign N2481 = N2416 & 1'b0;
  assign N2482 = N2418 & N2445;
  assign N2483 = N2418 & 1'b0;
  assign N2484 = N2420 & N2445;
  assign N2485 = N2420 & 1'b0;
  assign N2486 = N2422 & N2445;
  assign N2487 = N2422 & 1'b0;
  assign N2488 = N2424 & N2445;
  assign N2489 = N2424 & 1'b0;
  assign N2490 = N2426 & N2445;
  assign N2491 = N2426 & 1'b0;
  assign N2492 = N2428 & N2445;
  assign N2493 = N2428 & 1'b0;
  assign N2494 = N2430 & N2445;
  assign N2495 = N2430 & 1'b0;
  assign N2496 = N2432 & N2445;
  assign N2497 = N2432 & 1'b0;
  assign N2498 = N2434 & N2445;
  assign N2499 = N2434 & 1'b0;
  assign N2500 = N2436 & N2445;
  assign N2501 = N2436 & 1'b0;
  assign N2502 = N2438 & N2445;
  assign N2503 = N2438 & 1'b0;
  assign N2504 = N2440 & N2445;
  assign N2505 = N2440 & 1'b0;
  assign N2506 = N2442 & N2445;
  assign N2507 = N2442 & 1'b0;
  assign N2508 = N2444 & N2445;
  assign pe_i_1__62_ = mask[62] ^ 1'b0;
  assign pe_i_1__61_ = mask[61] ^ 1'b0;
  assign pe_i_1__60_ = mask[60] ^ 1'b0;
  assign pe_i_1__59_ = mask[59] ^ 1'b0;
  assign pe_i_1__58_ = mask[58] ^ 1'b0;
  assign pe_i_1__57_ = mask[57] ^ 1'b0;
  assign pe_i_1__56_ = mask[56] ^ 1'b0;
  assign pe_i_1__55_ = mask[55] ^ 1'b0;
  assign pe_i_1__54_ = mask[54] ^ 1'b0;
  assign pe_i_1__53_ = mask[53] ^ 1'b0;
  assign pe_i_1__52_ = mask[52] ^ 1'b0;
  assign pe_i_1__51_ = mask[51] ^ 1'b0;
  assign pe_i_1__50_ = mask[50] ^ 1'b0;
  assign pe_i_1__49_ = mask[49] ^ 1'b0;
  assign pe_i_1__48_ = mask[48] ^ 1'b0;
  assign pe_i_1__47_ = mask[47] ^ 1'b0;
  assign pe_i_1__46_ = mask[46] ^ 1'b0;
  assign pe_i_1__45_ = mask[45] ^ 1'b0;
  assign pe_i_1__44_ = mask[44] ^ 1'b0;
  assign pe_i_1__43_ = mask[43] ^ 1'b0;
  assign pe_i_1__42_ = mask[42] ^ 1'b0;
  assign pe_i_1__41_ = mask[41] ^ 1'b0;
  assign pe_i_1__40_ = mask[40] ^ 1'b0;
  assign pe_i_1__39_ = mask[39] ^ 1'b0;
  assign pe_i_1__38_ = mask[38] ^ 1'b0;
  assign pe_i_1__37_ = mask[37] ^ 1'b0;
  assign pe_i_1__36_ = mask[36] ^ 1'b0;
  assign pe_i_1__35_ = mask[35] ^ 1'b0;
  assign pe_i_1__34_ = mask[34] ^ 1'b0;
  assign pe_i_1__33_ = mask[33] ^ 1'b0;
  assign pe_i_1__32_ = mask[32] ^ 1'b0;
  assign pe_i_1__31_ = mask[31] ^ 1'b0;
  assign pe_i_1__30_ = mask[30] ^ 1'b0;
  assign pe_i_1__29_ = mask[29] ^ 1'b0;
  assign pe_i_1__28_ = mask[28] ^ 1'b0;
  assign pe_i_1__27_ = mask[27] ^ 1'b0;
  assign pe_i_1__26_ = mask[26] ^ 1'b0;
  assign pe_i_1__25_ = mask[25] ^ 1'b0;
  assign pe_i_1__24_ = mask[24] ^ 1'b0;
  assign pe_i_1__23_ = mask[23] ^ 1'b0;
  assign pe_i_1__22_ = mask[22] ^ 1'b0;
  assign pe_i_1__21_ = mask[21] ^ 1'b0;
  assign pe_i_1__20_ = mask[20] ^ 1'b0;
  assign pe_i_1__19_ = mask[19] ^ 1'b0;
  assign pe_i_1__18_ = mask[18] ^ 1'b0;
  assign pe_i_1__17_ = mask[17] ^ 1'b0;
  assign pe_i_1__16_ = mask[16] ^ 1'b0;
  assign pe_i_1__15_ = mask[15] ^ 1'b0;
  assign pe_i_1__14_ = mask[14] ^ 1'b0;
  assign pe_i_1__13_ = mask[13] ^ 1'b0;
  assign pe_i_1__12_ = mask[12] ^ 1'b0;
  assign pe_i_1__11_ = mask[11] ^ 1'b0;
  assign pe_i_1__10_ = mask[10] ^ 1'b0;
  assign pe_i_1__9_ = mask[9] ^ 1'b0;
  assign pe_i_1__8_ = mask[8] ^ 1'b0;
  assign pe_i_1__7_ = mask[7] ^ 1'b0;
  assign pe_i_1__6_ = mask[6] ^ 1'b0;
  assign pe_i_1__5_ = mask[5] ^ 1'b0;
  assign pe_i_1__4_ = mask[4] ^ 1'b0;
  assign pe_i_1__3_ = mask[3] ^ 1'b0;
  assign pe_i_1__2_ = mask[2] ^ 1'b0;
  assign pe_i_1__1_ = mask[1] ^ 1'b0;
  assign pe_i_1__0_ = 1'b1 ^ 1'b1;
  assign pe_i_2__62_ = pe_i_1__62_ ^ N2697;
  assign pe_i_2__61_ = pe_i_1__61_ ^ N2696;
  assign pe_i_2__60_ = pe_i_1__60_ ^ N2695;
  assign pe_i_2__59_ = pe_i_1__59_ ^ N2694;
  assign pe_i_2__58_ = pe_i_1__58_ ^ N2693;
  assign pe_i_2__57_ = pe_i_1__57_ ^ N2692;
  assign pe_i_2__56_ = pe_i_1__56_ ^ N2691;
  assign pe_i_2__55_ = pe_i_1__55_ ^ N2690;
  assign pe_i_2__54_ = pe_i_1__54_ ^ N2689;
  assign pe_i_2__53_ = pe_i_1__53_ ^ N2688;
  assign pe_i_2__52_ = pe_i_1__52_ ^ N2687;
  assign pe_i_2__51_ = pe_i_1__51_ ^ N2686;
  assign pe_i_2__50_ = pe_i_1__50_ ^ N2685;
  assign pe_i_2__49_ = pe_i_1__49_ ^ N2684;
  assign pe_i_2__48_ = pe_i_1__48_ ^ N2683;
  assign pe_i_2__47_ = pe_i_1__47_ ^ N2682;
  assign pe_i_2__46_ = pe_i_1__46_ ^ N2681;
  assign pe_i_2__45_ = pe_i_1__45_ ^ N2680;
  assign pe_i_2__44_ = pe_i_1__44_ ^ N2679;
  assign pe_i_2__43_ = pe_i_1__43_ ^ N2678;
  assign pe_i_2__42_ = pe_i_1__42_ ^ N2677;
  assign pe_i_2__41_ = pe_i_1__41_ ^ N2676;
  assign pe_i_2__40_ = pe_i_1__40_ ^ N2675;
  assign pe_i_2__39_ = pe_i_1__39_ ^ N2674;
  assign pe_i_2__38_ = pe_i_1__38_ ^ N2673;
  assign pe_i_2__37_ = pe_i_1__37_ ^ N2672;
  assign pe_i_2__36_ = pe_i_1__36_ ^ N2671;
  assign pe_i_2__35_ = pe_i_1__35_ ^ N2670;
  assign pe_i_2__34_ = pe_i_1__34_ ^ N2669;
  assign pe_i_2__33_ = pe_i_1__33_ ^ N2668;
  assign pe_i_2__32_ = pe_i_1__32_ ^ N2667;
  assign pe_i_2__31_ = pe_i_1__31_ ^ N2666;
  assign pe_i_2__30_ = pe_i_1__30_ ^ N2665;
  assign pe_i_2__29_ = pe_i_1__29_ ^ N2664;
  assign pe_i_2__28_ = pe_i_1__28_ ^ N2663;
  assign pe_i_2__27_ = pe_i_1__27_ ^ N2662;
  assign pe_i_2__26_ = pe_i_1__26_ ^ N2661;
  assign pe_i_2__25_ = pe_i_1__25_ ^ N2660;
  assign pe_i_2__24_ = pe_i_1__24_ ^ N2659;
  assign pe_i_2__23_ = pe_i_1__23_ ^ N2658;
  assign pe_i_2__22_ = pe_i_1__22_ ^ N2657;
  assign pe_i_2__21_ = pe_i_1__21_ ^ N2656;
  assign pe_i_2__20_ = pe_i_1__20_ ^ N2655;
  assign pe_i_2__19_ = pe_i_1__19_ ^ N2654;
  assign pe_i_2__18_ = pe_i_1__18_ ^ N2653;
  assign pe_i_2__17_ = pe_i_1__17_ ^ N2652;
  assign pe_i_2__16_ = pe_i_1__16_ ^ N2651;
  assign pe_i_2__15_ = pe_i_1__15_ ^ N2650;
  assign pe_i_2__14_ = pe_i_1__14_ ^ N2649;
  assign pe_i_2__13_ = pe_i_1__13_ ^ N2648;
  assign pe_i_2__12_ = pe_i_1__12_ ^ N2647;
  assign pe_i_2__11_ = pe_i_1__11_ ^ N2646;
  assign pe_i_2__10_ = pe_i_1__10_ ^ N2645;
  assign pe_i_2__9_ = pe_i_1__9_ ^ N2644;
  assign pe_i_2__8_ = pe_i_1__8_ ^ N2643;
  assign pe_i_2__7_ = pe_i_1__7_ ^ N2642;
  assign pe_i_2__6_ = pe_i_1__6_ ^ N2641;
  assign pe_i_2__5_ = pe_i_1__5_ ^ N2640;
  assign pe_i_2__4_ = pe_i_1__4_ ^ N2639;
  assign pe_i_2__3_ = pe_i_1__3_ ^ N2638;
  assign pe_i_2__2_ = pe_i_1__2_ ^ N2637;
  assign pe_i_2__1_ = pe_i_1__1_ ^ N2636;
  assign pe_i_2__0_ = pe_i_1__0_ ^ N2635;
  assign pe_i_3__62_ = pe_i_2__62_ ^ N2823;
  assign pe_i_3__61_ = pe_i_2__61_ ^ N2822;
  assign pe_i_3__60_ = pe_i_2__60_ ^ N2821;
  assign pe_i_3__59_ = pe_i_2__59_ ^ N2820;
  assign pe_i_3__58_ = pe_i_2__58_ ^ N2819;
  assign pe_i_3__57_ = pe_i_2__57_ ^ N2818;
  assign pe_i_3__56_ = pe_i_2__56_ ^ N2817;
  assign pe_i_3__55_ = pe_i_2__55_ ^ N2816;
  assign pe_i_3__54_ = pe_i_2__54_ ^ N2815;
  assign pe_i_3__53_ = pe_i_2__53_ ^ N2814;
  assign pe_i_3__52_ = pe_i_2__52_ ^ N2813;
  assign pe_i_3__51_ = pe_i_2__51_ ^ N2812;
  assign pe_i_3__50_ = pe_i_2__50_ ^ N2811;
  assign pe_i_3__49_ = pe_i_2__49_ ^ N2810;
  assign pe_i_3__48_ = pe_i_2__48_ ^ N2809;
  assign pe_i_3__47_ = pe_i_2__47_ ^ N2808;
  assign pe_i_3__46_ = pe_i_2__46_ ^ N2807;
  assign pe_i_3__45_ = pe_i_2__45_ ^ N2806;
  assign pe_i_3__44_ = pe_i_2__44_ ^ N2805;
  assign pe_i_3__43_ = pe_i_2__43_ ^ N2804;
  assign pe_i_3__42_ = pe_i_2__42_ ^ N2803;
  assign pe_i_3__41_ = pe_i_2__41_ ^ N2802;
  assign pe_i_3__40_ = pe_i_2__40_ ^ N2801;
  assign pe_i_3__39_ = pe_i_2__39_ ^ N2800;
  assign pe_i_3__38_ = pe_i_2__38_ ^ N2799;
  assign pe_i_3__37_ = pe_i_2__37_ ^ N2798;
  assign pe_i_3__36_ = pe_i_2__36_ ^ N2797;
  assign pe_i_3__35_ = pe_i_2__35_ ^ N2796;
  assign pe_i_3__34_ = pe_i_2__34_ ^ N2795;
  assign pe_i_3__33_ = pe_i_2__33_ ^ N2794;
  assign pe_i_3__32_ = pe_i_2__32_ ^ N2793;
  assign pe_i_3__31_ = pe_i_2__31_ ^ N2792;
  assign pe_i_3__30_ = pe_i_2__30_ ^ N2791;
  assign pe_i_3__29_ = pe_i_2__29_ ^ N2790;
  assign pe_i_3__28_ = pe_i_2__28_ ^ N2789;
  assign pe_i_3__27_ = pe_i_2__27_ ^ N2788;
  assign pe_i_3__26_ = pe_i_2__26_ ^ N2787;
  assign pe_i_3__25_ = pe_i_2__25_ ^ N2786;
  assign pe_i_3__24_ = pe_i_2__24_ ^ N2785;
  assign pe_i_3__23_ = pe_i_2__23_ ^ N2784;
  assign pe_i_3__22_ = pe_i_2__22_ ^ N2783;
  assign pe_i_3__21_ = pe_i_2__21_ ^ N2782;
  assign pe_i_3__20_ = pe_i_2__20_ ^ N2781;
  assign pe_i_3__19_ = pe_i_2__19_ ^ N2780;
  assign pe_i_3__18_ = pe_i_2__18_ ^ N2779;
  assign pe_i_3__17_ = pe_i_2__17_ ^ N2778;
  assign pe_i_3__16_ = pe_i_2__16_ ^ N2777;
  assign pe_i_3__15_ = pe_i_2__15_ ^ N2776;
  assign pe_i_3__14_ = pe_i_2__14_ ^ N2775;
  assign pe_i_3__13_ = pe_i_2__13_ ^ N2774;
  assign pe_i_3__12_ = pe_i_2__12_ ^ N2773;
  assign pe_i_3__11_ = pe_i_2__11_ ^ N2772;
  assign pe_i_3__10_ = pe_i_2__10_ ^ N2771;
  assign pe_i_3__9_ = pe_i_2__9_ ^ N2770;
  assign pe_i_3__8_ = pe_i_2__8_ ^ N2769;
  assign pe_i_3__7_ = pe_i_2__7_ ^ N2768;
  assign pe_i_3__6_ = pe_i_2__6_ ^ N2767;
  assign pe_i_3__5_ = pe_i_2__5_ ^ N2766;
  assign pe_i_3__4_ = pe_i_2__4_ ^ N2765;
  assign pe_i_3__3_ = pe_i_2__3_ ^ N2764;
  assign pe_i_3__2_ = pe_i_2__2_ ^ N2763;
  assign pe_i_3__1_ = pe_i_2__1_ ^ N2762;
  assign pe_i_3__0_ = pe_i_2__0_ ^ N2761;
  assign pe_i_4__62_ = pe_i_3__62_ ^ N2949;
  assign pe_i_4__61_ = pe_i_3__61_ ^ N2948;
  assign pe_i_4__60_ = pe_i_3__60_ ^ N2947;
  assign pe_i_4__59_ = pe_i_3__59_ ^ N2946;
  assign pe_i_4__58_ = pe_i_3__58_ ^ N2945;
  assign pe_i_4__57_ = pe_i_3__57_ ^ N2944;
  assign pe_i_4__56_ = pe_i_3__56_ ^ N2943;
  assign pe_i_4__55_ = pe_i_3__55_ ^ N2942;
  assign pe_i_4__54_ = pe_i_3__54_ ^ N2941;
  assign pe_i_4__53_ = pe_i_3__53_ ^ N2940;
  assign pe_i_4__52_ = pe_i_3__52_ ^ N2939;
  assign pe_i_4__51_ = pe_i_3__51_ ^ N2938;
  assign pe_i_4__50_ = pe_i_3__50_ ^ N2937;
  assign pe_i_4__49_ = pe_i_3__49_ ^ N2936;
  assign pe_i_4__48_ = pe_i_3__48_ ^ N2935;
  assign pe_i_4__47_ = pe_i_3__47_ ^ N2934;
  assign pe_i_4__46_ = pe_i_3__46_ ^ N2933;
  assign pe_i_4__45_ = pe_i_3__45_ ^ N2932;
  assign pe_i_4__44_ = pe_i_3__44_ ^ N2931;
  assign pe_i_4__43_ = pe_i_3__43_ ^ N2930;
  assign pe_i_4__42_ = pe_i_3__42_ ^ N2929;
  assign pe_i_4__41_ = pe_i_3__41_ ^ N2928;
  assign pe_i_4__40_ = pe_i_3__40_ ^ N2927;
  assign pe_i_4__39_ = pe_i_3__39_ ^ N2926;
  assign pe_i_4__38_ = pe_i_3__38_ ^ N2925;
  assign pe_i_4__37_ = pe_i_3__37_ ^ N2924;
  assign pe_i_4__36_ = pe_i_3__36_ ^ N2923;
  assign pe_i_4__35_ = pe_i_3__35_ ^ N2922;
  assign pe_i_4__34_ = pe_i_3__34_ ^ N2921;
  assign pe_i_4__33_ = pe_i_3__33_ ^ N2920;
  assign pe_i_4__32_ = pe_i_3__32_ ^ N2919;
  assign pe_i_4__31_ = pe_i_3__31_ ^ N2918;
  assign pe_i_4__30_ = pe_i_3__30_ ^ N2917;
  assign pe_i_4__29_ = pe_i_3__29_ ^ N2916;
  assign pe_i_4__28_ = pe_i_3__28_ ^ N2915;
  assign pe_i_4__27_ = pe_i_3__27_ ^ N2914;
  assign pe_i_4__26_ = pe_i_3__26_ ^ N2913;
  assign pe_i_4__25_ = pe_i_3__25_ ^ N2912;
  assign pe_i_4__24_ = pe_i_3__24_ ^ N2911;
  assign pe_i_4__23_ = pe_i_3__23_ ^ N2910;
  assign pe_i_4__22_ = pe_i_3__22_ ^ N2909;
  assign pe_i_4__21_ = pe_i_3__21_ ^ N2908;
  assign pe_i_4__20_ = pe_i_3__20_ ^ N2907;
  assign pe_i_4__19_ = pe_i_3__19_ ^ N2906;
  assign pe_i_4__18_ = pe_i_3__18_ ^ N2905;
  assign pe_i_4__17_ = pe_i_3__17_ ^ N2904;
  assign pe_i_4__16_ = pe_i_3__16_ ^ N2903;
  assign pe_i_4__15_ = pe_i_3__15_ ^ N2902;
  assign pe_i_4__14_ = pe_i_3__14_ ^ N2901;
  assign pe_i_4__13_ = pe_i_3__13_ ^ N2900;
  assign pe_i_4__12_ = pe_i_3__12_ ^ N2899;
  assign pe_i_4__11_ = pe_i_3__11_ ^ N2898;
  assign pe_i_4__10_ = pe_i_3__10_ ^ N2897;
  assign pe_i_4__9_ = pe_i_3__9_ ^ N2896;
  assign pe_i_4__8_ = pe_i_3__8_ ^ N2895;
  assign pe_i_4__7_ = pe_i_3__7_ ^ N2894;
  assign pe_i_4__6_ = pe_i_3__6_ ^ N2893;
  assign pe_i_4__5_ = pe_i_3__5_ ^ N2892;
  assign pe_i_4__4_ = pe_i_3__4_ ^ N2891;
  assign pe_i_4__3_ = pe_i_3__3_ ^ N2890;
  assign pe_i_4__2_ = pe_i_3__2_ ^ N2889;
  assign pe_i_4__1_ = pe_i_3__1_ ^ N2888;
  assign pe_i_4__0_ = pe_i_3__0_ ^ N2887;
  assign pe_i_5__62_ = pe_i_4__62_ ^ N3075;
  assign pe_i_5__61_ = pe_i_4__61_ ^ N3074;
  assign pe_i_5__60_ = pe_i_4__60_ ^ N3073;
  assign pe_i_5__59_ = pe_i_4__59_ ^ N3072;
  assign pe_i_5__58_ = pe_i_4__58_ ^ N3071;
  assign pe_i_5__57_ = pe_i_4__57_ ^ N3070;
  assign pe_i_5__56_ = pe_i_4__56_ ^ N3069;
  assign pe_i_5__55_ = pe_i_4__55_ ^ N3068;
  assign pe_i_5__54_ = pe_i_4__54_ ^ N3067;
  assign pe_i_5__53_ = pe_i_4__53_ ^ N3066;
  assign pe_i_5__52_ = pe_i_4__52_ ^ N3065;
  assign pe_i_5__51_ = pe_i_4__51_ ^ N3064;
  assign pe_i_5__50_ = pe_i_4__50_ ^ N3063;
  assign pe_i_5__49_ = pe_i_4__49_ ^ N3062;
  assign pe_i_5__48_ = pe_i_4__48_ ^ N3061;
  assign pe_i_5__47_ = pe_i_4__47_ ^ N3060;
  assign pe_i_5__46_ = pe_i_4__46_ ^ N3059;
  assign pe_i_5__45_ = pe_i_4__45_ ^ N3058;
  assign pe_i_5__44_ = pe_i_4__44_ ^ N3057;
  assign pe_i_5__43_ = pe_i_4__43_ ^ N3056;
  assign pe_i_5__42_ = pe_i_4__42_ ^ N3055;
  assign pe_i_5__41_ = pe_i_4__41_ ^ N3054;
  assign pe_i_5__40_ = pe_i_4__40_ ^ N3053;
  assign pe_i_5__39_ = pe_i_4__39_ ^ N3052;
  assign pe_i_5__38_ = pe_i_4__38_ ^ N3051;
  assign pe_i_5__37_ = pe_i_4__37_ ^ N3050;
  assign pe_i_5__36_ = pe_i_4__36_ ^ N3049;
  assign pe_i_5__35_ = pe_i_4__35_ ^ N3048;
  assign pe_i_5__34_ = pe_i_4__34_ ^ N3047;
  assign pe_i_5__33_ = pe_i_4__33_ ^ N3046;
  assign pe_i_5__32_ = pe_i_4__32_ ^ N3045;
  assign pe_i_5__31_ = pe_i_4__31_ ^ N3044;
  assign pe_i_5__30_ = pe_i_4__30_ ^ N3043;
  assign pe_i_5__29_ = pe_i_4__29_ ^ N3042;
  assign pe_i_5__28_ = pe_i_4__28_ ^ N3041;
  assign pe_i_5__27_ = pe_i_4__27_ ^ N3040;
  assign pe_i_5__26_ = pe_i_4__26_ ^ N3039;
  assign pe_i_5__25_ = pe_i_4__25_ ^ N3038;
  assign pe_i_5__24_ = pe_i_4__24_ ^ N3037;
  assign pe_i_5__23_ = pe_i_4__23_ ^ N3036;
  assign pe_i_5__22_ = pe_i_4__22_ ^ N3035;
  assign pe_i_5__21_ = pe_i_4__21_ ^ N3034;
  assign pe_i_5__20_ = pe_i_4__20_ ^ N3033;
  assign pe_i_5__19_ = pe_i_4__19_ ^ N3032;
  assign pe_i_5__18_ = pe_i_4__18_ ^ N3031;
  assign pe_i_5__17_ = pe_i_4__17_ ^ N3030;
  assign pe_i_5__16_ = pe_i_4__16_ ^ N3029;
  assign pe_i_5__15_ = pe_i_4__15_ ^ N3028;
  assign pe_i_5__14_ = pe_i_4__14_ ^ N3027;
  assign pe_i_5__13_ = pe_i_4__13_ ^ N3026;
  assign pe_i_5__12_ = pe_i_4__12_ ^ N3025;
  assign pe_i_5__11_ = pe_i_4__11_ ^ N3024;
  assign pe_i_5__10_ = pe_i_4__10_ ^ N3023;
  assign pe_i_5__9_ = pe_i_4__9_ ^ N3022;
  assign pe_i_5__8_ = pe_i_4__8_ ^ N3021;
  assign pe_i_5__7_ = pe_i_4__7_ ^ N3020;
  assign pe_i_5__6_ = pe_i_4__6_ ^ N3019;
  assign pe_i_5__5_ = pe_i_4__5_ ^ N3018;
  assign pe_i_5__4_ = pe_i_4__4_ ^ N3017;
  assign pe_i_5__3_ = pe_i_4__3_ ^ N3016;
  assign pe_i_5__2_ = pe_i_4__2_ ^ N3015;
  assign pe_i_5__1_ = pe_i_4__1_ ^ N3014;
  assign pe_i_5__0_ = pe_i_4__0_ ^ N3013;

endmodule

