

module top
(
  data_i,
  sel_i,
  data_o
);

  input [4095:0] data_i;
  input [5:0] sel_i;
  output [4095:0] data_o;

  bsg_mux_butterfly
  wrapper
  (
    .data_i(data_i),
    .sel_i(sel_i),
    .data_o(data_o)
  );


endmodule



module bsg_swap_width_p64
(
  data_i,
  swap_i,
  data_o
);

  input [127:0] data_i;
  output [127:0] data_o;
  input swap_i;
  wire [127:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[63:0], data_i[127:64] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p128
(
  data_i,
  swap_i,
  data_o
);

  input [255:0] data_i;
  output [255:0] data_o;
  input swap_i;
  wire [255:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[127:0], data_i[255:128] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p256
(
  data_i,
  swap_i,
  data_o
);

  input [511:0] data_i;
  output [511:0] data_o;
  input swap_i;
  wire [511:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[255:0], data_i[511:256] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p512
(
  data_i,
  swap_i,
  data_o
);

  input [1023:0] data_i;
  output [1023:0] data_o;
  input swap_i;
  wire [1023:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[511:0], data_i[1023:512] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p1024
(
  data_i,
  swap_i,
  data_o
);

  input [2047:0] data_i;
  output [2047:0] data_o;
  input swap_i;
  wire [2047:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[1023:0], data_i[2047:1024] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p2048
(
  data_i,
  swap_i,
  data_o
);

  input [4095:0] data_i;
  output [4095:0] data_o;
  input swap_i;
  wire [4095:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[2047:0], data_i[4095:2048] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_mux_butterfly
(
  data_i,
  sel_i,
  data_o
);

  input [4095:0] data_i;
  input [5:0] sel_i;
  output [4095:0] data_o;
  wire [4095:0] data_o;
  wire data_stage_1__4095_,data_stage_1__4094_,data_stage_1__4093_,data_stage_1__4092_,
  data_stage_1__4091_,data_stage_1__4090_,data_stage_1__4089_,data_stage_1__4088_,
  data_stage_1__4087_,data_stage_1__4086_,data_stage_1__4085_,data_stage_1__4084_,
  data_stage_1__4083_,data_stage_1__4082_,data_stage_1__4081_,data_stage_1__4080_,
  data_stage_1__4079_,data_stage_1__4078_,data_stage_1__4077_,data_stage_1__4076_,
  data_stage_1__4075_,data_stage_1__4074_,data_stage_1__4073_,data_stage_1__4072_,
  data_stage_1__4071_,data_stage_1__4070_,data_stage_1__4069_,data_stage_1__4068_,
  data_stage_1__4067_,data_stage_1__4066_,data_stage_1__4065_,data_stage_1__4064_,
  data_stage_1__4063_,data_stage_1__4062_,data_stage_1__4061_,data_stage_1__4060_,
  data_stage_1__4059_,data_stage_1__4058_,data_stage_1__4057_,data_stage_1__4056_,
  data_stage_1__4055_,data_stage_1__4054_,data_stage_1__4053_,data_stage_1__4052_,
  data_stage_1__4051_,data_stage_1__4050_,data_stage_1__4049_,data_stage_1__4048_,
  data_stage_1__4047_,data_stage_1__4046_,data_stage_1__4045_,data_stage_1__4044_,
  data_stage_1__4043_,data_stage_1__4042_,data_stage_1__4041_,data_stage_1__4040_,
  data_stage_1__4039_,data_stage_1__4038_,data_stage_1__4037_,data_stage_1__4036_,
  data_stage_1__4035_,data_stage_1__4034_,data_stage_1__4033_,data_stage_1__4032_,
  data_stage_1__4031_,data_stage_1__4030_,data_stage_1__4029_,data_stage_1__4028_,
  data_stage_1__4027_,data_stage_1__4026_,data_stage_1__4025_,data_stage_1__4024_,
  data_stage_1__4023_,data_stage_1__4022_,data_stage_1__4021_,data_stage_1__4020_,
  data_stage_1__4019_,data_stage_1__4018_,data_stage_1__4017_,data_stage_1__4016_,
  data_stage_1__4015_,data_stage_1__4014_,data_stage_1__4013_,data_stage_1__4012_,
  data_stage_1__4011_,data_stage_1__4010_,data_stage_1__4009_,data_stage_1__4008_,
  data_stage_1__4007_,data_stage_1__4006_,data_stage_1__4005_,data_stage_1__4004_,
  data_stage_1__4003_,data_stage_1__4002_,data_stage_1__4001_,data_stage_1__4000_,
  data_stage_1__3999_,data_stage_1__3998_,data_stage_1__3997_,data_stage_1__3996_,
  data_stage_1__3995_,data_stage_1__3994_,data_stage_1__3993_,data_stage_1__3992_,
  data_stage_1__3991_,data_stage_1__3990_,data_stage_1__3989_,data_stage_1__3988_,
  data_stage_1__3987_,data_stage_1__3986_,data_stage_1__3985_,data_stage_1__3984_,
  data_stage_1__3983_,data_stage_1__3982_,data_stage_1__3981_,data_stage_1__3980_,
  data_stage_1__3979_,data_stage_1__3978_,data_stage_1__3977_,data_stage_1__3976_,
  data_stage_1__3975_,data_stage_1__3974_,data_stage_1__3973_,data_stage_1__3972_,
  data_stage_1__3971_,data_stage_1__3970_,data_stage_1__3969_,data_stage_1__3968_,
  data_stage_1__3967_,data_stage_1__3966_,data_stage_1__3965_,data_stage_1__3964_,
  data_stage_1__3963_,data_stage_1__3962_,data_stage_1__3961_,data_stage_1__3960_,
  data_stage_1__3959_,data_stage_1__3958_,data_stage_1__3957_,data_stage_1__3956_,
  data_stage_1__3955_,data_stage_1__3954_,data_stage_1__3953_,data_stage_1__3952_,
  data_stage_1__3951_,data_stage_1__3950_,data_stage_1__3949_,data_stage_1__3948_,
  data_stage_1__3947_,data_stage_1__3946_,data_stage_1__3945_,data_stage_1__3944_,
  data_stage_1__3943_,data_stage_1__3942_,data_stage_1__3941_,data_stage_1__3940_,
  data_stage_1__3939_,data_stage_1__3938_,data_stage_1__3937_,data_stage_1__3936_,
  data_stage_1__3935_,data_stage_1__3934_,data_stage_1__3933_,data_stage_1__3932_,
  data_stage_1__3931_,data_stage_1__3930_,data_stage_1__3929_,data_stage_1__3928_,
  data_stage_1__3927_,data_stage_1__3926_,data_stage_1__3925_,data_stage_1__3924_,
  data_stage_1__3923_,data_stage_1__3922_,data_stage_1__3921_,data_stage_1__3920_,
  data_stage_1__3919_,data_stage_1__3918_,data_stage_1__3917_,data_stage_1__3916_,
  data_stage_1__3915_,data_stage_1__3914_,data_stage_1__3913_,data_stage_1__3912_,
  data_stage_1__3911_,data_stage_1__3910_,data_stage_1__3909_,data_stage_1__3908_,
  data_stage_1__3907_,data_stage_1__3906_,data_stage_1__3905_,data_stage_1__3904_,
  data_stage_1__3903_,data_stage_1__3902_,data_stage_1__3901_,data_stage_1__3900_,
  data_stage_1__3899_,data_stage_1__3898_,data_stage_1__3897_,data_stage_1__3896_,
  data_stage_1__3895_,data_stage_1__3894_,data_stage_1__3893_,data_stage_1__3892_,
  data_stage_1__3891_,data_stage_1__3890_,data_stage_1__3889_,data_stage_1__3888_,
  data_stage_1__3887_,data_stage_1__3886_,data_stage_1__3885_,data_stage_1__3884_,
  data_stage_1__3883_,data_stage_1__3882_,data_stage_1__3881_,data_stage_1__3880_,
  data_stage_1__3879_,data_stage_1__3878_,data_stage_1__3877_,data_stage_1__3876_,
  data_stage_1__3875_,data_stage_1__3874_,data_stage_1__3873_,data_stage_1__3872_,
  data_stage_1__3871_,data_stage_1__3870_,data_stage_1__3869_,data_stage_1__3868_,
  data_stage_1__3867_,data_stage_1__3866_,data_stage_1__3865_,data_stage_1__3864_,
  data_stage_1__3863_,data_stage_1__3862_,data_stage_1__3861_,data_stage_1__3860_,
  data_stage_1__3859_,data_stage_1__3858_,data_stage_1__3857_,data_stage_1__3856_,
  data_stage_1__3855_,data_stage_1__3854_,data_stage_1__3853_,data_stage_1__3852_,
  data_stage_1__3851_,data_stage_1__3850_,data_stage_1__3849_,data_stage_1__3848_,
  data_stage_1__3847_,data_stage_1__3846_,data_stage_1__3845_,data_stage_1__3844_,
  data_stage_1__3843_,data_stage_1__3842_,data_stage_1__3841_,data_stage_1__3840_,
  data_stage_1__3839_,data_stage_1__3838_,data_stage_1__3837_,data_stage_1__3836_,
  data_stage_1__3835_,data_stage_1__3834_,data_stage_1__3833_,data_stage_1__3832_,
  data_stage_1__3831_,data_stage_1__3830_,data_stage_1__3829_,data_stage_1__3828_,
  data_stage_1__3827_,data_stage_1__3826_,data_stage_1__3825_,data_stage_1__3824_,
  data_stage_1__3823_,data_stage_1__3822_,data_stage_1__3821_,data_stage_1__3820_,
  data_stage_1__3819_,data_stage_1__3818_,data_stage_1__3817_,data_stage_1__3816_,
  data_stage_1__3815_,data_stage_1__3814_,data_stage_1__3813_,data_stage_1__3812_,
  data_stage_1__3811_,data_stage_1__3810_,data_stage_1__3809_,data_stage_1__3808_,
  data_stage_1__3807_,data_stage_1__3806_,data_stage_1__3805_,data_stage_1__3804_,
  data_stage_1__3803_,data_stage_1__3802_,data_stage_1__3801_,data_stage_1__3800_,
  data_stage_1__3799_,data_stage_1__3798_,data_stage_1__3797_,data_stage_1__3796_,
  data_stage_1__3795_,data_stage_1__3794_,data_stage_1__3793_,data_stage_1__3792_,
  data_stage_1__3791_,data_stage_1__3790_,data_stage_1__3789_,data_stage_1__3788_,
  data_stage_1__3787_,data_stage_1__3786_,data_stage_1__3785_,data_stage_1__3784_,
  data_stage_1__3783_,data_stage_1__3782_,data_stage_1__3781_,data_stage_1__3780_,
  data_stage_1__3779_,data_stage_1__3778_,data_stage_1__3777_,data_stage_1__3776_,
  data_stage_1__3775_,data_stage_1__3774_,data_stage_1__3773_,data_stage_1__3772_,
  data_stage_1__3771_,data_stage_1__3770_,data_stage_1__3769_,data_stage_1__3768_,
  data_stage_1__3767_,data_stage_1__3766_,data_stage_1__3765_,data_stage_1__3764_,
  data_stage_1__3763_,data_stage_1__3762_,data_stage_1__3761_,data_stage_1__3760_,
  data_stage_1__3759_,data_stage_1__3758_,data_stage_1__3757_,data_stage_1__3756_,
  data_stage_1__3755_,data_stage_1__3754_,data_stage_1__3753_,data_stage_1__3752_,
  data_stage_1__3751_,data_stage_1__3750_,data_stage_1__3749_,data_stage_1__3748_,
  data_stage_1__3747_,data_stage_1__3746_,data_stage_1__3745_,data_stage_1__3744_,
  data_stage_1__3743_,data_stage_1__3742_,data_stage_1__3741_,data_stage_1__3740_,
  data_stage_1__3739_,data_stage_1__3738_,data_stage_1__3737_,data_stage_1__3736_,
  data_stage_1__3735_,data_stage_1__3734_,data_stage_1__3733_,data_stage_1__3732_,
  data_stage_1__3731_,data_stage_1__3730_,data_stage_1__3729_,data_stage_1__3728_,
  data_stage_1__3727_,data_stage_1__3726_,data_stage_1__3725_,data_stage_1__3724_,
  data_stage_1__3723_,data_stage_1__3722_,data_stage_1__3721_,data_stage_1__3720_,
  data_stage_1__3719_,data_stage_1__3718_,data_stage_1__3717_,data_stage_1__3716_,
  data_stage_1__3715_,data_stage_1__3714_,data_stage_1__3713_,data_stage_1__3712_,
  data_stage_1__3711_,data_stage_1__3710_,data_stage_1__3709_,data_stage_1__3708_,
  data_stage_1__3707_,data_stage_1__3706_,data_stage_1__3705_,data_stage_1__3704_,
  data_stage_1__3703_,data_stage_1__3702_,data_stage_1__3701_,data_stage_1__3700_,
  data_stage_1__3699_,data_stage_1__3698_,data_stage_1__3697_,data_stage_1__3696_,
  data_stage_1__3695_,data_stage_1__3694_,data_stage_1__3693_,data_stage_1__3692_,
  data_stage_1__3691_,data_stage_1__3690_,data_stage_1__3689_,data_stage_1__3688_,
  data_stage_1__3687_,data_stage_1__3686_,data_stage_1__3685_,data_stage_1__3684_,
  data_stage_1__3683_,data_stage_1__3682_,data_stage_1__3681_,data_stage_1__3680_,
  data_stage_1__3679_,data_stage_1__3678_,data_stage_1__3677_,data_stage_1__3676_,
  data_stage_1__3675_,data_stage_1__3674_,data_stage_1__3673_,data_stage_1__3672_,
  data_stage_1__3671_,data_stage_1__3670_,data_stage_1__3669_,data_stage_1__3668_,
  data_stage_1__3667_,data_stage_1__3666_,data_stage_1__3665_,data_stage_1__3664_,
  data_stage_1__3663_,data_stage_1__3662_,data_stage_1__3661_,data_stage_1__3660_,
  data_stage_1__3659_,data_stage_1__3658_,data_stage_1__3657_,data_stage_1__3656_,
  data_stage_1__3655_,data_stage_1__3654_,data_stage_1__3653_,data_stage_1__3652_,
  data_stage_1__3651_,data_stage_1__3650_,data_stage_1__3649_,data_stage_1__3648_,
  data_stage_1__3647_,data_stage_1__3646_,data_stage_1__3645_,data_stage_1__3644_,
  data_stage_1__3643_,data_stage_1__3642_,data_stage_1__3641_,data_stage_1__3640_,
  data_stage_1__3639_,data_stage_1__3638_,data_stage_1__3637_,data_stage_1__3636_,
  data_stage_1__3635_,data_stage_1__3634_,data_stage_1__3633_,data_stage_1__3632_,
  data_stage_1__3631_,data_stage_1__3630_,data_stage_1__3629_,data_stage_1__3628_,
  data_stage_1__3627_,data_stage_1__3626_,data_stage_1__3625_,data_stage_1__3624_,
  data_stage_1__3623_,data_stage_1__3622_,data_stage_1__3621_,data_stage_1__3620_,
  data_stage_1__3619_,data_stage_1__3618_,data_stage_1__3617_,data_stage_1__3616_,
  data_stage_1__3615_,data_stage_1__3614_,data_stage_1__3613_,data_stage_1__3612_,
  data_stage_1__3611_,data_stage_1__3610_,data_stage_1__3609_,data_stage_1__3608_,
  data_stage_1__3607_,data_stage_1__3606_,data_stage_1__3605_,data_stage_1__3604_,
  data_stage_1__3603_,data_stage_1__3602_,data_stage_1__3601_,data_stage_1__3600_,
  data_stage_1__3599_,data_stage_1__3598_,data_stage_1__3597_,data_stage_1__3596_,
  data_stage_1__3595_,data_stage_1__3594_,data_stage_1__3593_,data_stage_1__3592_,
  data_stage_1__3591_,data_stage_1__3590_,data_stage_1__3589_,data_stage_1__3588_,
  data_stage_1__3587_,data_stage_1__3586_,data_stage_1__3585_,data_stage_1__3584_,
  data_stage_1__3583_,data_stage_1__3582_,data_stage_1__3581_,data_stage_1__3580_,
  data_stage_1__3579_,data_stage_1__3578_,data_stage_1__3577_,data_stage_1__3576_,
  data_stage_1__3575_,data_stage_1__3574_,data_stage_1__3573_,data_stage_1__3572_,
  data_stage_1__3571_,data_stage_1__3570_,data_stage_1__3569_,data_stage_1__3568_,
  data_stage_1__3567_,data_stage_1__3566_,data_stage_1__3565_,data_stage_1__3564_,
  data_stage_1__3563_,data_stage_1__3562_,data_stage_1__3561_,data_stage_1__3560_,
  data_stage_1__3559_,data_stage_1__3558_,data_stage_1__3557_,data_stage_1__3556_,
  data_stage_1__3555_,data_stage_1__3554_,data_stage_1__3553_,data_stage_1__3552_,
  data_stage_1__3551_,data_stage_1__3550_,data_stage_1__3549_,data_stage_1__3548_,
  data_stage_1__3547_,data_stage_1__3546_,data_stage_1__3545_,data_stage_1__3544_,
  data_stage_1__3543_,data_stage_1__3542_,data_stage_1__3541_,data_stage_1__3540_,
  data_stage_1__3539_,data_stage_1__3538_,data_stage_1__3537_,data_stage_1__3536_,
  data_stage_1__3535_,data_stage_1__3534_,data_stage_1__3533_,data_stage_1__3532_,
  data_stage_1__3531_,data_stage_1__3530_,data_stage_1__3529_,data_stage_1__3528_,
  data_stage_1__3527_,data_stage_1__3526_,data_stage_1__3525_,data_stage_1__3524_,
  data_stage_1__3523_,data_stage_1__3522_,data_stage_1__3521_,data_stage_1__3520_,
  data_stage_1__3519_,data_stage_1__3518_,data_stage_1__3517_,data_stage_1__3516_,
  data_stage_1__3515_,data_stage_1__3514_,data_stage_1__3513_,data_stage_1__3512_,
  data_stage_1__3511_,data_stage_1__3510_,data_stage_1__3509_,data_stage_1__3508_,
  data_stage_1__3507_,data_stage_1__3506_,data_stage_1__3505_,data_stage_1__3504_,
  data_stage_1__3503_,data_stage_1__3502_,data_stage_1__3501_,data_stage_1__3500_,
  data_stage_1__3499_,data_stage_1__3498_,data_stage_1__3497_,data_stage_1__3496_,
  data_stage_1__3495_,data_stage_1__3494_,data_stage_1__3493_,data_stage_1__3492_,
  data_stage_1__3491_,data_stage_1__3490_,data_stage_1__3489_,data_stage_1__3488_,
  data_stage_1__3487_,data_stage_1__3486_,data_stage_1__3485_,data_stage_1__3484_,
  data_stage_1__3483_,data_stage_1__3482_,data_stage_1__3481_,data_stage_1__3480_,
  data_stage_1__3479_,data_stage_1__3478_,data_stage_1__3477_,data_stage_1__3476_,
  data_stage_1__3475_,data_stage_1__3474_,data_stage_1__3473_,data_stage_1__3472_,
  data_stage_1__3471_,data_stage_1__3470_,data_stage_1__3469_,data_stage_1__3468_,
  data_stage_1__3467_,data_stage_1__3466_,data_stage_1__3465_,data_stage_1__3464_,
  data_stage_1__3463_,data_stage_1__3462_,data_stage_1__3461_,data_stage_1__3460_,
  data_stage_1__3459_,data_stage_1__3458_,data_stage_1__3457_,data_stage_1__3456_,
  data_stage_1__3455_,data_stage_1__3454_,data_stage_1__3453_,data_stage_1__3452_,
  data_stage_1__3451_,data_stage_1__3450_,data_stage_1__3449_,data_stage_1__3448_,
  data_stage_1__3447_,data_stage_1__3446_,data_stage_1__3445_,data_stage_1__3444_,
  data_stage_1__3443_,data_stage_1__3442_,data_stage_1__3441_,data_stage_1__3440_,
  data_stage_1__3439_,data_stage_1__3438_,data_stage_1__3437_,data_stage_1__3436_,
  data_stage_1__3435_,data_stage_1__3434_,data_stage_1__3433_,data_stage_1__3432_,
  data_stage_1__3431_,data_stage_1__3430_,data_stage_1__3429_,data_stage_1__3428_,
  data_stage_1__3427_,data_stage_1__3426_,data_stage_1__3425_,data_stage_1__3424_,
  data_stage_1__3423_,data_stage_1__3422_,data_stage_1__3421_,data_stage_1__3420_,
  data_stage_1__3419_,data_stage_1__3418_,data_stage_1__3417_,data_stage_1__3416_,
  data_stage_1__3415_,data_stage_1__3414_,data_stage_1__3413_,data_stage_1__3412_,
  data_stage_1__3411_,data_stage_1__3410_,data_stage_1__3409_,data_stage_1__3408_,
  data_stage_1__3407_,data_stage_1__3406_,data_stage_1__3405_,data_stage_1__3404_,
  data_stage_1__3403_,data_stage_1__3402_,data_stage_1__3401_,data_stage_1__3400_,
  data_stage_1__3399_,data_stage_1__3398_,data_stage_1__3397_,data_stage_1__3396_,
  data_stage_1__3395_,data_stage_1__3394_,data_stage_1__3393_,data_stage_1__3392_,
  data_stage_1__3391_,data_stage_1__3390_,data_stage_1__3389_,data_stage_1__3388_,
  data_stage_1__3387_,data_stage_1__3386_,data_stage_1__3385_,data_stage_1__3384_,
  data_stage_1__3383_,data_stage_1__3382_,data_stage_1__3381_,data_stage_1__3380_,
  data_stage_1__3379_,data_stage_1__3378_,data_stage_1__3377_,data_stage_1__3376_,
  data_stage_1__3375_,data_stage_1__3374_,data_stage_1__3373_,data_stage_1__3372_,
  data_stage_1__3371_,data_stage_1__3370_,data_stage_1__3369_,data_stage_1__3368_,
  data_stage_1__3367_,data_stage_1__3366_,data_stage_1__3365_,data_stage_1__3364_,
  data_stage_1__3363_,data_stage_1__3362_,data_stage_1__3361_,data_stage_1__3360_,
  data_stage_1__3359_,data_stage_1__3358_,data_stage_1__3357_,data_stage_1__3356_,
  data_stage_1__3355_,data_stage_1__3354_,data_stage_1__3353_,data_stage_1__3352_,
  data_stage_1__3351_,data_stage_1__3350_,data_stage_1__3349_,data_stage_1__3348_,
  data_stage_1__3347_,data_stage_1__3346_,data_stage_1__3345_,data_stage_1__3344_,
  data_stage_1__3343_,data_stage_1__3342_,data_stage_1__3341_,data_stage_1__3340_,
  data_stage_1__3339_,data_stage_1__3338_,data_stage_1__3337_,data_stage_1__3336_,
  data_stage_1__3335_,data_stage_1__3334_,data_stage_1__3333_,data_stage_1__3332_,
  data_stage_1__3331_,data_stage_1__3330_,data_stage_1__3329_,data_stage_1__3328_,
  data_stage_1__3327_,data_stage_1__3326_,data_stage_1__3325_,data_stage_1__3324_,
  data_stage_1__3323_,data_stage_1__3322_,data_stage_1__3321_,data_stage_1__3320_,
  data_stage_1__3319_,data_stage_1__3318_,data_stage_1__3317_,data_stage_1__3316_,
  data_stage_1__3315_,data_stage_1__3314_,data_stage_1__3313_,data_stage_1__3312_,
  data_stage_1__3311_,data_stage_1__3310_,data_stage_1__3309_,data_stage_1__3308_,
  data_stage_1__3307_,data_stage_1__3306_,data_stage_1__3305_,data_stage_1__3304_,
  data_stage_1__3303_,data_stage_1__3302_,data_stage_1__3301_,data_stage_1__3300_,
  data_stage_1__3299_,data_stage_1__3298_,data_stage_1__3297_,data_stage_1__3296_,
  data_stage_1__3295_,data_stage_1__3294_,data_stage_1__3293_,data_stage_1__3292_,
  data_stage_1__3291_,data_stage_1__3290_,data_stage_1__3289_,data_stage_1__3288_,
  data_stage_1__3287_,data_stage_1__3286_,data_stage_1__3285_,data_stage_1__3284_,
  data_stage_1__3283_,data_stage_1__3282_,data_stage_1__3281_,data_stage_1__3280_,
  data_stage_1__3279_,data_stage_1__3278_,data_stage_1__3277_,data_stage_1__3276_,
  data_stage_1__3275_,data_stage_1__3274_,data_stage_1__3273_,data_stage_1__3272_,
  data_stage_1__3271_,data_stage_1__3270_,data_stage_1__3269_,data_stage_1__3268_,
  data_stage_1__3267_,data_stage_1__3266_,data_stage_1__3265_,data_stage_1__3264_,
  data_stage_1__3263_,data_stage_1__3262_,data_stage_1__3261_,data_stage_1__3260_,
  data_stage_1__3259_,data_stage_1__3258_,data_stage_1__3257_,data_stage_1__3256_,
  data_stage_1__3255_,data_stage_1__3254_,data_stage_1__3253_,data_stage_1__3252_,
  data_stage_1__3251_,data_stage_1__3250_,data_stage_1__3249_,data_stage_1__3248_,
  data_stage_1__3247_,data_stage_1__3246_,data_stage_1__3245_,data_stage_1__3244_,
  data_stage_1__3243_,data_stage_1__3242_,data_stage_1__3241_,data_stage_1__3240_,
  data_stage_1__3239_,data_stage_1__3238_,data_stage_1__3237_,data_stage_1__3236_,
  data_stage_1__3235_,data_stage_1__3234_,data_stage_1__3233_,data_stage_1__3232_,
  data_stage_1__3231_,data_stage_1__3230_,data_stage_1__3229_,data_stage_1__3228_,
  data_stage_1__3227_,data_stage_1__3226_,data_stage_1__3225_,data_stage_1__3224_,
  data_stage_1__3223_,data_stage_1__3222_,data_stage_1__3221_,data_stage_1__3220_,
  data_stage_1__3219_,data_stage_1__3218_,data_stage_1__3217_,data_stage_1__3216_,
  data_stage_1__3215_,data_stage_1__3214_,data_stage_1__3213_,data_stage_1__3212_,
  data_stage_1__3211_,data_stage_1__3210_,data_stage_1__3209_,data_stage_1__3208_,
  data_stage_1__3207_,data_stage_1__3206_,data_stage_1__3205_,data_stage_1__3204_,
  data_stage_1__3203_,data_stage_1__3202_,data_stage_1__3201_,data_stage_1__3200_,
  data_stage_1__3199_,data_stage_1__3198_,data_stage_1__3197_,data_stage_1__3196_,
  data_stage_1__3195_,data_stage_1__3194_,data_stage_1__3193_,data_stage_1__3192_,
  data_stage_1__3191_,data_stage_1__3190_,data_stage_1__3189_,data_stage_1__3188_,
  data_stage_1__3187_,data_stage_1__3186_,data_stage_1__3185_,data_stage_1__3184_,
  data_stage_1__3183_,data_stage_1__3182_,data_stage_1__3181_,data_stage_1__3180_,
  data_stage_1__3179_,data_stage_1__3178_,data_stage_1__3177_,data_stage_1__3176_,
  data_stage_1__3175_,data_stage_1__3174_,data_stage_1__3173_,data_stage_1__3172_,
  data_stage_1__3171_,data_stage_1__3170_,data_stage_1__3169_,data_stage_1__3168_,
  data_stage_1__3167_,data_stage_1__3166_,data_stage_1__3165_,data_stage_1__3164_,
  data_stage_1__3163_,data_stage_1__3162_,data_stage_1__3161_,data_stage_1__3160_,
  data_stage_1__3159_,data_stage_1__3158_,data_stage_1__3157_,data_stage_1__3156_,
  data_stage_1__3155_,data_stage_1__3154_,data_stage_1__3153_,data_stage_1__3152_,
  data_stage_1__3151_,data_stage_1__3150_,data_stage_1__3149_,data_stage_1__3148_,
  data_stage_1__3147_,data_stage_1__3146_,data_stage_1__3145_,data_stage_1__3144_,
  data_stage_1__3143_,data_stage_1__3142_,data_stage_1__3141_,data_stage_1__3140_,
  data_stage_1__3139_,data_stage_1__3138_,data_stage_1__3137_,data_stage_1__3136_,
  data_stage_1__3135_,data_stage_1__3134_,data_stage_1__3133_,data_stage_1__3132_,
  data_stage_1__3131_,data_stage_1__3130_,data_stage_1__3129_,data_stage_1__3128_,
  data_stage_1__3127_,data_stage_1__3126_,data_stage_1__3125_,data_stage_1__3124_,
  data_stage_1__3123_,data_stage_1__3122_,data_stage_1__3121_,data_stage_1__3120_,
  data_stage_1__3119_,data_stage_1__3118_,data_stage_1__3117_,data_stage_1__3116_,
  data_stage_1__3115_,data_stage_1__3114_,data_stage_1__3113_,data_stage_1__3112_,
  data_stage_1__3111_,data_stage_1__3110_,data_stage_1__3109_,data_stage_1__3108_,
  data_stage_1__3107_,data_stage_1__3106_,data_stage_1__3105_,data_stage_1__3104_,
  data_stage_1__3103_,data_stage_1__3102_,data_stage_1__3101_,data_stage_1__3100_,
  data_stage_1__3099_,data_stage_1__3098_,data_stage_1__3097_,data_stage_1__3096_,
  data_stage_1__3095_,data_stage_1__3094_,data_stage_1__3093_,data_stage_1__3092_,
  data_stage_1__3091_,data_stage_1__3090_,data_stage_1__3089_,data_stage_1__3088_,
  data_stage_1__3087_,data_stage_1__3086_,data_stage_1__3085_,data_stage_1__3084_,
  data_stage_1__3083_,data_stage_1__3082_,data_stage_1__3081_,data_stage_1__3080_,
  data_stage_1__3079_,data_stage_1__3078_,data_stage_1__3077_,data_stage_1__3076_,
  data_stage_1__3075_,data_stage_1__3074_,data_stage_1__3073_,data_stage_1__3072_,
  data_stage_1__3071_,data_stage_1__3070_,data_stage_1__3069_,data_stage_1__3068_,
  data_stage_1__3067_,data_stage_1__3066_,data_stage_1__3065_,data_stage_1__3064_,
  data_stage_1__3063_,data_stage_1__3062_,data_stage_1__3061_,data_stage_1__3060_,
  data_stage_1__3059_,data_stage_1__3058_,data_stage_1__3057_,data_stage_1__3056_,
  data_stage_1__3055_,data_stage_1__3054_,data_stage_1__3053_,data_stage_1__3052_,
  data_stage_1__3051_,data_stage_1__3050_,data_stage_1__3049_,data_stage_1__3048_,
  data_stage_1__3047_,data_stage_1__3046_,data_stage_1__3045_,data_stage_1__3044_,
  data_stage_1__3043_,data_stage_1__3042_,data_stage_1__3041_,data_stage_1__3040_,
  data_stage_1__3039_,data_stage_1__3038_,data_stage_1__3037_,data_stage_1__3036_,
  data_stage_1__3035_,data_stage_1__3034_,data_stage_1__3033_,data_stage_1__3032_,
  data_stage_1__3031_,data_stage_1__3030_,data_stage_1__3029_,data_stage_1__3028_,
  data_stage_1__3027_,data_stage_1__3026_,data_stage_1__3025_,data_stage_1__3024_,
  data_stage_1__3023_,data_stage_1__3022_,data_stage_1__3021_,data_stage_1__3020_,
  data_stage_1__3019_,data_stage_1__3018_,data_stage_1__3017_,data_stage_1__3016_,
  data_stage_1__3015_,data_stage_1__3014_,data_stage_1__3013_,data_stage_1__3012_,
  data_stage_1__3011_,data_stage_1__3010_,data_stage_1__3009_,data_stage_1__3008_,
  data_stage_1__3007_,data_stage_1__3006_,data_stage_1__3005_,data_stage_1__3004_,
  data_stage_1__3003_,data_stage_1__3002_,data_stage_1__3001_,data_stage_1__3000_,
  data_stage_1__2999_,data_stage_1__2998_,data_stage_1__2997_,data_stage_1__2996_,
  data_stage_1__2995_,data_stage_1__2994_,data_stage_1__2993_,data_stage_1__2992_,
  data_stage_1__2991_,data_stage_1__2990_,data_stage_1__2989_,data_stage_1__2988_,
  data_stage_1__2987_,data_stage_1__2986_,data_stage_1__2985_,data_stage_1__2984_,
  data_stage_1__2983_,data_stage_1__2982_,data_stage_1__2981_,data_stage_1__2980_,
  data_stage_1__2979_,data_stage_1__2978_,data_stage_1__2977_,data_stage_1__2976_,
  data_stage_1__2975_,data_stage_1__2974_,data_stage_1__2973_,data_stage_1__2972_,
  data_stage_1__2971_,data_stage_1__2970_,data_stage_1__2969_,data_stage_1__2968_,
  data_stage_1__2967_,data_stage_1__2966_,data_stage_1__2965_,data_stage_1__2964_,
  data_stage_1__2963_,data_stage_1__2962_,data_stage_1__2961_,data_stage_1__2960_,
  data_stage_1__2959_,data_stage_1__2958_,data_stage_1__2957_,data_stage_1__2956_,
  data_stage_1__2955_,data_stage_1__2954_,data_stage_1__2953_,data_stage_1__2952_,
  data_stage_1__2951_,data_stage_1__2950_,data_stage_1__2949_,data_stage_1__2948_,
  data_stage_1__2947_,data_stage_1__2946_,data_stage_1__2945_,data_stage_1__2944_,
  data_stage_1__2943_,data_stage_1__2942_,data_stage_1__2941_,data_stage_1__2940_,
  data_stage_1__2939_,data_stage_1__2938_,data_stage_1__2937_,data_stage_1__2936_,
  data_stage_1__2935_,data_stage_1__2934_,data_stage_1__2933_,data_stage_1__2932_,
  data_stage_1__2931_,data_stage_1__2930_,data_stage_1__2929_,data_stage_1__2928_,
  data_stage_1__2927_,data_stage_1__2926_,data_stage_1__2925_,data_stage_1__2924_,
  data_stage_1__2923_,data_stage_1__2922_,data_stage_1__2921_,data_stage_1__2920_,
  data_stage_1__2919_,data_stage_1__2918_,data_stage_1__2917_,data_stage_1__2916_,
  data_stage_1__2915_,data_stage_1__2914_,data_stage_1__2913_,data_stage_1__2912_,
  data_stage_1__2911_,data_stage_1__2910_,data_stage_1__2909_,data_stage_1__2908_,
  data_stage_1__2907_,data_stage_1__2906_,data_stage_1__2905_,data_stage_1__2904_,
  data_stage_1__2903_,data_stage_1__2902_,data_stage_1__2901_,data_stage_1__2900_,
  data_stage_1__2899_,data_stage_1__2898_,data_stage_1__2897_,data_stage_1__2896_,
  data_stage_1__2895_,data_stage_1__2894_,data_stage_1__2893_,data_stage_1__2892_,
  data_stage_1__2891_,data_stage_1__2890_,data_stage_1__2889_,data_stage_1__2888_,
  data_stage_1__2887_,data_stage_1__2886_,data_stage_1__2885_,data_stage_1__2884_,
  data_stage_1__2883_,data_stage_1__2882_,data_stage_1__2881_,data_stage_1__2880_,
  data_stage_1__2879_,data_stage_1__2878_,data_stage_1__2877_,data_stage_1__2876_,
  data_stage_1__2875_,data_stage_1__2874_,data_stage_1__2873_,data_stage_1__2872_,
  data_stage_1__2871_,data_stage_1__2870_,data_stage_1__2869_,data_stage_1__2868_,
  data_stage_1__2867_,data_stage_1__2866_,data_stage_1__2865_,data_stage_1__2864_,
  data_stage_1__2863_,data_stage_1__2862_,data_stage_1__2861_,data_stage_1__2860_,
  data_stage_1__2859_,data_stage_1__2858_,data_stage_1__2857_,data_stage_1__2856_,
  data_stage_1__2855_,data_stage_1__2854_,data_stage_1__2853_,data_stage_1__2852_,
  data_stage_1__2851_,data_stage_1__2850_,data_stage_1__2849_,data_stage_1__2848_,
  data_stage_1__2847_,data_stage_1__2846_,data_stage_1__2845_,data_stage_1__2844_,
  data_stage_1__2843_,data_stage_1__2842_,data_stage_1__2841_,data_stage_1__2840_,
  data_stage_1__2839_,data_stage_1__2838_,data_stage_1__2837_,data_stage_1__2836_,
  data_stage_1__2835_,data_stage_1__2834_,data_stage_1__2833_,data_stage_1__2832_,
  data_stage_1__2831_,data_stage_1__2830_,data_stage_1__2829_,data_stage_1__2828_,
  data_stage_1__2827_,data_stage_1__2826_,data_stage_1__2825_,data_stage_1__2824_,
  data_stage_1__2823_,data_stage_1__2822_,data_stage_1__2821_,data_stage_1__2820_,
  data_stage_1__2819_,data_stage_1__2818_,data_stage_1__2817_,data_stage_1__2816_,
  data_stage_1__2815_,data_stage_1__2814_,data_stage_1__2813_,data_stage_1__2812_,
  data_stage_1__2811_,data_stage_1__2810_,data_stage_1__2809_,data_stage_1__2808_,
  data_stage_1__2807_,data_stage_1__2806_,data_stage_1__2805_,data_stage_1__2804_,
  data_stage_1__2803_,data_stage_1__2802_,data_stage_1__2801_,data_stage_1__2800_,
  data_stage_1__2799_,data_stage_1__2798_,data_stage_1__2797_,data_stage_1__2796_,
  data_stage_1__2795_,data_stage_1__2794_,data_stage_1__2793_,data_stage_1__2792_,
  data_stage_1__2791_,data_stage_1__2790_,data_stage_1__2789_,data_stage_1__2788_,
  data_stage_1__2787_,data_stage_1__2786_,data_stage_1__2785_,data_stage_1__2784_,
  data_stage_1__2783_,data_stage_1__2782_,data_stage_1__2781_,data_stage_1__2780_,
  data_stage_1__2779_,data_stage_1__2778_,data_stage_1__2777_,data_stage_1__2776_,
  data_stage_1__2775_,data_stage_1__2774_,data_stage_1__2773_,data_stage_1__2772_,
  data_stage_1__2771_,data_stage_1__2770_,data_stage_1__2769_,data_stage_1__2768_,
  data_stage_1__2767_,data_stage_1__2766_,data_stage_1__2765_,data_stage_1__2764_,
  data_stage_1__2763_,data_stage_1__2762_,data_stage_1__2761_,data_stage_1__2760_,
  data_stage_1__2759_,data_stage_1__2758_,data_stage_1__2757_,data_stage_1__2756_,
  data_stage_1__2755_,data_stage_1__2754_,data_stage_1__2753_,data_stage_1__2752_,
  data_stage_1__2751_,data_stage_1__2750_,data_stage_1__2749_,data_stage_1__2748_,
  data_stage_1__2747_,data_stage_1__2746_,data_stage_1__2745_,data_stage_1__2744_,
  data_stage_1__2743_,data_stage_1__2742_,data_stage_1__2741_,data_stage_1__2740_,
  data_stage_1__2739_,data_stage_1__2738_,data_stage_1__2737_,data_stage_1__2736_,
  data_stage_1__2735_,data_stage_1__2734_,data_stage_1__2733_,data_stage_1__2732_,
  data_stage_1__2731_,data_stage_1__2730_,data_stage_1__2729_,data_stage_1__2728_,
  data_stage_1__2727_,data_stage_1__2726_,data_stage_1__2725_,data_stage_1__2724_,
  data_stage_1__2723_,data_stage_1__2722_,data_stage_1__2721_,data_stage_1__2720_,
  data_stage_1__2719_,data_stage_1__2718_,data_stage_1__2717_,data_stage_1__2716_,
  data_stage_1__2715_,data_stage_1__2714_,data_stage_1__2713_,data_stage_1__2712_,
  data_stage_1__2711_,data_stage_1__2710_,data_stage_1__2709_,data_stage_1__2708_,
  data_stage_1__2707_,data_stage_1__2706_,data_stage_1__2705_,data_stage_1__2704_,
  data_stage_1__2703_,data_stage_1__2702_,data_stage_1__2701_,data_stage_1__2700_,
  data_stage_1__2699_,data_stage_1__2698_,data_stage_1__2697_,data_stage_1__2696_,
  data_stage_1__2695_,data_stage_1__2694_,data_stage_1__2693_,data_stage_1__2692_,
  data_stage_1__2691_,data_stage_1__2690_,data_stage_1__2689_,data_stage_1__2688_,
  data_stage_1__2687_,data_stage_1__2686_,data_stage_1__2685_,data_stage_1__2684_,
  data_stage_1__2683_,data_stage_1__2682_,data_stage_1__2681_,data_stage_1__2680_,
  data_stage_1__2679_,data_stage_1__2678_,data_stage_1__2677_,data_stage_1__2676_,
  data_stage_1__2675_,data_stage_1__2674_,data_stage_1__2673_,data_stage_1__2672_,
  data_stage_1__2671_,data_stage_1__2670_,data_stage_1__2669_,data_stage_1__2668_,
  data_stage_1__2667_,data_stage_1__2666_,data_stage_1__2665_,data_stage_1__2664_,
  data_stage_1__2663_,data_stage_1__2662_,data_stage_1__2661_,data_stage_1__2660_,
  data_stage_1__2659_,data_stage_1__2658_,data_stage_1__2657_,data_stage_1__2656_,
  data_stage_1__2655_,data_stage_1__2654_,data_stage_1__2653_,data_stage_1__2652_,
  data_stage_1__2651_,data_stage_1__2650_,data_stage_1__2649_,data_stage_1__2648_,
  data_stage_1__2647_,data_stage_1__2646_,data_stage_1__2645_,data_stage_1__2644_,
  data_stage_1__2643_,data_stage_1__2642_,data_stage_1__2641_,data_stage_1__2640_,
  data_stage_1__2639_,data_stage_1__2638_,data_stage_1__2637_,data_stage_1__2636_,
  data_stage_1__2635_,data_stage_1__2634_,data_stage_1__2633_,data_stage_1__2632_,
  data_stage_1__2631_,data_stage_1__2630_,data_stage_1__2629_,data_stage_1__2628_,
  data_stage_1__2627_,data_stage_1__2626_,data_stage_1__2625_,data_stage_1__2624_,
  data_stage_1__2623_,data_stage_1__2622_,data_stage_1__2621_,data_stage_1__2620_,
  data_stage_1__2619_,data_stage_1__2618_,data_stage_1__2617_,data_stage_1__2616_,
  data_stage_1__2615_,data_stage_1__2614_,data_stage_1__2613_,data_stage_1__2612_,
  data_stage_1__2611_,data_stage_1__2610_,data_stage_1__2609_,data_stage_1__2608_,
  data_stage_1__2607_,data_stage_1__2606_,data_stage_1__2605_,data_stage_1__2604_,
  data_stage_1__2603_,data_stage_1__2602_,data_stage_1__2601_,data_stage_1__2600_,
  data_stage_1__2599_,data_stage_1__2598_,data_stage_1__2597_,data_stage_1__2596_,
  data_stage_1__2595_,data_stage_1__2594_,data_stage_1__2593_,data_stage_1__2592_,
  data_stage_1__2591_,data_stage_1__2590_,data_stage_1__2589_,data_stage_1__2588_,
  data_stage_1__2587_,data_stage_1__2586_,data_stage_1__2585_,data_stage_1__2584_,
  data_stage_1__2583_,data_stage_1__2582_,data_stage_1__2581_,data_stage_1__2580_,
  data_stage_1__2579_,data_stage_1__2578_,data_stage_1__2577_,data_stage_1__2576_,
  data_stage_1__2575_,data_stage_1__2574_,data_stage_1__2573_,data_stage_1__2572_,
  data_stage_1__2571_,data_stage_1__2570_,data_stage_1__2569_,data_stage_1__2568_,
  data_stage_1__2567_,data_stage_1__2566_,data_stage_1__2565_,data_stage_1__2564_,
  data_stage_1__2563_,data_stage_1__2562_,data_stage_1__2561_,data_stage_1__2560_,
  data_stage_1__2559_,data_stage_1__2558_,data_stage_1__2557_,data_stage_1__2556_,
  data_stage_1__2555_,data_stage_1__2554_,data_stage_1__2553_,data_stage_1__2552_,
  data_stage_1__2551_,data_stage_1__2550_,data_stage_1__2549_,data_stage_1__2548_,
  data_stage_1__2547_,data_stage_1__2546_,data_stage_1__2545_,data_stage_1__2544_,
  data_stage_1__2543_,data_stage_1__2542_,data_stage_1__2541_,data_stage_1__2540_,
  data_stage_1__2539_,data_stage_1__2538_,data_stage_1__2537_,data_stage_1__2536_,
  data_stage_1__2535_,data_stage_1__2534_,data_stage_1__2533_,data_stage_1__2532_,
  data_stage_1__2531_,data_stage_1__2530_,data_stage_1__2529_,data_stage_1__2528_,
  data_stage_1__2527_,data_stage_1__2526_,data_stage_1__2525_,data_stage_1__2524_,
  data_stage_1__2523_,data_stage_1__2522_,data_stage_1__2521_,data_stage_1__2520_,
  data_stage_1__2519_,data_stage_1__2518_,data_stage_1__2517_,data_stage_1__2516_,
  data_stage_1__2515_,data_stage_1__2514_,data_stage_1__2513_,data_stage_1__2512_,
  data_stage_1__2511_,data_stage_1__2510_,data_stage_1__2509_,data_stage_1__2508_,
  data_stage_1__2507_,data_stage_1__2506_,data_stage_1__2505_,data_stage_1__2504_,
  data_stage_1__2503_,data_stage_1__2502_,data_stage_1__2501_,data_stage_1__2500_,
  data_stage_1__2499_,data_stage_1__2498_,data_stage_1__2497_,data_stage_1__2496_,
  data_stage_1__2495_,data_stage_1__2494_,data_stage_1__2493_,data_stage_1__2492_,
  data_stage_1__2491_,data_stage_1__2490_,data_stage_1__2489_,data_stage_1__2488_,
  data_stage_1__2487_,data_stage_1__2486_,data_stage_1__2485_,data_stage_1__2484_,
  data_stage_1__2483_,data_stage_1__2482_,data_stage_1__2481_,data_stage_1__2480_,
  data_stage_1__2479_,data_stage_1__2478_,data_stage_1__2477_,data_stage_1__2476_,
  data_stage_1__2475_,data_stage_1__2474_,data_stage_1__2473_,data_stage_1__2472_,
  data_stage_1__2471_,data_stage_1__2470_,data_stage_1__2469_,data_stage_1__2468_,
  data_stage_1__2467_,data_stage_1__2466_,data_stage_1__2465_,data_stage_1__2464_,
  data_stage_1__2463_,data_stage_1__2462_,data_stage_1__2461_,data_stage_1__2460_,
  data_stage_1__2459_,data_stage_1__2458_,data_stage_1__2457_,data_stage_1__2456_,
  data_stage_1__2455_,data_stage_1__2454_,data_stage_1__2453_,data_stage_1__2452_,
  data_stage_1__2451_,data_stage_1__2450_,data_stage_1__2449_,data_stage_1__2448_,
  data_stage_1__2447_,data_stage_1__2446_,data_stage_1__2445_,data_stage_1__2444_,
  data_stage_1__2443_,data_stage_1__2442_,data_stage_1__2441_,data_stage_1__2440_,
  data_stage_1__2439_,data_stage_1__2438_,data_stage_1__2437_,data_stage_1__2436_,
  data_stage_1__2435_,data_stage_1__2434_,data_stage_1__2433_,data_stage_1__2432_,
  data_stage_1__2431_,data_stage_1__2430_,data_stage_1__2429_,data_stage_1__2428_,
  data_stage_1__2427_,data_stage_1__2426_,data_stage_1__2425_,data_stage_1__2424_,
  data_stage_1__2423_,data_stage_1__2422_,data_stage_1__2421_,data_stage_1__2420_,
  data_stage_1__2419_,data_stage_1__2418_,data_stage_1__2417_,data_stage_1__2416_,
  data_stage_1__2415_,data_stage_1__2414_,data_stage_1__2413_,data_stage_1__2412_,
  data_stage_1__2411_,data_stage_1__2410_,data_stage_1__2409_,data_stage_1__2408_,
  data_stage_1__2407_,data_stage_1__2406_,data_stage_1__2405_,data_stage_1__2404_,
  data_stage_1__2403_,data_stage_1__2402_,data_stage_1__2401_,data_stage_1__2400_,
  data_stage_1__2399_,data_stage_1__2398_,data_stage_1__2397_,data_stage_1__2396_,
  data_stage_1__2395_,data_stage_1__2394_,data_stage_1__2393_,data_stage_1__2392_,
  data_stage_1__2391_,data_stage_1__2390_,data_stage_1__2389_,data_stage_1__2388_,
  data_stage_1__2387_,data_stage_1__2386_,data_stage_1__2385_,data_stage_1__2384_,
  data_stage_1__2383_,data_stage_1__2382_,data_stage_1__2381_,data_stage_1__2380_,
  data_stage_1__2379_,data_stage_1__2378_,data_stage_1__2377_,data_stage_1__2376_,
  data_stage_1__2375_,data_stage_1__2374_,data_stage_1__2373_,data_stage_1__2372_,
  data_stage_1__2371_,data_stage_1__2370_,data_stage_1__2369_,data_stage_1__2368_,
  data_stage_1__2367_,data_stage_1__2366_,data_stage_1__2365_,data_stage_1__2364_,
  data_stage_1__2363_,data_stage_1__2362_,data_stage_1__2361_,data_stage_1__2360_,
  data_stage_1__2359_,data_stage_1__2358_,data_stage_1__2357_,data_stage_1__2356_,
  data_stage_1__2355_,data_stage_1__2354_,data_stage_1__2353_,data_stage_1__2352_,
  data_stage_1__2351_,data_stage_1__2350_,data_stage_1__2349_,data_stage_1__2348_,
  data_stage_1__2347_,data_stage_1__2346_,data_stage_1__2345_,data_stage_1__2344_,
  data_stage_1__2343_,data_stage_1__2342_,data_stage_1__2341_,data_stage_1__2340_,
  data_stage_1__2339_,data_stage_1__2338_,data_stage_1__2337_,data_stage_1__2336_,
  data_stage_1__2335_,data_stage_1__2334_,data_stage_1__2333_,data_stage_1__2332_,
  data_stage_1__2331_,data_stage_1__2330_,data_stage_1__2329_,data_stage_1__2328_,
  data_stage_1__2327_,data_stage_1__2326_,data_stage_1__2325_,data_stage_1__2324_,
  data_stage_1__2323_,data_stage_1__2322_,data_stage_1__2321_,data_stage_1__2320_,
  data_stage_1__2319_,data_stage_1__2318_,data_stage_1__2317_,data_stage_1__2316_,
  data_stage_1__2315_,data_stage_1__2314_,data_stage_1__2313_,data_stage_1__2312_,
  data_stage_1__2311_,data_stage_1__2310_,data_stage_1__2309_,data_stage_1__2308_,
  data_stage_1__2307_,data_stage_1__2306_,data_stage_1__2305_,data_stage_1__2304_,
  data_stage_1__2303_,data_stage_1__2302_,data_stage_1__2301_,data_stage_1__2300_,
  data_stage_1__2299_,data_stage_1__2298_,data_stage_1__2297_,data_stage_1__2296_,
  data_stage_1__2295_,data_stage_1__2294_,data_stage_1__2293_,data_stage_1__2292_,
  data_stage_1__2291_,data_stage_1__2290_,data_stage_1__2289_,data_stage_1__2288_,
  data_stage_1__2287_,data_stage_1__2286_,data_stage_1__2285_,data_stage_1__2284_,
  data_stage_1__2283_,data_stage_1__2282_,data_stage_1__2281_,data_stage_1__2280_,
  data_stage_1__2279_,data_stage_1__2278_,data_stage_1__2277_,data_stage_1__2276_,
  data_stage_1__2275_,data_stage_1__2274_,data_stage_1__2273_,data_stage_1__2272_,
  data_stage_1__2271_,data_stage_1__2270_,data_stage_1__2269_,data_stage_1__2268_,
  data_stage_1__2267_,data_stage_1__2266_,data_stage_1__2265_,data_stage_1__2264_,
  data_stage_1__2263_,data_stage_1__2262_,data_stage_1__2261_,data_stage_1__2260_,
  data_stage_1__2259_,data_stage_1__2258_,data_stage_1__2257_,data_stage_1__2256_,
  data_stage_1__2255_,data_stage_1__2254_,data_stage_1__2253_,data_stage_1__2252_,
  data_stage_1__2251_,data_stage_1__2250_,data_stage_1__2249_,data_stage_1__2248_,
  data_stage_1__2247_,data_stage_1__2246_,data_stage_1__2245_,data_stage_1__2244_,
  data_stage_1__2243_,data_stage_1__2242_,data_stage_1__2241_,data_stage_1__2240_,
  data_stage_1__2239_,data_stage_1__2238_,data_stage_1__2237_,data_stage_1__2236_,
  data_stage_1__2235_,data_stage_1__2234_,data_stage_1__2233_,data_stage_1__2232_,
  data_stage_1__2231_,data_stage_1__2230_,data_stage_1__2229_,data_stage_1__2228_,
  data_stage_1__2227_,data_stage_1__2226_,data_stage_1__2225_,data_stage_1__2224_,
  data_stage_1__2223_,data_stage_1__2222_,data_stage_1__2221_,data_stage_1__2220_,
  data_stage_1__2219_,data_stage_1__2218_,data_stage_1__2217_,data_stage_1__2216_,
  data_stage_1__2215_,data_stage_1__2214_,data_stage_1__2213_,data_stage_1__2212_,
  data_stage_1__2211_,data_stage_1__2210_,data_stage_1__2209_,data_stage_1__2208_,
  data_stage_1__2207_,data_stage_1__2206_,data_stage_1__2205_,data_stage_1__2204_,
  data_stage_1__2203_,data_stage_1__2202_,data_stage_1__2201_,data_stage_1__2200_,
  data_stage_1__2199_,data_stage_1__2198_,data_stage_1__2197_,data_stage_1__2196_,
  data_stage_1__2195_,data_stage_1__2194_,data_stage_1__2193_,data_stage_1__2192_,
  data_stage_1__2191_,data_stage_1__2190_,data_stage_1__2189_,data_stage_1__2188_,
  data_stage_1__2187_,data_stage_1__2186_,data_stage_1__2185_,data_stage_1__2184_,
  data_stage_1__2183_,data_stage_1__2182_,data_stage_1__2181_,data_stage_1__2180_,
  data_stage_1__2179_,data_stage_1__2178_,data_stage_1__2177_,data_stage_1__2176_,
  data_stage_1__2175_,data_stage_1__2174_,data_stage_1__2173_,data_stage_1__2172_,
  data_stage_1__2171_,data_stage_1__2170_,data_stage_1__2169_,data_stage_1__2168_,
  data_stage_1__2167_,data_stage_1__2166_,data_stage_1__2165_,data_stage_1__2164_,
  data_stage_1__2163_,data_stage_1__2162_,data_stage_1__2161_,data_stage_1__2160_,
  data_stage_1__2159_,data_stage_1__2158_,data_stage_1__2157_,data_stage_1__2156_,
  data_stage_1__2155_,data_stage_1__2154_,data_stage_1__2153_,data_stage_1__2152_,
  data_stage_1__2151_,data_stage_1__2150_,data_stage_1__2149_,data_stage_1__2148_,
  data_stage_1__2147_,data_stage_1__2146_,data_stage_1__2145_,data_stage_1__2144_,
  data_stage_1__2143_,data_stage_1__2142_,data_stage_1__2141_,data_stage_1__2140_,
  data_stage_1__2139_,data_stage_1__2138_,data_stage_1__2137_,data_stage_1__2136_,
  data_stage_1__2135_,data_stage_1__2134_,data_stage_1__2133_,data_stage_1__2132_,
  data_stage_1__2131_,data_stage_1__2130_,data_stage_1__2129_,data_stage_1__2128_,
  data_stage_1__2127_,data_stage_1__2126_,data_stage_1__2125_,data_stage_1__2124_,
  data_stage_1__2123_,data_stage_1__2122_,data_stage_1__2121_,data_stage_1__2120_,
  data_stage_1__2119_,data_stage_1__2118_,data_stage_1__2117_,data_stage_1__2116_,
  data_stage_1__2115_,data_stage_1__2114_,data_stage_1__2113_,data_stage_1__2112_,
  data_stage_1__2111_,data_stage_1__2110_,data_stage_1__2109_,data_stage_1__2108_,
  data_stage_1__2107_,data_stage_1__2106_,data_stage_1__2105_,data_stage_1__2104_,
  data_stage_1__2103_,data_stage_1__2102_,data_stage_1__2101_,data_stage_1__2100_,
  data_stage_1__2099_,data_stage_1__2098_,data_stage_1__2097_,data_stage_1__2096_,
  data_stage_1__2095_,data_stage_1__2094_,data_stage_1__2093_,data_stage_1__2092_,
  data_stage_1__2091_,data_stage_1__2090_,data_stage_1__2089_,data_stage_1__2088_,
  data_stage_1__2087_,data_stage_1__2086_,data_stage_1__2085_,data_stage_1__2084_,
  data_stage_1__2083_,data_stage_1__2082_,data_stage_1__2081_,data_stage_1__2080_,
  data_stage_1__2079_,data_stage_1__2078_,data_stage_1__2077_,data_stage_1__2076_,
  data_stage_1__2075_,data_stage_1__2074_,data_stage_1__2073_,data_stage_1__2072_,
  data_stage_1__2071_,data_stage_1__2070_,data_stage_1__2069_,data_stage_1__2068_,
  data_stage_1__2067_,data_stage_1__2066_,data_stage_1__2065_,data_stage_1__2064_,
  data_stage_1__2063_,data_stage_1__2062_,data_stage_1__2061_,data_stage_1__2060_,
  data_stage_1__2059_,data_stage_1__2058_,data_stage_1__2057_,data_stage_1__2056_,
  data_stage_1__2055_,data_stage_1__2054_,data_stage_1__2053_,data_stage_1__2052_,
  data_stage_1__2051_,data_stage_1__2050_,data_stage_1__2049_,data_stage_1__2048_,
  data_stage_1__2047_,data_stage_1__2046_,data_stage_1__2045_,data_stage_1__2044_,
  data_stage_1__2043_,data_stage_1__2042_,data_stage_1__2041_,data_stage_1__2040_,
  data_stage_1__2039_,data_stage_1__2038_,data_stage_1__2037_,data_stage_1__2036_,
  data_stage_1__2035_,data_stage_1__2034_,data_stage_1__2033_,data_stage_1__2032_,
  data_stage_1__2031_,data_stage_1__2030_,data_stage_1__2029_,data_stage_1__2028_,
  data_stage_1__2027_,data_stage_1__2026_,data_stage_1__2025_,data_stage_1__2024_,
  data_stage_1__2023_,data_stage_1__2022_,data_stage_1__2021_,data_stage_1__2020_,
  data_stage_1__2019_,data_stage_1__2018_,data_stage_1__2017_,data_stage_1__2016_,
  data_stage_1__2015_,data_stage_1__2014_,data_stage_1__2013_,data_stage_1__2012_,
  data_stage_1__2011_,data_stage_1__2010_,data_stage_1__2009_,data_stage_1__2008_,
  data_stage_1__2007_,data_stage_1__2006_,data_stage_1__2005_,data_stage_1__2004_,
  data_stage_1__2003_,data_stage_1__2002_,data_stage_1__2001_,data_stage_1__2000_,
  data_stage_1__1999_,data_stage_1__1998_,data_stage_1__1997_,data_stage_1__1996_,
  data_stage_1__1995_,data_stage_1__1994_,data_stage_1__1993_,data_stage_1__1992_,
  data_stage_1__1991_,data_stage_1__1990_,data_stage_1__1989_,data_stage_1__1988_,
  data_stage_1__1987_,data_stage_1__1986_,data_stage_1__1985_,data_stage_1__1984_,
  data_stage_1__1983_,data_stage_1__1982_,data_stage_1__1981_,data_stage_1__1980_,
  data_stage_1__1979_,data_stage_1__1978_,data_stage_1__1977_,data_stage_1__1976_,
  data_stage_1__1975_,data_stage_1__1974_,data_stage_1__1973_,data_stage_1__1972_,
  data_stage_1__1971_,data_stage_1__1970_,data_stage_1__1969_,data_stage_1__1968_,
  data_stage_1__1967_,data_stage_1__1966_,data_stage_1__1965_,data_stage_1__1964_,
  data_stage_1__1963_,data_stage_1__1962_,data_stage_1__1961_,data_stage_1__1960_,
  data_stage_1__1959_,data_stage_1__1958_,data_stage_1__1957_,data_stage_1__1956_,
  data_stage_1__1955_,data_stage_1__1954_,data_stage_1__1953_,data_stage_1__1952_,
  data_stage_1__1951_,data_stage_1__1950_,data_stage_1__1949_,data_stage_1__1948_,
  data_stage_1__1947_,data_stage_1__1946_,data_stage_1__1945_,data_stage_1__1944_,
  data_stage_1__1943_,data_stage_1__1942_,data_stage_1__1941_,data_stage_1__1940_,
  data_stage_1__1939_,data_stage_1__1938_,data_stage_1__1937_,data_stage_1__1936_,
  data_stage_1__1935_,data_stage_1__1934_,data_stage_1__1933_,data_stage_1__1932_,
  data_stage_1__1931_,data_stage_1__1930_,data_stage_1__1929_,data_stage_1__1928_,
  data_stage_1__1927_,data_stage_1__1926_,data_stage_1__1925_,data_stage_1__1924_,
  data_stage_1__1923_,data_stage_1__1922_,data_stage_1__1921_,data_stage_1__1920_,
  data_stage_1__1919_,data_stage_1__1918_,data_stage_1__1917_,data_stage_1__1916_,
  data_stage_1__1915_,data_stage_1__1914_,data_stage_1__1913_,data_stage_1__1912_,
  data_stage_1__1911_,data_stage_1__1910_,data_stage_1__1909_,data_stage_1__1908_,
  data_stage_1__1907_,data_stage_1__1906_,data_stage_1__1905_,data_stage_1__1904_,
  data_stage_1__1903_,data_stage_1__1902_,data_stage_1__1901_,data_stage_1__1900_,
  data_stage_1__1899_,data_stage_1__1898_,data_stage_1__1897_,data_stage_1__1896_,
  data_stage_1__1895_,data_stage_1__1894_,data_stage_1__1893_,data_stage_1__1892_,
  data_stage_1__1891_,data_stage_1__1890_,data_stage_1__1889_,data_stage_1__1888_,
  data_stage_1__1887_,data_stage_1__1886_,data_stage_1__1885_,data_stage_1__1884_,
  data_stage_1__1883_,data_stage_1__1882_,data_stage_1__1881_,data_stage_1__1880_,
  data_stage_1__1879_,data_stage_1__1878_,data_stage_1__1877_,data_stage_1__1876_,
  data_stage_1__1875_,data_stage_1__1874_,data_stage_1__1873_,data_stage_1__1872_,
  data_stage_1__1871_,data_stage_1__1870_,data_stage_1__1869_,data_stage_1__1868_,
  data_stage_1__1867_,data_stage_1__1866_,data_stage_1__1865_,data_stage_1__1864_,
  data_stage_1__1863_,data_stage_1__1862_,data_stage_1__1861_,data_stage_1__1860_,
  data_stage_1__1859_,data_stage_1__1858_,data_stage_1__1857_,data_stage_1__1856_,
  data_stage_1__1855_,data_stage_1__1854_,data_stage_1__1853_,data_stage_1__1852_,
  data_stage_1__1851_,data_stage_1__1850_,data_stage_1__1849_,data_stage_1__1848_,
  data_stage_1__1847_,data_stage_1__1846_,data_stage_1__1845_,data_stage_1__1844_,
  data_stage_1__1843_,data_stage_1__1842_,data_stage_1__1841_,data_stage_1__1840_,
  data_stage_1__1839_,data_stage_1__1838_,data_stage_1__1837_,data_stage_1__1836_,
  data_stage_1__1835_,data_stage_1__1834_,data_stage_1__1833_,data_stage_1__1832_,
  data_stage_1__1831_,data_stage_1__1830_,data_stage_1__1829_,data_stage_1__1828_,
  data_stage_1__1827_,data_stage_1__1826_,data_stage_1__1825_,data_stage_1__1824_,
  data_stage_1__1823_,data_stage_1__1822_,data_stage_1__1821_,data_stage_1__1820_,
  data_stage_1__1819_,data_stage_1__1818_,data_stage_1__1817_,data_stage_1__1816_,
  data_stage_1__1815_,data_stage_1__1814_,data_stage_1__1813_,data_stage_1__1812_,
  data_stage_1__1811_,data_stage_1__1810_,data_stage_1__1809_,data_stage_1__1808_,
  data_stage_1__1807_,data_stage_1__1806_,data_stage_1__1805_,data_stage_1__1804_,
  data_stage_1__1803_,data_stage_1__1802_,data_stage_1__1801_,data_stage_1__1800_,
  data_stage_1__1799_,data_stage_1__1798_,data_stage_1__1797_,data_stage_1__1796_,
  data_stage_1__1795_,data_stage_1__1794_,data_stage_1__1793_,data_stage_1__1792_,
  data_stage_1__1791_,data_stage_1__1790_,data_stage_1__1789_,data_stage_1__1788_,
  data_stage_1__1787_,data_stage_1__1786_,data_stage_1__1785_,data_stage_1__1784_,
  data_stage_1__1783_,data_stage_1__1782_,data_stage_1__1781_,data_stage_1__1780_,
  data_stage_1__1779_,data_stage_1__1778_,data_stage_1__1777_,data_stage_1__1776_,
  data_stage_1__1775_,data_stage_1__1774_,data_stage_1__1773_,data_stage_1__1772_,
  data_stage_1__1771_,data_stage_1__1770_,data_stage_1__1769_,data_stage_1__1768_,
  data_stage_1__1767_,data_stage_1__1766_,data_stage_1__1765_,data_stage_1__1764_,
  data_stage_1__1763_,data_stage_1__1762_,data_stage_1__1761_,data_stage_1__1760_,
  data_stage_1__1759_,data_stage_1__1758_,data_stage_1__1757_,data_stage_1__1756_,
  data_stage_1__1755_,data_stage_1__1754_,data_stage_1__1753_,data_stage_1__1752_,
  data_stage_1__1751_,data_stage_1__1750_,data_stage_1__1749_,data_stage_1__1748_,
  data_stage_1__1747_,data_stage_1__1746_,data_stage_1__1745_,data_stage_1__1744_,
  data_stage_1__1743_,data_stage_1__1742_,data_stage_1__1741_,data_stage_1__1740_,
  data_stage_1__1739_,data_stage_1__1738_,data_stage_1__1737_,data_stage_1__1736_,
  data_stage_1__1735_,data_stage_1__1734_,data_stage_1__1733_,data_stage_1__1732_,
  data_stage_1__1731_,data_stage_1__1730_,data_stage_1__1729_,data_stage_1__1728_,
  data_stage_1__1727_,data_stage_1__1726_,data_stage_1__1725_,data_stage_1__1724_,
  data_stage_1__1723_,data_stage_1__1722_,data_stage_1__1721_,data_stage_1__1720_,
  data_stage_1__1719_,data_stage_1__1718_,data_stage_1__1717_,data_stage_1__1716_,
  data_stage_1__1715_,data_stage_1__1714_,data_stage_1__1713_,data_stage_1__1712_,
  data_stage_1__1711_,data_stage_1__1710_,data_stage_1__1709_,data_stage_1__1708_,
  data_stage_1__1707_,data_stage_1__1706_,data_stage_1__1705_,data_stage_1__1704_,
  data_stage_1__1703_,data_stage_1__1702_,data_stage_1__1701_,data_stage_1__1700_,
  data_stage_1__1699_,data_stage_1__1698_,data_stage_1__1697_,data_stage_1__1696_,
  data_stage_1__1695_,data_stage_1__1694_,data_stage_1__1693_,data_stage_1__1692_,
  data_stage_1__1691_,data_stage_1__1690_,data_stage_1__1689_,data_stage_1__1688_,
  data_stage_1__1687_,data_stage_1__1686_,data_stage_1__1685_,data_stage_1__1684_,
  data_stage_1__1683_,data_stage_1__1682_,data_stage_1__1681_,data_stage_1__1680_,
  data_stage_1__1679_,data_stage_1__1678_,data_stage_1__1677_,data_stage_1__1676_,
  data_stage_1__1675_,data_stage_1__1674_,data_stage_1__1673_,data_stage_1__1672_,
  data_stage_1__1671_,data_stage_1__1670_,data_stage_1__1669_,data_stage_1__1668_,
  data_stage_1__1667_,data_stage_1__1666_,data_stage_1__1665_,data_stage_1__1664_,
  data_stage_1__1663_,data_stage_1__1662_,data_stage_1__1661_,data_stage_1__1660_,
  data_stage_1__1659_,data_stage_1__1658_,data_stage_1__1657_,data_stage_1__1656_,
  data_stage_1__1655_,data_stage_1__1654_,data_stage_1__1653_,data_stage_1__1652_,
  data_stage_1__1651_,data_stage_1__1650_,data_stage_1__1649_,data_stage_1__1648_,
  data_stage_1__1647_,data_stage_1__1646_,data_stage_1__1645_,data_stage_1__1644_,
  data_stage_1__1643_,data_stage_1__1642_,data_stage_1__1641_,data_stage_1__1640_,
  data_stage_1__1639_,data_stage_1__1638_,data_stage_1__1637_,data_stage_1__1636_,
  data_stage_1__1635_,data_stage_1__1634_,data_stage_1__1633_,data_stage_1__1632_,
  data_stage_1__1631_,data_stage_1__1630_,data_stage_1__1629_,data_stage_1__1628_,
  data_stage_1__1627_,data_stage_1__1626_,data_stage_1__1625_,data_stage_1__1624_,
  data_stage_1__1623_,data_stage_1__1622_,data_stage_1__1621_,data_stage_1__1620_,
  data_stage_1__1619_,data_stage_1__1618_,data_stage_1__1617_,data_stage_1__1616_,
  data_stage_1__1615_,data_stage_1__1614_,data_stage_1__1613_,data_stage_1__1612_,
  data_stage_1__1611_,data_stage_1__1610_,data_stage_1__1609_,data_stage_1__1608_,
  data_stage_1__1607_,data_stage_1__1606_,data_stage_1__1605_,data_stage_1__1604_,
  data_stage_1__1603_,data_stage_1__1602_,data_stage_1__1601_,data_stage_1__1600_,
  data_stage_1__1599_,data_stage_1__1598_,data_stage_1__1597_,data_stage_1__1596_,
  data_stage_1__1595_,data_stage_1__1594_,data_stage_1__1593_,data_stage_1__1592_,
  data_stage_1__1591_,data_stage_1__1590_,data_stage_1__1589_,data_stage_1__1588_,
  data_stage_1__1587_,data_stage_1__1586_,data_stage_1__1585_,data_stage_1__1584_,
  data_stage_1__1583_,data_stage_1__1582_,data_stage_1__1581_,data_stage_1__1580_,
  data_stage_1__1579_,data_stage_1__1578_,data_stage_1__1577_,data_stage_1__1576_,
  data_stage_1__1575_,data_stage_1__1574_,data_stage_1__1573_,data_stage_1__1572_,
  data_stage_1__1571_,data_stage_1__1570_,data_stage_1__1569_,data_stage_1__1568_,
  data_stage_1__1567_,data_stage_1__1566_,data_stage_1__1565_,data_stage_1__1564_,
  data_stage_1__1563_,data_stage_1__1562_,data_stage_1__1561_,data_stage_1__1560_,
  data_stage_1__1559_,data_stage_1__1558_,data_stage_1__1557_,data_stage_1__1556_,
  data_stage_1__1555_,data_stage_1__1554_,data_stage_1__1553_,data_stage_1__1552_,
  data_stage_1__1551_,data_stage_1__1550_,data_stage_1__1549_,data_stage_1__1548_,
  data_stage_1__1547_,data_stage_1__1546_,data_stage_1__1545_,data_stage_1__1544_,
  data_stage_1__1543_,data_stage_1__1542_,data_stage_1__1541_,data_stage_1__1540_,
  data_stage_1__1539_,data_stage_1__1538_,data_stage_1__1537_,data_stage_1__1536_,
  data_stage_1__1535_,data_stage_1__1534_,data_stage_1__1533_,data_stage_1__1532_,
  data_stage_1__1531_,data_stage_1__1530_,data_stage_1__1529_,data_stage_1__1528_,
  data_stage_1__1527_,data_stage_1__1526_,data_stage_1__1525_,data_stage_1__1524_,
  data_stage_1__1523_,data_stage_1__1522_,data_stage_1__1521_,data_stage_1__1520_,
  data_stage_1__1519_,data_stage_1__1518_,data_stage_1__1517_,data_stage_1__1516_,
  data_stage_1__1515_,data_stage_1__1514_,data_stage_1__1513_,data_stage_1__1512_,
  data_stage_1__1511_,data_stage_1__1510_,data_stage_1__1509_,data_stage_1__1508_,
  data_stage_1__1507_,data_stage_1__1506_,data_stage_1__1505_,data_stage_1__1504_,
  data_stage_1__1503_,data_stage_1__1502_,data_stage_1__1501_,data_stage_1__1500_,
  data_stage_1__1499_,data_stage_1__1498_,data_stage_1__1497_,data_stage_1__1496_,
  data_stage_1__1495_,data_stage_1__1494_,data_stage_1__1493_,data_stage_1__1492_,
  data_stage_1__1491_,data_stage_1__1490_,data_stage_1__1489_,data_stage_1__1488_,
  data_stage_1__1487_,data_stage_1__1486_,data_stage_1__1485_,data_stage_1__1484_,
  data_stage_1__1483_,data_stage_1__1482_,data_stage_1__1481_,data_stage_1__1480_,
  data_stage_1__1479_,data_stage_1__1478_,data_stage_1__1477_,data_stage_1__1476_,
  data_stage_1__1475_,data_stage_1__1474_,data_stage_1__1473_,data_stage_1__1472_,
  data_stage_1__1471_,data_stage_1__1470_,data_stage_1__1469_,data_stage_1__1468_,
  data_stage_1__1467_,data_stage_1__1466_,data_stage_1__1465_,data_stage_1__1464_,
  data_stage_1__1463_,data_stage_1__1462_,data_stage_1__1461_,data_stage_1__1460_,
  data_stage_1__1459_,data_stage_1__1458_,data_stage_1__1457_,data_stage_1__1456_,
  data_stage_1__1455_,data_stage_1__1454_,data_stage_1__1453_,data_stage_1__1452_,
  data_stage_1__1451_,data_stage_1__1450_,data_stage_1__1449_,data_stage_1__1448_,
  data_stage_1__1447_,data_stage_1__1446_,data_stage_1__1445_,data_stage_1__1444_,
  data_stage_1__1443_,data_stage_1__1442_,data_stage_1__1441_,data_stage_1__1440_,
  data_stage_1__1439_,data_stage_1__1438_,data_stage_1__1437_,data_stage_1__1436_,
  data_stage_1__1435_,data_stage_1__1434_,data_stage_1__1433_,data_stage_1__1432_,
  data_stage_1__1431_,data_stage_1__1430_,data_stage_1__1429_,data_stage_1__1428_,
  data_stage_1__1427_,data_stage_1__1426_,data_stage_1__1425_,data_stage_1__1424_,
  data_stage_1__1423_,data_stage_1__1422_,data_stage_1__1421_,data_stage_1__1420_,
  data_stage_1__1419_,data_stage_1__1418_,data_stage_1__1417_,data_stage_1__1416_,
  data_stage_1__1415_,data_stage_1__1414_,data_stage_1__1413_,data_stage_1__1412_,
  data_stage_1__1411_,data_stage_1__1410_,data_stage_1__1409_,data_stage_1__1408_,
  data_stage_1__1407_,data_stage_1__1406_,data_stage_1__1405_,data_stage_1__1404_,
  data_stage_1__1403_,data_stage_1__1402_,data_stage_1__1401_,data_stage_1__1400_,
  data_stage_1__1399_,data_stage_1__1398_,data_stage_1__1397_,data_stage_1__1396_,
  data_stage_1__1395_,data_stage_1__1394_,data_stage_1__1393_,data_stage_1__1392_,
  data_stage_1__1391_,data_stage_1__1390_,data_stage_1__1389_,data_stage_1__1388_,
  data_stage_1__1387_,data_stage_1__1386_,data_stage_1__1385_,data_stage_1__1384_,
  data_stage_1__1383_,data_stage_1__1382_,data_stage_1__1381_,data_stage_1__1380_,
  data_stage_1__1379_,data_stage_1__1378_,data_stage_1__1377_,data_stage_1__1376_,
  data_stage_1__1375_,data_stage_1__1374_,data_stage_1__1373_,data_stage_1__1372_,
  data_stage_1__1371_,data_stage_1__1370_,data_stage_1__1369_,data_stage_1__1368_,
  data_stage_1__1367_,data_stage_1__1366_,data_stage_1__1365_,data_stage_1__1364_,
  data_stage_1__1363_,data_stage_1__1362_,data_stage_1__1361_,data_stage_1__1360_,
  data_stage_1__1359_,data_stage_1__1358_,data_stage_1__1357_,data_stage_1__1356_,
  data_stage_1__1355_,data_stage_1__1354_,data_stage_1__1353_,data_stage_1__1352_,
  data_stage_1__1351_,data_stage_1__1350_,data_stage_1__1349_,data_stage_1__1348_,
  data_stage_1__1347_,data_stage_1__1346_,data_stage_1__1345_,data_stage_1__1344_,
  data_stage_1__1343_,data_stage_1__1342_,data_stage_1__1341_,data_stage_1__1340_,
  data_stage_1__1339_,data_stage_1__1338_,data_stage_1__1337_,data_stage_1__1336_,
  data_stage_1__1335_,data_stage_1__1334_,data_stage_1__1333_,data_stage_1__1332_,
  data_stage_1__1331_,data_stage_1__1330_,data_stage_1__1329_,data_stage_1__1328_,
  data_stage_1__1327_,data_stage_1__1326_,data_stage_1__1325_,data_stage_1__1324_,
  data_stage_1__1323_,data_stage_1__1322_,data_stage_1__1321_,data_stage_1__1320_,
  data_stage_1__1319_,data_stage_1__1318_,data_stage_1__1317_,data_stage_1__1316_,
  data_stage_1__1315_,data_stage_1__1314_,data_stage_1__1313_,data_stage_1__1312_,
  data_stage_1__1311_,data_stage_1__1310_,data_stage_1__1309_,data_stage_1__1308_,
  data_stage_1__1307_,data_stage_1__1306_,data_stage_1__1305_,data_stage_1__1304_,
  data_stage_1__1303_,data_stage_1__1302_,data_stage_1__1301_,data_stage_1__1300_,
  data_stage_1__1299_,data_stage_1__1298_,data_stage_1__1297_,data_stage_1__1296_,
  data_stage_1__1295_,data_stage_1__1294_,data_stage_1__1293_,data_stage_1__1292_,
  data_stage_1__1291_,data_stage_1__1290_,data_stage_1__1289_,data_stage_1__1288_,
  data_stage_1__1287_,data_stage_1__1286_,data_stage_1__1285_,data_stage_1__1284_,
  data_stage_1__1283_,data_stage_1__1282_,data_stage_1__1281_,data_stage_1__1280_,
  data_stage_1__1279_,data_stage_1__1278_,data_stage_1__1277_,data_stage_1__1276_,
  data_stage_1__1275_,data_stage_1__1274_,data_stage_1__1273_,data_stage_1__1272_,
  data_stage_1__1271_,data_stage_1__1270_,data_stage_1__1269_,data_stage_1__1268_,
  data_stage_1__1267_,data_stage_1__1266_,data_stage_1__1265_,data_stage_1__1264_,
  data_stage_1__1263_,data_stage_1__1262_,data_stage_1__1261_,data_stage_1__1260_,
  data_stage_1__1259_,data_stage_1__1258_,data_stage_1__1257_,data_stage_1__1256_,
  data_stage_1__1255_,data_stage_1__1254_,data_stage_1__1253_,data_stage_1__1252_,
  data_stage_1__1251_,data_stage_1__1250_,data_stage_1__1249_,data_stage_1__1248_,
  data_stage_1__1247_,data_stage_1__1246_,data_stage_1__1245_,data_stage_1__1244_,
  data_stage_1__1243_,data_stage_1__1242_,data_stage_1__1241_,data_stage_1__1240_,
  data_stage_1__1239_,data_stage_1__1238_,data_stage_1__1237_,data_stage_1__1236_,
  data_stage_1__1235_,data_stage_1__1234_,data_stage_1__1233_,data_stage_1__1232_,
  data_stage_1__1231_,data_stage_1__1230_,data_stage_1__1229_,data_stage_1__1228_,
  data_stage_1__1227_,data_stage_1__1226_,data_stage_1__1225_,data_stage_1__1224_,
  data_stage_1__1223_,data_stage_1__1222_,data_stage_1__1221_,data_stage_1__1220_,
  data_stage_1__1219_,data_stage_1__1218_,data_stage_1__1217_,data_stage_1__1216_,
  data_stage_1__1215_,data_stage_1__1214_,data_stage_1__1213_,data_stage_1__1212_,
  data_stage_1__1211_,data_stage_1__1210_,data_stage_1__1209_,data_stage_1__1208_,
  data_stage_1__1207_,data_stage_1__1206_,data_stage_1__1205_,data_stage_1__1204_,
  data_stage_1__1203_,data_stage_1__1202_,data_stage_1__1201_,data_stage_1__1200_,
  data_stage_1__1199_,data_stage_1__1198_,data_stage_1__1197_,data_stage_1__1196_,
  data_stage_1__1195_,data_stage_1__1194_,data_stage_1__1193_,data_stage_1__1192_,
  data_stage_1__1191_,data_stage_1__1190_,data_stage_1__1189_,data_stage_1__1188_,
  data_stage_1__1187_,data_stage_1__1186_,data_stage_1__1185_,data_stage_1__1184_,
  data_stage_1__1183_,data_stage_1__1182_,data_stage_1__1181_,data_stage_1__1180_,
  data_stage_1__1179_,data_stage_1__1178_,data_stage_1__1177_,data_stage_1__1176_,
  data_stage_1__1175_,data_stage_1__1174_,data_stage_1__1173_,data_stage_1__1172_,
  data_stage_1__1171_,data_stage_1__1170_,data_stage_1__1169_,data_stage_1__1168_,
  data_stage_1__1167_,data_stage_1__1166_,data_stage_1__1165_,data_stage_1__1164_,
  data_stage_1__1163_,data_stage_1__1162_,data_stage_1__1161_,data_stage_1__1160_,
  data_stage_1__1159_,data_stage_1__1158_,data_stage_1__1157_,data_stage_1__1156_,
  data_stage_1__1155_,data_stage_1__1154_,data_stage_1__1153_,data_stage_1__1152_,
  data_stage_1__1151_,data_stage_1__1150_,data_stage_1__1149_,data_stage_1__1148_,
  data_stage_1__1147_,data_stage_1__1146_,data_stage_1__1145_,data_stage_1__1144_,
  data_stage_1__1143_,data_stage_1__1142_,data_stage_1__1141_,data_stage_1__1140_,
  data_stage_1__1139_,data_stage_1__1138_,data_stage_1__1137_,data_stage_1__1136_,
  data_stage_1__1135_,data_stage_1__1134_,data_stage_1__1133_,data_stage_1__1132_,
  data_stage_1__1131_,data_stage_1__1130_,data_stage_1__1129_,data_stage_1__1128_,
  data_stage_1__1127_,data_stage_1__1126_,data_stage_1__1125_,data_stage_1__1124_,
  data_stage_1__1123_,data_stage_1__1122_,data_stage_1__1121_,data_stage_1__1120_,
  data_stage_1__1119_,data_stage_1__1118_,data_stage_1__1117_,data_stage_1__1116_,
  data_stage_1__1115_,data_stage_1__1114_,data_stage_1__1113_,data_stage_1__1112_,
  data_stage_1__1111_,data_stage_1__1110_,data_stage_1__1109_,data_stage_1__1108_,
  data_stage_1__1107_,data_stage_1__1106_,data_stage_1__1105_,data_stage_1__1104_,
  data_stage_1__1103_,data_stage_1__1102_,data_stage_1__1101_,data_stage_1__1100_,
  data_stage_1__1099_,data_stage_1__1098_,data_stage_1__1097_,data_stage_1__1096_,
  data_stage_1__1095_,data_stage_1__1094_,data_stage_1__1093_,data_stage_1__1092_,
  data_stage_1__1091_,data_stage_1__1090_,data_stage_1__1089_,data_stage_1__1088_,
  data_stage_1__1087_,data_stage_1__1086_,data_stage_1__1085_,data_stage_1__1084_,
  data_stage_1__1083_,data_stage_1__1082_,data_stage_1__1081_,data_stage_1__1080_,
  data_stage_1__1079_,data_stage_1__1078_,data_stage_1__1077_,data_stage_1__1076_,
  data_stage_1__1075_,data_stage_1__1074_,data_stage_1__1073_,data_stage_1__1072_,
  data_stage_1__1071_,data_stage_1__1070_,data_stage_1__1069_,data_stage_1__1068_,
  data_stage_1__1067_,data_stage_1__1066_,data_stage_1__1065_,data_stage_1__1064_,
  data_stage_1__1063_,data_stage_1__1062_,data_stage_1__1061_,data_stage_1__1060_,
  data_stage_1__1059_,data_stage_1__1058_,data_stage_1__1057_,data_stage_1__1056_,
  data_stage_1__1055_,data_stage_1__1054_,data_stage_1__1053_,data_stage_1__1052_,
  data_stage_1__1051_,data_stage_1__1050_,data_stage_1__1049_,data_stage_1__1048_,
  data_stage_1__1047_,data_stage_1__1046_,data_stage_1__1045_,data_stage_1__1044_,
  data_stage_1__1043_,data_stage_1__1042_,data_stage_1__1041_,data_stage_1__1040_,
  data_stage_1__1039_,data_stage_1__1038_,data_stage_1__1037_,data_stage_1__1036_,
  data_stage_1__1035_,data_stage_1__1034_,data_stage_1__1033_,data_stage_1__1032_,
  data_stage_1__1031_,data_stage_1__1030_,data_stage_1__1029_,data_stage_1__1028_,
  data_stage_1__1027_,data_stage_1__1026_,data_stage_1__1025_,data_stage_1__1024_,
  data_stage_1__1023_,data_stage_1__1022_,data_stage_1__1021_,data_stage_1__1020_,
  data_stage_1__1019_,data_stage_1__1018_,data_stage_1__1017_,data_stage_1__1016_,
  data_stage_1__1015_,data_stage_1__1014_,data_stage_1__1013_,data_stage_1__1012_,
  data_stage_1__1011_,data_stage_1__1010_,data_stage_1__1009_,data_stage_1__1008_,
  data_stage_1__1007_,data_stage_1__1006_,data_stage_1__1005_,data_stage_1__1004_,
  data_stage_1__1003_,data_stage_1__1002_,data_stage_1__1001_,data_stage_1__1000_,
  data_stage_1__999_,data_stage_1__998_,data_stage_1__997_,data_stage_1__996_,
  data_stage_1__995_,data_stage_1__994_,data_stage_1__993_,data_stage_1__992_,
  data_stage_1__991_,data_stage_1__990_,data_stage_1__989_,data_stage_1__988_,
  data_stage_1__987_,data_stage_1__986_,data_stage_1__985_,data_stage_1__984_,
  data_stage_1__983_,data_stage_1__982_,data_stage_1__981_,data_stage_1__980_,data_stage_1__979_,
  data_stage_1__978_,data_stage_1__977_,data_stage_1__976_,data_stage_1__975_,
  data_stage_1__974_,data_stage_1__973_,data_stage_1__972_,data_stage_1__971_,
  data_stage_1__970_,data_stage_1__969_,data_stage_1__968_,data_stage_1__967_,
  data_stage_1__966_,data_stage_1__965_,data_stage_1__964_,data_stage_1__963_,
  data_stage_1__962_,data_stage_1__961_,data_stage_1__960_,data_stage_1__959_,data_stage_1__958_,
  data_stage_1__957_,data_stage_1__956_,data_stage_1__955_,data_stage_1__954_,
  data_stage_1__953_,data_stage_1__952_,data_stage_1__951_,data_stage_1__950_,
  data_stage_1__949_,data_stage_1__948_,data_stage_1__947_,data_stage_1__946_,
  data_stage_1__945_,data_stage_1__944_,data_stage_1__943_,data_stage_1__942_,
  data_stage_1__941_,data_stage_1__940_,data_stage_1__939_,data_stage_1__938_,data_stage_1__937_,
  data_stage_1__936_,data_stage_1__935_,data_stage_1__934_,data_stage_1__933_,
  data_stage_1__932_,data_stage_1__931_,data_stage_1__930_,data_stage_1__929_,
  data_stage_1__928_,data_stage_1__927_,data_stage_1__926_,data_stage_1__925_,
  data_stage_1__924_,data_stage_1__923_,data_stage_1__922_,data_stage_1__921_,data_stage_1__920_,
  data_stage_1__919_,data_stage_1__918_,data_stage_1__917_,data_stage_1__916_,
  data_stage_1__915_,data_stage_1__914_,data_stage_1__913_,data_stage_1__912_,
  data_stage_1__911_,data_stage_1__910_,data_stage_1__909_,data_stage_1__908_,
  data_stage_1__907_,data_stage_1__906_,data_stage_1__905_,data_stage_1__904_,
  data_stage_1__903_,data_stage_1__902_,data_stage_1__901_,data_stage_1__900_,data_stage_1__899_,
  data_stage_1__898_,data_stage_1__897_,data_stage_1__896_,data_stage_1__895_,
  data_stage_1__894_,data_stage_1__893_,data_stage_1__892_,data_stage_1__891_,
  data_stage_1__890_,data_stage_1__889_,data_stage_1__888_,data_stage_1__887_,
  data_stage_1__886_,data_stage_1__885_,data_stage_1__884_,data_stage_1__883_,
  data_stage_1__882_,data_stage_1__881_,data_stage_1__880_,data_stage_1__879_,data_stage_1__878_,
  data_stage_1__877_,data_stage_1__876_,data_stage_1__875_,data_stage_1__874_,
  data_stage_1__873_,data_stage_1__872_,data_stage_1__871_,data_stage_1__870_,
  data_stage_1__869_,data_stage_1__868_,data_stage_1__867_,data_stage_1__866_,
  data_stage_1__865_,data_stage_1__864_,data_stage_1__863_,data_stage_1__862_,
  data_stage_1__861_,data_stage_1__860_,data_stage_1__859_,data_stage_1__858_,data_stage_1__857_,
  data_stage_1__856_,data_stage_1__855_,data_stage_1__854_,data_stage_1__853_,
  data_stage_1__852_,data_stage_1__851_,data_stage_1__850_,data_stage_1__849_,
  data_stage_1__848_,data_stage_1__847_,data_stage_1__846_,data_stage_1__845_,
  data_stage_1__844_,data_stage_1__843_,data_stage_1__842_,data_stage_1__841_,data_stage_1__840_,
  data_stage_1__839_,data_stage_1__838_,data_stage_1__837_,data_stage_1__836_,
  data_stage_1__835_,data_stage_1__834_,data_stage_1__833_,data_stage_1__832_,
  data_stage_1__831_,data_stage_1__830_,data_stage_1__829_,data_stage_1__828_,
  data_stage_1__827_,data_stage_1__826_,data_stage_1__825_,data_stage_1__824_,
  data_stage_1__823_,data_stage_1__822_,data_stage_1__821_,data_stage_1__820_,data_stage_1__819_,
  data_stage_1__818_,data_stage_1__817_,data_stage_1__816_,data_stage_1__815_,
  data_stage_1__814_,data_stage_1__813_,data_stage_1__812_,data_stage_1__811_,
  data_stage_1__810_,data_stage_1__809_,data_stage_1__808_,data_stage_1__807_,
  data_stage_1__806_,data_stage_1__805_,data_stage_1__804_,data_stage_1__803_,
  data_stage_1__802_,data_stage_1__801_,data_stage_1__800_,data_stage_1__799_,data_stage_1__798_,
  data_stage_1__797_,data_stage_1__796_,data_stage_1__795_,data_stage_1__794_,
  data_stage_1__793_,data_stage_1__792_,data_stage_1__791_,data_stage_1__790_,
  data_stage_1__789_,data_stage_1__788_,data_stage_1__787_,data_stage_1__786_,
  data_stage_1__785_,data_stage_1__784_,data_stage_1__783_,data_stage_1__782_,
  data_stage_1__781_,data_stage_1__780_,data_stage_1__779_,data_stage_1__778_,data_stage_1__777_,
  data_stage_1__776_,data_stage_1__775_,data_stage_1__774_,data_stage_1__773_,
  data_stage_1__772_,data_stage_1__771_,data_stage_1__770_,data_stage_1__769_,
  data_stage_1__768_,data_stage_1__767_,data_stage_1__766_,data_stage_1__765_,
  data_stage_1__764_,data_stage_1__763_,data_stage_1__762_,data_stage_1__761_,data_stage_1__760_,
  data_stage_1__759_,data_stage_1__758_,data_stage_1__757_,data_stage_1__756_,
  data_stage_1__755_,data_stage_1__754_,data_stage_1__753_,data_stage_1__752_,
  data_stage_1__751_,data_stage_1__750_,data_stage_1__749_,data_stage_1__748_,
  data_stage_1__747_,data_stage_1__746_,data_stage_1__745_,data_stage_1__744_,
  data_stage_1__743_,data_stage_1__742_,data_stage_1__741_,data_stage_1__740_,data_stage_1__739_,
  data_stage_1__738_,data_stage_1__737_,data_stage_1__736_,data_stage_1__735_,
  data_stage_1__734_,data_stage_1__733_,data_stage_1__732_,data_stage_1__731_,
  data_stage_1__730_,data_stage_1__729_,data_stage_1__728_,data_stage_1__727_,
  data_stage_1__726_,data_stage_1__725_,data_stage_1__724_,data_stage_1__723_,
  data_stage_1__722_,data_stage_1__721_,data_stage_1__720_,data_stage_1__719_,data_stage_1__718_,
  data_stage_1__717_,data_stage_1__716_,data_stage_1__715_,data_stage_1__714_,
  data_stage_1__713_,data_stage_1__712_,data_stage_1__711_,data_stage_1__710_,
  data_stage_1__709_,data_stage_1__708_,data_stage_1__707_,data_stage_1__706_,
  data_stage_1__705_,data_stage_1__704_,data_stage_1__703_,data_stage_1__702_,
  data_stage_1__701_,data_stage_1__700_,data_stage_1__699_,data_stage_1__698_,data_stage_1__697_,
  data_stage_1__696_,data_stage_1__695_,data_stage_1__694_,data_stage_1__693_,
  data_stage_1__692_,data_stage_1__691_,data_stage_1__690_,data_stage_1__689_,
  data_stage_1__688_,data_stage_1__687_,data_stage_1__686_,data_stage_1__685_,
  data_stage_1__684_,data_stage_1__683_,data_stage_1__682_,data_stage_1__681_,data_stage_1__680_,
  data_stage_1__679_,data_stage_1__678_,data_stage_1__677_,data_stage_1__676_,
  data_stage_1__675_,data_stage_1__674_,data_stage_1__673_,data_stage_1__672_,
  data_stage_1__671_,data_stage_1__670_,data_stage_1__669_,data_stage_1__668_,
  data_stage_1__667_,data_stage_1__666_,data_stage_1__665_,data_stage_1__664_,
  data_stage_1__663_,data_stage_1__662_,data_stage_1__661_,data_stage_1__660_,data_stage_1__659_,
  data_stage_1__658_,data_stage_1__657_,data_stage_1__656_,data_stage_1__655_,
  data_stage_1__654_,data_stage_1__653_,data_stage_1__652_,data_stage_1__651_,
  data_stage_1__650_,data_stage_1__649_,data_stage_1__648_,data_stage_1__647_,
  data_stage_1__646_,data_stage_1__645_,data_stage_1__644_,data_stage_1__643_,
  data_stage_1__642_,data_stage_1__641_,data_stage_1__640_,data_stage_1__639_,data_stage_1__638_,
  data_stage_1__637_,data_stage_1__636_,data_stage_1__635_,data_stage_1__634_,
  data_stage_1__633_,data_stage_1__632_,data_stage_1__631_,data_stage_1__630_,
  data_stage_1__629_,data_stage_1__628_,data_stage_1__627_,data_stage_1__626_,
  data_stage_1__625_,data_stage_1__624_,data_stage_1__623_,data_stage_1__622_,
  data_stage_1__621_,data_stage_1__620_,data_stage_1__619_,data_stage_1__618_,data_stage_1__617_,
  data_stage_1__616_,data_stage_1__615_,data_stage_1__614_,data_stage_1__613_,
  data_stage_1__612_,data_stage_1__611_,data_stage_1__610_,data_stage_1__609_,
  data_stage_1__608_,data_stage_1__607_,data_stage_1__606_,data_stage_1__605_,
  data_stage_1__604_,data_stage_1__603_,data_stage_1__602_,data_stage_1__601_,data_stage_1__600_,
  data_stage_1__599_,data_stage_1__598_,data_stage_1__597_,data_stage_1__596_,
  data_stage_1__595_,data_stage_1__594_,data_stage_1__593_,data_stage_1__592_,
  data_stage_1__591_,data_stage_1__590_,data_stage_1__589_,data_stage_1__588_,
  data_stage_1__587_,data_stage_1__586_,data_stage_1__585_,data_stage_1__584_,
  data_stage_1__583_,data_stage_1__582_,data_stage_1__581_,data_stage_1__580_,data_stage_1__579_,
  data_stage_1__578_,data_stage_1__577_,data_stage_1__576_,data_stage_1__575_,
  data_stage_1__574_,data_stage_1__573_,data_stage_1__572_,data_stage_1__571_,
  data_stage_1__570_,data_stage_1__569_,data_stage_1__568_,data_stage_1__567_,
  data_stage_1__566_,data_stage_1__565_,data_stage_1__564_,data_stage_1__563_,
  data_stage_1__562_,data_stage_1__561_,data_stage_1__560_,data_stage_1__559_,data_stage_1__558_,
  data_stage_1__557_,data_stage_1__556_,data_stage_1__555_,data_stage_1__554_,
  data_stage_1__553_,data_stage_1__552_,data_stage_1__551_,data_stage_1__550_,
  data_stage_1__549_,data_stage_1__548_,data_stage_1__547_,data_stage_1__546_,
  data_stage_1__545_,data_stage_1__544_,data_stage_1__543_,data_stage_1__542_,
  data_stage_1__541_,data_stage_1__540_,data_stage_1__539_,data_stage_1__538_,data_stage_1__537_,
  data_stage_1__536_,data_stage_1__535_,data_stage_1__534_,data_stage_1__533_,
  data_stage_1__532_,data_stage_1__531_,data_stage_1__530_,data_stage_1__529_,
  data_stage_1__528_,data_stage_1__527_,data_stage_1__526_,data_stage_1__525_,
  data_stage_1__524_,data_stage_1__523_,data_stage_1__522_,data_stage_1__521_,data_stage_1__520_,
  data_stage_1__519_,data_stage_1__518_,data_stage_1__517_,data_stage_1__516_,
  data_stage_1__515_,data_stage_1__514_,data_stage_1__513_,data_stage_1__512_,
  data_stage_1__511_,data_stage_1__510_,data_stage_1__509_,data_stage_1__508_,
  data_stage_1__507_,data_stage_1__506_,data_stage_1__505_,data_stage_1__504_,
  data_stage_1__503_,data_stage_1__502_,data_stage_1__501_,data_stage_1__500_,data_stage_1__499_,
  data_stage_1__498_,data_stage_1__497_,data_stage_1__496_,data_stage_1__495_,
  data_stage_1__494_,data_stage_1__493_,data_stage_1__492_,data_stage_1__491_,
  data_stage_1__490_,data_stage_1__489_,data_stage_1__488_,data_stage_1__487_,
  data_stage_1__486_,data_stage_1__485_,data_stage_1__484_,data_stage_1__483_,
  data_stage_1__482_,data_stage_1__481_,data_stage_1__480_,data_stage_1__479_,data_stage_1__478_,
  data_stage_1__477_,data_stage_1__476_,data_stage_1__475_,data_stage_1__474_,
  data_stage_1__473_,data_stage_1__472_,data_stage_1__471_,data_stage_1__470_,
  data_stage_1__469_,data_stage_1__468_,data_stage_1__467_,data_stage_1__466_,
  data_stage_1__465_,data_stage_1__464_,data_stage_1__463_,data_stage_1__462_,
  data_stage_1__461_,data_stage_1__460_,data_stage_1__459_,data_stage_1__458_,data_stage_1__457_,
  data_stage_1__456_,data_stage_1__455_,data_stage_1__454_,data_stage_1__453_,
  data_stage_1__452_,data_stage_1__451_,data_stage_1__450_,data_stage_1__449_,
  data_stage_1__448_,data_stage_1__447_,data_stage_1__446_,data_stage_1__445_,
  data_stage_1__444_,data_stage_1__443_,data_stage_1__442_,data_stage_1__441_,data_stage_1__440_,
  data_stage_1__439_,data_stage_1__438_,data_stage_1__437_,data_stage_1__436_,
  data_stage_1__435_,data_stage_1__434_,data_stage_1__433_,data_stage_1__432_,
  data_stage_1__431_,data_stage_1__430_,data_stage_1__429_,data_stage_1__428_,
  data_stage_1__427_,data_stage_1__426_,data_stage_1__425_,data_stage_1__424_,
  data_stage_1__423_,data_stage_1__422_,data_stage_1__421_,data_stage_1__420_,data_stage_1__419_,
  data_stage_1__418_,data_stage_1__417_,data_stage_1__416_,data_stage_1__415_,
  data_stage_1__414_,data_stage_1__413_,data_stage_1__412_,data_stage_1__411_,
  data_stage_1__410_,data_stage_1__409_,data_stage_1__408_,data_stage_1__407_,
  data_stage_1__406_,data_stage_1__405_,data_stage_1__404_,data_stage_1__403_,
  data_stage_1__402_,data_stage_1__401_,data_stage_1__400_,data_stage_1__399_,data_stage_1__398_,
  data_stage_1__397_,data_stage_1__396_,data_stage_1__395_,data_stage_1__394_,
  data_stage_1__393_,data_stage_1__392_,data_stage_1__391_,data_stage_1__390_,
  data_stage_1__389_,data_stage_1__388_,data_stage_1__387_,data_stage_1__386_,
  data_stage_1__385_,data_stage_1__384_,data_stage_1__383_,data_stage_1__382_,
  data_stage_1__381_,data_stage_1__380_,data_stage_1__379_,data_stage_1__378_,data_stage_1__377_,
  data_stage_1__376_,data_stage_1__375_,data_stage_1__374_,data_stage_1__373_,
  data_stage_1__372_,data_stage_1__371_,data_stage_1__370_,data_stage_1__369_,
  data_stage_1__368_,data_stage_1__367_,data_stage_1__366_,data_stage_1__365_,
  data_stage_1__364_,data_stage_1__363_,data_stage_1__362_,data_stage_1__361_,data_stage_1__360_,
  data_stage_1__359_,data_stage_1__358_,data_stage_1__357_,data_stage_1__356_,
  data_stage_1__355_,data_stage_1__354_,data_stage_1__353_,data_stage_1__352_,
  data_stage_1__351_,data_stage_1__350_,data_stage_1__349_,data_stage_1__348_,
  data_stage_1__347_,data_stage_1__346_,data_stage_1__345_,data_stage_1__344_,
  data_stage_1__343_,data_stage_1__342_,data_stage_1__341_,data_stage_1__340_,data_stage_1__339_,
  data_stage_1__338_,data_stage_1__337_,data_stage_1__336_,data_stage_1__335_,
  data_stage_1__334_,data_stage_1__333_,data_stage_1__332_,data_stage_1__331_,
  data_stage_1__330_,data_stage_1__329_,data_stage_1__328_,data_stage_1__327_,
  data_stage_1__326_,data_stage_1__325_,data_stage_1__324_,data_stage_1__323_,
  data_stage_1__322_,data_stage_1__321_,data_stage_1__320_,data_stage_1__319_,data_stage_1__318_,
  data_stage_1__317_,data_stage_1__316_,data_stage_1__315_,data_stage_1__314_,
  data_stage_1__313_,data_stage_1__312_,data_stage_1__311_,data_stage_1__310_,
  data_stage_1__309_,data_stage_1__308_,data_stage_1__307_,data_stage_1__306_,
  data_stage_1__305_,data_stage_1__304_,data_stage_1__303_,data_stage_1__302_,
  data_stage_1__301_,data_stage_1__300_,data_stage_1__299_,data_stage_1__298_,data_stage_1__297_,
  data_stage_1__296_,data_stage_1__295_,data_stage_1__294_,data_stage_1__293_,
  data_stage_1__292_,data_stage_1__291_,data_stage_1__290_,data_stage_1__289_,
  data_stage_1__288_,data_stage_1__287_,data_stage_1__286_,data_stage_1__285_,
  data_stage_1__284_,data_stage_1__283_,data_stage_1__282_,data_stage_1__281_,data_stage_1__280_,
  data_stage_1__279_,data_stage_1__278_,data_stage_1__277_,data_stage_1__276_,
  data_stage_1__275_,data_stage_1__274_,data_stage_1__273_,data_stage_1__272_,
  data_stage_1__271_,data_stage_1__270_,data_stage_1__269_,data_stage_1__268_,
  data_stage_1__267_,data_stage_1__266_,data_stage_1__265_,data_stage_1__264_,
  data_stage_1__263_,data_stage_1__262_,data_stage_1__261_,data_stage_1__260_,data_stage_1__259_,
  data_stage_1__258_,data_stage_1__257_,data_stage_1__256_,data_stage_1__255_,
  data_stage_1__254_,data_stage_1__253_,data_stage_1__252_,data_stage_1__251_,
  data_stage_1__250_,data_stage_1__249_,data_stage_1__248_,data_stage_1__247_,
  data_stage_1__246_,data_stage_1__245_,data_stage_1__244_,data_stage_1__243_,
  data_stage_1__242_,data_stage_1__241_,data_stage_1__240_,data_stage_1__239_,data_stage_1__238_,
  data_stage_1__237_,data_stage_1__236_,data_stage_1__235_,data_stage_1__234_,
  data_stage_1__233_,data_stage_1__232_,data_stage_1__231_,data_stage_1__230_,
  data_stage_1__229_,data_stage_1__228_,data_stage_1__227_,data_stage_1__226_,
  data_stage_1__225_,data_stage_1__224_,data_stage_1__223_,data_stage_1__222_,
  data_stage_1__221_,data_stage_1__220_,data_stage_1__219_,data_stage_1__218_,data_stage_1__217_,
  data_stage_1__216_,data_stage_1__215_,data_stage_1__214_,data_stage_1__213_,
  data_stage_1__212_,data_stage_1__211_,data_stage_1__210_,data_stage_1__209_,
  data_stage_1__208_,data_stage_1__207_,data_stage_1__206_,data_stage_1__205_,
  data_stage_1__204_,data_stage_1__203_,data_stage_1__202_,data_stage_1__201_,data_stage_1__200_,
  data_stage_1__199_,data_stage_1__198_,data_stage_1__197_,data_stage_1__196_,
  data_stage_1__195_,data_stage_1__194_,data_stage_1__193_,data_stage_1__192_,
  data_stage_1__191_,data_stage_1__190_,data_stage_1__189_,data_stage_1__188_,
  data_stage_1__187_,data_stage_1__186_,data_stage_1__185_,data_stage_1__184_,
  data_stage_1__183_,data_stage_1__182_,data_stage_1__181_,data_stage_1__180_,data_stage_1__179_,
  data_stage_1__178_,data_stage_1__177_,data_stage_1__176_,data_stage_1__175_,
  data_stage_1__174_,data_stage_1__173_,data_stage_1__172_,data_stage_1__171_,
  data_stage_1__170_,data_stage_1__169_,data_stage_1__168_,data_stage_1__167_,
  data_stage_1__166_,data_stage_1__165_,data_stage_1__164_,data_stage_1__163_,
  data_stage_1__162_,data_stage_1__161_,data_stage_1__160_,data_stage_1__159_,data_stage_1__158_,
  data_stage_1__157_,data_stage_1__156_,data_stage_1__155_,data_stage_1__154_,
  data_stage_1__153_,data_stage_1__152_,data_stage_1__151_,data_stage_1__150_,
  data_stage_1__149_,data_stage_1__148_,data_stage_1__147_,data_stage_1__146_,
  data_stage_1__145_,data_stage_1__144_,data_stage_1__143_,data_stage_1__142_,
  data_stage_1__141_,data_stage_1__140_,data_stage_1__139_,data_stage_1__138_,data_stage_1__137_,
  data_stage_1__136_,data_stage_1__135_,data_stage_1__134_,data_stage_1__133_,
  data_stage_1__132_,data_stage_1__131_,data_stage_1__130_,data_stage_1__129_,
  data_stage_1__128_,data_stage_1__127_,data_stage_1__126_,data_stage_1__125_,
  data_stage_1__124_,data_stage_1__123_,data_stage_1__122_,data_stage_1__121_,data_stage_1__120_,
  data_stage_1__119_,data_stage_1__118_,data_stage_1__117_,data_stage_1__116_,
  data_stage_1__115_,data_stage_1__114_,data_stage_1__113_,data_stage_1__112_,
  data_stage_1__111_,data_stage_1__110_,data_stage_1__109_,data_stage_1__108_,
  data_stage_1__107_,data_stage_1__106_,data_stage_1__105_,data_stage_1__104_,
  data_stage_1__103_,data_stage_1__102_,data_stage_1__101_,data_stage_1__100_,data_stage_1__99_,
  data_stage_1__98_,data_stage_1__97_,data_stage_1__96_,data_stage_1__95_,
  data_stage_1__94_,data_stage_1__93_,data_stage_1__92_,data_stage_1__91_,data_stage_1__90_,
  data_stage_1__89_,data_stage_1__88_,data_stage_1__87_,data_stage_1__86_,
  data_stage_1__85_,data_stage_1__84_,data_stage_1__83_,data_stage_1__82_,
  data_stage_1__81_,data_stage_1__80_,data_stage_1__79_,data_stage_1__78_,data_stage_1__77_,
  data_stage_1__76_,data_stage_1__75_,data_stage_1__74_,data_stage_1__73_,
  data_stage_1__72_,data_stage_1__71_,data_stage_1__70_,data_stage_1__69_,data_stage_1__68_,
  data_stage_1__67_,data_stage_1__66_,data_stage_1__65_,data_stage_1__64_,
  data_stage_1__63_,data_stage_1__62_,data_stage_1__61_,data_stage_1__60_,data_stage_1__59_,
  data_stage_1__58_,data_stage_1__57_,data_stage_1__56_,data_stage_1__55_,
  data_stage_1__54_,data_stage_1__53_,data_stage_1__52_,data_stage_1__51_,data_stage_1__50_,
  data_stage_1__49_,data_stage_1__48_,data_stage_1__47_,data_stage_1__46_,
  data_stage_1__45_,data_stage_1__44_,data_stage_1__43_,data_stage_1__42_,
  data_stage_1__41_,data_stage_1__40_,data_stage_1__39_,data_stage_1__38_,data_stage_1__37_,
  data_stage_1__36_,data_stage_1__35_,data_stage_1__34_,data_stage_1__33_,
  data_stage_1__32_,data_stage_1__31_,data_stage_1__30_,data_stage_1__29_,data_stage_1__28_,
  data_stage_1__27_,data_stage_1__26_,data_stage_1__25_,data_stage_1__24_,
  data_stage_1__23_,data_stage_1__22_,data_stage_1__21_,data_stage_1__20_,data_stage_1__19_,
  data_stage_1__18_,data_stage_1__17_,data_stage_1__16_,data_stage_1__15_,
  data_stage_1__14_,data_stage_1__13_,data_stage_1__12_,data_stage_1__11_,data_stage_1__10_,
  data_stage_1__9_,data_stage_1__8_,data_stage_1__7_,data_stage_1__6_,
  data_stage_1__5_,data_stage_1__4_,data_stage_1__3_,data_stage_1__2_,data_stage_1__1_,
  data_stage_1__0_,data_stage_2__4095_,data_stage_2__4094_,data_stage_2__4093_,
  data_stage_2__4092_,data_stage_2__4091_,data_stage_2__4090_,data_stage_2__4089_,
  data_stage_2__4088_,data_stage_2__4087_,data_stage_2__4086_,data_stage_2__4085_,
  data_stage_2__4084_,data_stage_2__4083_,data_stage_2__4082_,data_stage_2__4081_,
  data_stage_2__4080_,data_stage_2__4079_,data_stage_2__4078_,data_stage_2__4077_,
  data_stage_2__4076_,data_stage_2__4075_,data_stage_2__4074_,data_stage_2__4073_,
  data_stage_2__4072_,data_stage_2__4071_,data_stage_2__4070_,data_stage_2__4069_,
  data_stage_2__4068_,data_stage_2__4067_,data_stage_2__4066_,data_stage_2__4065_,
  data_stage_2__4064_,data_stage_2__4063_,data_stage_2__4062_,data_stage_2__4061_,
  data_stage_2__4060_,data_stage_2__4059_,data_stage_2__4058_,data_stage_2__4057_,
  data_stage_2__4056_,data_stage_2__4055_,data_stage_2__4054_,data_stage_2__4053_,
  data_stage_2__4052_,data_stage_2__4051_,data_stage_2__4050_,data_stage_2__4049_,
  data_stage_2__4048_,data_stage_2__4047_,data_stage_2__4046_,data_stage_2__4045_,
  data_stage_2__4044_,data_stage_2__4043_,data_stage_2__4042_,data_stage_2__4041_,
  data_stage_2__4040_,data_stage_2__4039_,data_stage_2__4038_,data_stage_2__4037_,
  data_stage_2__4036_,data_stage_2__4035_,data_stage_2__4034_,data_stage_2__4033_,
  data_stage_2__4032_,data_stage_2__4031_,data_stage_2__4030_,data_stage_2__4029_,
  data_stage_2__4028_,data_stage_2__4027_,data_stage_2__4026_,data_stage_2__4025_,
  data_stage_2__4024_,data_stage_2__4023_,data_stage_2__4022_,data_stage_2__4021_,
  data_stage_2__4020_,data_stage_2__4019_,data_stage_2__4018_,data_stage_2__4017_,
  data_stage_2__4016_,data_stage_2__4015_,data_stage_2__4014_,data_stage_2__4013_,
  data_stage_2__4012_,data_stage_2__4011_,data_stage_2__4010_,data_stage_2__4009_,
  data_stage_2__4008_,data_stage_2__4007_,data_stage_2__4006_,data_stage_2__4005_,
  data_stage_2__4004_,data_stage_2__4003_,data_stage_2__4002_,data_stage_2__4001_,
  data_stage_2__4000_,data_stage_2__3999_,data_stage_2__3998_,data_stage_2__3997_,
  data_stage_2__3996_,data_stage_2__3995_,data_stage_2__3994_,data_stage_2__3993_,
  data_stage_2__3992_,data_stage_2__3991_,data_stage_2__3990_,data_stage_2__3989_,
  data_stage_2__3988_,data_stage_2__3987_,data_stage_2__3986_,data_stage_2__3985_,
  data_stage_2__3984_,data_stage_2__3983_,data_stage_2__3982_,data_stage_2__3981_,
  data_stage_2__3980_,data_stage_2__3979_,data_stage_2__3978_,data_stage_2__3977_,
  data_stage_2__3976_,data_stage_2__3975_,data_stage_2__3974_,data_stage_2__3973_,
  data_stage_2__3972_,data_stage_2__3971_,data_stage_2__3970_,data_stage_2__3969_,
  data_stage_2__3968_,data_stage_2__3967_,data_stage_2__3966_,data_stage_2__3965_,
  data_stage_2__3964_,data_stage_2__3963_,data_stage_2__3962_,data_stage_2__3961_,
  data_stage_2__3960_,data_stage_2__3959_,data_stage_2__3958_,data_stage_2__3957_,
  data_stage_2__3956_,data_stage_2__3955_,data_stage_2__3954_,data_stage_2__3953_,
  data_stage_2__3952_,data_stage_2__3951_,data_stage_2__3950_,data_stage_2__3949_,
  data_stage_2__3948_,data_stage_2__3947_,data_stage_2__3946_,data_stage_2__3945_,
  data_stage_2__3944_,data_stage_2__3943_,data_stage_2__3942_,data_stage_2__3941_,
  data_stage_2__3940_,data_stage_2__3939_,data_stage_2__3938_,data_stage_2__3937_,
  data_stage_2__3936_,data_stage_2__3935_,data_stage_2__3934_,data_stage_2__3933_,
  data_stage_2__3932_,data_stage_2__3931_,data_stage_2__3930_,data_stage_2__3929_,
  data_stage_2__3928_,data_stage_2__3927_,data_stage_2__3926_,data_stage_2__3925_,
  data_stage_2__3924_,data_stage_2__3923_,data_stage_2__3922_,data_stage_2__3921_,
  data_stage_2__3920_,data_stage_2__3919_,data_stage_2__3918_,data_stage_2__3917_,
  data_stage_2__3916_,data_stage_2__3915_,data_stage_2__3914_,data_stage_2__3913_,
  data_stage_2__3912_,data_stage_2__3911_,data_stage_2__3910_,data_stage_2__3909_,
  data_stage_2__3908_,data_stage_2__3907_,data_stage_2__3906_,data_stage_2__3905_,
  data_stage_2__3904_,data_stage_2__3903_,data_stage_2__3902_,data_stage_2__3901_,
  data_stage_2__3900_,data_stage_2__3899_,data_stage_2__3898_,data_stage_2__3897_,
  data_stage_2__3896_,data_stage_2__3895_,data_stage_2__3894_,data_stage_2__3893_,
  data_stage_2__3892_,data_stage_2__3891_,data_stage_2__3890_,data_stage_2__3889_,
  data_stage_2__3888_,data_stage_2__3887_,data_stage_2__3886_,data_stage_2__3885_,
  data_stage_2__3884_,data_stage_2__3883_,data_stage_2__3882_,data_stage_2__3881_,
  data_stage_2__3880_,data_stage_2__3879_,data_stage_2__3878_,data_stage_2__3877_,
  data_stage_2__3876_,data_stage_2__3875_,data_stage_2__3874_,data_stage_2__3873_,
  data_stage_2__3872_,data_stage_2__3871_,data_stage_2__3870_,data_stage_2__3869_,
  data_stage_2__3868_,data_stage_2__3867_,data_stage_2__3866_,data_stage_2__3865_,
  data_stage_2__3864_,data_stage_2__3863_,data_stage_2__3862_,data_stage_2__3861_,
  data_stage_2__3860_,data_stage_2__3859_,data_stage_2__3858_,data_stage_2__3857_,
  data_stage_2__3856_,data_stage_2__3855_,data_stage_2__3854_,data_stage_2__3853_,
  data_stage_2__3852_,data_stage_2__3851_,data_stage_2__3850_,data_stage_2__3849_,
  data_stage_2__3848_,data_stage_2__3847_,data_stage_2__3846_,data_stage_2__3845_,
  data_stage_2__3844_,data_stage_2__3843_,data_stage_2__3842_,data_stage_2__3841_,
  data_stage_2__3840_,data_stage_2__3839_,data_stage_2__3838_,data_stage_2__3837_,
  data_stage_2__3836_,data_stage_2__3835_,data_stage_2__3834_,data_stage_2__3833_,
  data_stage_2__3832_,data_stage_2__3831_,data_stage_2__3830_,data_stage_2__3829_,
  data_stage_2__3828_,data_stage_2__3827_,data_stage_2__3826_,data_stage_2__3825_,
  data_stage_2__3824_,data_stage_2__3823_,data_stage_2__3822_,data_stage_2__3821_,
  data_stage_2__3820_,data_stage_2__3819_,data_stage_2__3818_,data_stage_2__3817_,
  data_stage_2__3816_,data_stage_2__3815_,data_stage_2__3814_,data_stage_2__3813_,
  data_stage_2__3812_,data_stage_2__3811_,data_stage_2__3810_,data_stage_2__3809_,
  data_stage_2__3808_,data_stage_2__3807_,data_stage_2__3806_,data_stage_2__3805_,
  data_stage_2__3804_,data_stage_2__3803_,data_stage_2__3802_,data_stage_2__3801_,
  data_stage_2__3800_,data_stage_2__3799_,data_stage_2__3798_,data_stage_2__3797_,
  data_stage_2__3796_,data_stage_2__3795_,data_stage_2__3794_,data_stage_2__3793_,
  data_stage_2__3792_,data_stage_2__3791_,data_stage_2__3790_,data_stage_2__3789_,
  data_stage_2__3788_,data_stage_2__3787_,data_stage_2__3786_,data_stage_2__3785_,
  data_stage_2__3784_,data_stage_2__3783_,data_stage_2__3782_,data_stage_2__3781_,
  data_stage_2__3780_,data_stage_2__3779_,data_stage_2__3778_,data_stage_2__3777_,
  data_stage_2__3776_,data_stage_2__3775_,data_stage_2__3774_,data_stage_2__3773_,
  data_stage_2__3772_,data_stage_2__3771_,data_stage_2__3770_,data_stage_2__3769_,
  data_stage_2__3768_,data_stage_2__3767_,data_stage_2__3766_,data_stage_2__3765_,
  data_stage_2__3764_,data_stage_2__3763_,data_stage_2__3762_,data_stage_2__3761_,
  data_stage_2__3760_,data_stage_2__3759_,data_stage_2__3758_,data_stage_2__3757_,
  data_stage_2__3756_,data_stage_2__3755_,data_stage_2__3754_,data_stage_2__3753_,
  data_stage_2__3752_,data_stage_2__3751_,data_stage_2__3750_,data_stage_2__3749_,
  data_stage_2__3748_,data_stage_2__3747_,data_stage_2__3746_,data_stage_2__3745_,
  data_stage_2__3744_,data_stage_2__3743_,data_stage_2__3742_,data_stage_2__3741_,
  data_stage_2__3740_,data_stage_2__3739_,data_stage_2__3738_,data_stage_2__3737_,
  data_stage_2__3736_,data_stage_2__3735_,data_stage_2__3734_,data_stage_2__3733_,
  data_stage_2__3732_,data_stage_2__3731_,data_stage_2__3730_,data_stage_2__3729_,
  data_stage_2__3728_,data_stage_2__3727_,data_stage_2__3726_,data_stage_2__3725_,
  data_stage_2__3724_,data_stage_2__3723_,data_stage_2__3722_,data_stage_2__3721_,
  data_stage_2__3720_,data_stage_2__3719_,data_stage_2__3718_,data_stage_2__3717_,
  data_stage_2__3716_,data_stage_2__3715_,data_stage_2__3714_,data_stage_2__3713_,
  data_stage_2__3712_,data_stage_2__3711_,data_stage_2__3710_,data_stage_2__3709_,
  data_stage_2__3708_,data_stage_2__3707_,data_stage_2__3706_,data_stage_2__3705_,
  data_stage_2__3704_,data_stage_2__3703_,data_stage_2__3702_,data_stage_2__3701_,
  data_stage_2__3700_,data_stage_2__3699_,data_stage_2__3698_,data_stage_2__3697_,
  data_stage_2__3696_,data_stage_2__3695_,data_stage_2__3694_,data_stage_2__3693_,
  data_stage_2__3692_,data_stage_2__3691_,data_stage_2__3690_,data_stage_2__3689_,
  data_stage_2__3688_,data_stage_2__3687_,data_stage_2__3686_,data_stage_2__3685_,
  data_stage_2__3684_,data_stage_2__3683_,data_stage_2__3682_,data_stage_2__3681_,
  data_stage_2__3680_,data_stage_2__3679_,data_stage_2__3678_,data_stage_2__3677_,
  data_stage_2__3676_,data_stage_2__3675_,data_stage_2__3674_,data_stage_2__3673_,
  data_stage_2__3672_,data_stage_2__3671_,data_stage_2__3670_,data_stage_2__3669_,
  data_stage_2__3668_,data_stage_2__3667_,data_stage_2__3666_,data_stage_2__3665_,
  data_stage_2__3664_,data_stage_2__3663_,data_stage_2__3662_,data_stage_2__3661_,
  data_stage_2__3660_,data_stage_2__3659_,data_stage_2__3658_,data_stage_2__3657_,
  data_stage_2__3656_,data_stage_2__3655_,data_stage_2__3654_,data_stage_2__3653_,
  data_stage_2__3652_,data_stage_2__3651_,data_stage_2__3650_,data_stage_2__3649_,
  data_stage_2__3648_,data_stage_2__3647_,data_stage_2__3646_,data_stage_2__3645_,
  data_stage_2__3644_,data_stage_2__3643_,data_stage_2__3642_,data_stage_2__3641_,
  data_stage_2__3640_,data_stage_2__3639_,data_stage_2__3638_,data_stage_2__3637_,
  data_stage_2__3636_,data_stage_2__3635_,data_stage_2__3634_,data_stage_2__3633_,
  data_stage_2__3632_,data_stage_2__3631_,data_stage_2__3630_,data_stage_2__3629_,
  data_stage_2__3628_,data_stage_2__3627_,data_stage_2__3626_,data_stage_2__3625_,
  data_stage_2__3624_,data_stage_2__3623_,data_stage_2__3622_,data_stage_2__3621_,
  data_stage_2__3620_,data_stage_2__3619_,data_stage_2__3618_,data_stage_2__3617_,
  data_stage_2__3616_,data_stage_2__3615_,data_stage_2__3614_,data_stage_2__3613_,
  data_stage_2__3612_,data_stage_2__3611_,data_stage_2__3610_,data_stage_2__3609_,
  data_stage_2__3608_,data_stage_2__3607_,data_stage_2__3606_,data_stage_2__3605_,
  data_stage_2__3604_,data_stage_2__3603_,data_stage_2__3602_,data_stage_2__3601_,
  data_stage_2__3600_,data_stage_2__3599_,data_stage_2__3598_,data_stage_2__3597_,
  data_stage_2__3596_,data_stage_2__3595_,data_stage_2__3594_,data_stage_2__3593_,
  data_stage_2__3592_,data_stage_2__3591_,data_stage_2__3590_,data_stage_2__3589_,
  data_stage_2__3588_,data_stage_2__3587_,data_stage_2__3586_,data_stage_2__3585_,
  data_stage_2__3584_,data_stage_2__3583_,data_stage_2__3582_,data_stage_2__3581_,
  data_stage_2__3580_,data_stage_2__3579_,data_stage_2__3578_,data_stage_2__3577_,
  data_stage_2__3576_,data_stage_2__3575_,data_stage_2__3574_,data_stage_2__3573_,
  data_stage_2__3572_,data_stage_2__3571_,data_stage_2__3570_,data_stage_2__3569_,
  data_stage_2__3568_,data_stage_2__3567_,data_stage_2__3566_,data_stage_2__3565_,
  data_stage_2__3564_,data_stage_2__3563_,data_stage_2__3562_,data_stage_2__3561_,
  data_stage_2__3560_,data_stage_2__3559_,data_stage_2__3558_,data_stage_2__3557_,
  data_stage_2__3556_,data_stage_2__3555_,data_stage_2__3554_,data_stage_2__3553_,
  data_stage_2__3552_,data_stage_2__3551_,data_stage_2__3550_,data_stage_2__3549_,
  data_stage_2__3548_,data_stage_2__3547_,data_stage_2__3546_,data_stage_2__3545_,
  data_stage_2__3544_,data_stage_2__3543_,data_stage_2__3542_,data_stage_2__3541_,
  data_stage_2__3540_,data_stage_2__3539_,data_stage_2__3538_,data_stage_2__3537_,
  data_stage_2__3536_,data_stage_2__3535_,data_stage_2__3534_,data_stage_2__3533_,
  data_stage_2__3532_,data_stage_2__3531_,data_stage_2__3530_,data_stage_2__3529_,
  data_stage_2__3528_,data_stage_2__3527_,data_stage_2__3526_,data_stage_2__3525_,
  data_stage_2__3524_,data_stage_2__3523_,data_stage_2__3522_,data_stage_2__3521_,
  data_stage_2__3520_,data_stage_2__3519_,data_stage_2__3518_,data_stage_2__3517_,
  data_stage_2__3516_,data_stage_2__3515_,data_stage_2__3514_,data_stage_2__3513_,
  data_stage_2__3512_,data_stage_2__3511_,data_stage_2__3510_,data_stage_2__3509_,
  data_stage_2__3508_,data_stage_2__3507_,data_stage_2__3506_,data_stage_2__3505_,
  data_stage_2__3504_,data_stage_2__3503_,data_stage_2__3502_,data_stage_2__3501_,
  data_stage_2__3500_,data_stage_2__3499_,data_stage_2__3498_,data_stage_2__3497_,
  data_stage_2__3496_,data_stage_2__3495_,data_stage_2__3494_,data_stage_2__3493_,
  data_stage_2__3492_,data_stage_2__3491_,data_stage_2__3490_,data_stage_2__3489_,
  data_stage_2__3488_,data_stage_2__3487_,data_stage_2__3486_,data_stage_2__3485_,
  data_stage_2__3484_,data_stage_2__3483_,data_stage_2__3482_,data_stage_2__3481_,
  data_stage_2__3480_,data_stage_2__3479_,data_stage_2__3478_,data_stage_2__3477_,
  data_stage_2__3476_,data_stage_2__3475_,data_stage_2__3474_,data_stage_2__3473_,
  data_stage_2__3472_,data_stage_2__3471_,data_stage_2__3470_,data_stage_2__3469_,
  data_stage_2__3468_,data_stage_2__3467_,data_stage_2__3466_,data_stage_2__3465_,
  data_stage_2__3464_,data_stage_2__3463_,data_stage_2__3462_,data_stage_2__3461_,
  data_stage_2__3460_,data_stage_2__3459_,data_stage_2__3458_,data_stage_2__3457_,
  data_stage_2__3456_,data_stage_2__3455_,data_stage_2__3454_,data_stage_2__3453_,
  data_stage_2__3452_,data_stage_2__3451_,data_stage_2__3450_,data_stage_2__3449_,
  data_stage_2__3448_,data_stage_2__3447_,data_stage_2__3446_,data_stage_2__3445_,
  data_stage_2__3444_,data_stage_2__3443_,data_stage_2__3442_,data_stage_2__3441_,
  data_stage_2__3440_,data_stage_2__3439_,data_stage_2__3438_,data_stage_2__3437_,
  data_stage_2__3436_,data_stage_2__3435_,data_stage_2__3434_,data_stage_2__3433_,
  data_stage_2__3432_,data_stage_2__3431_,data_stage_2__3430_,data_stage_2__3429_,
  data_stage_2__3428_,data_stage_2__3427_,data_stage_2__3426_,data_stage_2__3425_,
  data_stage_2__3424_,data_stage_2__3423_,data_stage_2__3422_,data_stage_2__3421_,
  data_stage_2__3420_,data_stage_2__3419_,data_stage_2__3418_,data_stage_2__3417_,
  data_stage_2__3416_,data_stage_2__3415_,data_stage_2__3414_,data_stage_2__3413_,
  data_stage_2__3412_,data_stage_2__3411_,data_stage_2__3410_,data_stage_2__3409_,
  data_stage_2__3408_,data_stage_2__3407_,data_stage_2__3406_,data_stage_2__3405_,
  data_stage_2__3404_,data_stage_2__3403_,data_stage_2__3402_,data_stage_2__3401_,
  data_stage_2__3400_,data_stage_2__3399_,data_stage_2__3398_,data_stage_2__3397_,
  data_stage_2__3396_,data_stage_2__3395_,data_stage_2__3394_,data_stage_2__3393_,
  data_stage_2__3392_,data_stage_2__3391_,data_stage_2__3390_,data_stage_2__3389_,
  data_stage_2__3388_,data_stage_2__3387_,data_stage_2__3386_,data_stage_2__3385_,
  data_stage_2__3384_,data_stage_2__3383_,data_stage_2__3382_,data_stage_2__3381_,
  data_stage_2__3380_,data_stage_2__3379_,data_stage_2__3378_,data_stage_2__3377_,
  data_stage_2__3376_,data_stage_2__3375_,data_stage_2__3374_,data_stage_2__3373_,
  data_stage_2__3372_,data_stage_2__3371_,data_stage_2__3370_,data_stage_2__3369_,
  data_stage_2__3368_,data_stage_2__3367_,data_stage_2__3366_,data_stage_2__3365_,
  data_stage_2__3364_,data_stage_2__3363_,data_stage_2__3362_,data_stage_2__3361_,
  data_stage_2__3360_,data_stage_2__3359_,data_stage_2__3358_,data_stage_2__3357_,
  data_stage_2__3356_,data_stage_2__3355_,data_stage_2__3354_,data_stage_2__3353_,
  data_stage_2__3352_,data_stage_2__3351_,data_stage_2__3350_,data_stage_2__3349_,
  data_stage_2__3348_,data_stage_2__3347_,data_stage_2__3346_,data_stage_2__3345_,
  data_stage_2__3344_,data_stage_2__3343_,data_stage_2__3342_,data_stage_2__3341_,
  data_stage_2__3340_,data_stage_2__3339_,data_stage_2__3338_,data_stage_2__3337_,
  data_stage_2__3336_,data_stage_2__3335_,data_stage_2__3334_,data_stage_2__3333_,
  data_stage_2__3332_,data_stage_2__3331_,data_stage_2__3330_,data_stage_2__3329_,
  data_stage_2__3328_,data_stage_2__3327_,data_stage_2__3326_,data_stage_2__3325_,
  data_stage_2__3324_,data_stage_2__3323_,data_stage_2__3322_,data_stage_2__3321_,
  data_stage_2__3320_,data_stage_2__3319_,data_stage_2__3318_,data_stage_2__3317_,
  data_stage_2__3316_,data_stage_2__3315_,data_stage_2__3314_,data_stage_2__3313_,
  data_stage_2__3312_,data_stage_2__3311_,data_stage_2__3310_,data_stage_2__3309_,
  data_stage_2__3308_,data_stage_2__3307_,data_stage_2__3306_,data_stage_2__3305_,
  data_stage_2__3304_,data_stage_2__3303_,data_stage_2__3302_,data_stage_2__3301_,
  data_stage_2__3300_,data_stage_2__3299_,data_stage_2__3298_,data_stage_2__3297_,
  data_stage_2__3296_,data_stage_2__3295_,data_stage_2__3294_,data_stage_2__3293_,
  data_stage_2__3292_,data_stage_2__3291_,data_stage_2__3290_,data_stage_2__3289_,
  data_stage_2__3288_,data_stage_2__3287_,data_stage_2__3286_,data_stage_2__3285_,
  data_stage_2__3284_,data_stage_2__3283_,data_stage_2__3282_,data_stage_2__3281_,
  data_stage_2__3280_,data_stage_2__3279_,data_stage_2__3278_,data_stage_2__3277_,
  data_stage_2__3276_,data_stage_2__3275_,data_stage_2__3274_,data_stage_2__3273_,
  data_stage_2__3272_,data_stage_2__3271_,data_stage_2__3270_,data_stage_2__3269_,
  data_stage_2__3268_,data_stage_2__3267_,data_stage_2__3266_,data_stage_2__3265_,
  data_stage_2__3264_,data_stage_2__3263_,data_stage_2__3262_,data_stage_2__3261_,
  data_stage_2__3260_,data_stage_2__3259_,data_stage_2__3258_,data_stage_2__3257_,
  data_stage_2__3256_,data_stage_2__3255_,data_stage_2__3254_,data_stage_2__3253_,
  data_stage_2__3252_,data_stage_2__3251_,data_stage_2__3250_,data_stage_2__3249_,
  data_stage_2__3248_,data_stage_2__3247_,data_stage_2__3246_,data_stage_2__3245_,
  data_stage_2__3244_,data_stage_2__3243_,data_stage_2__3242_,data_stage_2__3241_,
  data_stage_2__3240_,data_stage_2__3239_,data_stage_2__3238_,data_stage_2__3237_,
  data_stage_2__3236_,data_stage_2__3235_,data_stage_2__3234_,data_stage_2__3233_,
  data_stage_2__3232_,data_stage_2__3231_,data_stage_2__3230_,data_stage_2__3229_,
  data_stage_2__3228_,data_stage_2__3227_,data_stage_2__3226_,data_stage_2__3225_,
  data_stage_2__3224_,data_stage_2__3223_,data_stage_2__3222_,data_stage_2__3221_,
  data_stage_2__3220_,data_stage_2__3219_,data_stage_2__3218_,data_stage_2__3217_,
  data_stage_2__3216_,data_stage_2__3215_,data_stage_2__3214_,data_stage_2__3213_,
  data_stage_2__3212_,data_stage_2__3211_,data_stage_2__3210_,data_stage_2__3209_,
  data_stage_2__3208_,data_stage_2__3207_,data_stage_2__3206_,data_stage_2__3205_,
  data_stage_2__3204_,data_stage_2__3203_,data_stage_2__3202_,data_stage_2__3201_,
  data_stage_2__3200_,data_stage_2__3199_,data_stage_2__3198_,data_stage_2__3197_,
  data_stage_2__3196_,data_stage_2__3195_,data_stage_2__3194_,data_stage_2__3193_,
  data_stage_2__3192_,data_stage_2__3191_,data_stage_2__3190_,data_stage_2__3189_,
  data_stage_2__3188_,data_stage_2__3187_,data_stage_2__3186_,data_stage_2__3185_,
  data_stage_2__3184_,data_stage_2__3183_,data_stage_2__3182_,data_stage_2__3181_,
  data_stage_2__3180_,data_stage_2__3179_,data_stage_2__3178_,data_stage_2__3177_,
  data_stage_2__3176_,data_stage_2__3175_,data_stage_2__3174_,data_stage_2__3173_,
  data_stage_2__3172_,data_stage_2__3171_,data_stage_2__3170_,data_stage_2__3169_,
  data_stage_2__3168_,data_stage_2__3167_,data_stage_2__3166_,data_stage_2__3165_,
  data_stage_2__3164_,data_stage_2__3163_,data_stage_2__3162_,data_stage_2__3161_,
  data_stage_2__3160_,data_stage_2__3159_,data_stage_2__3158_,data_stage_2__3157_,
  data_stage_2__3156_,data_stage_2__3155_,data_stage_2__3154_,data_stage_2__3153_,
  data_stage_2__3152_,data_stage_2__3151_,data_stage_2__3150_,data_stage_2__3149_,
  data_stage_2__3148_,data_stage_2__3147_,data_stage_2__3146_,data_stage_2__3145_,
  data_stage_2__3144_,data_stage_2__3143_,data_stage_2__3142_,data_stage_2__3141_,
  data_stage_2__3140_,data_stage_2__3139_,data_stage_2__3138_,data_stage_2__3137_,
  data_stage_2__3136_,data_stage_2__3135_,data_stage_2__3134_,data_stage_2__3133_,
  data_stage_2__3132_,data_stage_2__3131_,data_stage_2__3130_,data_stage_2__3129_,
  data_stage_2__3128_,data_stage_2__3127_,data_stage_2__3126_,data_stage_2__3125_,
  data_stage_2__3124_,data_stage_2__3123_,data_stage_2__3122_,data_stage_2__3121_,
  data_stage_2__3120_,data_stage_2__3119_,data_stage_2__3118_,data_stage_2__3117_,
  data_stage_2__3116_,data_stage_2__3115_,data_stage_2__3114_,data_stage_2__3113_,
  data_stage_2__3112_,data_stage_2__3111_,data_stage_2__3110_,data_stage_2__3109_,
  data_stage_2__3108_,data_stage_2__3107_,data_stage_2__3106_,data_stage_2__3105_,
  data_stage_2__3104_,data_stage_2__3103_,data_stage_2__3102_,data_stage_2__3101_,
  data_stage_2__3100_,data_stage_2__3099_,data_stage_2__3098_,data_stage_2__3097_,
  data_stage_2__3096_,data_stage_2__3095_,data_stage_2__3094_,data_stage_2__3093_,
  data_stage_2__3092_,data_stage_2__3091_,data_stage_2__3090_,data_stage_2__3089_,
  data_stage_2__3088_,data_stage_2__3087_,data_stage_2__3086_,data_stage_2__3085_,
  data_stage_2__3084_,data_stage_2__3083_,data_stage_2__3082_,data_stage_2__3081_,
  data_stage_2__3080_,data_stage_2__3079_,data_stage_2__3078_,data_stage_2__3077_,
  data_stage_2__3076_,data_stage_2__3075_,data_stage_2__3074_,data_stage_2__3073_,
  data_stage_2__3072_,data_stage_2__3071_,data_stage_2__3070_,data_stage_2__3069_,
  data_stage_2__3068_,data_stage_2__3067_,data_stage_2__3066_,data_stage_2__3065_,
  data_stage_2__3064_,data_stage_2__3063_,data_stage_2__3062_,data_stage_2__3061_,
  data_stage_2__3060_,data_stage_2__3059_,data_stage_2__3058_,data_stage_2__3057_,
  data_stage_2__3056_,data_stage_2__3055_,data_stage_2__3054_,data_stage_2__3053_,
  data_stage_2__3052_,data_stage_2__3051_,data_stage_2__3050_,data_stage_2__3049_,
  data_stage_2__3048_,data_stage_2__3047_,data_stage_2__3046_,data_stage_2__3045_,
  data_stage_2__3044_,data_stage_2__3043_,data_stage_2__3042_,data_stage_2__3041_,
  data_stage_2__3040_,data_stage_2__3039_,data_stage_2__3038_,data_stage_2__3037_,
  data_stage_2__3036_,data_stage_2__3035_,data_stage_2__3034_,data_stage_2__3033_,
  data_stage_2__3032_,data_stage_2__3031_,data_stage_2__3030_,data_stage_2__3029_,
  data_stage_2__3028_,data_stage_2__3027_,data_stage_2__3026_,data_stage_2__3025_,
  data_stage_2__3024_,data_stage_2__3023_,data_stage_2__3022_,data_stage_2__3021_,
  data_stage_2__3020_,data_stage_2__3019_,data_stage_2__3018_,data_stage_2__3017_,
  data_stage_2__3016_,data_stage_2__3015_,data_stage_2__3014_,data_stage_2__3013_,
  data_stage_2__3012_,data_stage_2__3011_,data_stage_2__3010_,data_stage_2__3009_,
  data_stage_2__3008_,data_stage_2__3007_,data_stage_2__3006_,data_stage_2__3005_,
  data_stage_2__3004_,data_stage_2__3003_,data_stage_2__3002_,data_stage_2__3001_,
  data_stage_2__3000_,data_stage_2__2999_,data_stage_2__2998_,data_stage_2__2997_,
  data_stage_2__2996_,data_stage_2__2995_,data_stage_2__2994_,data_stage_2__2993_,
  data_stage_2__2992_,data_stage_2__2991_,data_stage_2__2990_,data_stage_2__2989_,
  data_stage_2__2988_,data_stage_2__2987_,data_stage_2__2986_,data_stage_2__2985_,
  data_stage_2__2984_,data_stage_2__2983_,data_stage_2__2982_,data_stage_2__2981_,
  data_stage_2__2980_,data_stage_2__2979_,data_stage_2__2978_,data_stage_2__2977_,
  data_stage_2__2976_,data_stage_2__2975_,data_stage_2__2974_,data_stage_2__2973_,
  data_stage_2__2972_,data_stage_2__2971_,data_stage_2__2970_,data_stage_2__2969_,
  data_stage_2__2968_,data_stage_2__2967_,data_stage_2__2966_,data_stage_2__2965_,
  data_stage_2__2964_,data_stage_2__2963_,data_stage_2__2962_,data_stage_2__2961_,
  data_stage_2__2960_,data_stage_2__2959_,data_stage_2__2958_,data_stage_2__2957_,
  data_stage_2__2956_,data_stage_2__2955_,data_stage_2__2954_,data_stage_2__2953_,
  data_stage_2__2952_,data_stage_2__2951_,data_stage_2__2950_,data_stage_2__2949_,
  data_stage_2__2948_,data_stage_2__2947_,data_stage_2__2946_,data_stage_2__2945_,
  data_stage_2__2944_,data_stage_2__2943_,data_stage_2__2942_,data_stage_2__2941_,
  data_stage_2__2940_,data_stage_2__2939_,data_stage_2__2938_,data_stage_2__2937_,
  data_stage_2__2936_,data_stage_2__2935_,data_stage_2__2934_,data_stage_2__2933_,
  data_stage_2__2932_,data_stage_2__2931_,data_stage_2__2930_,data_stage_2__2929_,
  data_stage_2__2928_,data_stage_2__2927_,data_stage_2__2926_,data_stage_2__2925_,
  data_stage_2__2924_,data_stage_2__2923_,data_stage_2__2922_,data_stage_2__2921_,
  data_stage_2__2920_,data_stage_2__2919_,data_stage_2__2918_,data_stage_2__2917_,
  data_stage_2__2916_,data_stage_2__2915_,data_stage_2__2914_,data_stage_2__2913_,
  data_stage_2__2912_,data_stage_2__2911_,data_stage_2__2910_,data_stage_2__2909_,
  data_stage_2__2908_,data_stage_2__2907_,data_stage_2__2906_,data_stage_2__2905_,
  data_stage_2__2904_,data_stage_2__2903_,data_stage_2__2902_,data_stage_2__2901_,
  data_stage_2__2900_,data_stage_2__2899_,data_stage_2__2898_,data_stage_2__2897_,
  data_stage_2__2896_,data_stage_2__2895_,data_stage_2__2894_,data_stage_2__2893_,
  data_stage_2__2892_,data_stage_2__2891_,data_stage_2__2890_,data_stage_2__2889_,
  data_stage_2__2888_,data_stage_2__2887_,data_stage_2__2886_,data_stage_2__2885_,
  data_stage_2__2884_,data_stage_2__2883_,data_stage_2__2882_,data_stage_2__2881_,
  data_stage_2__2880_,data_stage_2__2879_,data_stage_2__2878_,data_stage_2__2877_,
  data_stage_2__2876_,data_stage_2__2875_,data_stage_2__2874_,data_stage_2__2873_,
  data_stage_2__2872_,data_stage_2__2871_,data_stage_2__2870_,data_stage_2__2869_,
  data_stage_2__2868_,data_stage_2__2867_,data_stage_2__2866_,data_stage_2__2865_,
  data_stage_2__2864_,data_stage_2__2863_,data_stage_2__2862_,data_stage_2__2861_,
  data_stage_2__2860_,data_stage_2__2859_,data_stage_2__2858_,data_stage_2__2857_,
  data_stage_2__2856_,data_stage_2__2855_,data_stage_2__2854_,data_stage_2__2853_,
  data_stage_2__2852_,data_stage_2__2851_,data_stage_2__2850_,data_stage_2__2849_,
  data_stage_2__2848_,data_stage_2__2847_,data_stage_2__2846_,data_stage_2__2845_,
  data_stage_2__2844_,data_stage_2__2843_,data_stage_2__2842_,data_stage_2__2841_,
  data_stage_2__2840_,data_stage_2__2839_,data_stage_2__2838_,data_stage_2__2837_,
  data_stage_2__2836_,data_stage_2__2835_,data_stage_2__2834_,data_stage_2__2833_,
  data_stage_2__2832_,data_stage_2__2831_,data_stage_2__2830_,data_stage_2__2829_,
  data_stage_2__2828_,data_stage_2__2827_,data_stage_2__2826_,data_stage_2__2825_,
  data_stage_2__2824_,data_stage_2__2823_,data_stage_2__2822_,data_stage_2__2821_,
  data_stage_2__2820_,data_stage_2__2819_,data_stage_2__2818_,data_stage_2__2817_,
  data_stage_2__2816_,data_stage_2__2815_,data_stage_2__2814_,data_stage_2__2813_,
  data_stage_2__2812_,data_stage_2__2811_,data_stage_2__2810_,data_stage_2__2809_,
  data_stage_2__2808_,data_stage_2__2807_,data_stage_2__2806_,data_stage_2__2805_,
  data_stage_2__2804_,data_stage_2__2803_,data_stage_2__2802_,data_stage_2__2801_,
  data_stage_2__2800_,data_stage_2__2799_,data_stage_2__2798_,data_stage_2__2797_,
  data_stage_2__2796_,data_stage_2__2795_,data_stage_2__2794_,data_stage_2__2793_,
  data_stage_2__2792_,data_stage_2__2791_,data_stage_2__2790_,data_stage_2__2789_,
  data_stage_2__2788_,data_stage_2__2787_,data_stage_2__2786_,data_stage_2__2785_,
  data_stage_2__2784_,data_stage_2__2783_,data_stage_2__2782_,data_stage_2__2781_,
  data_stage_2__2780_,data_stage_2__2779_,data_stage_2__2778_,data_stage_2__2777_,
  data_stage_2__2776_,data_stage_2__2775_,data_stage_2__2774_,data_stage_2__2773_,
  data_stage_2__2772_,data_stage_2__2771_,data_stage_2__2770_,data_stage_2__2769_,
  data_stage_2__2768_,data_stage_2__2767_,data_stage_2__2766_,data_stage_2__2765_,
  data_stage_2__2764_,data_stage_2__2763_,data_stage_2__2762_,data_stage_2__2761_,
  data_stage_2__2760_,data_stage_2__2759_,data_stage_2__2758_,data_stage_2__2757_,
  data_stage_2__2756_,data_stage_2__2755_,data_stage_2__2754_,data_stage_2__2753_,
  data_stage_2__2752_,data_stage_2__2751_,data_stage_2__2750_,data_stage_2__2749_,
  data_stage_2__2748_,data_stage_2__2747_,data_stage_2__2746_,data_stage_2__2745_,
  data_stage_2__2744_,data_stage_2__2743_,data_stage_2__2742_,data_stage_2__2741_,
  data_stage_2__2740_,data_stage_2__2739_,data_stage_2__2738_,data_stage_2__2737_,
  data_stage_2__2736_,data_stage_2__2735_,data_stage_2__2734_,data_stage_2__2733_,
  data_stage_2__2732_,data_stage_2__2731_,data_stage_2__2730_,data_stage_2__2729_,
  data_stage_2__2728_,data_stage_2__2727_,data_stage_2__2726_,data_stage_2__2725_,
  data_stage_2__2724_,data_stage_2__2723_,data_stage_2__2722_,data_stage_2__2721_,
  data_stage_2__2720_,data_stage_2__2719_,data_stage_2__2718_,data_stage_2__2717_,
  data_stage_2__2716_,data_stage_2__2715_,data_stage_2__2714_,data_stage_2__2713_,
  data_stage_2__2712_,data_stage_2__2711_,data_stage_2__2710_,data_stage_2__2709_,
  data_stage_2__2708_,data_stage_2__2707_,data_stage_2__2706_,data_stage_2__2705_,
  data_stage_2__2704_,data_stage_2__2703_,data_stage_2__2702_,data_stage_2__2701_,
  data_stage_2__2700_,data_stage_2__2699_,data_stage_2__2698_,data_stage_2__2697_,
  data_stage_2__2696_,data_stage_2__2695_,data_stage_2__2694_,data_stage_2__2693_,
  data_stage_2__2692_,data_stage_2__2691_,data_stage_2__2690_,data_stage_2__2689_,
  data_stage_2__2688_,data_stage_2__2687_,data_stage_2__2686_,data_stage_2__2685_,
  data_stage_2__2684_,data_stage_2__2683_,data_stage_2__2682_,data_stage_2__2681_,
  data_stage_2__2680_,data_stage_2__2679_,data_stage_2__2678_,data_stage_2__2677_,
  data_stage_2__2676_,data_stage_2__2675_,data_stage_2__2674_,data_stage_2__2673_,
  data_stage_2__2672_,data_stage_2__2671_,data_stage_2__2670_,data_stage_2__2669_,
  data_stage_2__2668_,data_stage_2__2667_,data_stage_2__2666_,data_stage_2__2665_,
  data_stage_2__2664_,data_stage_2__2663_,data_stage_2__2662_,data_stage_2__2661_,
  data_stage_2__2660_,data_stage_2__2659_,data_stage_2__2658_,data_stage_2__2657_,
  data_stage_2__2656_,data_stage_2__2655_,data_stage_2__2654_,data_stage_2__2653_,
  data_stage_2__2652_,data_stage_2__2651_,data_stage_2__2650_,data_stage_2__2649_,
  data_stage_2__2648_,data_stage_2__2647_,data_stage_2__2646_,data_stage_2__2645_,
  data_stage_2__2644_,data_stage_2__2643_,data_stage_2__2642_,data_stage_2__2641_,
  data_stage_2__2640_,data_stage_2__2639_,data_stage_2__2638_,data_stage_2__2637_,
  data_stage_2__2636_,data_stage_2__2635_,data_stage_2__2634_,data_stage_2__2633_,
  data_stage_2__2632_,data_stage_2__2631_,data_stage_2__2630_,data_stage_2__2629_,
  data_stage_2__2628_,data_stage_2__2627_,data_stage_2__2626_,data_stage_2__2625_,
  data_stage_2__2624_,data_stage_2__2623_,data_stage_2__2622_,data_stage_2__2621_,
  data_stage_2__2620_,data_stage_2__2619_,data_stage_2__2618_,data_stage_2__2617_,
  data_stage_2__2616_,data_stage_2__2615_,data_stage_2__2614_,data_stage_2__2613_,
  data_stage_2__2612_,data_stage_2__2611_,data_stage_2__2610_,data_stage_2__2609_,
  data_stage_2__2608_,data_stage_2__2607_,data_stage_2__2606_,data_stage_2__2605_,
  data_stage_2__2604_,data_stage_2__2603_,data_stage_2__2602_,data_stage_2__2601_,
  data_stage_2__2600_,data_stage_2__2599_,data_stage_2__2598_,data_stage_2__2597_,
  data_stage_2__2596_,data_stage_2__2595_,data_stage_2__2594_,data_stage_2__2593_,
  data_stage_2__2592_,data_stage_2__2591_,data_stage_2__2590_,data_stage_2__2589_,
  data_stage_2__2588_,data_stage_2__2587_,data_stage_2__2586_,data_stage_2__2585_,
  data_stage_2__2584_,data_stage_2__2583_,data_stage_2__2582_,data_stage_2__2581_,
  data_stage_2__2580_,data_stage_2__2579_,data_stage_2__2578_,data_stage_2__2577_,
  data_stage_2__2576_,data_stage_2__2575_,data_stage_2__2574_,data_stage_2__2573_,
  data_stage_2__2572_,data_stage_2__2571_,data_stage_2__2570_,data_stage_2__2569_,
  data_stage_2__2568_,data_stage_2__2567_,data_stage_2__2566_,data_stage_2__2565_,
  data_stage_2__2564_,data_stage_2__2563_,data_stage_2__2562_,data_stage_2__2561_,
  data_stage_2__2560_,data_stage_2__2559_,data_stage_2__2558_,data_stage_2__2557_,
  data_stage_2__2556_,data_stage_2__2555_,data_stage_2__2554_,data_stage_2__2553_,
  data_stage_2__2552_,data_stage_2__2551_,data_stage_2__2550_,data_stage_2__2549_,
  data_stage_2__2548_,data_stage_2__2547_,data_stage_2__2546_,data_stage_2__2545_,
  data_stage_2__2544_,data_stage_2__2543_,data_stage_2__2542_,data_stage_2__2541_,
  data_stage_2__2540_,data_stage_2__2539_,data_stage_2__2538_,data_stage_2__2537_,
  data_stage_2__2536_,data_stage_2__2535_,data_stage_2__2534_,data_stage_2__2533_,
  data_stage_2__2532_,data_stage_2__2531_,data_stage_2__2530_,data_stage_2__2529_,
  data_stage_2__2528_,data_stage_2__2527_,data_stage_2__2526_,data_stage_2__2525_,
  data_stage_2__2524_,data_stage_2__2523_,data_stage_2__2522_,data_stage_2__2521_,
  data_stage_2__2520_,data_stage_2__2519_,data_stage_2__2518_,data_stage_2__2517_,
  data_stage_2__2516_,data_stage_2__2515_,data_stage_2__2514_,data_stage_2__2513_,
  data_stage_2__2512_,data_stage_2__2511_,data_stage_2__2510_,data_stage_2__2509_,
  data_stage_2__2508_,data_stage_2__2507_,data_stage_2__2506_,data_stage_2__2505_,
  data_stage_2__2504_,data_stage_2__2503_,data_stage_2__2502_,data_stage_2__2501_,
  data_stage_2__2500_,data_stage_2__2499_,data_stage_2__2498_,data_stage_2__2497_,
  data_stage_2__2496_,data_stage_2__2495_,data_stage_2__2494_,data_stage_2__2493_,
  data_stage_2__2492_,data_stage_2__2491_,data_stage_2__2490_,data_stage_2__2489_,
  data_stage_2__2488_,data_stage_2__2487_,data_stage_2__2486_,data_stage_2__2485_,
  data_stage_2__2484_,data_stage_2__2483_,data_stage_2__2482_,data_stage_2__2481_,
  data_stage_2__2480_,data_stage_2__2479_,data_stage_2__2478_,data_stage_2__2477_,
  data_stage_2__2476_,data_stage_2__2475_,data_stage_2__2474_,data_stage_2__2473_,
  data_stage_2__2472_,data_stage_2__2471_,data_stage_2__2470_,data_stage_2__2469_,
  data_stage_2__2468_,data_stage_2__2467_,data_stage_2__2466_,data_stage_2__2465_,
  data_stage_2__2464_,data_stage_2__2463_,data_stage_2__2462_,data_stage_2__2461_,
  data_stage_2__2460_,data_stage_2__2459_,data_stage_2__2458_,data_stage_2__2457_,
  data_stage_2__2456_,data_stage_2__2455_,data_stage_2__2454_,data_stage_2__2453_,
  data_stage_2__2452_,data_stage_2__2451_,data_stage_2__2450_,data_stage_2__2449_,
  data_stage_2__2448_,data_stage_2__2447_,data_stage_2__2446_,data_stage_2__2445_,
  data_stage_2__2444_,data_stage_2__2443_,data_stage_2__2442_,data_stage_2__2441_,
  data_stage_2__2440_,data_stage_2__2439_,data_stage_2__2438_,data_stage_2__2437_,
  data_stage_2__2436_,data_stage_2__2435_,data_stage_2__2434_,data_stage_2__2433_,
  data_stage_2__2432_,data_stage_2__2431_,data_stage_2__2430_,data_stage_2__2429_,
  data_stage_2__2428_,data_stage_2__2427_,data_stage_2__2426_,data_stage_2__2425_,
  data_stage_2__2424_,data_stage_2__2423_,data_stage_2__2422_,data_stage_2__2421_,
  data_stage_2__2420_,data_stage_2__2419_,data_stage_2__2418_,data_stage_2__2417_,
  data_stage_2__2416_,data_stage_2__2415_,data_stage_2__2414_,data_stage_2__2413_,
  data_stage_2__2412_,data_stage_2__2411_,data_stage_2__2410_,data_stage_2__2409_,
  data_stage_2__2408_,data_stage_2__2407_,data_stage_2__2406_,data_stage_2__2405_,
  data_stage_2__2404_,data_stage_2__2403_,data_stage_2__2402_,data_stage_2__2401_,
  data_stage_2__2400_,data_stage_2__2399_,data_stage_2__2398_,data_stage_2__2397_,
  data_stage_2__2396_,data_stage_2__2395_,data_stage_2__2394_,data_stage_2__2393_,
  data_stage_2__2392_,data_stage_2__2391_,data_stage_2__2390_,data_stage_2__2389_,
  data_stage_2__2388_,data_stage_2__2387_,data_stage_2__2386_,data_stage_2__2385_,
  data_stage_2__2384_,data_stage_2__2383_,data_stage_2__2382_,data_stage_2__2381_,
  data_stage_2__2380_,data_stage_2__2379_,data_stage_2__2378_,data_stage_2__2377_,
  data_stage_2__2376_,data_stage_2__2375_,data_stage_2__2374_,data_stage_2__2373_,
  data_stage_2__2372_,data_stage_2__2371_,data_stage_2__2370_,data_stage_2__2369_,
  data_stage_2__2368_,data_stage_2__2367_,data_stage_2__2366_,data_stage_2__2365_,
  data_stage_2__2364_,data_stage_2__2363_,data_stage_2__2362_,data_stage_2__2361_,
  data_stage_2__2360_,data_stage_2__2359_,data_stage_2__2358_,data_stage_2__2357_,
  data_stage_2__2356_,data_stage_2__2355_,data_stage_2__2354_,data_stage_2__2353_,
  data_stage_2__2352_,data_stage_2__2351_,data_stage_2__2350_,data_stage_2__2349_,
  data_stage_2__2348_,data_stage_2__2347_,data_stage_2__2346_,data_stage_2__2345_,
  data_stage_2__2344_,data_stage_2__2343_,data_stage_2__2342_,data_stage_2__2341_,
  data_stage_2__2340_,data_stage_2__2339_,data_stage_2__2338_,data_stage_2__2337_,
  data_stage_2__2336_,data_stage_2__2335_,data_stage_2__2334_,data_stage_2__2333_,
  data_stage_2__2332_,data_stage_2__2331_,data_stage_2__2330_,data_stage_2__2329_,
  data_stage_2__2328_,data_stage_2__2327_,data_stage_2__2326_,data_stage_2__2325_,
  data_stage_2__2324_,data_stage_2__2323_,data_stage_2__2322_,data_stage_2__2321_,
  data_stage_2__2320_,data_stage_2__2319_,data_stage_2__2318_,data_stage_2__2317_,
  data_stage_2__2316_,data_stage_2__2315_,data_stage_2__2314_,data_stage_2__2313_,
  data_stage_2__2312_,data_stage_2__2311_,data_stage_2__2310_,data_stage_2__2309_,
  data_stage_2__2308_,data_stage_2__2307_,data_stage_2__2306_,data_stage_2__2305_,
  data_stage_2__2304_,data_stage_2__2303_,data_stage_2__2302_,data_stage_2__2301_,
  data_stage_2__2300_,data_stage_2__2299_,data_stage_2__2298_,data_stage_2__2297_,
  data_stage_2__2296_,data_stage_2__2295_,data_stage_2__2294_,data_stage_2__2293_,
  data_stage_2__2292_,data_stage_2__2291_,data_stage_2__2290_,data_stage_2__2289_,
  data_stage_2__2288_,data_stage_2__2287_,data_stage_2__2286_,data_stage_2__2285_,
  data_stage_2__2284_,data_stage_2__2283_,data_stage_2__2282_,data_stage_2__2281_,
  data_stage_2__2280_,data_stage_2__2279_,data_stage_2__2278_,data_stage_2__2277_,
  data_stage_2__2276_,data_stage_2__2275_,data_stage_2__2274_,data_stage_2__2273_,
  data_stage_2__2272_,data_stage_2__2271_,data_stage_2__2270_,data_stage_2__2269_,
  data_stage_2__2268_,data_stage_2__2267_,data_stage_2__2266_,data_stage_2__2265_,
  data_stage_2__2264_,data_stage_2__2263_,data_stage_2__2262_,data_stage_2__2261_,
  data_stage_2__2260_,data_stage_2__2259_,data_stage_2__2258_,data_stage_2__2257_,
  data_stage_2__2256_,data_stage_2__2255_,data_stage_2__2254_,data_stage_2__2253_,
  data_stage_2__2252_,data_stage_2__2251_,data_stage_2__2250_,data_stage_2__2249_,
  data_stage_2__2248_,data_stage_2__2247_,data_stage_2__2246_,data_stage_2__2245_,
  data_stage_2__2244_,data_stage_2__2243_,data_stage_2__2242_,data_stage_2__2241_,
  data_stage_2__2240_,data_stage_2__2239_,data_stage_2__2238_,data_stage_2__2237_,
  data_stage_2__2236_,data_stage_2__2235_,data_stage_2__2234_,data_stage_2__2233_,
  data_stage_2__2232_,data_stage_2__2231_,data_stage_2__2230_,data_stage_2__2229_,
  data_stage_2__2228_,data_stage_2__2227_,data_stage_2__2226_,data_stage_2__2225_,
  data_stage_2__2224_,data_stage_2__2223_,data_stage_2__2222_,data_stage_2__2221_,
  data_stage_2__2220_,data_stage_2__2219_,data_stage_2__2218_,data_stage_2__2217_,
  data_stage_2__2216_,data_stage_2__2215_,data_stage_2__2214_,data_stage_2__2213_,
  data_stage_2__2212_,data_stage_2__2211_,data_stage_2__2210_,data_stage_2__2209_,
  data_stage_2__2208_,data_stage_2__2207_,data_stage_2__2206_,data_stage_2__2205_,
  data_stage_2__2204_,data_stage_2__2203_,data_stage_2__2202_,data_stage_2__2201_,
  data_stage_2__2200_,data_stage_2__2199_,data_stage_2__2198_,data_stage_2__2197_,
  data_stage_2__2196_,data_stage_2__2195_,data_stage_2__2194_,data_stage_2__2193_,
  data_stage_2__2192_,data_stage_2__2191_,data_stage_2__2190_,data_stage_2__2189_,
  data_stage_2__2188_,data_stage_2__2187_,data_stage_2__2186_,data_stage_2__2185_,
  data_stage_2__2184_,data_stage_2__2183_,data_stage_2__2182_,data_stage_2__2181_,
  data_stage_2__2180_,data_stage_2__2179_,data_stage_2__2178_,data_stage_2__2177_,
  data_stage_2__2176_,data_stage_2__2175_,data_stage_2__2174_,data_stage_2__2173_,
  data_stage_2__2172_,data_stage_2__2171_,data_stage_2__2170_,data_stage_2__2169_,
  data_stage_2__2168_,data_stage_2__2167_,data_stage_2__2166_,data_stage_2__2165_,
  data_stage_2__2164_,data_stage_2__2163_,data_stage_2__2162_,data_stage_2__2161_,
  data_stage_2__2160_,data_stage_2__2159_,data_stage_2__2158_,data_stage_2__2157_,
  data_stage_2__2156_,data_stage_2__2155_,data_stage_2__2154_,data_stage_2__2153_,
  data_stage_2__2152_,data_stage_2__2151_,data_stage_2__2150_,data_stage_2__2149_,
  data_stage_2__2148_,data_stage_2__2147_,data_stage_2__2146_,data_stage_2__2145_,
  data_stage_2__2144_,data_stage_2__2143_,data_stage_2__2142_,data_stage_2__2141_,
  data_stage_2__2140_,data_stage_2__2139_,data_stage_2__2138_,data_stage_2__2137_,
  data_stage_2__2136_,data_stage_2__2135_,data_stage_2__2134_,data_stage_2__2133_,
  data_stage_2__2132_,data_stage_2__2131_,data_stage_2__2130_,data_stage_2__2129_,
  data_stage_2__2128_,data_stage_2__2127_,data_stage_2__2126_,data_stage_2__2125_,
  data_stage_2__2124_,data_stage_2__2123_,data_stage_2__2122_,data_stage_2__2121_,
  data_stage_2__2120_,data_stage_2__2119_,data_stage_2__2118_,data_stage_2__2117_,
  data_stage_2__2116_,data_stage_2__2115_,data_stage_2__2114_,data_stage_2__2113_,
  data_stage_2__2112_,data_stage_2__2111_,data_stage_2__2110_,data_stage_2__2109_,
  data_stage_2__2108_,data_stage_2__2107_,data_stage_2__2106_,data_stage_2__2105_,
  data_stage_2__2104_,data_stage_2__2103_,data_stage_2__2102_,data_stage_2__2101_,
  data_stage_2__2100_,data_stage_2__2099_,data_stage_2__2098_,data_stage_2__2097_,
  data_stage_2__2096_,data_stage_2__2095_,data_stage_2__2094_,data_stage_2__2093_,
  data_stage_2__2092_,data_stage_2__2091_,data_stage_2__2090_,data_stage_2__2089_,
  data_stage_2__2088_,data_stage_2__2087_,data_stage_2__2086_,data_stage_2__2085_,
  data_stage_2__2084_,data_stage_2__2083_,data_stage_2__2082_,data_stage_2__2081_,
  data_stage_2__2080_,data_stage_2__2079_,data_stage_2__2078_,data_stage_2__2077_,
  data_stage_2__2076_,data_stage_2__2075_,data_stage_2__2074_,data_stage_2__2073_,
  data_stage_2__2072_,data_stage_2__2071_,data_stage_2__2070_,data_stage_2__2069_,
  data_stage_2__2068_,data_stage_2__2067_,data_stage_2__2066_,data_stage_2__2065_,
  data_stage_2__2064_,data_stage_2__2063_,data_stage_2__2062_,data_stage_2__2061_,
  data_stage_2__2060_,data_stage_2__2059_,data_stage_2__2058_,data_stage_2__2057_,
  data_stage_2__2056_,data_stage_2__2055_,data_stage_2__2054_,data_stage_2__2053_,
  data_stage_2__2052_,data_stage_2__2051_,data_stage_2__2050_,data_stage_2__2049_,
  data_stage_2__2048_,data_stage_2__2047_,data_stage_2__2046_,data_stage_2__2045_,
  data_stage_2__2044_,data_stage_2__2043_,data_stage_2__2042_,data_stage_2__2041_,
  data_stage_2__2040_,data_stage_2__2039_,data_stage_2__2038_,data_stage_2__2037_,
  data_stage_2__2036_,data_stage_2__2035_,data_stage_2__2034_,data_stage_2__2033_,
  data_stage_2__2032_,data_stage_2__2031_,data_stage_2__2030_,data_stage_2__2029_,
  data_stage_2__2028_,data_stage_2__2027_,data_stage_2__2026_,data_stage_2__2025_,
  data_stage_2__2024_,data_stage_2__2023_,data_stage_2__2022_,data_stage_2__2021_,
  data_stage_2__2020_,data_stage_2__2019_,data_stage_2__2018_,data_stage_2__2017_,
  data_stage_2__2016_,data_stage_2__2015_,data_stage_2__2014_,data_stage_2__2013_,
  data_stage_2__2012_,data_stage_2__2011_,data_stage_2__2010_,data_stage_2__2009_,
  data_stage_2__2008_,data_stage_2__2007_,data_stage_2__2006_,data_stage_2__2005_,
  data_stage_2__2004_,data_stage_2__2003_,data_stage_2__2002_,data_stage_2__2001_,
  data_stage_2__2000_,data_stage_2__1999_,data_stage_2__1998_,data_stage_2__1997_,
  data_stage_2__1996_,data_stage_2__1995_,data_stage_2__1994_,data_stage_2__1993_,
  data_stage_2__1992_,data_stage_2__1991_,data_stage_2__1990_,data_stage_2__1989_,
  data_stage_2__1988_,data_stage_2__1987_,data_stage_2__1986_,data_stage_2__1985_,
  data_stage_2__1984_,data_stage_2__1983_,data_stage_2__1982_,data_stage_2__1981_,
  data_stage_2__1980_,data_stage_2__1979_,data_stage_2__1978_,data_stage_2__1977_,
  data_stage_2__1976_,data_stage_2__1975_,data_stage_2__1974_,data_stage_2__1973_,
  data_stage_2__1972_,data_stage_2__1971_,data_stage_2__1970_,data_stage_2__1969_,
  data_stage_2__1968_,data_stage_2__1967_,data_stage_2__1966_,data_stage_2__1965_,
  data_stage_2__1964_,data_stage_2__1963_,data_stage_2__1962_,data_stage_2__1961_,
  data_stage_2__1960_,data_stage_2__1959_,data_stage_2__1958_,data_stage_2__1957_,
  data_stage_2__1956_,data_stage_2__1955_,data_stage_2__1954_,data_stage_2__1953_,
  data_stage_2__1952_,data_stage_2__1951_,data_stage_2__1950_,data_stage_2__1949_,
  data_stage_2__1948_,data_stage_2__1947_,data_stage_2__1946_,data_stage_2__1945_,
  data_stage_2__1944_,data_stage_2__1943_,data_stage_2__1942_,data_stage_2__1941_,
  data_stage_2__1940_,data_stage_2__1939_,data_stage_2__1938_,data_stage_2__1937_,
  data_stage_2__1936_,data_stage_2__1935_,data_stage_2__1934_,data_stage_2__1933_,
  data_stage_2__1932_,data_stage_2__1931_,data_stage_2__1930_,data_stage_2__1929_,
  data_stage_2__1928_,data_stage_2__1927_,data_stage_2__1926_,data_stage_2__1925_,
  data_stage_2__1924_,data_stage_2__1923_,data_stage_2__1922_,data_stage_2__1921_,
  data_stage_2__1920_,data_stage_2__1919_,data_stage_2__1918_,data_stage_2__1917_,
  data_stage_2__1916_,data_stage_2__1915_,data_stage_2__1914_,data_stage_2__1913_,
  data_stage_2__1912_,data_stage_2__1911_,data_stage_2__1910_,data_stage_2__1909_,
  data_stage_2__1908_,data_stage_2__1907_,data_stage_2__1906_,data_stage_2__1905_,
  data_stage_2__1904_,data_stage_2__1903_,data_stage_2__1902_,data_stage_2__1901_,
  data_stage_2__1900_,data_stage_2__1899_,data_stage_2__1898_,data_stage_2__1897_,
  data_stage_2__1896_,data_stage_2__1895_,data_stage_2__1894_,data_stage_2__1893_,
  data_stage_2__1892_,data_stage_2__1891_,data_stage_2__1890_,data_stage_2__1889_,
  data_stage_2__1888_,data_stage_2__1887_,data_stage_2__1886_,data_stage_2__1885_,
  data_stage_2__1884_,data_stage_2__1883_,data_stage_2__1882_,data_stage_2__1881_,
  data_stage_2__1880_,data_stage_2__1879_,data_stage_2__1878_,data_stage_2__1877_,
  data_stage_2__1876_,data_stage_2__1875_,data_stage_2__1874_,data_stage_2__1873_,
  data_stage_2__1872_,data_stage_2__1871_,data_stage_2__1870_,data_stage_2__1869_,
  data_stage_2__1868_,data_stage_2__1867_,data_stage_2__1866_,data_stage_2__1865_,
  data_stage_2__1864_,data_stage_2__1863_,data_stage_2__1862_,data_stage_2__1861_,
  data_stage_2__1860_,data_stage_2__1859_,data_stage_2__1858_,data_stage_2__1857_,
  data_stage_2__1856_,data_stage_2__1855_,data_stage_2__1854_,data_stage_2__1853_,
  data_stage_2__1852_,data_stage_2__1851_,data_stage_2__1850_,data_stage_2__1849_,
  data_stage_2__1848_,data_stage_2__1847_,data_stage_2__1846_,data_stage_2__1845_,
  data_stage_2__1844_,data_stage_2__1843_,data_stage_2__1842_,data_stage_2__1841_,
  data_stage_2__1840_,data_stage_2__1839_,data_stage_2__1838_,data_stage_2__1837_,
  data_stage_2__1836_,data_stage_2__1835_,data_stage_2__1834_,data_stage_2__1833_,
  data_stage_2__1832_,data_stage_2__1831_,data_stage_2__1830_,data_stage_2__1829_,
  data_stage_2__1828_,data_stage_2__1827_,data_stage_2__1826_,data_stage_2__1825_,
  data_stage_2__1824_,data_stage_2__1823_,data_stage_2__1822_,data_stage_2__1821_,
  data_stage_2__1820_,data_stage_2__1819_,data_stage_2__1818_,data_stage_2__1817_,
  data_stage_2__1816_,data_stage_2__1815_,data_stage_2__1814_,data_stage_2__1813_,
  data_stage_2__1812_,data_stage_2__1811_,data_stage_2__1810_,data_stage_2__1809_,
  data_stage_2__1808_,data_stage_2__1807_,data_stage_2__1806_,data_stage_2__1805_,
  data_stage_2__1804_,data_stage_2__1803_,data_stage_2__1802_,data_stage_2__1801_,
  data_stage_2__1800_,data_stage_2__1799_,data_stage_2__1798_,data_stage_2__1797_,
  data_stage_2__1796_,data_stage_2__1795_,data_stage_2__1794_,data_stage_2__1793_,
  data_stage_2__1792_,data_stage_2__1791_,data_stage_2__1790_,data_stage_2__1789_,
  data_stage_2__1788_,data_stage_2__1787_,data_stage_2__1786_,data_stage_2__1785_,
  data_stage_2__1784_,data_stage_2__1783_,data_stage_2__1782_,data_stage_2__1781_,
  data_stage_2__1780_,data_stage_2__1779_,data_stage_2__1778_,data_stage_2__1777_,
  data_stage_2__1776_,data_stage_2__1775_,data_stage_2__1774_,data_stage_2__1773_,
  data_stage_2__1772_,data_stage_2__1771_,data_stage_2__1770_,data_stage_2__1769_,
  data_stage_2__1768_,data_stage_2__1767_,data_stage_2__1766_,data_stage_2__1765_,
  data_stage_2__1764_,data_stage_2__1763_,data_stage_2__1762_,data_stage_2__1761_,
  data_stage_2__1760_,data_stage_2__1759_,data_stage_2__1758_,data_stage_2__1757_,
  data_stage_2__1756_,data_stage_2__1755_,data_stage_2__1754_,data_stage_2__1753_,
  data_stage_2__1752_,data_stage_2__1751_,data_stage_2__1750_,data_stage_2__1749_,
  data_stage_2__1748_,data_stage_2__1747_,data_stage_2__1746_,data_stage_2__1745_,
  data_stage_2__1744_,data_stage_2__1743_,data_stage_2__1742_,data_stage_2__1741_,
  data_stage_2__1740_,data_stage_2__1739_,data_stage_2__1738_,data_stage_2__1737_,
  data_stage_2__1736_,data_stage_2__1735_,data_stage_2__1734_,data_stage_2__1733_,
  data_stage_2__1732_,data_stage_2__1731_,data_stage_2__1730_,data_stage_2__1729_,
  data_stage_2__1728_,data_stage_2__1727_,data_stage_2__1726_,data_stage_2__1725_,
  data_stage_2__1724_,data_stage_2__1723_,data_stage_2__1722_,data_stage_2__1721_,
  data_stage_2__1720_,data_stage_2__1719_,data_stage_2__1718_,data_stage_2__1717_,
  data_stage_2__1716_,data_stage_2__1715_,data_stage_2__1714_,data_stage_2__1713_,
  data_stage_2__1712_,data_stage_2__1711_,data_stage_2__1710_,data_stage_2__1709_,
  data_stage_2__1708_,data_stage_2__1707_,data_stage_2__1706_,data_stage_2__1705_,
  data_stage_2__1704_,data_stage_2__1703_,data_stage_2__1702_,data_stage_2__1701_,
  data_stage_2__1700_,data_stage_2__1699_,data_stage_2__1698_,data_stage_2__1697_,
  data_stage_2__1696_,data_stage_2__1695_,data_stage_2__1694_,data_stage_2__1693_,
  data_stage_2__1692_,data_stage_2__1691_,data_stage_2__1690_,data_stage_2__1689_,
  data_stage_2__1688_,data_stage_2__1687_,data_stage_2__1686_,data_stage_2__1685_,
  data_stage_2__1684_,data_stage_2__1683_,data_stage_2__1682_,data_stage_2__1681_,
  data_stage_2__1680_,data_stage_2__1679_,data_stage_2__1678_,data_stage_2__1677_,
  data_stage_2__1676_,data_stage_2__1675_,data_stage_2__1674_,data_stage_2__1673_,
  data_stage_2__1672_,data_stage_2__1671_,data_stage_2__1670_,data_stage_2__1669_,
  data_stage_2__1668_,data_stage_2__1667_,data_stage_2__1666_,data_stage_2__1665_,
  data_stage_2__1664_,data_stage_2__1663_,data_stage_2__1662_,data_stage_2__1661_,
  data_stage_2__1660_,data_stage_2__1659_,data_stage_2__1658_,data_stage_2__1657_,
  data_stage_2__1656_,data_stage_2__1655_,data_stage_2__1654_,data_stage_2__1653_,
  data_stage_2__1652_,data_stage_2__1651_,data_stage_2__1650_,data_stage_2__1649_,
  data_stage_2__1648_,data_stage_2__1647_,data_stage_2__1646_,data_stage_2__1645_,
  data_stage_2__1644_,data_stage_2__1643_,data_stage_2__1642_,data_stage_2__1641_,
  data_stage_2__1640_,data_stage_2__1639_,data_stage_2__1638_,data_stage_2__1637_,
  data_stage_2__1636_,data_stage_2__1635_,data_stage_2__1634_,data_stage_2__1633_,
  data_stage_2__1632_,data_stage_2__1631_,data_stage_2__1630_,data_stage_2__1629_,
  data_stage_2__1628_,data_stage_2__1627_,data_stage_2__1626_,data_stage_2__1625_,
  data_stage_2__1624_,data_stage_2__1623_,data_stage_2__1622_,data_stage_2__1621_,
  data_stage_2__1620_,data_stage_2__1619_,data_stage_2__1618_,data_stage_2__1617_,
  data_stage_2__1616_,data_stage_2__1615_,data_stage_2__1614_,data_stage_2__1613_,
  data_stage_2__1612_,data_stage_2__1611_,data_stage_2__1610_,data_stage_2__1609_,
  data_stage_2__1608_,data_stage_2__1607_,data_stage_2__1606_,data_stage_2__1605_,
  data_stage_2__1604_,data_stage_2__1603_,data_stage_2__1602_,data_stage_2__1601_,
  data_stage_2__1600_,data_stage_2__1599_,data_stage_2__1598_,data_stage_2__1597_,
  data_stage_2__1596_,data_stage_2__1595_,data_stage_2__1594_,data_stage_2__1593_,
  data_stage_2__1592_,data_stage_2__1591_,data_stage_2__1590_,data_stage_2__1589_,
  data_stage_2__1588_,data_stage_2__1587_,data_stage_2__1586_,data_stage_2__1585_,
  data_stage_2__1584_,data_stage_2__1583_,data_stage_2__1582_,data_stage_2__1581_,
  data_stage_2__1580_,data_stage_2__1579_,data_stage_2__1578_,data_stage_2__1577_,
  data_stage_2__1576_,data_stage_2__1575_,data_stage_2__1574_,data_stage_2__1573_,
  data_stage_2__1572_,data_stage_2__1571_,data_stage_2__1570_,data_stage_2__1569_,
  data_stage_2__1568_,data_stage_2__1567_,data_stage_2__1566_,data_stage_2__1565_,
  data_stage_2__1564_,data_stage_2__1563_,data_stage_2__1562_,data_stage_2__1561_,
  data_stage_2__1560_,data_stage_2__1559_,data_stage_2__1558_,data_stage_2__1557_,
  data_stage_2__1556_,data_stage_2__1555_,data_stage_2__1554_,data_stage_2__1553_,
  data_stage_2__1552_,data_stage_2__1551_,data_stage_2__1550_,data_stage_2__1549_,
  data_stage_2__1548_,data_stage_2__1547_,data_stage_2__1546_,data_stage_2__1545_,
  data_stage_2__1544_,data_stage_2__1543_,data_stage_2__1542_,data_stage_2__1541_,
  data_stage_2__1540_,data_stage_2__1539_,data_stage_2__1538_,data_stage_2__1537_,
  data_stage_2__1536_,data_stage_2__1535_,data_stage_2__1534_,data_stage_2__1533_,
  data_stage_2__1532_,data_stage_2__1531_,data_stage_2__1530_,data_stage_2__1529_,
  data_stage_2__1528_,data_stage_2__1527_,data_stage_2__1526_,data_stage_2__1525_,
  data_stage_2__1524_,data_stage_2__1523_,data_stage_2__1522_,data_stage_2__1521_,
  data_stage_2__1520_,data_stage_2__1519_,data_stage_2__1518_,data_stage_2__1517_,
  data_stage_2__1516_,data_stage_2__1515_,data_stage_2__1514_,data_stage_2__1513_,
  data_stage_2__1512_,data_stage_2__1511_,data_stage_2__1510_,data_stage_2__1509_,
  data_stage_2__1508_,data_stage_2__1507_,data_stage_2__1506_,data_stage_2__1505_,
  data_stage_2__1504_,data_stage_2__1503_,data_stage_2__1502_,data_stage_2__1501_,
  data_stage_2__1500_,data_stage_2__1499_,data_stage_2__1498_,data_stage_2__1497_,
  data_stage_2__1496_,data_stage_2__1495_,data_stage_2__1494_,data_stage_2__1493_,
  data_stage_2__1492_,data_stage_2__1491_,data_stage_2__1490_,data_stage_2__1489_,
  data_stage_2__1488_,data_stage_2__1487_,data_stage_2__1486_,data_stage_2__1485_,
  data_stage_2__1484_,data_stage_2__1483_,data_stage_2__1482_,data_stage_2__1481_,
  data_stage_2__1480_,data_stage_2__1479_,data_stage_2__1478_,data_stage_2__1477_,
  data_stage_2__1476_,data_stage_2__1475_,data_stage_2__1474_,data_stage_2__1473_,
  data_stage_2__1472_,data_stage_2__1471_,data_stage_2__1470_,data_stage_2__1469_,
  data_stage_2__1468_,data_stage_2__1467_,data_stage_2__1466_,data_stage_2__1465_,
  data_stage_2__1464_,data_stage_2__1463_,data_stage_2__1462_,data_stage_2__1461_,
  data_stage_2__1460_,data_stage_2__1459_,data_stage_2__1458_,data_stage_2__1457_,
  data_stage_2__1456_,data_stage_2__1455_,data_stage_2__1454_,data_stage_2__1453_,
  data_stage_2__1452_,data_stage_2__1451_,data_stage_2__1450_,data_stage_2__1449_,
  data_stage_2__1448_,data_stage_2__1447_,data_stage_2__1446_,data_stage_2__1445_,
  data_stage_2__1444_,data_stage_2__1443_,data_stage_2__1442_,data_stage_2__1441_,
  data_stage_2__1440_,data_stage_2__1439_,data_stage_2__1438_,data_stage_2__1437_,
  data_stage_2__1436_,data_stage_2__1435_,data_stage_2__1434_,data_stage_2__1433_,
  data_stage_2__1432_,data_stage_2__1431_,data_stage_2__1430_,data_stage_2__1429_,
  data_stage_2__1428_,data_stage_2__1427_,data_stage_2__1426_,data_stage_2__1425_,
  data_stage_2__1424_,data_stage_2__1423_,data_stage_2__1422_,data_stage_2__1421_,
  data_stage_2__1420_,data_stage_2__1419_,data_stage_2__1418_,data_stage_2__1417_,
  data_stage_2__1416_,data_stage_2__1415_,data_stage_2__1414_,data_stage_2__1413_,
  data_stage_2__1412_,data_stage_2__1411_,data_stage_2__1410_,data_stage_2__1409_,
  data_stage_2__1408_,data_stage_2__1407_,data_stage_2__1406_,data_stage_2__1405_,
  data_stage_2__1404_,data_stage_2__1403_,data_stage_2__1402_,data_stage_2__1401_,
  data_stage_2__1400_,data_stage_2__1399_,data_stage_2__1398_,data_stage_2__1397_,
  data_stage_2__1396_,data_stage_2__1395_,data_stage_2__1394_,data_stage_2__1393_,
  data_stage_2__1392_,data_stage_2__1391_,data_stage_2__1390_,data_stage_2__1389_,
  data_stage_2__1388_,data_stage_2__1387_,data_stage_2__1386_,data_stage_2__1385_,
  data_stage_2__1384_,data_stage_2__1383_,data_stage_2__1382_,data_stage_2__1381_,
  data_stage_2__1380_,data_stage_2__1379_,data_stage_2__1378_,data_stage_2__1377_,
  data_stage_2__1376_,data_stage_2__1375_,data_stage_2__1374_,data_stage_2__1373_,
  data_stage_2__1372_,data_stage_2__1371_,data_stage_2__1370_,data_stage_2__1369_,
  data_stage_2__1368_,data_stage_2__1367_,data_stage_2__1366_,data_stage_2__1365_,
  data_stage_2__1364_,data_stage_2__1363_,data_stage_2__1362_,data_stage_2__1361_,
  data_stage_2__1360_,data_stage_2__1359_,data_stage_2__1358_,data_stage_2__1357_,
  data_stage_2__1356_,data_stage_2__1355_,data_stage_2__1354_,data_stage_2__1353_,
  data_stage_2__1352_,data_stage_2__1351_,data_stage_2__1350_,data_stage_2__1349_,
  data_stage_2__1348_,data_stage_2__1347_,data_stage_2__1346_,data_stage_2__1345_,
  data_stage_2__1344_,data_stage_2__1343_,data_stage_2__1342_,data_stage_2__1341_,
  data_stage_2__1340_,data_stage_2__1339_,data_stage_2__1338_,data_stage_2__1337_,
  data_stage_2__1336_,data_stage_2__1335_,data_stage_2__1334_,data_stage_2__1333_,
  data_stage_2__1332_,data_stage_2__1331_,data_stage_2__1330_,data_stage_2__1329_,
  data_stage_2__1328_,data_stage_2__1327_,data_stage_2__1326_,data_stage_2__1325_,
  data_stage_2__1324_,data_stage_2__1323_,data_stage_2__1322_,data_stage_2__1321_,
  data_stage_2__1320_,data_stage_2__1319_,data_stage_2__1318_,data_stage_2__1317_,
  data_stage_2__1316_,data_stage_2__1315_,data_stage_2__1314_,data_stage_2__1313_,
  data_stage_2__1312_,data_stage_2__1311_,data_stage_2__1310_,data_stage_2__1309_,
  data_stage_2__1308_,data_stage_2__1307_,data_stage_2__1306_,data_stage_2__1305_,
  data_stage_2__1304_,data_stage_2__1303_,data_stage_2__1302_,data_stage_2__1301_,
  data_stage_2__1300_,data_stage_2__1299_,data_stage_2__1298_,data_stage_2__1297_,
  data_stage_2__1296_,data_stage_2__1295_,data_stage_2__1294_,data_stage_2__1293_,
  data_stage_2__1292_,data_stage_2__1291_,data_stage_2__1290_,data_stage_2__1289_,
  data_stage_2__1288_,data_stage_2__1287_,data_stage_2__1286_,data_stage_2__1285_,
  data_stage_2__1284_,data_stage_2__1283_,data_stage_2__1282_,data_stage_2__1281_,
  data_stage_2__1280_,data_stage_2__1279_,data_stage_2__1278_,data_stage_2__1277_,
  data_stage_2__1276_,data_stage_2__1275_,data_stage_2__1274_,data_stage_2__1273_,
  data_stage_2__1272_,data_stage_2__1271_,data_stage_2__1270_,data_stage_2__1269_,
  data_stage_2__1268_,data_stage_2__1267_,data_stage_2__1266_,data_stage_2__1265_,
  data_stage_2__1264_,data_stage_2__1263_,data_stage_2__1262_,data_stage_2__1261_,
  data_stage_2__1260_,data_stage_2__1259_,data_stage_2__1258_,data_stage_2__1257_,
  data_stage_2__1256_,data_stage_2__1255_,data_stage_2__1254_,data_stage_2__1253_,
  data_stage_2__1252_,data_stage_2__1251_,data_stage_2__1250_,data_stage_2__1249_,
  data_stage_2__1248_,data_stage_2__1247_,data_stage_2__1246_,data_stage_2__1245_,
  data_stage_2__1244_,data_stage_2__1243_,data_stage_2__1242_,data_stage_2__1241_,
  data_stage_2__1240_,data_stage_2__1239_,data_stage_2__1238_,data_stage_2__1237_,
  data_stage_2__1236_,data_stage_2__1235_,data_stage_2__1234_,data_stage_2__1233_,
  data_stage_2__1232_,data_stage_2__1231_,data_stage_2__1230_,data_stage_2__1229_,
  data_stage_2__1228_,data_stage_2__1227_,data_stage_2__1226_,data_stage_2__1225_,
  data_stage_2__1224_,data_stage_2__1223_,data_stage_2__1222_,data_stage_2__1221_,
  data_stage_2__1220_,data_stage_2__1219_,data_stage_2__1218_,data_stage_2__1217_,
  data_stage_2__1216_,data_stage_2__1215_,data_stage_2__1214_,data_stage_2__1213_,
  data_stage_2__1212_,data_stage_2__1211_,data_stage_2__1210_,data_stage_2__1209_,
  data_stage_2__1208_,data_stage_2__1207_,data_stage_2__1206_,data_stage_2__1205_,
  data_stage_2__1204_,data_stage_2__1203_,data_stage_2__1202_,data_stage_2__1201_,
  data_stage_2__1200_,data_stage_2__1199_,data_stage_2__1198_,data_stage_2__1197_,
  data_stage_2__1196_,data_stage_2__1195_,data_stage_2__1194_,data_stage_2__1193_,
  data_stage_2__1192_,data_stage_2__1191_,data_stage_2__1190_,data_stage_2__1189_,
  data_stage_2__1188_,data_stage_2__1187_,data_stage_2__1186_,data_stage_2__1185_,
  data_stage_2__1184_,data_stage_2__1183_,data_stage_2__1182_,data_stage_2__1181_,
  data_stage_2__1180_,data_stage_2__1179_,data_stage_2__1178_,data_stage_2__1177_,
  data_stage_2__1176_,data_stage_2__1175_,data_stage_2__1174_,data_stage_2__1173_,
  data_stage_2__1172_,data_stage_2__1171_,data_stage_2__1170_,data_stage_2__1169_,
  data_stage_2__1168_,data_stage_2__1167_,data_stage_2__1166_,data_stage_2__1165_,
  data_stage_2__1164_,data_stage_2__1163_,data_stage_2__1162_,data_stage_2__1161_,
  data_stage_2__1160_,data_stage_2__1159_,data_stage_2__1158_,data_stage_2__1157_,
  data_stage_2__1156_,data_stage_2__1155_,data_stage_2__1154_,data_stage_2__1153_,
  data_stage_2__1152_,data_stage_2__1151_,data_stage_2__1150_,data_stage_2__1149_,
  data_stage_2__1148_,data_stage_2__1147_,data_stage_2__1146_,data_stage_2__1145_,
  data_stage_2__1144_,data_stage_2__1143_,data_stage_2__1142_,data_stage_2__1141_,
  data_stage_2__1140_,data_stage_2__1139_,data_stage_2__1138_,data_stage_2__1137_,
  data_stage_2__1136_,data_stage_2__1135_,data_stage_2__1134_,data_stage_2__1133_,
  data_stage_2__1132_,data_stage_2__1131_,data_stage_2__1130_,data_stage_2__1129_,
  data_stage_2__1128_,data_stage_2__1127_,data_stage_2__1126_,data_stage_2__1125_,
  data_stage_2__1124_,data_stage_2__1123_,data_stage_2__1122_,data_stage_2__1121_,
  data_stage_2__1120_,data_stage_2__1119_,data_stage_2__1118_,data_stage_2__1117_,
  data_stage_2__1116_,data_stage_2__1115_,data_stage_2__1114_,data_stage_2__1113_,
  data_stage_2__1112_,data_stage_2__1111_,data_stage_2__1110_,data_stage_2__1109_,
  data_stage_2__1108_,data_stage_2__1107_,data_stage_2__1106_,data_stage_2__1105_,
  data_stage_2__1104_,data_stage_2__1103_,data_stage_2__1102_,data_stage_2__1101_,
  data_stage_2__1100_,data_stage_2__1099_,data_stage_2__1098_,data_stage_2__1097_,
  data_stage_2__1096_,data_stage_2__1095_,data_stage_2__1094_,data_stage_2__1093_,
  data_stage_2__1092_,data_stage_2__1091_,data_stage_2__1090_,data_stage_2__1089_,
  data_stage_2__1088_,data_stage_2__1087_,data_stage_2__1086_,data_stage_2__1085_,
  data_stage_2__1084_,data_stage_2__1083_,data_stage_2__1082_,data_stage_2__1081_,
  data_stage_2__1080_,data_stage_2__1079_,data_stage_2__1078_,data_stage_2__1077_,
  data_stage_2__1076_,data_stage_2__1075_,data_stage_2__1074_,data_stage_2__1073_,
  data_stage_2__1072_,data_stage_2__1071_,data_stage_2__1070_,data_stage_2__1069_,
  data_stage_2__1068_,data_stage_2__1067_,data_stage_2__1066_,data_stage_2__1065_,
  data_stage_2__1064_,data_stage_2__1063_,data_stage_2__1062_,data_stage_2__1061_,
  data_stage_2__1060_,data_stage_2__1059_,data_stage_2__1058_,data_stage_2__1057_,
  data_stage_2__1056_,data_stage_2__1055_,data_stage_2__1054_,data_stage_2__1053_,
  data_stage_2__1052_,data_stage_2__1051_,data_stage_2__1050_,data_stage_2__1049_,
  data_stage_2__1048_,data_stage_2__1047_,data_stage_2__1046_,data_stage_2__1045_,
  data_stage_2__1044_,data_stage_2__1043_,data_stage_2__1042_,data_stage_2__1041_,
  data_stage_2__1040_,data_stage_2__1039_,data_stage_2__1038_,data_stage_2__1037_,
  data_stage_2__1036_,data_stage_2__1035_,data_stage_2__1034_,data_stage_2__1033_,
  data_stage_2__1032_,data_stage_2__1031_,data_stage_2__1030_,data_stage_2__1029_,
  data_stage_2__1028_,data_stage_2__1027_,data_stage_2__1026_,data_stage_2__1025_,
  data_stage_2__1024_,data_stage_2__1023_,data_stage_2__1022_,data_stage_2__1021_,
  data_stage_2__1020_,data_stage_2__1019_,data_stage_2__1018_,data_stage_2__1017_,
  data_stage_2__1016_,data_stage_2__1015_,data_stage_2__1014_,data_stage_2__1013_,
  data_stage_2__1012_,data_stage_2__1011_,data_stage_2__1010_,data_stage_2__1009_,
  data_stage_2__1008_,data_stage_2__1007_,data_stage_2__1006_,data_stage_2__1005_,
  data_stage_2__1004_,data_stage_2__1003_,data_stage_2__1002_,data_stage_2__1001_,
  data_stage_2__1000_,data_stage_2__999_,data_stage_2__998_,data_stage_2__997_,
  data_stage_2__996_,data_stage_2__995_,data_stage_2__994_,data_stage_2__993_,
  data_stage_2__992_,data_stage_2__991_,data_stage_2__990_,data_stage_2__989_,data_stage_2__988_,
  data_stage_2__987_,data_stage_2__986_,data_stage_2__985_,data_stage_2__984_,
  data_stage_2__983_,data_stage_2__982_,data_stage_2__981_,data_stage_2__980_,
  data_stage_2__979_,data_stage_2__978_,data_stage_2__977_,data_stage_2__976_,
  data_stage_2__975_,data_stage_2__974_,data_stage_2__973_,data_stage_2__972_,
  data_stage_2__971_,data_stage_2__970_,data_stage_2__969_,data_stage_2__968_,data_stage_2__967_,
  data_stage_2__966_,data_stage_2__965_,data_stage_2__964_,data_stage_2__963_,
  data_stage_2__962_,data_stage_2__961_,data_stage_2__960_,data_stage_2__959_,
  data_stage_2__958_,data_stage_2__957_,data_stage_2__956_,data_stage_2__955_,
  data_stage_2__954_,data_stage_2__953_,data_stage_2__952_,data_stage_2__951_,data_stage_2__950_,
  data_stage_2__949_,data_stage_2__948_,data_stage_2__947_,data_stage_2__946_,
  data_stage_2__945_,data_stage_2__944_,data_stage_2__943_,data_stage_2__942_,
  data_stage_2__941_,data_stage_2__940_,data_stage_2__939_,data_stage_2__938_,
  data_stage_2__937_,data_stage_2__936_,data_stage_2__935_,data_stage_2__934_,
  data_stage_2__933_,data_stage_2__932_,data_stage_2__931_,data_stage_2__930_,data_stage_2__929_,
  data_stage_2__928_,data_stage_2__927_,data_stage_2__926_,data_stage_2__925_,
  data_stage_2__924_,data_stage_2__923_,data_stage_2__922_,data_stage_2__921_,
  data_stage_2__920_,data_stage_2__919_,data_stage_2__918_,data_stage_2__917_,
  data_stage_2__916_,data_stage_2__915_,data_stage_2__914_,data_stage_2__913_,
  data_stage_2__912_,data_stage_2__911_,data_stage_2__910_,data_stage_2__909_,data_stage_2__908_,
  data_stage_2__907_,data_stage_2__906_,data_stage_2__905_,data_stage_2__904_,
  data_stage_2__903_,data_stage_2__902_,data_stage_2__901_,data_stage_2__900_,
  data_stage_2__899_,data_stage_2__898_,data_stage_2__897_,data_stage_2__896_,
  data_stage_2__895_,data_stage_2__894_,data_stage_2__893_,data_stage_2__892_,
  data_stage_2__891_,data_stage_2__890_,data_stage_2__889_,data_stage_2__888_,data_stage_2__887_,
  data_stage_2__886_,data_stage_2__885_,data_stage_2__884_,data_stage_2__883_,
  data_stage_2__882_,data_stage_2__881_,data_stage_2__880_,data_stage_2__879_,
  data_stage_2__878_,data_stage_2__877_,data_stage_2__876_,data_stage_2__875_,
  data_stage_2__874_,data_stage_2__873_,data_stage_2__872_,data_stage_2__871_,data_stage_2__870_,
  data_stage_2__869_,data_stage_2__868_,data_stage_2__867_,data_stage_2__866_,
  data_stage_2__865_,data_stage_2__864_,data_stage_2__863_,data_stage_2__862_,
  data_stage_2__861_,data_stage_2__860_,data_stage_2__859_,data_stage_2__858_,
  data_stage_2__857_,data_stage_2__856_,data_stage_2__855_,data_stage_2__854_,
  data_stage_2__853_,data_stage_2__852_,data_stage_2__851_,data_stage_2__850_,data_stage_2__849_,
  data_stage_2__848_,data_stage_2__847_,data_stage_2__846_,data_stage_2__845_,
  data_stage_2__844_,data_stage_2__843_,data_stage_2__842_,data_stage_2__841_,
  data_stage_2__840_,data_stage_2__839_,data_stage_2__838_,data_stage_2__837_,
  data_stage_2__836_,data_stage_2__835_,data_stage_2__834_,data_stage_2__833_,
  data_stage_2__832_,data_stage_2__831_,data_stage_2__830_,data_stage_2__829_,data_stage_2__828_,
  data_stage_2__827_,data_stage_2__826_,data_stage_2__825_,data_stage_2__824_,
  data_stage_2__823_,data_stage_2__822_,data_stage_2__821_,data_stage_2__820_,
  data_stage_2__819_,data_stage_2__818_,data_stage_2__817_,data_stage_2__816_,
  data_stage_2__815_,data_stage_2__814_,data_stage_2__813_,data_stage_2__812_,
  data_stage_2__811_,data_stage_2__810_,data_stage_2__809_,data_stage_2__808_,data_stage_2__807_,
  data_stage_2__806_,data_stage_2__805_,data_stage_2__804_,data_stage_2__803_,
  data_stage_2__802_,data_stage_2__801_,data_stage_2__800_,data_stage_2__799_,
  data_stage_2__798_,data_stage_2__797_,data_stage_2__796_,data_stage_2__795_,
  data_stage_2__794_,data_stage_2__793_,data_stage_2__792_,data_stage_2__791_,data_stage_2__790_,
  data_stage_2__789_,data_stage_2__788_,data_stage_2__787_,data_stage_2__786_,
  data_stage_2__785_,data_stage_2__784_,data_stage_2__783_,data_stage_2__782_,
  data_stage_2__781_,data_stage_2__780_,data_stage_2__779_,data_stage_2__778_,
  data_stage_2__777_,data_stage_2__776_,data_stage_2__775_,data_stage_2__774_,
  data_stage_2__773_,data_stage_2__772_,data_stage_2__771_,data_stage_2__770_,data_stage_2__769_,
  data_stage_2__768_,data_stage_2__767_,data_stage_2__766_,data_stage_2__765_,
  data_stage_2__764_,data_stage_2__763_,data_stage_2__762_,data_stage_2__761_,
  data_stage_2__760_,data_stage_2__759_,data_stage_2__758_,data_stage_2__757_,
  data_stage_2__756_,data_stage_2__755_,data_stage_2__754_,data_stage_2__753_,
  data_stage_2__752_,data_stage_2__751_,data_stage_2__750_,data_stage_2__749_,data_stage_2__748_,
  data_stage_2__747_,data_stage_2__746_,data_stage_2__745_,data_stage_2__744_,
  data_stage_2__743_,data_stage_2__742_,data_stage_2__741_,data_stage_2__740_,
  data_stage_2__739_,data_stage_2__738_,data_stage_2__737_,data_stage_2__736_,
  data_stage_2__735_,data_stage_2__734_,data_stage_2__733_,data_stage_2__732_,
  data_stage_2__731_,data_stage_2__730_,data_stage_2__729_,data_stage_2__728_,data_stage_2__727_,
  data_stage_2__726_,data_stage_2__725_,data_stage_2__724_,data_stage_2__723_,
  data_stage_2__722_,data_stage_2__721_,data_stage_2__720_,data_stage_2__719_,
  data_stage_2__718_,data_stage_2__717_,data_stage_2__716_,data_stage_2__715_,
  data_stage_2__714_,data_stage_2__713_,data_stage_2__712_,data_stage_2__711_,data_stage_2__710_,
  data_stage_2__709_,data_stage_2__708_,data_stage_2__707_,data_stage_2__706_,
  data_stage_2__705_,data_stage_2__704_,data_stage_2__703_,data_stage_2__702_,
  data_stage_2__701_,data_stage_2__700_,data_stage_2__699_,data_stage_2__698_,
  data_stage_2__697_,data_stage_2__696_,data_stage_2__695_,data_stage_2__694_,
  data_stage_2__693_,data_stage_2__692_,data_stage_2__691_,data_stage_2__690_,data_stage_2__689_,
  data_stage_2__688_,data_stage_2__687_,data_stage_2__686_,data_stage_2__685_,
  data_stage_2__684_,data_stage_2__683_,data_stage_2__682_,data_stage_2__681_,
  data_stage_2__680_,data_stage_2__679_,data_stage_2__678_,data_stage_2__677_,
  data_stage_2__676_,data_stage_2__675_,data_stage_2__674_,data_stage_2__673_,
  data_stage_2__672_,data_stage_2__671_,data_stage_2__670_,data_stage_2__669_,data_stage_2__668_,
  data_stage_2__667_,data_stage_2__666_,data_stage_2__665_,data_stage_2__664_,
  data_stage_2__663_,data_stage_2__662_,data_stage_2__661_,data_stage_2__660_,
  data_stage_2__659_,data_stage_2__658_,data_stage_2__657_,data_stage_2__656_,
  data_stage_2__655_,data_stage_2__654_,data_stage_2__653_,data_stage_2__652_,
  data_stage_2__651_,data_stage_2__650_,data_stage_2__649_,data_stage_2__648_,data_stage_2__647_,
  data_stage_2__646_,data_stage_2__645_,data_stage_2__644_,data_stage_2__643_,
  data_stage_2__642_,data_stage_2__641_,data_stage_2__640_,data_stage_2__639_,
  data_stage_2__638_,data_stage_2__637_,data_stage_2__636_,data_stage_2__635_,
  data_stage_2__634_,data_stage_2__633_,data_stage_2__632_,data_stage_2__631_,data_stage_2__630_,
  data_stage_2__629_,data_stage_2__628_,data_stage_2__627_,data_stage_2__626_,
  data_stage_2__625_,data_stage_2__624_,data_stage_2__623_,data_stage_2__622_,
  data_stage_2__621_,data_stage_2__620_,data_stage_2__619_,data_stage_2__618_,
  data_stage_2__617_,data_stage_2__616_,data_stage_2__615_,data_stage_2__614_,
  data_stage_2__613_,data_stage_2__612_,data_stage_2__611_,data_stage_2__610_,data_stage_2__609_,
  data_stage_2__608_,data_stage_2__607_,data_stage_2__606_,data_stage_2__605_,
  data_stage_2__604_,data_stage_2__603_,data_stage_2__602_,data_stage_2__601_,
  data_stage_2__600_,data_stage_2__599_,data_stage_2__598_,data_stage_2__597_,
  data_stage_2__596_,data_stage_2__595_,data_stage_2__594_,data_stage_2__593_,
  data_stage_2__592_,data_stage_2__591_,data_stage_2__590_,data_stage_2__589_,data_stage_2__588_,
  data_stage_2__587_,data_stage_2__586_,data_stage_2__585_,data_stage_2__584_,
  data_stage_2__583_,data_stage_2__582_,data_stage_2__581_,data_stage_2__580_,
  data_stage_2__579_,data_stage_2__578_,data_stage_2__577_,data_stage_2__576_,
  data_stage_2__575_,data_stage_2__574_,data_stage_2__573_,data_stage_2__572_,
  data_stage_2__571_,data_stage_2__570_,data_stage_2__569_,data_stage_2__568_,data_stage_2__567_,
  data_stage_2__566_,data_stage_2__565_,data_stage_2__564_,data_stage_2__563_,
  data_stage_2__562_,data_stage_2__561_,data_stage_2__560_,data_stage_2__559_,
  data_stage_2__558_,data_stage_2__557_,data_stage_2__556_,data_stage_2__555_,
  data_stage_2__554_,data_stage_2__553_,data_stage_2__552_,data_stage_2__551_,data_stage_2__550_,
  data_stage_2__549_,data_stage_2__548_,data_stage_2__547_,data_stage_2__546_,
  data_stage_2__545_,data_stage_2__544_,data_stage_2__543_,data_stage_2__542_,
  data_stage_2__541_,data_stage_2__540_,data_stage_2__539_,data_stage_2__538_,
  data_stage_2__537_,data_stage_2__536_,data_stage_2__535_,data_stage_2__534_,
  data_stage_2__533_,data_stage_2__532_,data_stage_2__531_,data_stage_2__530_,data_stage_2__529_,
  data_stage_2__528_,data_stage_2__527_,data_stage_2__526_,data_stage_2__525_,
  data_stage_2__524_,data_stage_2__523_,data_stage_2__522_,data_stage_2__521_,
  data_stage_2__520_,data_stage_2__519_,data_stage_2__518_,data_stage_2__517_,
  data_stage_2__516_,data_stage_2__515_,data_stage_2__514_,data_stage_2__513_,
  data_stage_2__512_,data_stage_2__511_,data_stage_2__510_,data_stage_2__509_,data_stage_2__508_,
  data_stage_2__507_,data_stage_2__506_,data_stage_2__505_,data_stage_2__504_,
  data_stage_2__503_,data_stage_2__502_,data_stage_2__501_,data_stage_2__500_,
  data_stage_2__499_,data_stage_2__498_,data_stage_2__497_,data_stage_2__496_,
  data_stage_2__495_,data_stage_2__494_,data_stage_2__493_,data_stage_2__492_,
  data_stage_2__491_,data_stage_2__490_,data_stage_2__489_,data_stage_2__488_,data_stage_2__487_,
  data_stage_2__486_,data_stage_2__485_,data_stage_2__484_,data_stage_2__483_,
  data_stage_2__482_,data_stage_2__481_,data_stage_2__480_,data_stage_2__479_,
  data_stage_2__478_,data_stage_2__477_,data_stage_2__476_,data_stage_2__475_,
  data_stage_2__474_,data_stage_2__473_,data_stage_2__472_,data_stage_2__471_,data_stage_2__470_,
  data_stage_2__469_,data_stage_2__468_,data_stage_2__467_,data_stage_2__466_,
  data_stage_2__465_,data_stage_2__464_,data_stage_2__463_,data_stage_2__462_,
  data_stage_2__461_,data_stage_2__460_,data_stage_2__459_,data_stage_2__458_,
  data_stage_2__457_,data_stage_2__456_,data_stage_2__455_,data_stage_2__454_,
  data_stage_2__453_,data_stage_2__452_,data_stage_2__451_,data_stage_2__450_,data_stage_2__449_,
  data_stage_2__448_,data_stage_2__447_,data_stage_2__446_,data_stage_2__445_,
  data_stage_2__444_,data_stage_2__443_,data_stage_2__442_,data_stage_2__441_,
  data_stage_2__440_,data_stage_2__439_,data_stage_2__438_,data_stage_2__437_,
  data_stage_2__436_,data_stage_2__435_,data_stage_2__434_,data_stage_2__433_,
  data_stage_2__432_,data_stage_2__431_,data_stage_2__430_,data_stage_2__429_,data_stage_2__428_,
  data_stage_2__427_,data_stage_2__426_,data_stage_2__425_,data_stage_2__424_,
  data_stage_2__423_,data_stage_2__422_,data_stage_2__421_,data_stage_2__420_,
  data_stage_2__419_,data_stage_2__418_,data_stage_2__417_,data_stage_2__416_,
  data_stage_2__415_,data_stage_2__414_,data_stage_2__413_,data_stage_2__412_,
  data_stage_2__411_,data_stage_2__410_,data_stage_2__409_,data_stage_2__408_,data_stage_2__407_,
  data_stage_2__406_,data_stage_2__405_,data_stage_2__404_,data_stage_2__403_,
  data_stage_2__402_,data_stage_2__401_,data_stage_2__400_,data_stage_2__399_,
  data_stage_2__398_,data_stage_2__397_,data_stage_2__396_,data_stage_2__395_,
  data_stage_2__394_,data_stage_2__393_,data_stage_2__392_,data_stage_2__391_,data_stage_2__390_,
  data_stage_2__389_,data_stage_2__388_,data_stage_2__387_,data_stage_2__386_,
  data_stage_2__385_,data_stage_2__384_,data_stage_2__383_,data_stage_2__382_,
  data_stage_2__381_,data_stage_2__380_,data_stage_2__379_,data_stage_2__378_,
  data_stage_2__377_,data_stage_2__376_,data_stage_2__375_,data_stage_2__374_,
  data_stage_2__373_,data_stage_2__372_,data_stage_2__371_,data_stage_2__370_,data_stage_2__369_,
  data_stage_2__368_,data_stage_2__367_,data_stage_2__366_,data_stage_2__365_,
  data_stage_2__364_,data_stage_2__363_,data_stage_2__362_,data_stage_2__361_,
  data_stage_2__360_,data_stage_2__359_,data_stage_2__358_,data_stage_2__357_,
  data_stage_2__356_,data_stage_2__355_,data_stage_2__354_,data_stage_2__353_,
  data_stage_2__352_,data_stage_2__351_,data_stage_2__350_,data_stage_2__349_,data_stage_2__348_,
  data_stage_2__347_,data_stage_2__346_,data_stage_2__345_,data_stage_2__344_,
  data_stage_2__343_,data_stage_2__342_,data_stage_2__341_,data_stage_2__340_,
  data_stage_2__339_,data_stage_2__338_,data_stage_2__337_,data_stage_2__336_,
  data_stage_2__335_,data_stage_2__334_,data_stage_2__333_,data_stage_2__332_,
  data_stage_2__331_,data_stage_2__330_,data_stage_2__329_,data_stage_2__328_,data_stage_2__327_,
  data_stage_2__326_,data_stage_2__325_,data_stage_2__324_,data_stage_2__323_,
  data_stage_2__322_,data_stage_2__321_,data_stage_2__320_,data_stage_2__319_,
  data_stage_2__318_,data_stage_2__317_,data_stage_2__316_,data_stage_2__315_,
  data_stage_2__314_,data_stage_2__313_,data_stage_2__312_,data_stage_2__311_,data_stage_2__310_,
  data_stage_2__309_,data_stage_2__308_,data_stage_2__307_,data_stage_2__306_,
  data_stage_2__305_,data_stage_2__304_,data_stage_2__303_,data_stage_2__302_,
  data_stage_2__301_,data_stage_2__300_,data_stage_2__299_,data_stage_2__298_,
  data_stage_2__297_,data_stage_2__296_,data_stage_2__295_,data_stage_2__294_,
  data_stage_2__293_,data_stage_2__292_,data_stage_2__291_,data_stage_2__290_,data_stage_2__289_,
  data_stage_2__288_,data_stage_2__287_,data_stage_2__286_,data_stage_2__285_,
  data_stage_2__284_,data_stage_2__283_,data_stage_2__282_,data_stage_2__281_,
  data_stage_2__280_,data_stage_2__279_,data_stage_2__278_,data_stage_2__277_,
  data_stage_2__276_,data_stage_2__275_,data_stage_2__274_,data_stage_2__273_,
  data_stage_2__272_,data_stage_2__271_,data_stage_2__270_,data_stage_2__269_,data_stage_2__268_,
  data_stage_2__267_,data_stage_2__266_,data_stage_2__265_,data_stage_2__264_,
  data_stage_2__263_,data_stage_2__262_,data_stage_2__261_,data_stage_2__260_,
  data_stage_2__259_,data_stage_2__258_,data_stage_2__257_,data_stage_2__256_,
  data_stage_2__255_,data_stage_2__254_,data_stage_2__253_,data_stage_2__252_,
  data_stage_2__251_,data_stage_2__250_,data_stage_2__249_,data_stage_2__248_,data_stage_2__247_,
  data_stage_2__246_,data_stage_2__245_,data_stage_2__244_,data_stage_2__243_,
  data_stage_2__242_,data_stage_2__241_,data_stage_2__240_,data_stage_2__239_,
  data_stage_2__238_,data_stage_2__237_,data_stage_2__236_,data_stage_2__235_,
  data_stage_2__234_,data_stage_2__233_,data_stage_2__232_,data_stage_2__231_,data_stage_2__230_,
  data_stage_2__229_,data_stage_2__228_,data_stage_2__227_,data_stage_2__226_,
  data_stage_2__225_,data_stage_2__224_,data_stage_2__223_,data_stage_2__222_,
  data_stage_2__221_,data_stage_2__220_,data_stage_2__219_,data_stage_2__218_,
  data_stage_2__217_,data_stage_2__216_,data_stage_2__215_,data_stage_2__214_,
  data_stage_2__213_,data_stage_2__212_,data_stage_2__211_,data_stage_2__210_,data_stage_2__209_,
  data_stage_2__208_,data_stage_2__207_,data_stage_2__206_,data_stage_2__205_,
  data_stage_2__204_,data_stage_2__203_,data_stage_2__202_,data_stage_2__201_,
  data_stage_2__200_,data_stage_2__199_,data_stage_2__198_,data_stage_2__197_,
  data_stage_2__196_,data_stage_2__195_,data_stage_2__194_,data_stage_2__193_,
  data_stage_2__192_,data_stage_2__191_,data_stage_2__190_,data_stage_2__189_,data_stage_2__188_,
  data_stage_2__187_,data_stage_2__186_,data_stage_2__185_,data_stage_2__184_,
  data_stage_2__183_,data_stage_2__182_,data_stage_2__181_,data_stage_2__180_,
  data_stage_2__179_,data_stage_2__178_,data_stage_2__177_,data_stage_2__176_,
  data_stage_2__175_,data_stage_2__174_,data_stage_2__173_,data_stage_2__172_,
  data_stage_2__171_,data_stage_2__170_,data_stage_2__169_,data_stage_2__168_,data_stage_2__167_,
  data_stage_2__166_,data_stage_2__165_,data_stage_2__164_,data_stage_2__163_,
  data_stage_2__162_,data_stage_2__161_,data_stage_2__160_,data_stage_2__159_,
  data_stage_2__158_,data_stage_2__157_,data_stage_2__156_,data_stage_2__155_,
  data_stage_2__154_,data_stage_2__153_,data_stage_2__152_,data_stage_2__151_,data_stage_2__150_,
  data_stage_2__149_,data_stage_2__148_,data_stage_2__147_,data_stage_2__146_,
  data_stage_2__145_,data_stage_2__144_,data_stage_2__143_,data_stage_2__142_,
  data_stage_2__141_,data_stage_2__140_,data_stage_2__139_,data_stage_2__138_,
  data_stage_2__137_,data_stage_2__136_,data_stage_2__135_,data_stage_2__134_,
  data_stage_2__133_,data_stage_2__132_,data_stage_2__131_,data_stage_2__130_,data_stage_2__129_,
  data_stage_2__128_,data_stage_2__127_,data_stage_2__126_,data_stage_2__125_,
  data_stage_2__124_,data_stage_2__123_,data_stage_2__122_,data_stage_2__121_,
  data_stage_2__120_,data_stage_2__119_,data_stage_2__118_,data_stage_2__117_,
  data_stage_2__116_,data_stage_2__115_,data_stage_2__114_,data_stage_2__113_,
  data_stage_2__112_,data_stage_2__111_,data_stage_2__110_,data_stage_2__109_,data_stage_2__108_,
  data_stage_2__107_,data_stage_2__106_,data_stage_2__105_,data_stage_2__104_,
  data_stage_2__103_,data_stage_2__102_,data_stage_2__101_,data_stage_2__100_,
  data_stage_2__99_,data_stage_2__98_,data_stage_2__97_,data_stage_2__96_,data_stage_2__95_,
  data_stage_2__94_,data_stage_2__93_,data_stage_2__92_,data_stage_2__91_,
  data_stage_2__90_,data_stage_2__89_,data_stage_2__88_,data_stage_2__87_,
  data_stage_2__86_,data_stage_2__85_,data_stage_2__84_,data_stage_2__83_,data_stage_2__82_,
  data_stage_2__81_,data_stage_2__80_,data_stage_2__79_,data_stage_2__78_,
  data_stage_2__77_,data_stage_2__76_,data_stage_2__75_,data_stage_2__74_,data_stage_2__73_,
  data_stage_2__72_,data_stage_2__71_,data_stage_2__70_,data_stage_2__69_,
  data_stage_2__68_,data_stage_2__67_,data_stage_2__66_,data_stage_2__65_,data_stage_2__64_,
  data_stage_2__63_,data_stage_2__62_,data_stage_2__61_,data_stage_2__60_,
  data_stage_2__59_,data_stage_2__58_,data_stage_2__57_,data_stage_2__56_,data_stage_2__55_,
  data_stage_2__54_,data_stage_2__53_,data_stage_2__52_,data_stage_2__51_,
  data_stage_2__50_,data_stage_2__49_,data_stage_2__48_,data_stage_2__47_,
  data_stage_2__46_,data_stage_2__45_,data_stage_2__44_,data_stage_2__43_,data_stage_2__42_,
  data_stage_2__41_,data_stage_2__40_,data_stage_2__39_,data_stage_2__38_,
  data_stage_2__37_,data_stage_2__36_,data_stage_2__35_,data_stage_2__34_,data_stage_2__33_,
  data_stage_2__32_,data_stage_2__31_,data_stage_2__30_,data_stage_2__29_,
  data_stage_2__28_,data_stage_2__27_,data_stage_2__26_,data_stage_2__25_,data_stage_2__24_,
  data_stage_2__23_,data_stage_2__22_,data_stage_2__21_,data_stage_2__20_,
  data_stage_2__19_,data_stage_2__18_,data_stage_2__17_,data_stage_2__16_,data_stage_2__15_,
  data_stage_2__14_,data_stage_2__13_,data_stage_2__12_,data_stage_2__11_,
  data_stage_2__10_,data_stage_2__9_,data_stage_2__8_,data_stage_2__7_,data_stage_2__6_,
  data_stage_2__5_,data_stage_2__4_,data_stage_2__3_,data_stage_2__2_,
  data_stage_2__1_,data_stage_2__0_,data_stage_3__4095_,data_stage_3__4094_,data_stage_3__4093_,
  data_stage_3__4092_,data_stage_3__4091_,data_stage_3__4090_,data_stage_3__4089_,
  data_stage_3__4088_,data_stage_3__4087_,data_stage_3__4086_,data_stage_3__4085_,
  data_stage_3__4084_,data_stage_3__4083_,data_stage_3__4082_,data_stage_3__4081_,
  data_stage_3__4080_,data_stage_3__4079_,data_stage_3__4078_,data_stage_3__4077_,
  data_stage_3__4076_,data_stage_3__4075_,data_stage_3__4074_,data_stage_3__4073_,
  data_stage_3__4072_,data_stage_3__4071_,data_stage_3__4070_,data_stage_3__4069_,
  data_stage_3__4068_,data_stage_3__4067_,data_stage_3__4066_,data_stage_3__4065_,
  data_stage_3__4064_,data_stage_3__4063_,data_stage_3__4062_,data_stage_3__4061_,
  data_stage_3__4060_,data_stage_3__4059_,data_stage_3__4058_,data_stage_3__4057_,
  data_stage_3__4056_,data_stage_3__4055_,data_stage_3__4054_,data_stage_3__4053_,
  data_stage_3__4052_,data_stage_3__4051_,data_stage_3__4050_,data_stage_3__4049_,
  data_stage_3__4048_,data_stage_3__4047_,data_stage_3__4046_,data_stage_3__4045_,
  data_stage_3__4044_,data_stage_3__4043_,data_stage_3__4042_,data_stage_3__4041_,
  data_stage_3__4040_,data_stage_3__4039_,data_stage_3__4038_,data_stage_3__4037_,
  data_stage_3__4036_,data_stage_3__4035_,data_stage_3__4034_,data_stage_3__4033_,
  data_stage_3__4032_,data_stage_3__4031_,data_stage_3__4030_,data_stage_3__4029_,
  data_stage_3__4028_,data_stage_3__4027_,data_stage_3__4026_,data_stage_3__4025_,
  data_stage_3__4024_,data_stage_3__4023_,data_stage_3__4022_,data_stage_3__4021_,
  data_stage_3__4020_,data_stage_3__4019_,data_stage_3__4018_,data_stage_3__4017_,
  data_stage_3__4016_,data_stage_3__4015_,data_stage_3__4014_,data_stage_3__4013_,
  data_stage_3__4012_,data_stage_3__4011_,data_stage_3__4010_,data_stage_3__4009_,
  data_stage_3__4008_,data_stage_3__4007_,data_stage_3__4006_,data_stage_3__4005_,
  data_stage_3__4004_,data_stage_3__4003_,data_stage_3__4002_,data_stage_3__4001_,
  data_stage_3__4000_,data_stage_3__3999_,data_stage_3__3998_,data_stage_3__3997_,
  data_stage_3__3996_,data_stage_3__3995_,data_stage_3__3994_,data_stage_3__3993_,
  data_stage_3__3992_,data_stage_3__3991_,data_stage_3__3990_,data_stage_3__3989_,
  data_stage_3__3988_,data_stage_3__3987_,data_stage_3__3986_,data_stage_3__3985_,
  data_stage_3__3984_,data_stage_3__3983_,data_stage_3__3982_,data_stage_3__3981_,
  data_stage_3__3980_,data_stage_3__3979_,data_stage_3__3978_,data_stage_3__3977_,
  data_stage_3__3976_,data_stage_3__3975_,data_stage_3__3974_,data_stage_3__3973_,
  data_stage_3__3972_,data_stage_3__3971_,data_stage_3__3970_,data_stage_3__3969_,
  data_stage_3__3968_,data_stage_3__3967_,data_stage_3__3966_,data_stage_3__3965_,
  data_stage_3__3964_,data_stage_3__3963_,data_stage_3__3962_,data_stage_3__3961_,
  data_stage_3__3960_,data_stage_3__3959_,data_stage_3__3958_,data_stage_3__3957_,
  data_stage_3__3956_,data_stage_3__3955_,data_stage_3__3954_,data_stage_3__3953_,
  data_stage_3__3952_,data_stage_3__3951_,data_stage_3__3950_,data_stage_3__3949_,
  data_stage_3__3948_,data_stage_3__3947_,data_stage_3__3946_,data_stage_3__3945_,
  data_stage_3__3944_,data_stage_3__3943_,data_stage_3__3942_,data_stage_3__3941_,
  data_stage_3__3940_,data_stage_3__3939_,data_stage_3__3938_,data_stage_3__3937_,
  data_stage_3__3936_,data_stage_3__3935_,data_stage_3__3934_,data_stage_3__3933_,
  data_stage_3__3932_,data_stage_3__3931_,data_stage_3__3930_,data_stage_3__3929_,
  data_stage_3__3928_,data_stage_3__3927_,data_stage_3__3926_,data_stage_3__3925_,
  data_stage_3__3924_,data_stage_3__3923_,data_stage_3__3922_,data_stage_3__3921_,
  data_stage_3__3920_,data_stage_3__3919_,data_stage_3__3918_,data_stage_3__3917_,
  data_stage_3__3916_,data_stage_3__3915_,data_stage_3__3914_,data_stage_3__3913_,
  data_stage_3__3912_,data_stage_3__3911_,data_stage_3__3910_,data_stage_3__3909_,
  data_stage_3__3908_,data_stage_3__3907_,data_stage_3__3906_,data_stage_3__3905_,
  data_stage_3__3904_,data_stage_3__3903_,data_stage_3__3902_,data_stage_3__3901_,
  data_stage_3__3900_,data_stage_3__3899_,data_stage_3__3898_,data_stage_3__3897_,
  data_stage_3__3896_,data_stage_3__3895_,data_stage_3__3894_,data_stage_3__3893_,
  data_stage_3__3892_,data_stage_3__3891_,data_stage_3__3890_,data_stage_3__3889_,
  data_stage_3__3888_,data_stage_3__3887_,data_stage_3__3886_,data_stage_3__3885_,
  data_stage_3__3884_,data_stage_3__3883_,data_stage_3__3882_,data_stage_3__3881_,
  data_stage_3__3880_,data_stage_3__3879_,data_stage_3__3878_,data_stage_3__3877_,
  data_stage_3__3876_,data_stage_3__3875_,data_stage_3__3874_,data_stage_3__3873_,
  data_stage_3__3872_,data_stage_3__3871_,data_stage_3__3870_,data_stage_3__3869_,
  data_stage_3__3868_,data_stage_3__3867_,data_stage_3__3866_,data_stage_3__3865_,
  data_stage_3__3864_,data_stage_3__3863_,data_stage_3__3862_,data_stage_3__3861_,
  data_stage_3__3860_,data_stage_3__3859_,data_stage_3__3858_,data_stage_3__3857_,
  data_stage_3__3856_,data_stage_3__3855_,data_stage_3__3854_,data_stage_3__3853_,
  data_stage_3__3852_,data_stage_3__3851_,data_stage_3__3850_,data_stage_3__3849_,
  data_stage_3__3848_,data_stage_3__3847_,data_stage_3__3846_,data_stage_3__3845_,
  data_stage_3__3844_,data_stage_3__3843_,data_stage_3__3842_,data_stage_3__3841_,
  data_stage_3__3840_,data_stage_3__3839_,data_stage_3__3838_,data_stage_3__3837_,
  data_stage_3__3836_,data_stage_3__3835_,data_stage_3__3834_,data_stage_3__3833_,
  data_stage_3__3832_,data_stage_3__3831_,data_stage_3__3830_,data_stage_3__3829_,
  data_stage_3__3828_,data_stage_3__3827_,data_stage_3__3826_,data_stage_3__3825_,
  data_stage_3__3824_,data_stage_3__3823_,data_stage_3__3822_,data_stage_3__3821_,
  data_stage_3__3820_,data_stage_3__3819_,data_stage_3__3818_,data_stage_3__3817_,
  data_stage_3__3816_,data_stage_3__3815_,data_stage_3__3814_,data_stage_3__3813_,
  data_stage_3__3812_,data_stage_3__3811_,data_stage_3__3810_,data_stage_3__3809_,
  data_stage_3__3808_,data_stage_3__3807_,data_stage_3__3806_,data_stage_3__3805_,
  data_stage_3__3804_,data_stage_3__3803_,data_stage_3__3802_,data_stage_3__3801_,
  data_stage_3__3800_,data_stage_3__3799_,data_stage_3__3798_,data_stage_3__3797_,
  data_stage_3__3796_,data_stage_3__3795_,data_stage_3__3794_,data_stage_3__3793_,
  data_stage_3__3792_,data_stage_3__3791_,data_stage_3__3790_,data_stage_3__3789_,
  data_stage_3__3788_,data_stage_3__3787_,data_stage_3__3786_,data_stage_3__3785_,
  data_stage_3__3784_,data_stage_3__3783_,data_stage_3__3782_,data_stage_3__3781_,
  data_stage_3__3780_,data_stage_3__3779_,data_stage_3__3778_,data_stage_3__3777_,
  data_stage_3__3776_,data_stage_3__3775_,data_stage_3__3774_,data_stage_3__3773_,
  data_stage_3__3772_,data_stage_3__3771_,data_stage_3__3770_,data_stage_3__3769_,
  data_stage_3__3768_,data_stage_3__3767_,data_stage_3__3766_,data_stage_3__3765_,
  data_stage_3__3764_,data_stage_3__3763_,data_stage_3__3762_,data_stage_3__3761_,
  data_stage_3__3760_,data_stage_3__3759_,data_stage_3__3758_,data_stage_3__3757_,
  data_stage_3__3756_,data_stage_3__3755_,data_stage_3__3754_,data_stage_3__3753_,
  data_stage_3__3752_,data_stage_3__3751_,data_stage_3__3750_,data_stage_3__3749_,
  data_stage_3__3748_,data_stage_3__3747_,data_stage_3__3746_,data_stage_3__3745_,
  data_stage_3__3744_,data_stage_3__3743_,data_stage_3__3742_,data_stage_3__3741_,
  data_stage_3__3740_,data_stage_3__3739_,data_stage_3__3738_,data_stage_3__3737_,
  data_stage_3__3736_,data_stage_3__3735_,data_stage_3__3734_,data_stage_3__3733_,
  data_stage_3__3732_,data_stage_3__3731_,data_stage_3__3730_,data_stage_3__3729_,
  data_stage_3__3728_,data_stage_3__3727_,data_stage_3__3726_,data_stage_3__3725_,
  data_stage_3__3724_,data_stage_3__3723_,data_stage_3__3722_,data_stage_3__3721_,
  data_stage_3__3720_,data_stage_3__3719_,data_stage_3__3718_,data_stage_3__3717_,
  data_stage_3__3716_,data_stage_3__3715_,data_stage_3__3714_,data_stage_3__3713_,
  data_stage_3__3712_,data_stage_3__3711_,data_stage_3__3710_,data_stage_3__3709_,
  data_stage_3__3708_,data_stage_3__3707_,data_stage_3__3706_,data_stage_3__3705_,
  data_stage_3__3704_,data_stage_3__3703_,data_stage_3__3702_,data_stage_3__3701_,
  data_stage_3__3700_,data_stage_3__3699_,data_stage_3__3698_,data_stage_3__3697_,
  data_stage_3__3696_,data_stage_3__3695_,data_stage_3__3694_,data_stage_3__3693_,
  data_stage_3__3692_,data_stage_3__3691_,data_stage_3__3690_,data_stage_3__3689_,
  data_stage_3__3688_,data_stage_3__3687_,data_stage_3__3686_,data_stage_3__3685_,
  data_stage_3__3684_,data_stage_3__3683_,data_stage_3__3682_,data_stage_3__3681_,
  data_stage_3__3680_,data_stage_3__3679_,data_stage_3__3678_,data_stage_3__3677_,
  data_stage_3__3676_,data_stage_3__3675_,data_stage_3__3674_,data_stage_3__3673_,
  data_stage_3__3672_,data_stage_3__3671_,data_stage_3__3670_,data_stage_3__3669_,
  data_stage_3__3668_,data_stage_3__3667_,data_stage_3__3666_,data_stage_3__3665_,
  data_stage_3__3664_,data_stage_3__3663_,data_stage_3__3662_,data_stage_3__3661_,
  data_stage_3__3660_,data_stage_3__3659_,data_stage_3__3658_,data_stage_3__3657_,
  data_stage_3__3656_,data_stage_3__3655_,data_stage_3__3654_,data_stage_3__3653_,
  data_stage_3__3652_,data_stage_3__3651_,data_stage_3__3650_,data_stage_3__3649_,
  data_stage_3__3648_,data_stage_3__3647_,data_stage_3__3646_,data_stage_3__3645_,
  data_stage_3__3644_,data_stage_3__3643_,data_stage_3__3642_,data_stage_3__3641_,
  data_stage_3__3640_,data_stage_3__3639_,data_stage_3__3638_,data_stage_3__3637_,
  data_stage_3__3636_,data_stage_3__3635_,data_stage_3__3634_,data_stage_3__3633_,
  data_stage_3__3632_,data_stage_3__3631_,data_stage_3__3630_,data_stage_3__3629_,
  data_stage_3__3628_,data_stage_3__3627_,data_stage_3__3626_,data_stage_3__3625_,
  data_stage_3__3624_,data_stage_3__3623_,data_stage_3__3622_,data_stage_3__3621_,
  data_stage_3__3620_,data_stage_3__3619_,data_stage_3__3618_,data_stage_3__3617_,
  data_stage_3__3616_,data_stage_3__3615_,data_stage_3__3614_,data_stage_3__3613_,
  data_stage_3__3612_,data_stage_3__3611_,data_stage_3__3610_,data_stage_3__3609_,
  data_stage_3__3608_,data_stage_3__3607_,data_stage_3__3606_,data_stage_3__3605_,
  data_stage_3__3604_,data_stage_3__3603_,data_stage_3__3602_,data_stage_3__3601_,
  data_stage_3__3600_,data_stage_3__3599_,data_stage_3__3598_,data_stage_3__3597_,
  data_stage_3__3596_,data_stage_3__3595_,data_stage_3__3594_,data_stage_3__3593_,
  data_stage_3__3592_,data_stage_3__3591_,data_stage_3__3590_,data_stage_3__3589_,
  data_stage_3__3588_,data_stage_3__3587_,data_stage_3__3586_,data_stage_3__3585_,
  data_stage_3__3584_,data_stage_3__3583_,data_stage_3__3582_,data_stage_3__3581_,
  data_stage_3__3580_,data_stage_3__3579_,data_stage_3__3578_,data_stage_3__3577_,
  data_stage_3__3576_,data_stage_3__3575_,data_stage_3__3574_,data_stage_3__3573_,
  data_stage_3__3572_,data_stage_3__3571_,data_stage_3__3570_,data_stage_3__3569_,
  data_stage_3__3568_,data_stage_3__3567_,data_stage_3__3566_,data_stage_3__3565_,
  data_stage_3__3564_,data_stage_3__3563_,data_stage_3__3562_,data_stage_3__3561_,
  data_stage_3__3560_,data_stage_3__3559_,data_stage_3__3558_,data_stage_3__3557_,
  data_stage_3__3556_,data_stage_3__3555_,data_stage_3__3554_,data_stage_3__3553_,
  data_stage_3__3552_,data_stage_3__3551_,data_stage_3__3550_,data_stage_3__3549_,
  data_stage_3__3548_,data_stage_3__3547_,data_stage_3__3546_,data_stage_3__3545_,
  data_stage_3__3544_,data_stage_3__3543_,data_stage_3__3542_,data_stage_3__3541_,
  data_stage_3__3540_,data_stage_3__3539_,data_stage_3__3538_,data_stage_3__3537_,
  data_stage_3__3536_,data_stage_3__3535_,data_stage_3__3534_,data_stage_3__3533_,
  data_stage_3__3532_,data_stage_3__3531_,data_stage_3__3530_,data_stage_3__3529_,
  data_stage_3__3528_,data_stage_3__3527_,data_stage_3__3526_,data_stage_3__3525_,
  data_stage_3__3524_,data_stage_3__3523_,data_stage_3__3522_,data_stage_3__3521_,
  data_stage_3__3520_,data_stage_3__3519_,data_stage_3__3518_,data_stage_3__3517_,
  data_stage_3__3516_,data_stage_3__3515_,data_stage_3__3514_,data_stage_3__3513_,
  data_stage_3__3512_,data_stage_3__3511_,data_stage_3__3510_,data_stage_3__3509_,
  data_stage_3__3508_,data_stage_3__3507_,data_stage_3__3506_,data_stage_3__3505_,
  data_stage_3__3504_,data_stage_3__3503_,data_stage_3__3502_,data_stage_3__3501_,
  data_stage_3__3500_,data_stage_3__3499_,data_stage_3__3498_,data_stage_3__3497_,
  data_stage_3__3496_,data_stage_3__3495_,data_stage_3__3494_,data_stage_3__3493_,
  data_stage_3__3492_,data_stage_3__3491_,data_stage_3__3490_,data_stage_3__3489_,
  data_stage_3__3488_,data_stage_3__3487_,data_stage_3__3486_,data_stage_3__3485_,
  data_stage_3__3484_,data_stage_3__3483_,data_stage_3__3482_,data_stage_3__3481_,
  data_stage_3__3480_,data_stage_3__3479_,data_stage_3__3478_,data_stage_3__3477_,
  data_stage_3__3476_,data_stage_3__3475_,data_stage_3__3474_,data_stage_3__3473_,
  data_stage_3__3472_,data_stage_3__3471_,data_stage_3__3470_,data_stage_3__3469_,
  data_stage_3__3468_,data_stage_3__3467_,data_stage_3__3466_,data_stage_3__3465_,
  data_stage_3__3464_,data_stage_3__3463_,data_stage_3__3462_,data_stage_3__3461_,
  data_stage_3__3460_,data_stage_3__3459_,data_stage_3__3458_,data_stage_3__3457_,
  data_stage_3__3456_,data_stage_3__3455_,data_stage_3__3454_,data_stage_3__3453_,
  data_stage_3__3452_,data_stage_3__3451_,data_stage_3__3450_,data_stage_3__3449_,
  data_stage_3__3448_,data_stage_3__3447_,data_stage_3__3446_,data_stage_3__3445_,
  data_stage_3__3444_,data_stage_3__3443_,data_stage_3__3442_,data_stage_3__3441_,
  data_stage_3__3440_,data_stage_3__3439_,data_stage_3__3438_,data_stage_3__3437_,
  data_stage_3__3436_,data_stage_3__3435_,data_stage_3__3434_,data_stage_3__3433_,
  data_stage_3__3432_,data_stage_3__3431_,data_stage_3__3430_,data_stage_3__3429_,
  data_stage_3__3428_,data_stage_3__3427_,data_stage_3__3426_,data_stage_3__3425_,
  data_stage_3__3424_,data_stage_3__3423_,data_stage_3__3422_,data_stage_3__3421_,
  data_stage_3__3420_,data_stage_3__3419_,data_stage_3__3418_,data_stage_3__3417_,
  data_stage_3__3416_,data_stage_3__3415_,data_stage_3__3414_,data_stage_3__3413_,
  data_stage_3__3412_,data_stage_3__3411_,data_stage_3__3410_,data_stage_3__3409_,
  data_stage_3__3408_,data_stage_3__3407_,data_stage_3__3406_,data_stage_3__3405_,
  data_stage_3__3404_,data_stage_3__3403_,data_stage_3__3402_,data_stage_3__3401_,
  data_stage_3__3400_,data_stage_3__3399_,data_stage_3__3398_,data_stage_3__3397_,
  data_stage_3__3396_,data_stage_3__3395_,data_stage_3__3394_,data_stage_3__3393_,
  data_stage_3__3392_,data_stage_3__3391_,data_stage_3__3390_,data_stage_3__3389_,
  data_stage_3__3388_,data_stage_3__3387_,data_stage_3__3386_,data_stage_3__3385_,
  data_stage_3__3384_,data_stage_3__3383_,data_stage_3__3382_,data_stage_3__3381_,
  data_stage_3__3380_,data_stage_3__3379_,data_stage_3__3378_,data_stage_3__3377_,
  data_stage_3__3376_,data_stage_3__3375_,data_stage_3__3374_,data_stage_3__3373_,
  data_stage_3__3372_,data_stage_3__3371_,data_stage_3__3370_,data_stage_3__3369_,
  data_stage_3__3368_,data_stage_3__3367_,data_stage_3__3366_,data_stage_3__3365_,
  data_stage_3__3364_,data_stage_3__3363_,data_stage_3__3362_,data_stage_3__3361_,
  data_stage_3__3360_,data_stage_3__3359_,data_stage_3__3358_,data_stage_3__3357_,
  data_stage_3__3356_,data_stage_3__3355_,data_stage_3__3354_,data_stage_3__3353_,
  data_stage_3__3352_,data_stage_3__3351_,data_stage_3__3350_,data_stage_3__3349_,
  data_stage_3__3348_,data_stage_3__3347_,data_stage_3__3346_,data_stage_3__3345_,
  data_stage_3__3344_,data_stage_3__3343_,data_stage_3__3342_,data_stage_3__3341_,
  data_stage_3__3340_,data_stage_3__3339_,data_stage_3__3338_,data_stage_3__3337_,
  data_stage_3__3336_,data_stage_3__3335_,data_stage_3__3334_,data_stage_3__3333_,
  data_stage_3__3332_,data_stage_3__3331_,data_stage_3__3330_,data_stage_3__3329_,
  data_stage_3__3328_,data_stage_3__3327_,data_stage_3__3326_,data_stage_3__3325_,
  data_stage_3__3324_,data_stage_3__3323_,data_stage_3__3322_,data_stage_3__3321_,
  data_stage_3__3320_,data_stage_3__3319_,data_stage_3__3318_,data_stage_3__3317_,
  data_stage_3__3316_,data_stage_3__3315_,data_stage_3__3314_,data_stage_3__3313_,
  data_stage_3__3312_,data_stage_3__3311_,data_stage_3__3310_,data_stage_3__3309_,
  data_stage_3__3308_,data_stage_3__3307_,data_stage_3__3306_,data_stage_3__3305_,
  data_stage_3__3304_,data_stage_3__3303_,data_stage_3__3302_,data_stage_3__3301_,
  data_stage_3__3300_,data_stage_3__3299_,data_stage_3__3298_,data_stage_3__3297_,
  data_stage_3__3296_,data_stage_3__3295_,data_stage_3__3294_,data_stage_3__3293_,
  data_stage_3__3292_,data_stage_3__3291_,data_stage_3__3290_,data_stage_3__3289_,
  data_stage_3__3288_,data_stage_3__3287_,data_stage_3__3286_,data_stage_3__3285_,
  data_stage_3__3284_,data_stage_3__3283_,data_stage_3__3282_,data_stage_3__3281_,
  data_stage_3__3280_,data_stage_3__3279_,data_stage_3__3278_,data_stage_3__3277_,
  data_stage_3__3276_,data_stage_3__3275_,data_stage_3__3274_,data_stage_3__3273_,
  data_stage_3__3272_,data_stage_3__3271_,data_stage_3__3270_,data_stage_3__3269_,
  data_stage_3__3268_,data_stage_3__3267_,data_stage_3__3266_,data_stage_3__3265_,
  data_stage_3__3264_,data_stage_3__3263_,data_stage_3__3262_,data_stage_3__3261_,
  data_stage_3__3260_,data_stage_3__3259_,data_stage_3__3258_,data_stage_3__3257_,
  data_stage_3__3256_,data_stage_3__3255_,data_stage_3__3254_,data_stage_3__3253_,
  data_stage_3__3252_,data_stage_3__3251_,data_stage_3__3250_,data_stage_3__3249_,
  data_stage_3__3248_,data_stage_3__3247_,data_stage_3__3246_,data_stage_3__3245_,
  data_stage_3__3244_,data_stage_3__3243_,data_stage_3__3242_,data_stage_3__3241_,
  data_stage_3__3240_,data_stage_3__3239_,data_stage_3__3238_,data_stage_3__3237_,
  data_stage_3__3236_,data_stage_3__3235_,data_stage_3__3234_,data_stage_3__3233_,
  data_stage_3__3232_,data_stage_3__3231_,data_stage_3__3230_,data_stage_3__3229_,
  data_stage_3__3228_,data_stage_3__3227_,data_stage_3__3226_,data_stage_3__3225_,
  data_stage_3__3224_,data_stage_3__3223_,data_stage_3__3222_,data_stage_3__3221_,
  data_stage_3__3220_,data_stage_3__3219_,data_stage_3__3218_,data_stage_3__3217_,
  data_stage_3__3216_,data_stage_3__3215_,data_stage_3__3214_,data_stage_3__3213_,
  data_stage_3__3212_,data_stage_3__3211_,data_stage_3__3210_,data_stage_3__3209_,
  data_stage_3__3208_,data_stage_3__3207_,data_stage_3__3206_,data_stage_3__3205_,
  data_stage_3__3204_,data_stage_3__3203_,data_stage_3__3202_,data_stage_3__3201_,
  data_stage_3__3200_,data_stage_3__3199_,data_stage_3__3198_,data_stage_3__3197_,
  data_stage_3__3196_,data_stage_3__3195_,data_stage_3__3194_,data_stage_3__3193_,
  data_stage_3__3192_,data_stage_3__3191_,data_stage_3__3190_,data_stage_3__3189_,
  data_stage_3__3188_,data_stage_3__3187_,data_stage_3__3186_,data_stage_3__3185_,
  data_stage_3__3184_,data_stage_3__3183_,data_stage_3__3182_,data_stage_3__3181_,
  data_stage_3__3180_,data_stage_3__3179_,data_stage_3__3178_,data_stage_3__3177_,
  data_stage_3__3176_,data_stage_3__3175_,data_stage_3__3174_,data_stage_3__3173_,
  data_stage_3__3172_,data_stage_3__3171_,data_stage_3__3170_,data_stage_3__3169_,
  data_stage_3__3168_,data_stage_3__3167_,data_stage_3__3166_,data_stage_3__3165_,
  data_stage_3__3164_,data_stage_3__3163_,data_stage_3__3162_,data_stage_3__3161_,
  data_stage_3__3160_,data_stage_3__3159_,data_stage_3__3158_,data_stage_3__3157_,
  data_stage_3__3156_,data_stage_3__3155_,data_stage_3__3154_,data_stage_3__3153_,
  data_stage_3__3152_,data_stage_3__3151_,data_stage_3__3150_,data_stage_3__3149_,
  data_stage_3__3148_,data_stage_3__3147_,data_stage_3__3146_,data_stage_3__3145_,
  data_stage_3__3144_,data_stage_3__3143_,data_stage_3__3142_,data_stage_3__3141_,
  data_stage_3__3140_,data_stage_3__3139_,data_stage_3__3138_,data_stage_3__3137_,
  data_stage_3__3136_,data_stage_3__3135_,data_stage_3__3134_,data_stage_3__3133_,
  data_stage_3__3132_,data_stage_3__3131_,data_stage_3__3130_,data_stage_3__3129_,
  data_stage_3__3128_,data_stage_3__3127_,data_stage_3__3126_,data_stage_3__3125_,
  data_stage_3__3124_,data_stage_3__3123_,data_stage_3__3122_,data_stage_3__3121_,
  data_stage_3__3120_,data_stage_3__3119_,data_stage_3__3118_,data_stage_3__3117_,
  data_stage_3__3116_,data_stage_3__3115_,data_stage_3__3114_,data_stage_3__3113_,
  data_stage_3__3112_,data_stage_3__3111_,data_stage_3__3110_,data_stage_3__3109_,
  data_stage_3__3108_,data_stage_3__3107_,data_stage_3__3106_,data_stage_3__3105_,
  data_stage_3__3104_,data_stage_3__3103_,data_stage_3__3102_,data_stage_3__3101_,
  data_stage_3__3100_,data_stage_3__3099_,data_stage_3__3098_,data_stage_3__3097_,
  data_stage_3__3096_,data_stage_3__3095_,data_stage_3__3094_,data_stage_3__3093_,
  data_stage_3__3092_,data_stage_3__3091_,data_stage_3__3090_,data_stage_3__3089_,
  data_stage_3__3088_,data_stage_3__3087_,data_stage_3__3086_,data_stage_3__3085_,
  data_stage_3__3084_,data_stage_3__3083_,data_stage_3__3082_,data_stage_3__3081_,
  data_stage_3__3080_,data_stage_3__3079_,data_stage_3__3078_,data_stage_3__3077_,
  data_stage_3__3076_,data_stage_3__3075_,data_stage_3__3074_,data_stage_3__3073_,
  data_stage_3__3072_,data_stage_3__3071_,data_stage_3__3070_,data_stage_3__3069_,
  data_stage_3__3068_,data_stage_3__3067_,data_stage_3__3066_,data_stage_3__3065_,
  data_stage_3__3064_,data_stage_3__3063_,data_stage_3__3062_,data_stage_3__3061_,
  data_stage_3__3060_,data_stage_3__3059_,data_stage_3__3058_,data_stage_3__3057_,
  data_stage_3__3056_,data_stage_3__3055_,data_stage_3__3054_,data_stage_3__3053_,
  data_stage_3__3052_,data_stage_3__3051_,data_stage_3__3050_,data_stage_3__3049_,
  data_stage_3__3048_,data_stage_3__3047_,data_stage_3__3046_,data_stage_3__3045_,
  data_stage_3__3044_,data_stage_3__3043_,data_stage_3__3042_,data_stage_3__3041_,
  data_stage_3__3040_,data_stage_3__3039_,data_stage_3__3038_,data_stage_3__3037_,
  data_stage_3__3036_,data_stage_3__3035_,data_stage_3__3034_,data_stage_3__3033_,
  data_stage_3__3032_,data_stage_3__3031_,data_stage_3__3030_,data_stage_3__3029_,
  data_stage_3__3028_,data_stage_3__3027_,data_stage_3__3026_,data_stage_3__3025_,
  data_stage_3__3024_,data_stage_3__3023_,data_stage_3__3022_,data_stage_3__3021_,
  data_stage_3__3020_,data_stage_3__3019_,data_stage_3__3018_,data_stage_3__3017_,
  data_stage_3__3016_,data_stage_3__3015_,data_stage_3__3014_,data_stage_3__3013_,
  data_stage_3__3012_,data_stage_3__3011_,data_stage_3__3010_,data_stage_3__3009_,
  data_stage_3__3008_,data_stage_3__3007_,data_stage_3__3006_,data_stage_3__3005_,
  data_stage_3__3004_,data_stage_3__3003_,data_stage_3__3002_,data_stage_3__3001_,
  data_stage_3__3000_,data_stage_3__2999_,data_stage_3__2998_,data_stage_3__2997_,
  data_stage_3__2996_,data_stage_3__2995_,data_stage_3__2994_,data_stage_3__2993_,
  data_stage_3__2992_,data_stage_3__2991_,data_stage_3__2990_,data_stage_3__2989_,
  data_stage_3__2988_,data_stage_3__2987_,data_stage_3__2986_,data_stage_3__2985_,
  data_stage_3__2984_,data_stage_3__2983_,data_stage_3__2982_,data_stage_3__2981_,
  data_stage_3__2980_,data_stage_3__2979_,data_stage_3__2978_,data_stage_3__2977_,
  data_stage_3__2976_,data_stage_3__2975_,data_stage_3__2974_,data_stage_3__2973_,
  data_stage_3__2972_,data_stage_3__2971_,data_stage_3__2970_,data_stage_3__2969_,
  data_stage_3__2968_,data_stage_3__2967_,data_stage_3__2966_,data_stage_3__2965_,
  data_stage_3__2964_,data_stage_3__2963_,data_stage_3__2962_,data_stage_3__2961_,
  data_stage_3__2960_,data_stage_3__2959_,data_stage_3__2958_,data_stage_3__2957_,
  data_stage_3__2956_,data_stage_3__2955_,data_stage_3__2954_,data_stage_3__2953_,
  data_stage_3__2952_,data_stage_3__2951_,data_stage_3__2950_,data_stage_3__2949_,
  data_stage_3__2948_,data_stage_3__2947_,data_stage_3__2946_,data_stage_3__2945_,
  data_stage_3__2944_,data_stage_3__2943_,data_stage_3__2942_,data_stage_3__2941_,
  data_stage_3__2940_,data_stage_3__2939_,data_stage_3__2938_,data_stage_3__2937_,
  data_stage_3__2936_,data_stage_3__2935_,data_stage_3__2934_,data_stage_3__2933_,
  data_stage_3__2932_,data_stage_3__2931_,data_stage_3__2930_,data_stage_3__2929_,
  data_stage_3__2928_,data_stage_3__2927_,data_stage_3__2926_,data_stage_3__2925_,
  data_stage_3__2924_,data_stage_3__2923_,data_stage_3__2922_,data_stage_3__2921_,
  data_stage_3__2920_,data_stage_3__2919_,data_stage_3__2918_,data_stage_3__2917_,
  data_stage_3__2916_,data_stage_3__2915_,data_stage_3__2914_,data_stage_3__2913_,
  data_stage_3__2912_,data_stage_3__2911_,data_stage_3__2910_,data_stage_3__2909_,
  data_stage_3__2908_,data_stage_3__2907_,data_stage_3__2906_,data_stage_3__2905_,
  data_stage_3__2904_,data_stage_3__2903_,data_stage_3__2902_,data_stage_3__2901_,
  data_stage_3__2900_,data_stage_3__2899_,data_stage_3__2898_,data_stage_3__2897_,
  data_stage_3__2896_,data_stage_3__2895_,data_stage_3__2894_,data_stage_3__2893_,
  data_stage_3__2892_,data_stage_3__2891_,data_stage_3__2890_,data_stage_3__2889_,
  data_stage_3__2888_,data_stage_3__2887_,data_stage_3__2886_,data_stage_3__2885_,
  data_stage_3__2884_,data_stage_3__2883_,data_stage_3__2882_,data_stage_3__2881_,
  data_stage_3__2880_,data_stage_3__2879_,data_stage_3__2878_,data_stage_3__2877_,
  data_stage_3__2876_,data_stage_3__2875_,data_stage_3__2874_,data_stage_3__2873_,
  data_stage_3__2872_,data_stage_3__2871_,data_stage_3__2870_,data_stage_3__2869_,
  data_stage_3__2868_,data_stage_3__2867_,data_stage_3__2866_,data_stage_3__2865_,
  data_stage_3__2864_,data_stage_3__2863_,data_stage_3__2862_,data_stage_3__2861_,
  data_stage_3__2860_,data_stage_3__2859_,data_stage_3__2858_,data_stage_3__2857_,
  data_stage_3__2856_,data_stage_3__2855_,data_stage_3__2854_,data_stage_3__2853_,
  data_stage_3__2852_,data_stage_3__2851_,data_stage_3__2850_,data_stage_3__2849_,
  data_stage_3__2848_,data_stage_3__2847_,data_stage_3__2846_,data_stage_3__2845_,
  data_stage_3__2844_,data_stage_3__2843_,data_stage_3__2842_,data_stage_3__2841_,
  data_stage_3__2840_,data_stage_3__2839_,data_stage_3__2838_,data_stage_3__2837_,
  data_stage_3__2836_,data_stage_3__2835_,data_stage_3__2834_,data_stage_3__2833_,
  data_stage_3__2832_,data_stage_3__2831_,data_stage_3__2830_,data_stage_3__2829_,
  data_stage_3__2828_,data_stage_3__2827_,data_stage_3__2826_,data_stage_3__2825_,
  data_stage_3__2824_,data_stage_3__2823_,data_stage_3__2822_,data_stage_3__2821_,
  data_stage_3__2820_,data_stage_3__2819_,data_stage_3__2818_,data_stage_3__2817_,
  data_stage_3__2816_,data_stage_3__2815_,data_stage_3__2814_,data_stage_3__2813_,
  data_stage_3__2812_,data_stage_3__2811_,data_stage_3__2810_,data_stage_3__2809_,
  data_stage_3__2808_,data_stage_3__2807_,data_stage_3__2806_,data_stage_3__2805_,
  data_stage_3__2804_,data_stage_3__2803_,data_stage_3__2802_,data_stage_3__2801_,
  data_stage_3__2800_,data_stage_3__2799_,data_stage_3__2798_,data_stage_3__2797_,
  data_stage_3__2796_,data_stage_3__2795_,data_stage_3__2794_,data_stage_3__2793_,
  data_stage_3__2792_,data_stage_3__2791_,data_stage_3__2790_,data_stage_3__2789_,
  data_stage_3__2788_,data_stage_3__2787_,data_stage_3__2786_,data_stage_3__2785_,
  data_stage_3__2784_,data_stage_3__2783_,data_stage_3__2782_,data_stage_3__2781_,
  data_stage_3__2780_,data_stage_3__2779_,data_stage_3__2778_,data_stage_3__2777_,
  data_stage_3__2776_,data_stage_3__2775_,data_stage_3__2774_,data_stage_3__2773_,
  data_stage_3__2772_,data_stage_3__2771_,data_stage_3__2770_,data_stage_3__2769_,
  data_stage_3__2768_,data_stage_3__2767_,data_stage_3__2766_,data_stage_3__2765_,
  data_stage_3__2764_,data_stage_3__2763_,data_stage_3__2762_,data_stage_3__2761_,
  data_stage_3__2760_,data_stage_3__2759_,data_stage_3__2758_,data_stage_3__2757_,
  data_stage_3__2756_,data_stage_3__2755_,data_stage_3__2754_,data_stage_3__2753_,
  data_stage_3__2752_,data_stage_3__2751_,data_stage_3__2750_,data_stage_3__2749_,
  data_stage_3__2748_,data_stage_3__2747_,data_stage_3__2746_,data_stage_3__2745_,
  data_stage_3__2744_,data_stage_3__2743_,data_stage_3__2742_,data_stage_3__2741_,
  data_stage_3__2740_,data_stage_3__2739_,data_stage_3__2738_,data_stage_3__2737_,
  data_stage_3__2736_,data_stage_3__2735_,data_stage_3__2734_,data_stage_3__2733_,
  data_stage_3__2732_,data_stage_3__2731_,data_stage_3__2730_,data_stage_3__2729_,
  data_stage_3__2728_,data_stage_3__2727_,data_stage_3__2726_,data_stage_3__2725_,
  data_stage_3__2724_,data_stage_3__2723_,data_stage_3__2722_,data_stage_3__2721_,
  data_stage_3__2720_,data_stage_3__2719_,data_stage_3__2718_,data_stage_3__2717_,
  data_stage_3__2716_,data_stage_3__2715_,data_stage_3__2714_,data_stage_3__2713_,
  data_stage_3__2712_,data_stage_3__2711_,data_stage_3__2710_,data_stage_3__2709_,
  data_stage_3__2708_,data_stage_3__2707_,data_stage_3__2706_,data_stage_3__2705_,
  data_stage_3__2704_,data_stage_3__2703_,data_stage_3__2702_,data_stage_3__2701_,
  data_stage_3__2700_,data_stage_3__2699_,data_stage_3__2698_,data_stage_3__2697_,
  data_stage_3__2696_,data_stage_3__2695_,data_stage_3__2694_,data_stage_3__2693_,
  data_stage_3__2692_,data_stage_3__2691_,data_stage_3__2690_,data_stage_3__2689_,
  data_stage_3__2688_,data_stage_3__2687_,data_stage_3__2686_,data_stage_3__2685_,
  data_stage_3__2684_,data_stage_3__2683_,data_stage_3__2682_,data_stage_3__2681_,
  data_stage_3__2680_,data_stage_3__2679_,data_stage_3__2678_,data_stage_3__2677_,
  data_stage_3__2676_,data_stage_3__2675_,data_stage_3__2674_,data_stage_3__2673_,
  data_stage_3__2672_,data_stage_3__2671_,data_stage_3__2670_,data_stage_3__2669_,
  data_stage_3__2668_,data_stage_3__2667_,data_stage_3__2666_,data_stage_3__2665_,
  data_stage_3__2664_,data_stage_3__2663_,data_stage_3__2662_,data_stage_3__2661_,
  data_stage_3__2660_,data_stage_3__2659_,data_stage_3__2658_,data_stage_3__2657_,
  data_stage_3__2656_,data_stage_3__2655_,data_stage_3__2654_,data_stage_3__2653_,
  data_stage_3__2652_,data_stage_3__2651_,data_stage_3__2650_,data_stage_3__2649_,
  data_stage_3__2648_,data_stage_3__2647_,data_stage_3__2646_,data_stage_3__2645_,
  data_stage_3__2644_,data_stage_3__2643_,data_stage_3__2642_,data_stage_3__2641_,
  data_stage_3__2640_,data_stage_3__2639_,data_stage_3__2638_,data_stage_3__2637_,
  data_stage_3__2636_,data_stage_3__2635_,data_stage_3__2634_,data_stage_3__2633_,
  data_stage_3__2632_,data_stage_3__2631_,data_stage_3__2630_,data_stage_3__2629_,
  data_stage_3__2628_,data_stage_3__2627_,data_stage_3__2626_,data_stage_3__2625_,
  data_stage_3__2624_,data_stage_3__2623_,data_stage_3__2622_,data_stage_3__2621_,
  data_stage_3__2620_,data_stage_3__2619_,data_stage_3__2618_,data_stage_3__2617_,
  data_stage_3__2616_,data_stage_3__2615_,data_stage_3__2614_,data_stage_3__2613_,
  data_stage_3__2612_,data_stage_3__2611_,data_stage_3__2610_,data_stage_3__2609_,
  data_stage_3__2608_,data_stage_3__2607_,data_stage_3__2606_,data_stage_3__2605_,
  data_stage_3__2604_,data_stage_3__2603_,data_stage_3__2602_,data_stage_3__2601_,
  data_stage_3__2600_,data_stage_3__2599_,data_stage_3__2598_,data_stage_3__2597_,
  data_stage_3__2596_,data_stage_3__2595_,data_stage_3__2594_,data_stage_3__2593_,
  data_stage_3__2592_,data_stage_3__2591_,data_stage_3__2590_,data_stage_3__2589_,
  data_stage_3__2588_,data_stage_3__2587_,data_stage_3__2586_,data_stage_3__2585_,
  data_stage_3__2584_,data_stage_3__2583_,data_stage_3__2582_,data_stage_3__2581_,
  data_stage_3__2580_,data_stage_3__2579_,data_stage_3__2578_,data_stage_3__2577_,
  data_stage_3__2576_,data_stage_3__2575_,data_stage_3__2574_,data_stage_3__2573_,
  data_stage_3__2572_,data_stage_3__2571_,data_stage_3__2570_,data_stage_3__2569_,
  data_stage_3__2568_,data_stage_3__2567_,data_stage_3__2566_,data_stage_3__2565_,
  data_stage_3__2564_,data_stage_3__2563_,data_stage_3__2562_,data_stage_3__2561_,
  data_stage_3__2560_,data_stage_3__2559_,data_stage_3__2558_,data_stage_3__2557_,
  data_stage_3__2556_,data_stage_3__2555_,data_stage_3__2554_,data_stage_3__2553_,
  data_stage_3__2552_,data_stage_3__2551_,data_stage_3__2550_,data_stage_3__2549_,
  data_stage_3__2548_,data_stage_3__2547_,data_stage_3__2546_,data_stage_3__2545_,
  data_stage_3__2544_,data_stage_3__2543_,data_stage_3__2542_,data_stage_3__2541_,
  data_stage_3__2540_,data_stage_3__2539_,data_stage_3__2538_,data_stage_3__2537_,
  data_stage_3__2536_,data_stage_3__2535_,data_stage_3__2534_,data_stage_3__2533_,
  data_stage_3__2532_,data_stage_3__2531_,data_stage_3__2530_,data_stage_3__2529_,
  data_stage_3__2528_,data_stage_3__2527_,data_stage_3__2526_,data_stage_3__2525_,
  data_stage_3__2524_,data_stage_3__2523_,data_stage_3__2522_,data_stage_3__2521_,
  data_stage_3__2520_,data_stage_3__2519_,data_stage_3__2518_,data_stage_3__2517_,
  data_stage_3__2516_,data_stage_3__2515_,data_stage_3__2514_,data_stage_3__2513_,
  data_stage_3__2512_,data_stage_3__2511_,data_stage_3__2510_,data_stage_3__2509_,
  data_stage_3__2508_,data_stage_3__2507_,data_stage_3__2506_,data_stage_3__2505_,
  data_stage_3__2504_,data_stage_3__2503_,data_stage_3__2502_,data_stage_3__2501_,
  data_stage_3__2500_,data_stage_3__2499_,data_stage_3__2498_,data_stage_3__2497_,
  data_stage_3__2496_,data_stage_3__2495_,data_stage_3__2494_,data_stage_3__2493_,
  data_stage_3__2492_,data_stage_3__2491_,data_stage_3__2490_,data_stage_3__2489_,
  data_stage_3__2488_,data_stage_3__2487_,data_stage_3__2486_,data_stage_3__2485_,
  data_stage_3__2484_,data_stage_3__2483_,data_stage_3__2482_,data_stage_3__2481_,
  data_stage_3__2480_,data_stage_3__2479_,data_stage_3__2478_,data_stage_3__2477_,
  data_stage_3__2476_,data_stage_3__2475_,data_stage_3__2474_,data_stage_3__2473_,
  data_stage_3__2472_,data_stage_3__2471_,data_stage_3__2470_,data_stage_3__2469_,
  data_stage_3__2468_,data_stage_3__2467_,data_stage_3__2466_,data_stage_3__2465_,
  data_stage_3__2464_,data_stage_3__2463_,data_stage_3__2462_,data_stage_3__2461_,
  data_stage_3__2460_,data_stage_3__2459_,data_stage_3__2458_,data_stage_3__2457_,
  data_stage_3__2456_,data_stage_3__2455_,data_stage_3__2454_,data_stage_3__2453_,
  data_stage_3__2452_,data_stage_3__2451_,data_stage_3__2450_,data_stage_3__2449_,
  data_stage_3__2448_,data_stage_3__2447_,data_stage_3__2446_,data_stage_3__2445_,
  data_stage_3__2444_,data_stage_3__2443_,data_stage_3__2442_,data_stage_3__2441_,
  data_stage_3__2440_,data_stage_3__2439_,data_stage_3__2438_,data_stage_3__2437_,
  data_stage_3__2436_,data_stage_3__2435_,data_stage_3__2434_,data_stage_3__2433_,
  data_stage_3__2432_,data_stage_3__2431_,data_stage_3__2430_,data_stage_3__2429_,
  data_stage_3__2428_,data_stage_3__2427_,data_stage_3__2426_,data_stage_3__2425_,
  data_stage_3__2424_,data_stage_3__2423_,data_stage_3__2422_,data_stage_3__2421_,
  data_stage_3__2420_,data_stage_3__2419_,data_stage_3__2418_,data_stage_3__2417_,
  data_stage_3__2416_,data_stage_3__2415_,data_stage_3__2414_,data_stage_3__2413_,
  data_stage_3__2412_,data_stage_3__2411_,data_stage_3__2410_,data_stage_3__2409_,
  data_stage_3__2408_,data_stage_3__2407_,data_stage_3__2406_,data_stage_3__2405_,
  data_stage_3__2404_,data_stage_3__2403_,data_stage_3__2402_,data_stage_3__2401_,
  data_stage_3__2400_,data_stage_3__2399_,data_stage_3__2398_,data_stage_3__2397_,
  data_stage_3__2396_,data_stage_3__2395_,data_stage_3__2394_,data_stage_3__2393_,
  data_stage_3__2392_,data_stage_3__2391_,data_stage_3__2390_,data_stage_3__2389_,
  data_stage_3__2388_,data_stage_3__2387_,data_stage_3__2386_,data_stage_3__2385_,
  data_stage_3__2384_,data_stage_3__2383_,data_stage_3__2382_,data_stage_3__2381_,
  data_stage_3__2380_,data_stage_3__2379_,data_stage_3__2378_,data_stage_3__2377_,
  data_stage_3__2376_,data_stage_3__2375_,data_stage_3__2374_,data_stage_3__2373_,
  data_stage_3__2372_,data_stage_3__2371_,data_stage_3__2370_,data_stage_3__2369_,
  data_stage_3__2368_,data_stage_3__2367_,data_stage_3__2366_,data_stage_3__2365_,
  data_stage_3__2364_,data_stage_3__2363_,data_stage_3__2362_,data_stage_3__2361_,
  data_stage_3__2360_,data_stage_3__2359_,data_stage_3__2358_,data_stage_3__2357_,
  data_stage_3__2356_,data_stage_3__2355_,data_stage_3__2354_,data_stage_3__2353_,
  data_stage_3__2352_,data_stage_3__2351_,data_stage_3__2350_,data_stage_3__2349_,
  data_stage_3__2348_,data_stage_3__2347_,data_stage_3__2346_,data_stage_3__2345_,
  data_stage_3__2344_,data_stage_3__2343_,data_stage_3__2342_,data_stage_3__2341_,
  data_stage_3__2340_,data_stage_3__2339_,data_stage_3__2338_,data_stage_3__2337_,
  data_stage_3__2336_,data_stage_3__2335_,data_stage_3__2334_,data_stage_3__2333_,
  data_stage_3__2332_,data_stage_3__2331_,data_stage_3__2330_,data_stage_3__2329_,
  data_stage_3__2328_,data_stage_3__2327_,data_stage_3__2326_,data_stage_3__2325_,
  data_stage_3__2324_,data_stage_3__2323_,data_stage_3__2322_,data_stage_3__2321_,
  data_stage_3__2320_,data_stage_3__2319_,data_stage_3__2318_,data_stage_3__2317_,
  data_stage_3__2316_,data_stage_3__2315_,data_stage_3__2314_,data_stage_3__2313_,
  data_stage_3__2312_,data_stage_3__2311_,data_stage_3__2310_,data_stage_3__2309_,
  data_stage_3__2308_,data_stage_3__2307_,data_stage_3__2306_,data_stage_3__2305_,
  data_stage_3__2304_,data_stage_3__2303_,data_stage_3__2302_,data_stage_3__2301_,
  data_stage_3__2300_,data_stage_3__2299_,data_stage_3__2298_,data_stage_3__2297_,
  data_stage_3__2296_,data_stage_3__2295_,data_stage_3__2294_,data_stage_3__2293_,
  data_stage_3__2292_,data_stage_3__2291_,data_stage_3__2290_,data_stage_3__2289_,
  data_stage_3__2288_,data_stage_3__2287_,data_stage_3__2286_,data_stage_3__2285_,
  data_stage_3__2284_,data_stage_3__2283_,data_stage_3__2282_,data_stage_3__2281_,
  data_stage_3__2280_,data_stage_3__2279_,data_stage_3__2278_,data_stage_3__2277_,
  data_stage_3__2276_,data_stage_3__2275_,data_stage_3__2274_,data_stage_3__2273_,
  data_stage_3__2272_,data_stage_3__2271_,data_stage_3__2270_,data_stage_3__2269_,
  data_stage_3__2268_,data_stage_3__2267_,data_stage_3__2266_,data_stage_3__2265_,
  data_stage_3__2264_,data_stage_3__2263_,data_stage_3__2262_,data_stage_3__2261_,
  data_stage_3__2260_,data_stage_3__2259_,data_stage_3__2258_,data_stage_3__2257_,
  data_stage_3__2256_,data_stage_3__2255_,data_stage_3__2254_,data_stage_3__2253_,
  data_stage_3__2252_,data_stage_3__2251_,data_stage_3__2250_,data_stage_3__2249_,
  data_stage_3__2248_,data_stage_3__2247_,data_stage_3__2246_,data_stage_3__2245_,
  data_stage_3__2244_,data_stage_3__2243_,data_stage_3__2242_,data_stage_3__2241_,
  data_stage_3__2240_,data_stage_3__2239_,data_stage_3__2238_,data_stage_3__2237_,
  data_stage_3__2236_,data_stage_3__2235_,data_stage_3__2234_,data_stage_3__2233_,
  data_stage_3__2232_,data_stage_3__2231_,data_stage_3__2230_,data_stage_3__2229_,
  data_stage_3__2228_,data_stage_3__2227_,data_stage_3__2226_,data_stage_3__2225_,
  data_stage_3__2224_,data_stage_3__2223_,data_stage_3__2222_,data_stage_3__2221_,
  data_stage_3__2220_,data_stage_3__2219_,data_stage_3__2218_,data_stage_3__2217_,
  data_stage_3__2216_,data_stage_3__2215_,data_stage_3__2214_,data_stage_3__2213_,
  data_stage_3__2212_,data_stage_3__2211_,data_stage_3__2210_,data_stage_3__2209_,
  data_stage_3__2208_,data_stage_3__2207_,data_stage_3__2206_,data_stage_3__2205_,
  data_stage_3__2204_,data_stage_3__2203_,data_stage_3__2202_,data_stage_3__2201_,
  data_stage_3__2200_,data_stage_3__2199_,data_stage_3__2198_,data_stage_3__2197_,
  data_stage_3__2196_,data_stage_3__2195_,data_stage_3__2194_,data_stage_3__2193_,
  data_stage_3__2192_,data_stage_3__2191_,data_stage_3__2190_,data_stage_3__2189_,
  data_stage_3__2188_,data_stage_3__2187_,data_stage_3__2186_,data_stage_3__2185_,
  data_stage_3__2184_,data_stage_3__2183_,data_stage_3__2182_,data_stage_3__2181_,
  data_stage_3__2180_,data_stage_3__2179_,data_stage_3__2178_,data_stage_3__2177_,
  data_stage_3__2176_,data_stage_3__2175_,data_stage_3__2174_,data_stage_3__2173_,
  data_stage_3__2172_,data_stage_3__2171_,data_stage_3__2170_,data_stage_3__2169_,
  data_stage_3__2168_,data_stage_3__2167_,data_stage_3__2166_,data_stage_3__2165_,
  data_stage_3__2164_,data_stage_3__2163_,data_stage_3__2162_,data_stage_3__2161_,
  data_stage_3__2160_,data_stage_3__2159_,data_stage_3__2158_,data_stage_3__2157_,
  data_stage_3__2156_,data_stage_3__2155_,data_stage_3__2154_,data_stage_3__2153_,
  data_stage_3__2152_,data_stage_3__2151_,data_stage_3__2150_,data_stage_3__2149_,
  data_stage_3__2148_,data_stage_3__2147_,data_stage_3__2146_,data_stage_3__2145_,
  data_stage_3__2144_,data_stage_3__2143_,data_stage_3__2142_,data_stage_3__2141_,
  data_stage_3__2140_,data_stage_3__2139_,data_stage_3__2138_,data_stage_3__2137_,
  data_stage_3__2136_,data_stage_3__2135_,data_stage_3__2134_,data_stage_3__2133_,
  data_stage_3__2132_,data_stage_3__2131_,data_stage_3__2130_,data_stage_3__2129_,
  data_stage_3__2128_,data_stage_3__2127_,data_stage_3__2126_,data_stage_3__2125_,
  data_stage_3__2124_,data_stage_3__2123_,data_stage_3__2122_,data_stage_3__2121_,
  data_stage_3__2120_,data_stage_3__2119_,data_stage_3__2118_,data_stage_3__2117_,
  data_stage_3__2116_,data_stage_3__2115_,data_stage_3__2114_,data_stage_3__2113_,
  data_stage_3__2112_,data_stage_3__2111_,data_stage_3__2110_,data_stage_3__2109_,
  data_stage_3__2108_,data_stage_3__2107_,data_stage_3__2106_,data_stage_3__2105_,
  data_stage_3__2104_,data_stage_3__2103_,data_stage_3__2102_,data_stage_3__2101_,
  data_stage_3__2100_,data_stage_3__2099_,data_stage_3__2098_,data_stage_3__2097_,
  data_stage_3__2096_,data_stage_3__2095_,data_stage_3__2094_,data_stage_3__2093_,
  data_stage_3__2092_,data_stage_3__2091_,data_stage_3__2090_,data_stage_3__2089_,
  data_stage_3__2088_,data_stage_3__2087_,data_stage_3__2086_,data_stage_3__2085_,
  data_stage_3__2084_,data_stage_3__2083_,data_stage_3__2082_,data_stage_3__2081_,
  data_stage_3__2080_,data_stage_3__2079_,data_stage_3__2078_,data_stage_3__2077_,
  data_stage_3__2076_,data_stage_3__2075_,data_stage_3__2074_,data_stage_3__2073_,
  data_stage_3__2072_,data_stage_3__2071_,data_stage_3__2070_,data_stage_3__2069_,
  data_stage_3__2068_,data_stage_3__2067_,data_stage_3__2066_,data_stage_3__2065_,
  data_stage_3__2064_,data_stage_3__2063_,data_stage_3__2062_,data_stage_3__2061_,
  data_stage_3__2060_,data_stage_3__2059_,data_stage_3__2058_,data_stage_3__2057_,
  data_stage_3__2056_,data_stage_3__2055_,data_stage_3__2054_,data_stage_3__2053_,
  data_stage_3__2052_,data_stage_3__2051_,data_stage_3__2050_,data_stage_3__2049_,
  data_stage_3__2048_,data_stage_3__2047_,data_stage_3__2046_,data_stage_3__2045_,
  data_stage_3__2044_,data_stage_3__2043_,data_stage_3__2042_,data_stage_3__2041_,
  data_stage_3__2040_,data_stage_3__2039_,data_stage_3__2038_,data_stage_3__2037_,
  data_stage_3__2036_,data_stage_3__2035_,data_stage_3__2034_,data_stage_3__2033_,
  data_stage_3__2032_,data_stage_3__2031_,data_stage_3__2030_,data_stage_3__2029_,
  data_stage_3__2028_,data_stage_3__2027_,data_stage_3__2026_,data_stage_3__2025_,
  data_stage_3__2024_,data_stage_3__2023_,data_stage_3__2022_,data_stage_3__2021_,
  data_stage_3__2020_,data_stage_3__2019_,data_stage_3__2018_,data_stage_3__2017_,
  data_stage_3__2016_,data_stage_3__2015_,data_stage_3__2014_,data_stage_3__2013_,
  data_stage_3__2012_,data_stage_3__2011_,data_stage_3__2010_,data_stage_3__2009_,
  data_stage_3__2008_,data_stage_3__2007_,data_stage_3__2006_,data_stage_3__2005_,
  data_stage_3__2004_,data_stage_3__2003_,data_stage_3__2002_,data_stage_3__2001_,
  data_stage_3__2000_,data_stage_3__1999_,data_stage_3__1998_,data_stage_3__1997_,
  data_stage_3__1996_,data_stage_3__1995_,data_stage_3__1994_,data_stage_3__1993_,
  data_stage_3__1992_,data_stage_3__1991_,data_stage_3__1990_,data_stage_3__1989_,
  data_stage_3__1988_,data_stage_3__1987_,data_stage_3__1986_,data_stage_3__1985_,
  data_stage_3__1984_,data_stage_3__1983_,data_stage_3__1982_,data_stage_3__1981_,
  data_stage_3__1980_,data_stage_3__1979_,data_stage_3__1978_,data_stage_3__1977_,
  data_stage_3__1976_,data_stage_3__1975_,data_stage_3__1974_,data_stage_3__1973_,
  data_stage_3__1972_,data_stage_3__1971_,data_stage_3__1970_,data_stage_3__1969_,
  data_stage_3__1968_,data_stage_3__1967_,data_stage_3__1966_,data_stage_3__1965_,
  data_stage_3__1964_,data_stage_3__1963_,data_stage_3__1962_,data_stage_3__1961_,
  data_stage_3__1960_,data_stage_3__1959_,data_stage_3__1958_,data_stage_3__1957_,
  data_stage_3__1956_,data_stage_3__1955_,data_stage_3__1954_,data_stage_3__1953_,
  data_stage_3__1952_,data_stage_3__1951_,data_stage_3__1950_,data_stage_3__1949_,
  data_stage_3__1948_,data_stage_3__1947_,data_stage_3__1946_,data_stage_3__1945_,
  data_stage_3__1944_,data_stage_3__1943_,data_stage_3__1942_,data_stage_3__1941_,
  data_stage_3__1940_,data_stage_3__1939_,data_stage_3__1938_,data_stage_3__1937_,
  data_stage_3__1936_,data_stage_3__1935_,data_stage_3__1934_,data_stage_3__1933_,
  data_stage_3__1932_,data_stage_3__1931_,data_stage_3__1930_,data_stage_3__1929_,
  data_stage_3__1928_,data_stage_3__1927_,data_stage_3__1926_,data_stage_3__1925_,
  data_stage_3__1924_,data_stage_3__1923_,data_stage_3__1922_,data_stage_3__1921_,
  data_stage_3__1920_,data_stage_3__1919_,data_stage_3__1918_,data_stage_3__1917_,
  data_stage_3__1916_,data_stage_3__1915_,data_stage_3__1914_,data_stage_3__1913_,
  data_stage_3__1912_,data_stage_3__1911_,data_stage_3__1910_,data_stage_3__1909_,
  data_stage_3__1908_,data_stage_3__1907_,data_stage_3__1906_,data_stage_3__1905_,
  data_stage_3__1904_,data_stage_3__1903_,data_stage_3__1902_,data_stage_3__1901_,
  data_stage_3__1900_,data_stage_3__1899_,data_stage_3__1898_,data_stage_3__1897_,
  data_stage_3__1896_,data_stage_3__1895_,data_stage_3__1894_,data_stage_3__1893_,
  data_stage_3__1892_,data_stage_3__1891_,data_stage_3__1890_,data_stage_3__1889_,
  data_stage_3__1888_,data_stage_3__1887_,data_stage_3__1886_,data_stage_3__1885_,
  data_stage_3__1884_,data_stage_3__1883_,data_stage_3__1882_,data_stage_3__1881_,
  data_stage_3__1880_,data_stage_3__1879_,data_stage_3__1878_,data_stage_3__1877_,
  data_stage_3__1876_,data_stage_3__1875_,data_stage_3__1874_,data_stage_3__1873_,
  data_stage_3__1872_,data_stage_3__1871_,data_stage_3__1870_,data_stage_3__1869_,
  data_stage_3__1868_,data_stage_3__1867_,data_stage_3__1866_,data_stage_3__1865_,
  data_stage_3__1864_,data_stage_3__1863_,data_stage_3__1862_,data_stage_3__1861_,
  data_stage_3__1860_,data_stage_3__1859_,data_stage_3__1858_,data_stage_3__1857_,
  data_stage_3__1856_,data_stage_3__1855_,data_stage_3__1854_,data_stage_3__1853_,
  data_stage_3__1852_,data_stage_3__1851_,data_stage_3__1850_,data_stage_3__1849_,
  data_stage_3__1848_,data_stage_3__1847_,data_stage_3__1846_,data_stage_3__1845_,
  data_stage_3__1844_,data_stage_3__1843_,data_stage_3__1842_,data_stage_3__1841_,
  data_stage_3__1840_,data_stage_3__1839_,data_stage_3__1838_,data_stage_3__1837_,
  data_stage_3__1836_,data_stage_3__1835_,data_stage_3__1834_,data_stage_3__1833_,
  data_stage_3__1832_,data_stage_3__1831_,data_stage_3__1830_,data_stage_3__1829_,
  data_stage_3__1828_,data_stage_3__1827_,data_stage_3__1826_,data_stage_3__1825_,
  data_stage_3__1824_,data_stage_3__1823_,data_stage_3__1822_,data_stage_3__1821_,
  data_stage_3__1820_,data_stage_3__1819_,data_stage_3__1818_,data_stage_3__1817_,
  data_stage_3__1816_,data_stage_3__1815_,data_stage_3__1814_,data_stage_3__1813_,
  data_stage_3__1812_,data_stage_3__1811_,data_stage_3__1810_,data_stage_3__1809_,
  data_stage_3__1808_,data_stage_3__1807_,data_stage_3__1806_,data_stage_3__1805_,
  data_stage_3__1804_,data_stage_3__1803_,data_stage_3__1802_,data_stage_3__1801_,
  data_stage_3__1800_,data_stage_3__1799_,data_stage_3__1798_,data_stage_3__1797_,
  data_stage_3__1796_,data_stage_3__1795_,data_stage_3__1794_,data_stage_3__1793_,
  data_stage_3__1792_,data_stage_3__1791_,data_stage_3__1790_,data_stage_3__1789_,
  data_stage_3__1788_,data_stage_3__1787_,data_stage_3__1786_,data_stage_3__1785_,
  data_stage_3__1784_,data_stage_3__1783_,data_stage_3__1782_,data_stage_3__1781_,
  data_stage_3__1780_,data_stage_3__1779_,data_stage_3__1778_,data_stage_3__1777_,
  data_stage_3__1776_,data_stage_3__1775_,data_stage_3__1774_,data_stage_3__1773_,
  data_stage_3__1772_,data_stage_3__1771_,data_stage_3__1770_,data_stage_3__1769_,
  data_stage_3__1768_,data_stage_3__1767_,data_stage_3__1766_,data_stage_3__1765_,
  data_stage_3__1764_,data_stage_3__1763_,data_stage_3__1762_,data_stage_3__1761_,
  data_stage_3__1760_,data_stage_3__1759_,data_stage_3__1758_,data_stage_3__1757_,
  data_stage_3__1756_,data_stage_3__1755_,data_stage_3__1754_,data_stage_3__1753_,
  data_stage_3__1752_,data_stage_3__1751_,data_stage_3__1750_,data_stage_3__1749_,
  data_stage_3__1748_,data_stage_3__1747_,data_stage_3__1746_,data_stage_3__1745_,
  data_stage_3__1744_,data_stage_3__1743_,data_stage_3__1742_,data_stage_3__1741_,
  data_stage_3__1740_,data_stage_3__1739_,data_stage_3__1738_,data_stage_3__1737_,
  data_stage_3__1736_,data_stage_3__1735_,data_stage_3__1734_,data_stage_3__1733_,
  data_stage_3__1732_,data_stage_3__1731_,data_stage_3__1730_,data_stage_3__1729_,
  data_stage_3__1728_,data_stage_3__1727_,data_stage_3__1726_,data_stage_3__1725_,
  data_stage_3__1724_,data_stage_3__1723_,data_stage_3__1722_,data_stage_3__1721_,
  data_stage_3__1720_,data_stage_3__1719_,data_stage_3__1718_,data_stage_3__1717_,
  data_stage_3__1716_,data_stage_3__1715_,data_stage_3__1714_,data_stage_3__1713_,
  data_stage_3__1712_,data_stage_3__1711_,data_stage_3__1710_,data_stage_3__1709_,
  data_stage_3__1708_,data_stage_3__1707_,data_stage_3__1706_,data_stage_3__1705_,
  data_stage_3__1704_,data_stage_3__1703_,data_stage_3__1702_,data_stage_3__1701_,
  data_stage_3__1700_,data_stage_3__1699_,data_stage_3__1698_,data_stage_3__1697_,
  data_stage_3__1696_,data_stage_3__1695_,data_stage_3__1694_,data_stage_3__1693_,
  data_stage_3__1692_,data_stage_3__1691_,data_stage_3__1690_,data_stage_3__1689_,
  data_stage_3__1688_,data_stage_3__1687_,data_stage_3__1686_,data_stage_3__1685_,
  data_stage_3__1684_,data_stage_3__1683_,data_stage_3__1682_,data_stage_3__1681_,
  data_stage_3__1680_,data_stage_3__1679_,data_stage_3__1678_,data_stage_3__1677_,
  data_stage_3__1676_,data_stage_3__1675_,data_stage_3__1674_,data_stage_3__1673_,
  data_stage_3__1672_,data_stage_3__1671_,data_stage_3__1670_,data_stage_3__1669_,
  data_stage_3__1668_,data_stage_3__1667_,data_stage_3__1666_,data_stage_3__1665_,
  data_stage_3__1664_,data_stage_3__1663_,data_stage_3__1662_,data_stage_3__1661_,
  data_stage_3__1660_,data_stage_3__1659_,data_stage_3__1658_,data_stage_3__1657_,
  data_stage_3__1656_,data_stage_3__1655_,data_stage_3__1654_,data_stage_3__1653_,
  data_stage_3__1652_,data_stage_3__1651_,data_stage_3__1650_,data_stage_3__1649_,
  data_stage_3__1648_,data_stage_3__1647_,data_stage_3__1646_,data_stage_3__1645_,
  data_stage_3__1644_,data_stage_3__1643_,data_stage_3__1642_,data_stage_3__1641_,
  data_stage_3__1640_,data_stage_3__1639_,data_stage_3__1638_,data_stage_3__1637_,
  data_stage_3__1636_,data_stage_3__1635_,data_stage_3__1634_,data_stage_3__1633_,
  data_stage_3__1632_,data_stage_3__1631_,data_stage_3__1630_,data_stage_3__1629_,
  data_stage_3__1628_,data_stage_3__1627_,data_stage_3__1626_,data_stage_3__1625_,
  data_stage_3__1624_,data_stage_3__1623_,data_stage_3__1622_,data_stage_3__1621_,
  data_stage_3__1620_,data_stage_3__1619_,data_stage_3__1618_,data_stage_3__1617_,
  data_stage_3__1616_,data_stage_3__1615_,data_stage_3__1614_,data_stage_3__1613_,
  data_stage_3__1612_,data_stage_3__1611_,data_stage_3__1610_,data_stage_3__1609_,
  data_stage_3__1608_,data_stage_3__1607_,data_stage_3__1606_,data_stage_3__1605_,
  data_stage_3__1604_,data_stage_3__1603_,data_stage_3__1602_,data_stage_3__1601_,
  data_stage_3__1600_,data_stage_3__1599_,data_stage_3__1598_,data_stage_3__1597_,
  data_stage_3__1596_,data_stage_3__1595_,data_stage_3__1594_,data_stage_3__1593_,
  data_stage_3__1592_,data_stage_3__1591_,data_stage_3__1590_,data_stage_3__1589_,
  data_stage_3__1588_,data_stage_3__1587_,data_stage_3__1586_,data_stage_3__1585_,
  data_stage_3__1584_,data_stage_3__1583_,data_stage_3__1582_,data_stage_3__1581_,
  data_stage_3__1580_,data_stage_3__1579_,data_stage_3__1578_,data_stage_3__1577_,
  data_stage_3__1576_,data_stage_3__1575_,data_stage_3__1574_,data_stage_3__1573_,
  data_stage_3__1572_,data_stage_3__1571_,data_stage_3__1570_,data_stage_3__1569_,
  data_stage_3__1568_,data_stage_3__1567_,data_stage_3__1566_,data_stage_3__1565_,
  data_stage_3__1564_,data_stage_3__1563_,data_stage_3__1562_,data_stage_3__1561_,
  data_stage_3__1560_,data_stage_3__1559_,data_stage_3__1558_,data_stage_3__1557_,
  data_stage_3__1556_,data_stage_3__1555_,data_stage_3__1554_,data_stage_3__1553_,
  data_stage_3__1552_,data_stage_3__1551_,data_stage_3__1550_,data_stage_3__1549_,
  data_stage_3__1548_,data_stage_3__1547_,data_stage_3__1546_,data_stage_3__1545_,
  data_stage_3__1544_,data_stage_3__1543_,data_stage_3__1542_,data_stage_3__1541_,
  data_stage_3__1540_,data_stage_3__1539_,data_stage_3__1538_,data_stage_3__1537_,
  data_stage_3__1536_,data_stage_3__1535_,data_stage_3__1534_,data_stage_3__1533_,
  data_stage_3__1532_,data_stage_3__1531_,data_stage_3__1530_,data_stage_3__1529_,
  data_stage_3__1528_,data_stage_3__1527_,data_stage_3__1526_,data_stage_3__1525_,
  data_stage_3__1524_,data_stage_3__1523_,data_stage_3__1522_,data_stage_3__1521_,
  data_stage_3__1520_,data_stage_3__1519_,data_stage_3__1518_,data_stage_3__1517_,
  data_stage_3__1516_,data_stage_3__1515_,data_stage_3__1514_,data_stage_3__1513_,
  data_stage_3__1512_,data_stage_3__1511_,data_stage_3__1510_,data_stage_3__1509_,
  data_stage_3__1508_,data_stage_3__1507_,data_stage_3__1506_,data_stage_3__1505_,
  data_stage_3__1504_,data_stage_3__1503_,data_stage_3__1502_,data_stage_3__1501_,
  data_stage_3__1500_,data_stage_3__1499_,data_stage_3__1498_,data_stage_3__1497_,
  data_stage_3__1496_,data_stage_3__1495_,data_stage_3__1494_,data_stage_3__1493_,
  data_stage_3__1492_,data_stage_3__1491_,data_stage_3__1490_,data_stage_3__1489_,
  data_stage_3__1488_,data_stage_3__1487_,data_stage_3__1486_,data_stage_3__1485_,
  data_stage_3__1484_,data_stage_3__1483_,data_stage_3__1482_,data_stage_3__1481_,
  data_stage_3__1480_,data_stage_3__1479_,data_stage_3__1478_,data_stage_3__1477_,
  data_stage_3__1476_,data_stage_3__1475_,data_stage_3__1474_,data_stage_3__1473_,
  data_stage_3__1472_,data_stage_3__1471_,data_stage_3__1470_,data_stage_3__1469_,
  data_stage_3__1468_,data_stage_3__1467_,data_stage_3__1466_,data_stage_3__1465_,
  data_stage_3__1464_,data_stage_3__1463_,data_stage_3__1462_,data_stage_3__1461_,
  data_stage_3__1460_,data_stage_3__1459_,data_stage_3__1458_,data_stage_3__1457_,
  data_stage_3__1456_,data_stage_3__1455_,data_stage_3__1454_,data_stage_3__1453_,
  data_stage_3__1452_,data_stage_3__1451_,data_stage_3__1450_,data_stage_3__1449_,
  data_stage_3__1448_,data_stage_3__1447_,data_stage_3__1446_,data_stage_3__1445_,
  data_stage_3__1444_,data_stage_3__1443_,data_stage_3__1442_,data_stage_3__1441_,
  data_stage_3__1440_,data_stage_3__1439_,data_stage_3__1438_,data_stage_3__1437_,
  data_stage_3__1436_,data_stage_3__1435_,data_stage_3__1434_,data_stage_3__1433_,
  data_stage_3__1432_,data_stage_3__1431_,data_stage_3__1430_,data_stage_3__1429_,
  data_stage_3__1428_,data_stage_3__1427_,data_stage_3__1426_,data_stage_3__1425_,
  data_stage_3__1424_,data_stage_3__1423_,data_stage_3__1422_,data_stage_3__1421_,
  data_stage_3__1420_,data_stage_3__1419_,data_stage_3__1418_,data_stage_3__1417_,
  data_stage_3__1416_,data_stage_3__1415_,data_stage_3__1414_,data_stage_3__1413_,
  data_stage_3__1412_,data_stage_3__1411_,data_stage_3__1410_,data_stage_3__1409_,
  data_stage_3__1408_,data_stage_3__1407_,data_stage_3__1406_,data_stage_3__1405_,
  data_stage_3__1404_,data_stage_3__1403_,data_stage_3__1402_,data_stage_3__1401_,
  data_stage_3__1400_,data_stage_3__1399_,data_stage_3__1398_,data_stage_3__1397_,
  data_stage_3__1396_,data_stage_3__1395_,data_stage_3__1394_,data_stage_3__1393_,
  data_stage_3__1392_,data_stage_3__1391_,data_stage_3__1390_,data_stage_3__1389_,
  data_stage_3__1388_,data_stage_3__1387_,data_stage_3__1386_,data_stage_3__1385_,
  data_stage_3__1384_,data_stage_3__1383_,data_stage_3__1382_,data_stage_3__1381_,
  data_stage_3__1380_,data_stage_3__1379_,data_stage_3__1378_,data_stage_3__1377_,
  data_stage_3__1376_,data_stage_3__1375_,data_stage_3__1374_,data_stage_3__1373_,
  data_stage_3__1372_,data_stage_3__1371_,data_stage_3__1370_,data_stage_3__1369_,
  data_stage_3__1368_,data_stage_3__1367_,data_stage_3__1366_,data_stage_3__1365_,
  data_stage_3__1364_,data_stage_3__1363_,data_stage_3__1362_,data_stage_3__1361_,
  data_stage_3__1360_,data_stage_3__1359_,data_stage_3__1358_,data_stage_3__1357_,
  data_stage_3__1356_,data_stage_3__1355_,data_stage_3__1354_,data_stage_3__1353_,
  data_stage_3__1352_,data_stage_3__1351_,data_stage_3__1350_,data_stage_3__1349_,
  data_stage_3__1348_,data_stage_3__1347_,data_stage_3__1346_,data_stage_3__1345_,
  data_stage_3__1344_,data_stage_3__1343_,data_stage_3__1342_,data_stage_3__1341_,
  data_stage_3__1340_,data_stage_3__1339_,data_stage_3__1338_,data_stage_3__1337_,
  data_stage_3__1336_,data_stage_3__1335_,data_stage_3__1334_,data_stage_3__1333_,
  data_stage_3__1332_,data_stage_3__1331_,data_stage_3__1330_,data_stage_3__1329_,
  data_stage_3__1328_,data_stage_3__1327_,data_stage_3__1326_,data_stage_3__1325_,
  data_stage_3__1324_,data_stage_3__1323_,data_stage_3__1322_,data_stage_3__1321_,
  data_stage_3__1320_,data_stage_3__1319_,data_stage_3__1318_,data_stage_3__1317_,
  data_stage_3__1316_,data_stage_3__1315_,data_stage_3__1314_,data_stage_3__1313_,
  data_stage_3__1312_,data_stage_3__1311_,data_stage_3__1310_,data_stage_3__1309_,
  data_stage_3__1308_,data_stage_3__1307_,data_stage_3__1306_,data_stage_3__1305_,
  data_stage_3__1304_,data_stage_3__1303_,data_stage_3__1302_,data_stage_3__1301_,
  data_stage_3__1300_,data_stage_3__1299_,data_stage_3__1298_,data_stage_3__1297_,
  data_stage_3__1296_,data_stage_3__1295_,data_stage_3__1294_,data_stage_3__1293_,
  data_stage_3__1292_,data_stage_3__1291_,data_stage_3__1290_,data_stage_3__1289_,
  data_stage_3__1288_,data_stage_3__1287_,data_stage_3__1286_,data_stage_3__1285_,
  data_stage_3__1284_,data_stage_3__1283_,data_stage_3__1282_,data_stage_3__1281_,
  data_stage_3__1280_,data_stage_3__1279_,data_stage_3__1278_,data_stage_3__1277_,
  data_stage_3__1276_,data_stage_3__1275_,data_stage_3__1274_,data_stage_3__1273_,
  data_stage_3__1272_,data_stage_3__1271_,data_stage_3__1270_,data_stage_3__1269_,
  data_stage_3__1268_,data_stage_3__1267_,data_stage_3__1266_,data_stage_3__1265_,
  data_stage_3__1264_,data_stage_3__1263_,data_stage_3__1262_,data_stage_3__1261_,
  data_stage_3__1260_,data_stage_3__1259_,data_stage_3__1258_,data_stage_3__1257_,
  data_stage_3__1256_,data_stage_3__1255_,data_stage_3__1254_,data_stage_3__1253_,
  data_stage_3__1252_,data_stage_3__1251_,data_stage_3__1250_,data_stage_3__1249_,
  data_stage_3__1248_,data_stage_3__1247_,data_stage_3__1246_,data_stage_3__1245_,
  data_stage_3__1244_,data_stage_3__1243_,data_stage_3__1242_,data_stage_3__1241_,
  data_stage_3__1240_,data_stage_3__1239_,data_stage_3__1238_,data_stage_3__1237_,
  data_stage_3__1236_,data_stage_3__1235_,data_stage_3__1234_,data_stage_3__1233_,
  data_stage_3__1232_,data_stage_3__1231_,data_stage_3__1230_,data_stage_3__1229_,
  data_stage_3__1228_,data_stage_3__1227_,data_stage_3__1226_,data_stage_3__1225_,
  data_stage_3__1224_,data_stage_3__1223_,data_stage_3__1222_,data_stage_3__1221_,
  data_stage_3__1220_,data_stage_3__1219_,data_stage_3__1218_,data_stage_3__1217_,
  data_stage_3__1216_,data_stage_3__1215_,data_stage_3__1214_,data_stage_3__1213_,
  data_stage_3__1212_,data_stage_3__1211_,data_stage_3__1210_,data_stage_3__1209_,
  data_stage_3__1208_,data_stage_3__1207_,data_stage_3__1206_,data_stage_3__1205_,
  data_stage_3__1204_,data_stage_3__1203_,data_stage_3__1202_,data_stage_3__1201_,
  data_stage_3__1200_,data_stage_3__1199_,data_stage_3__1198_,data_stage_3__1197_,
  data_stage_3__1196_,data_stage_3__1195_,data_stage_3__1194_,data_stage_3__1193_,
  data_stage_3__1192_,data_stage_3__1191_,data_stage_3__1190_,data_stage_3__1189_,
  data_stage_3__1188_,data_stage_3__1187_,data_stage_3__1186_,data_stage_3__1185_,
  data_stage_3__1184_,data_stage_3__1183_,data_stage_3__1182_,data_stage_3__1181_,
  data_stage_3__1180_,data_stage_3__1179_,data_stage_3__1178_,data_stage_3__1177_,
  data_stage_3__1176_,data_stage_3__1175_,data_stage_3__1174_,data_stage_3__1173_,
  data_stage_3__1172_,data_stage_3__1171_,data_stage_3__1170_,data_stage_3__1169_,
  data_stage_3__1168_,data_stage_3__1167_,data_stage_3__1166_,data_stage_3__1165_,
  data_stage_3__1164_,data_stage_3__1163_,data_stage_3__1162_,data_stage_3__1161_,
  data_stage_3__1160_,data_stage_3__1159_,data_stage_3__1158_,data_stage_3__1157_,
  data_stage_3__1156_,data_stage_3__1155_,data_stage_3__1154_,data_stage_3__1153_,
  data_stage_3__1152_,data_stage_3__1151_,data_stage_3__1150_,data_stage_3__1149_,
  data_stage_3__1148_,data_stage_3__1147_,data_stage_3__1146_,data_stage_3__1145_,
  data_stage_3__1144_,data_stage_3__1143_,data_stage_3__1142_,data_stage_3__1141_,
  data_stage_3__1140_,data_stage_3__1139_,data_stage_3__1138_,data_stage_3__1137_,
  data_stage_3__1136_,data_stage_3__1135_,data_stage_3__1134_,data_stage_3__1133_,
  data_stage_3__1132_,data_stage_3__1131_,data_stage_3__1130_,data_stage_3__1129_,
  data_stage_3__1128_,data_stage_3__1127_,data_stage_3__1126_,data_stage_3__1125_,
  data_stage_3__1124_,data_stage_3__1123_,data_stage_3__1122_,data_stage_3__1121_,
  data_stage_3__1120_,data_stage_3__1119_,data_stage_3__1118_,data_stage_3__1117_,
  data_stage_3__1116_,data_stage_3__1115_,data_stage_3__1114_,data_stage_3__1113_,
  data_stage_3__1112_,data_stage_3__1111_,data_stage_3__1110_,data_stage_3__1109_,
  data_stage_3__1108_,data_stage_3__1107_,data_stage_3__1106_,data_stage_3__1105_,
  data_stage_3__1104_,data_stage_3__1103_,data_stage_3__1102_,data_stage_3__1101_,
  data_stage_3__1100_,data_stage_3__1099_,data_stage_3__1098_,data_stage_3__1097_,
  data_stage_3__1096_,data_stage_3__1095_,data_stage_3__1094_,data_stage_3__1093_,
  data_stage_3__1092_,data_stage_3__1091_,data_stage_3__1090_,data_stage_3__1089_,
  data_stage_3__1088_,data_stage_3__1087_,data_stage_3__1086_,data_stage_3__1085_,
  data_stage_3__1084_,data_stage_3__1083_,data_stage_3__1082_,data_stage_3__1081_,
  data_stage_3__1080_,data_stage_3__1079_,data_stage_3__1078_,data_stage_3__1077_,
  data_stage_3__1076_,data_stage_3__1075_,data_stage_3__1074_,data_stage_3__1073_,
  data_stage_3__1072_,data_stage_3__1071_,data_stage_3__1070_,data_stage_3__1069_,
  data_stage_3__1068_,data_stage_3__1067_,data_stage_3__1066_,data_stage_3__1065_,
  data_stage_3__1064_,data_stage_3__1063_,data_stage_3__1062_,data_stage_3__1061_,
  data_stage_3__1060_,data_stage_3__1059_,data_stage_3__1058_,data_stage_3__1057_,
  data_stage_3__1056_,data_stage_3__1055_,data_stage_3__1054_,data_stage_3__1053_,
  data_stage_3__1052_,data_stage_3__1051_,data_stage_3__1050_,data_stage_3__1049_,
  data_stage_3__1048_,data_stage_3__1047_,data_stage_3__1046_,data_stage_3__1045_,
  data_stage_3__1044_,data_stage_3__1043_,data_stage_3__1042_,data_stage_3__1041_,
  data_stage_3__1040_,data_stage_3__1039_,data_stage_3__1038_,data_stage_3__1037_,
  data_stage_3__1036_,data_stage_3__1035_,data_stage_3__1034_,data_stage_3__1033_,
  data_stage_3__1032_,data_stage_3__1031_,data_stage_3__1030_,data_stage_3__1029_,
  data_stage_3__1028_,data_stage_3__1027_,data_stage_3__1026_,data_stage_3__1025_,
  data_stage_3__1024_,data_stage_3__1023_,data_stage_3__1022_,data_stage_3__1021_,
  data_stage_3__1020_,data_stage_3__1019_,data_stage_3__1018_,data_stage_3__1017_,
  data_stage_3__1016_,data_stage_3__1015_,data_stage_3__1014_,data_stage_3__1013_,
  data_stage_3__1012_,data_stage_3__1011_,data_stage_3__1010_,data_stage_3__1009_,
  data_stage_3__1008_,data_stage_3__1007_,data_stage_3__1006_,data_stage_3__1005_,
  data_stage_3__1004_,data_stage_3__1003_,data_stage_3__1002_,data_stage_3__1001_,
  data_stage_3__1000_,data_stage_3__999_,data_stage_3__998_,data_stage_3__997_,
  data_stage_3__996_,data_stage_3__995_,data_stage_3__994_,data_stage_3__993_,
  data_stage_3__992_,data_stage_3__991_,data_stage_3__990_,data_stage_3__989_,
  data_stage_3__988_,data_stage_3__987_,data_stage_3__986_,data_stage_3__985_,
  data_stage_3__984_,data_stage_3__983_,data_stage_3__982_,data_stage_3__981_,data_stage_3__980_,
  data_stage_3__979_,data_stage_3__978_,data_stage_3__977_,data_stage_3__976_,
  data_stage_3__975_,data_stage_3__974_,data_stage_3__973_,data_stage_3__972_,
  data_stage_3__971_,data_stage_3__970_,data_stage_3__969_,data_stage_3__968_,
  data_stage_3__967_,data_stage_3__966_,data_stage_3__965_,data_stage_3__964_,
  data_stage_3__963_,data_stage_3__962_,data_stage_3__961_,data_stage_3__960_,data_stage_3__959_,
  data_stage_3__958_,data_stage_3__957_,data_stage_3__956_,data_stage_3__955_,
  data_stage_3__954_,data_stage_3__953_,data_stage_3__952_,data_stage_3__951_,
  data_stage_3__950_,data_stage_3__949_,data_stage_3__948_,data_stage_3__947_,
  data_stage_3__946_,data_stage_3__945_,data_stage_3__944_,data_stage_3__943_,
  data_stage_3__942_,data_stage_3__941_,data_stage_3__940_,data_stage_3__939_,data_stage_3__938_,
  data_stage_3__937_,data_stage_3__936_,data_stage_3__935_,data_stage_3__934_,
  data_stage_3__933_,data_stage_3__932_,data_stage_3__931_,data_stage_3__930_,
  data_stage_3__929_,data_stage_3__928_,data_stage_3__927_,data_stage_3__926_,
  data_stage_3__925_,data_stage_3__924_,data_stage_3__923_,data_stage_3__922_,
  data_stage_3__921_,data_stage_3__920_,data_stage_3__919_,data_stage_3__918_,data_stage_3__917_,
  data_stage_3__916_,data_stage_3__915_,data_stage_3__914_,data_stage_3__913_,
  data_stage_3__912_,data_stage_3__911_,data_stage_3__910_,data_stage_3__909_,
  data_stage_3__908_,data_stage_3__907_,data_stage_3__906_,data_stage_3__905_,
  data_stage_3__904_,data_stage_3__903_,data_stage_3__902_,data_stage_3__901_,data_stage_3__900_,
  data_stage_3__899_,data_stage_3__898_,data_stage_3__897_,data_stage_3__896_,
  data_stage_3__895_,data_stage_3__894_,data_stage_3__893_,data_stage_3__892_,
  data_stage_3__891_,data_stage_3__890_,data_stage_3__889_,data_stage_3__888_,
  data_stage_3__887_,data_stage_3__886_,data_stage_3__885_,data_stage_3__884_,
  data_stage_3__883_,data_stage_3__882_,data_stage_3__881_,data_stage_3__880_,data_stage_3__879_,
  data_stage_3__878_,data_stage_3__877_,data_stage_3__876_,data_stage_3__875_,
  data_stage_3__874_,data_stage_3__873_,data_stage_3__872_,data_stage_3__871_,
  data_stage_3__870_,data_stage_3__869_,data_stage_3__868_,data_stage_3__867_,
  data_stage_3__866_,data_stage_3__865_,data_stage_3__864_,data_stage_3__863_,
  data_stage_3__862_,data_stage_3__861_,data_stage_3__860_,data_stage_3__859_,data_stage_3__858_,
  data_stage_3__857_,data_stage_3__856_,data_stage_3__855_,data_stage_3__854_,
  data_stage_3__853_,data_stage_3__852_,data_stage_3__851_,data_stage_3__850_,
  data_stage_3__849_,data_stage_3__848_,data_stage_3__847_,data_stage_3__846_,
  data_stage_3__845_,data_stage_3__844_,data_stage_3__843_,data_stage_3__842_,
  data_stage_3__841_,data_stage_3__840_,data_stage_3__839_,data_stage_3__838_,data_stage_3__837_,
  data_stage_3__836_,data_stage_3__835_,data_stage_3__834_,data_stage_3__833_,
  data_stage_3__832_,data_stage_3__831_,data_stage_3__830_,data_stage_3__829_,
  data_stage_3__828_,data_stage_3__827_,data_stage_3__826_,data_stage_3__825_,
  data_stage_3__824_,data_stage_3__823_,data_stage_3__822_,data_stage_3__821_,data_stage_3__820_,
  data_stage_3__819_,data_stage_3__818_,data_stage_3__817_,data_stage_3__816_,
  data_stage_3__815_,data_stage_3__814_,data_stage_3__813_,data_stage_3__812_,
  data_stage_3__811_,data_stage_3__810_,data_stage_3__809_,data_stage_3__808_,
  data_stage_3__807_,data_stage_3__806_,data_stage_3__805_,data_stage_3__804_,
  data_stage_3__803_,data_stage_3__802_,data_stage_3__801_,data_stage_3__800_,data_stage_3__799_,
  data_stage_3__798_,data_stage_3__797_,data_stage_3__796_,data_stage_3__795_,
  data_stage_3__794_,data_stage_3__793_,data_stage_3__792_,data_stage_3__791_,
  data_stage_3__790_,data_stage_3__789_,data_stage_3__788_,data_stage_3__787_,
  data_stage_3__786_,data_stage_3__785_,data_stage_3__784_,data_stage_3__783_,
  data_stage_3__782_,data_stage_3__781_,data_stage_3__780_,data_stage_3__779_,data_stage_3__778_,
  data_stage_3__777_,data_stage_3__776_,data_stage_3__775_,data_stage_3__774_,
  data_stage_3__773_,data_stage_3__772_,data_stage_3__771_,data_stage_3__770_,
  data_stage_3__769_,data_stage_3__768_,data_stage_3__767_,data_stage_3__766_,
  data_stage_3__765_,data_stage_3__764_,data_stage_3__763_,data_stage_3__762_,
  data_stage_3__761_,data_stage_3__760_,data_stage_3__759_,data_stage_3__758_,data_stage_3__757_,
  data_stage_3__756_,data_stage_3__755_,data_stage_3__754_,data_stage_3__753_,
  data_stage_3__752_,data_stage_3__751_,data_stage_3__750_,data_stage_3__749_,
  data_stage_3__748_,data_stage_3__747_,data_stage_3__746_,data_stage_3__745_,
  data_stage_3__744_,data_stage_3__743_,data_stage_3__742_,data_stage_3__741_,data_stage_3__740_,
  data_stage_3__739_,data_stage_3__738_,data_stage_3__737_,data_stage_3__736_,
  data_stage_3__735_,data_stage_3__734_,data_stage_3__733_,data_stage_3__732_,
  data_stage_3__731_,data_stage_3__730_,data_stage_3__729_,data_stage_3__728_,
  data_stage_3__727_,data_stage_3__726_,data_stage_3__725_,data_stage_3__724_,
  data_stage_3__723_,data_stage_3__722_,data_stage_3__721_,data_stage_3__720_,data_stage_3__719_,
  data_stage_3__718_,data_stage_3__717_,data_stage_3__716_,data_stage_3__715_,
  data_stage_3__714_,data_stage_3__713_,data_stage_3__712_,data_stage_3__711_,
  data_stage_3__710_,data_stage_3__709_,data_stage_3__708_,data_stage_3__707_,
  data_stage_3__706_,data_stage_3__705_,data_stage_3__704_,data_stage_3__703_,
  data_stage_3__702_,data_stage_3__701_,data_stage_3__700_,data_stage_3__699_,data_stage_3__698_,
  data_stage_3__697_,data_stage_3__696_,data_stage_3__695_,data_stage_3__694_,
  data_stage_3__693_,data_stage_3__692_,data_stage_3__691_,data_stage_3__690_,
  data_stage_3__689_,data_stage_3__688_,data_stage_3__687_,data_stage_3__686_,
  data_stage_3__685_,data_stage_3__684_,data_stage_3__683_,data_stage_3__682_,
  data_stage_3__681_,data_stage_3__680_,data_stage_3__679_,data_stage_3__678_,data_stage_3__677_,
  data_stage_3__676_,data_stage_3__675_,data_stage_3__674_,data_stage_3__673_,
  data_stage_3__672_,data_stage_3__671_,data_stage_3__670_,data_stage_3__669_,
  data_stage_3__668_,data_stage_3__667_,data_stage_3__666_,data_stage_3__665_,
  data_stage_3__664_,data_stage_3__663_,data_stage_3__662_,data_stage_3__661_,data_stage_3__660_,
  data_stage_3__659_,data_stage_3__658_,data_stage_3__657_,data_stage_3__656_,
  data_stage_3__655_,data_stage_3__654_,data_stage_3__653_,data_stage_3__652_,
  data_stage_3__651_,data_stage_3__650_,data_stage_3__649_,data_stage_3__648_,
  data_stage_3__647_,data_stage_3__646_,data_stage_3__645_,data_stage_3__644_,
  data_stage_3__643_,data_stage_3__642_,data_stage_3__641_,data_stage_3__640_,data_stage_3__639_,
  data_stage_3__638_,data_stage_3__637_,data_stage_3__636_,data_stage_3__635_,
  data_stage_3__634_,data_stage_3__633_,data_stage_3__632_,data_stage_3__631_,
  data_stage_3__630_,data_stage_3__629_,data_stage_3__628_,data_stage_3__627_,
  data_stage_3__626_,data_stage_3__625_,data_stage_3__624_,data_stage_3__623_,
  data_stage_3__622_,data_stage_3__621_,data_stage_3__620_,data_stage_3__619_,data_stage_3__618_,
  data_stage_3__617_,data_stage_3__616_,data_stage_3__615_,data_stage_3__614_,
  data_stage_3__613_,data_stage_3__612_,data_stage_3__611_,data_stage_3__610_,
  data_stage_3__609_,data_stage_3__608_,data_stage_3__607_,data_stage_3__606_,
  data_stage_3__605_,data_stage_3__604_,data_stage_3__603_,data_stage_3__602_,
  data_stage_3__601_,data_stage_3__600_,data_stage_3__599_,data_stage_3__598_,data_stage_3__597_,
  data_stage_3__596_,data_stage_3__595_,data_stage_3__594_,data_stage_3__593_,
  data_stage_3__592_,data_stage_3__591_,data_stage_3__590_,data_stage_3__589_,
  data_stage_3__588_,data_stage_3__587_,data_stage_3__586_,data_stage_3__585_,
  data_stage_3__584_,data_stage_3__583_,data_stage_3__582_,data_stage_3__581_,data_stage_3__580_,
  data_stage_3__579_,data_stage_3__578_,data_stage_3__577_,data_stage_3__576_,
  data_stage_3__575_,data_stage_3__574_,data_stage_3__573_,data_stage_3__572_,
  data_stage_3__571_,data_stage_3__570_,data_stage_3__569_,data_stage_3__568_,
  data_stage_3__567_,data_stage_3__566_,data_stage_3__565_,data_stage_3__564_,
  data_stage_3__563_,data_stage_3__562_,data_stage_3__561_,data_stage_3__560_,data_stage_3__559_,
  data_stage_3__558_,data_stage_3__557_,data_stage_3__556_,data_stage_3__555_,
  data_stage_3__554_,data_stage_3__553_,data_stage_3__552_,data_stage_3__551_,
  data_stage_3__550_,data_stage_3__549_,data_stage_3__548_,data_stage_3__547_,
  data_stage_3__546_,data_stage_3__545_,data_stage_3__544_,data_stage_3__543_,
  data_stage_3__542_,data_stage_3__541_,data_stage_3__540_,data_stage_3__539_,data_stage_3__538_,
  data_stage_3__537_,data_stage_3__536_,data_stage_3__535_,data_stage_3__534_,
  data_stage_3__533_,data_stage_3__532_,data_stage_3__531_,data_stage_3__530_,
  data_stage_3__529_,data_stage_3__528_,data_stage_3__527_,data_stage_3__526_,
  data_stage_3__525_,data_stage_3__524_,data_stage_3__523_,data_stage_3__522_,
  data_stage_3__521_,data_stage_3__520_,data_stage_3__519_,data_stage_3__518_,data_stage_3__517_,
  data_stage_3__516_,data_stage_3__515_,data_stage_3__514_,data_stage_3__513_,
  data_stage_3__512_,data_stage_3__511_,data_stage_3__510_,data_stage_3__509_,
  data_stage_3__508_,data_stage_3__507_,data_stage_3__506_,data_stage_3__505_,
  data_stage_3__504_,data_stage_3__503_,data_stage_3__502_,data_stage_3__501_,data_stage_3__500_,
  data_stage_3__499_,data_stage_3__498_,data_stage_3__497_,data_stage_3__496_,
  data_stage_3__495_,data_stage_3__494_,data_stage_3__493_,data_stage_3__492_,
  data_stage_3__491_,data_stage_3__490_,data_stage_3__489_,data_stage_3__488_,
  data_stage_3__487_,data_stage_3__486_,data_stage_3__485_,data_stage_3__484_,
  data_stage_3__483_,data_stage_3__482_,data_stage_3__481_,data_stage_3__480_,data_stage_3__479_,
  data_stage_3__478_,data_stage_3__477_,data_stage_3__476_,data_stage_3__475_,
  data_stage_3__474_,data_stage_3__473_,data_stage_3__472_,data_stage_3__471_,
  data_stage_3__470_,data_stage_3__469_,data_stage_3__468_,data_stage_3__467_,
  data_stage_3__466_,data_stage_3__465_,data_stage_3__464_,data_stage_3__463_,
  data_stage_3__462_,data_stage_3__461_,data_stage_3__460_,data_stage_3__459_,data_stage_3__458_,
  data_stage_3__457_,data_stage_3__456_,data_stage_3__455_,data_stage_3__454_,
  data_stage_3__453_,data_stage_3__452_,data_stage_3__451_,data_stage_3__450_,
  data_stage_3__449_,data_stage_3__448_,data_stage_3__447_,data_stage_3__446_,
  data_stage_3__445_,data_stage_3__444_,data_stage_3__443_,data_stage_3__442_,
  data_stage_3__441_,data_stage_3__440_,data_stage_3__439_,data_stage_3__438_,data_stage_3__437_,
  data_stage_3__436_,data_stage_3__435_,data_stage_3__434_,data_stage_3__433_,
  data_stage_3__432_,data_stage_3__431_,data_stage_3__430_,data_stage_3__429_,
  data_stage_3__428_,data_stage_3__427_,data_stage_3__426_,data_stage_3__425_,
  data_stage_3__424_,data_stage_3__423_,data_stage_3__422_,data_stage_3__421_,data_stage_3__420_,
  data_stage_3__419_,data_stage_3__418_,data_stage_3__417_,data_stage_3__416_,
  data_stage_3__415_,data_stage_3__414_,data_stage_3__413_,data_stage_3__412_,
  data_stage_3__411_,data_stage_3__410_,data_stage_3__409_,data_stage_3__408_,
  data_stage_3__407_,data_stage_3__406_,data_stage_3__405_,data_stage_3__404_,
  data_stage_3__403_,data_stage_3__402_,data_stage_3__401_,data_stage_3__400_,data_stage_3__399_,
  data_stage_3__398_,data_stage_3__397_,data_stage_3__396_,data_stage_3__395_,
  data_stage_3__394_,data_stage_3__393_,data_stage_3__392_,data_stage_3__391_,
  data_stage_3__390_,data_stage_3__389_,data_stage_3__388_,data_stage_3__387_,
  data_stage_3__386_,data_stage_3__385_,data_stage_3__384_,data_stage_3__383_,
  data_stage_3__382_,data_stage_3__381_,data_stage_3__380_,data_stage_3__379_,data_stage_3__378_,
  data_stage_3__377_,data_stage_3__376_,data_stage_3__375_,data_stage_3__374_,
  data_stage_3__373_,data_stage_3__372_,data_stage_3__371_,data_stage_3__370_,
  data_stage_3__369_,data_stage_3__368_,data_stage_3__367_,data_stage_3__366_,
  data_stage_3__365_,data_stage_3__364_,data_stage_3__363_,data_stage_3__362_,
  data_stage_3__361_,data_stage_3__360_,data_stage_3__359_,data_stage_3__358_,data_stage_3__357_,
  data_stage_3__356_,data_stage_3__355_,data_stage_3__354_,data_stage_3__353_,
  data_stage_3__352_,data_stage_3__351_,data_stage_3__350_,data_stage_3__349_,
  data_stage_3__348_,data_stage_3__347_,data_stage_3__346_,data_stage_3__345_,
  data_stage_3__344_,data_stage_3__343_,data_stage_3__342_,data_stage_3__341_,data_stage_3__340_,
  data_stage_3__339_,data_stage_3__338_,data_stage_3__337_,data_stage_3__336_,
  data_stage_3__335_,data_stage_3__334_,data_stage_3__333_,data_stage_3__332_,
  data_stage_3__331_,data_stage_3__330_,data_stage_3__329_,data_stage_3__328_,
  data_stage_3__327_,data_stage_3__326_,data_stage_3__325_,data_stage_3__324_,
  data_stage_3__323_,data_stage_3__322_,data_stage_3__321_,data_stage_3__320_,data_stage_3__319_,
  data_stage_3__318_,data_stage_3__317_,data_stage_3__316_,data_stage_3__315_,
  data_stage_3__314_,data_stage_3__313_,data_stage_3__312_,data_stage_3__311_,
  data_stage_3__310_,data_stage_3__309_,data_stage_3__308_,data_stage_3__307_,
  data_stage_3__306_,data_stage_3__305_,data_stage_3__304_,data_stage_3__303_,
  data_stage_3__302_,data_stage_3__301_,data_stage_3__300_,data_stage_3__299_,data_stage_3__298_,
  data_stage_3__297_,data_stage_3__296_,data_stage_3__295_,data_stage_3__294_,
  data_stage_3__293_,data_stage_3__292_,data_stage_3__291_,data_stage_3__290_,
  data_stage_3__289_,data_stage_3__288_,data_stage_3__287_,data_stage_3__286_,
  data_stage_3__285_,data_stage_3__284_,data_stage_3__283_,data_stage_3__282_,
  data_stage_3__281_,data_stage_3__280_,data_stage_3__279_,data_stage_3__278_,data_stage_3__277_,
  data_stage_3__276_,data_stage_3__275_,data_stage_3__274_,data_stage_3__273_,
  data_stage_3__272_,data_stage_3__271_,data_stage_3__270_,data_stage_3__269_,
  data_stage_3__268_,data_stage_3__267_,data_stage_3__266_,data_stage_3__265_,
  data_stage_3__264_,data_stage_3__263_,data_stage_3__262_,data_stage_3__261_,data_stage_3__260_,
  data_stage_3__259_,data_stage_3__258_,data_stage_3__257_,data_stage_3__256_,
  data_stage_3__255_,data_stage_3__254_,data_stage_3__253_,data_stage_3__252_,
  data_stage_3__251_,data_stage_3__250_,data_stage_3__249_,data_stage_3__248_,
  data_stage_3__247_,data_stage_3__246_,data_stage_3__245_,data_stage_3__244_,
  data_stage_3__243_,data_stage_3__242_,data_stage_3__241_,data_stage_3__240_,data_stage_3__239_,
  data_stage_3__238_,data_stage_3__237_,data_stage_3__236_,data_stage_3__235_,
  data_stage_3__234_,data_stage_3__233_,data_stage_3__232_,data_stage_3__231_,
  data_stage_3__230_,data_stage_3__229_,data_stage_3__228_,data_stage_3__227_,
  data_stage_3__226_,data_stage_3__225_,data_stage_3__224_,data_stage_3__223_,
  data_stage_3__222_,data_stage_3__221_,data_stage_3__220_,data_stage_3__219_,data_stage_3__218_,
  data_stage_3__217_,data_stage_3__216_,data_stage_3__215_,data_stage_3__214_,
  data_stage_3__213_,data_stage_3__212_,data_stage_3__211_,data_stage_3__210_,
  data_stage_3__209_,data_stage_3__208_,data_stage_3__207_,data_stage_3__206_,
  data_stage_3__205_,data_stage_3__204_,data_stage_3__203_,data_stage_3__202_,
  data_stage_3__201_,data_stage_3__200_,data_stage_3__199_,data_stage_3__198_,data_stage_3__197_,
  data_stage_3__196_,data_stage_3__195_,data_stage_3__194_,data_stage_3__193_,
  data_stage_3__192_,data_stage_3__191_,data_stage_3__190_,data_stage_3__189_,
  data_stage_3__188_,data_stage_3__187_,data_stage_3__186_,data_stage_3__185_,
  data_stage_3__184_,data_stage_3__183_,data_stage_3__182_,data_stage_3__181_,data_stage_3__180_,
  data_stage_3__179_,data_stage_3__178_,data_stage_3__177_,data_stage_3__176_,
  data_stage_3__175_,data_stage_3__174_,data_stage_3__173_,data_stage_3__172_,
  data_stage_3__171_,data_stage_3__170_,data_stage_3__169_,data_stage_3__168_,
  data_stage_3__167_,data_stage_3__166_,data_stage_3__165_,data_stage_3__164_,
  data_stage_3__163_,data_stage_3__162_,data_stage_3__161_,data_stage_3__160_,data_stage_3__159_,
  data_stage_3__158_,data_stage_3__157_,data_stage_3__156_,data_stage_3__155_,
  data_stage_3__154_,data_stage_3__153_,data_stage_3__152_,data_stage_3__151_,
  data_stage_3__150_,data_stage_3__149_,data_stage_3__148_,data_stage_3__147_,
  data_stage_3__146_,data_stage_3__145_,data_stage_3__144_,data_stage_3__143_,
  data_stage_3__142_,data_stage_3__141_,data_stage_3__140_,data_stage_3__139_,data_stage_3__138_,
  data_stage_3__137_,data_stage_3__136_,data_stage_3__135_,data_stage_3__134_,
  data_stage_3__133_,data_stage_3__132_,data_stage_3__131_,data_stage_3__130_,
  data_stage_3__129_,data_stage_3__128_,data_stage_3__127_,data_stage_3__126_,
  data_stage_3__125_,data_stage_3__124_,data_stage_3__123_,data_stage_3__122_,
  data_stage_3__121_,data_stage_3__120_,data_stage_3__119_,data_stage_3__118_,data_stage_3__117_,
  data_stage_3__116_,data_stage_3__115_,data_stage_3__114_,data_stage_3__113_,
  data_stage_3__112_,data_stage_3__111_,data_stage_3__110_,data_stage_3__109_,
  data_stage_3__108_,data_stage_3__107_,data_stage_3__106_,data_stage_3__105_,
  data_stage_3__104_,data_stage_3__103_,data_stage_3__102_,data_stage_3__101_,data_stage_3__100_,
  data_stage_3__99_,data_stage_3__98_,data_stage_3__97_,data_stage_3__96_,
  data_stage_3__95_,data_stage_3__94_,data_stage_3__93_,data_stage_3__92_,
  data_stage_3__91_,data_stage_3__90_,data_stage_3__89_,data_stage_3__88_,data_stage_3__87_,
  data_stage_3__86_,data_stage_3__85_,data_stage_3__84_,data_stage_3__83_,
  data_stage_3__82_,data_stage_3__81_,data_stage_3__80_,data_stage_3__79_,data_stage_3__78_,
  data_stage_3__77_,data_stage_3__76_,data_stage_3__75_,data_stage_3__74_,
  data_stage_3__73_,data_stage_3__72_,data_stage_3__71_,data_stage_3__70_,data_stage_3__69_,
  data_stage_3__68_,data_stage_3__67_,data_stage_3__66_,data_stage_3__65_,
  data_stage_3__64_,data_stage_3__63_,data_stage_3__62_,data_stage_3__61_,data_stage_3__60_,
  data_stage_3__59_,data_stage_3__58_,data_stage_3__57_,data_stage_3__56_,
  data_stage_3__55_,data_stage_3__54_,data_stage_3__53_,data_stage_3__52_,
  data_stage_3__51_,data_stage_3__50_,data_stage_3__49_,data_stage_3__48_,data_stage_3__47_,
  data_stage_3__46_,data_stage_3__45_,data_stage_3__44_,data_stage_3__43_,
  data_stage_3__42_,data_stage_3__41_,data_stage_3__40_,data_stage_3__39_,data_stage_3__38_,
  data_stage_3__37_,data_stage_3__36_,data_stage_3__35_,data_stage_3__34_,
  data_stage_3__33_,data_stage_3__32_,data_stage_3__31_,data_stage_3__30_,data_stage_3__29_,
  data_stage_3__28_,data_stage_3__27_,data_stage_3__26_,data_stage_3__25_,
  data_stage_3__24_,data_stage_3__23_,data_stage_3__22_,data_stage_3__21_,data_stage_3__20_,
  data_stage_3__19_,data_stage_3__18_,data_stage_3__17_,data_stage_3__16_,
  data_stage_3__15_,data_stage_3__14_,data_stage_3__13_,data_stage_3__12_,
  data_stage_3__11_,data_stage_3__10_,data_stage_3__9_,data_stage_3__8_,data_stage_3__7_,
  data_stage_3__6_,data_stage_3__5_,data_stage_3__4_,data_stage_3__3_,data_stage_3__2_,
  data_stage_3__1_,data_stage_3__0_,data_stage_4__4095_,data_stage_4__4094_,
  data_stage_4__4093_,data_stage_4__4092_,data_stage_4__4091_,data_stage_4__4090_,
  data_stage_4__4089_,data_stage_4__4088_,data_stage_4__4087_,data_stage_4__4086_,
  data_stage_4__4085_,data_stage_4__4084_,data_stage_4__4083_,data_stage_4__4082_,
  data_stage_4__4081_,data_stage_4__4080_,data_stage_4__4079_,data_stage_4__4078_,
  data_stage_4__4077_,data_stage_4__4076_,data_stage_4__4075_,data_stage_4__4074_,
  data_stage_4__4073_,data_stage_4__4072_,data_stage_4__4071_,data_stage_4__4070_,
  data_stage_4__4069_,data_stage_4__4068_,data_stage_4__4067_,data_stage_4__4066_,
  data_stage_4__4065_,data_stage_4__4064_,data_stage_4__4063_,data_stage_4__4062_,
  data_stage_4__4061_,data_stage_4__4060_,data_stage_4__4059_,data_stage_4__4058_,
  data_stage_4__4057_,data_stage_4__4056_,data_stage_4__4055_,data_stage_4__4054_,
  data_stage_4__4053_,data_stage_4__4052_,data_stage_4__4051_,data_stage_4__4050_,
  data_stage_4__4049_,data_stage_4__4048_,data_stage_4__4047_,data_stage_4__4046_,
  data_stage_4__4045_,data_stage_4__4044_,data_stage_4__4043_,data_stage_4__4042_,
  data_stage_4__4041_,data_stage_4__4040_,data_stage_4__4039_,data_stage_4__4038_,
  data_stage_4__4037_,data_stage_4__4036_,data_stage_4__4035_,data_stage_4__4034_,
  data_stage_4__4033_,data_stage_4__4032_,data_stage_4__4031_,data_stage_4__4030_,
  data_stage_4__4029_,data_stage_4__4028_,data_stage_4__4027_,data_stage_4__4026_,
  data_stage_4__4025_,data_stage_4__4024_,data_stage_4__4023_,data_stage_4__4022_,
  data_stage_4__4021_,data_stage_4__4020_,data_stage_4__4019_,data_stage_4__4018_,
  data_stage_4__4017_,data_stage_4__4016_,data_stage_4__4015_,data_stage_4__4014_,
  data_stage_4__4013_,data_stage_4__4012_,data_stage_4__4011_,data_stage_4__4010_,
  data_stage_4__4009_,data_stage_4__4008_,data_stage_4__4007_,data_stage_4__4006_,
  data_stage_4__4005_,data_stage_4__4004_,data_stage_4__4003_,data_stage_4__4002_,
  data_stage_4__4001_,data_stage_4__4000_,data_stage_4__3999_,data_stage_4__3998_,
  data_stage_4__3997_,data_stage_4__3996_,data_stage_4__3995_,data_stage_4__3994_,
  data_stage_4__3993_,data_stage_4__3992_,data_stage_4__3991_,data_stage_4__3990_,
  data_stage_4__3989_,data_stage_4__3988_,data_stage_4__3987_,data_stage_4__3986_,
  data_stage_4__3985_,data_stage_4__3984_,data_stage_4__3983_,data_stage_4__3982_,
  data_stage_4__3981_,data_stage_4__3980_,data_stage_4__3979_,data_stage_4__3978_,
  data_stage_4__3977_,data_stage_4__3976_,data_stage_4__3975_,data_stage_4__3974_,
  data_stage_4__3973_,data_stage_4__3972_,data_stage_4__3971_,data_stage_4__3970_,
  data_stage_4__3969_,data_stage_4__3968_,data_stage_4__3967_,data_stage_4__3966_,
  data_stage_4__3965_,data_stage_4__3964_,data_stage_4__3963_,data_stage_4__3962_,
  data_stage_4__3961_,data_stage_4__3960_,data_stage_4__3959_,data_stage_4__3958_,
  data_stage_4__3957_,data_stage_4__3956_,data_stage_4__3955_,data_stage_4__3954_,
  data_stage_4__3953_,data_stage_4__3952_,data_stage_4__3951_,data_stage_4__3950_,
  data_stage_4__3949_,data_stage_4__3948_,data_stage_4__3947_,data_stage_4__3946_,
  data_stage_4__3945_,data_stage_4__3944_,data_stage_4__3943_,data_stage_4__3942_,
  data_stage_4__3941_,data_stage_4__3940_,data_stage_4__3939_,data_stage_4__3938_,
  data_stage_4__3937_,data_stage_4__3936_,data_stage_4__3935_,data_stage_4__3934_,
  data_stage_4__3933_,data_stage_4__3932_,data_stage_4__3931_,data_stage_4__3930_,
  data_stage_4__3929_,data_stage_4__3928_,data_stage_4__3927_,data_stage_4__3926_,
  data_stage_4__3925_,data_stage_4__3924_,data_stage_4__3923_,data_stage_4__3922_,
  data_stage_4__3921_,data_stage_4__3920_,data_stage_4__3919_,data_stage_4__3918_,
  data_stage_4__3917_,data_stage_4__3916_,data_stage_4__3915_,data_stage_4__3914_,
  data_stage_4__3913_,data_stage_4__3912_,data_stage_4__3911_,data_stage_4__3910_,
  data_stage_4__3909_,data_stage_4__3908_,data_stage_4__3907_,data_stage_4__3906_,
  data_stage_4__3905_,data_stage_4__3904_,data_stage_4__3903_,data_stage_4__3902_,
  data_stage_4__3901_,data_stage_4__3900_,data_stage_4__3899_,data_stage_4__3898_,
  data_stage_4__3897_,data_stage_4__3896_,data_stage_4__3895_,data_stage_4__3894_,
  data_stage_4__3893_,data_stage_4__3892_,data_stage_4__3891_,data_stage_4__3890_,
  data_stage_4__3889_,data_stage_4__3888_,data_stage_4__3887_,data_stage_4__3886_,
  data_stage_4__3885_,data_stage_4__3884_,data_stage_4__3883_,data_stage_4__3882_,
  data_stage_4__3881_,data_stage_4__3880_,data_stage_4__3879_,data_stage_4__3878_,
  data_stage_4__3877_,data_stage_4__3876_,data_stage_4__3875_,data_stage_4__3874_,
  data_stage_4__3873_,data_stage_4__3872_,data_stage_4__3871_,data_stage_4__3870_,
  data_stage_4__3869_,data_stage_4__3868_,data_stage_4__3867_,data_stage_4__3866_,
  data_stage_4__3865_,data_stage_4__3864_,data_stage_4__3863_,data_stage_4__3862_,
  data_stage_4__3861_,data_stage_4__3860_,data_stage_4__3859_,data_stage_4__3858_,
  data_stage_4__3857_,data_stage_4__3856_,data_stage_4__3855_,data_stage_4__3854_,
  data_stage_4__3853_,data_stage_4__3852_,data_stage_4__3851_,data_stage_4__3850_,
  data_stage_4__3849_,data_stage_4__3848_,data_stage_4__3847_,data_stage_4__3846_,
  data_stage_4__3845_,data_stage_4__3844_,data_stage_4__3843_,data_stage_4__3842_,
  data_stage_4__3841_,data_stage_4__3840_,data_stage_4__3839_,data_stage_4__3838_,
  data_stage_4__3837_,data_stage_4__3836_,data_stage_4__3835_,data_stage_4__3834_,
  data_stage_4__3833_,data_stage_4__3832_,data_stage_4__3831_,data_stage_4__3830_,
  data_stage_4__3829_,data_stage_4__3828_,data_stage_4__3827_,data_stage_4__3826_,
  data_stage_4__3825_,data_stage_4__3824_,data_stage_4__3823_,data_stage_4__3822_,
  data_stage_4__3821_,data_stage_4__3820_,data_stage_4__3819_,data_stage_4__3818_,
  data_stage_4__3817_,data_stage_4__3816_,data_stage_4__3815_,data_stage_4__3814_,
  data_stage_4__3813_,data_stage_4__3812_,data_stage_4__3811_,data_stage_4__3810_,
  data_stage_4__3809_,data_stage_4__3808_,data_stage_4__3807_,data_stage_4__3806_,
  data_stage_4__3805_,data_stage_4__3804_,data_stage_4__3803_,data_stage_4__3802_,
  data_stage_4__3801_,data_stage_4__3800_,data_stage_4__3799_,data_stage_4__3798_,
  data_stage_4__3797_,data_stage_4__3796_,data_stage_4__3795_,data_stage_4__3794_,
  data_stage_4__3793_,data_stage_4__3792_,data_stage_4__3791_,data_stage_4__3790_,
  data_stage_4__3789_,data_stage_4__3788_,data_stage_4__3787_,data_stage_4__3786_,
  data_stage_4__3785_,data_stage_4__3784_,data_stage_4__3783_,data_stage_4__3782_,
  data_stage_4__3781_,data_stage_4__3780_,data_stage_4__3779_,data_stage_4__3778_,
  data_stage_4__3777_,data_stage_4__3776_,data_stage_4__3775_,data_stage_4__3774_,
  data_stage_4__3773_,data_stage_4__3772_,data_stage_4__3771_,data_stage_4__3770_,
  data_stage_4__3769_,data_stage_4__3768_,data_stage_4__3767_,data_stage_4__3766_,
  data_stage_4__3765_,data_stage_4__3764_,data_stage_4__3763_,data_stage_4__3762_,
  data_stage_4__3761_,data_stage_4__3760_,data_stage_4__3759_,data_stage_4__3758_,
  data_stage_4__3757_,data_stage_4__3756_,data_stage_4__3755_,data_stage_4__3754_,
  data_stage_4__3753_,data_stage_4__3752_,data_stage_4__3751_,data_stage_4__3750_,
  data_stage_4__3749_,data_stage_4__3748_,data_stage_4__3747_,data_stage_4__3746_,
  data_stage_4__3745_,data_stage_4__3744_,data_stage_4__3743_,data_stage_4__3742_,
  data_stage_4__3741_,data_stage_4__3740_,data_stage_4__3739_,data_stage_4__3738_,
  data_stage_4__3737_,data_stage_4__3736_,data_stage_4__3735_,data_stage_4__3734_,
  data_stage_4__3733_,data_stage_4__3732_,data_stage_4__3731_,data_stage_4__3730_,
  data_stage_4__3729_,data_stage_4__3728_,data_stage_4__3727_,data_stage_4__3726_,
  data_stage_4__3725_,data_stage_4__3724_,data_stage_4__3723_,data_stage_4__3722_,
  data_stage_4__3721_,data_stage_4__3720_,data_stage_4__3719_,data_stage_4__3718_,
  data_stage_4__3717_,data_stage_4__3716_,data_stage_4__3715_,data_stage_4__3714_,
  data_stage_4__3713_,data_stage_4__3712_,data_stage_4__3711_,data_stage_4__3710_,
  data_stage_4__3709_,data_stage_4__3708_,data_stage_4__3707_,data_stage_4__3706_,
  data_stage_4__3705_,data_stage_4__3704_,data_stage_4__3703_,data_stage_4__3702_,
  data_stage_4__3701_,data_stage_4__3700_,data_stage_4__3699_,data_stage_4__3698_,
  data_stage_4__3697_,data_stage_4__3696_,data_stage_4__3695_,data_stage_4__3694_,
  data_stage_4__3693_,data_stage_4__3692_,data_stage_4__3691_,data_stage_4__3690_,
  data_stage_4__3689_,data_stage_4__3688_,data_stage_4__3687_,data_stage_4__3686_,
  data_stage_4__3685_,data_stage_4__3684_,data_stage_4__3683_,data_stage_4__3682_,
  data_stage_4__3681_,data_stage_4__3680_,data_stage_4__3679_,data_stage_4__3678_,
  data_stage_4__3677_,data_stage_4__3676_,data_stage_4__3675_,data_stage_4__3674_,
  data_stage_4__3673_,data_stage_4__3672_,data_stage_4__3671_,data_stage_4__3670_,
  data_stage_4__3669_,data_stage_4__3668_,data_stage_4__3667_,data_stage_4__3666_,
  data_stage_4__3665_,data_stage_4__3664_,data_stage_4__3663_,data_stage_4__3662_,
  data_stage_4__3661_,data_stage_4__3660_,data_stage_4__3659_,data_stage_4__3658_,
  data_stage_4__3657_,data_stage_4__3656_,data_stage_4__3655_,data_stage_4__3654_,
  data_stage_4__3653_,data_stage_4__3652_,data_stage_4__3651_,data_stage_4__3650_,
  data_stage_4__3649_,data_stage_4__3648_,data_stage_4__3647_,data_stage_4__3646_,
  data_stage_4__3645_,data_stage_4__3644_,data_stage_4__3643_,data_stage_4__3642_,
  data_stage_4__3641_,data_stage_4__3640_,data_stage_4__3639_,data_stage_4__3638_,
  data_stage_4__3637_,data_stage_4__3636_,data_stage_4__3635_,data_stage_4__3634_,
  data_stage_4__3633_,data_stage_4__3632_,data_stage_4__3631_,data_stage_4__3630_,
  data_stage_4__3629_,data_stage_4__3628_,data_stage_4__3627_,data_stage_4__3626_,
  data_stage_4__3625_,data_stage_4__3624_,data_stage_4__3623_,data_stage_4__3622_,
  data_stage_4__3621_,data_stage_4__3620_,data_stage_4__3619_,data_stage_4__3618_,
  data_stage_4__3617_,data_stage_4__3616_,data_stage_4__3615_,data_stage_4__3614_,
  data_stage_4__3613_,data_stage_4__3612_,data_stage_4__3611_,data_stage_4__3610_,
  data_stage_4__3609_,data_stage_4__3608_,data_stage_4__3607_,data_stage_4__3606_,
  data_stage_4__3605_,data_stage_4__3604_,data_stage_4__3603_,data_stage_4__3602_,
  data_stage_4__3601_,data_stage_4__3600_,data_stage_4__3599_,data_stage_4__3598_,
  data_stage_4__3597_,data_stage_4__3596_,data_stage_4__3595_,data_stage_4__3594_,
  data_stage_4__3593_,data_stage_4__3592_,data_stage_4__3591_,data_stage_4__3590_,
  data_stage_4__3589_,data_stage_4__3588_,data_stage_4__3587_,data_stage_4__3586_,
  data_stage_4__3585_,data_stage_4__3584_,data_stage_4__3583_,data_stage_4__3582_,
  data_stage_4__3581_,data_stage_4__3580_,data_stage_4__3579_,data_stage_4__3578_,
  data_stage_4__3577_,data_stage_4__3576_,data_stage_4__3575_,data_stage_4__3574_,
  data_stage_4__3573_,data_stage_4__3572_,data_stage_4__3571_,data_stage_4__3570_,
  data_stage_4__3569_,data_stage_4__3568_,data_stage_4__3567_,data_stage_4__3566_,
  data_stage_4__3565_,data_stage_4__3564_,data_stage_4__3563_,data_stage_4__3562_,
  data_stage_4__3561_,data_stage_4__3560_,data_stage_4__3559_,data_stage_4__3558_,
  data_stage_4__3557_,data_stage_4__3556_,data_stage_4__3555_,data_stage_4__3554_,
  data_stage_4__3553_,data_stage_4__3552_,data_stage_4__3551_,data_stage_4__3550_,
  data_stage_4__3549_,data_stage_4__3548_,data_stage_4__3547_,data_stage_4__3546_,
  data_stage_4__3545_,data_stage_4__3544_,data_stage_4__3543_,data_stage_4__3542_,
  data_stage_4__3541_,data_stage_4__3540_,data_stage_4__3539_,data_stage_4__3538_,
  data_stage_4__3537_,data_stage_4__3536_,data_stage_4__3535_,data_stage_4__3534_,
  data_stage_4__3533_,data_stage_4__3532_,data_stage_4__3531_,data_stage_4__3530_,
  data_stage_4__3529_,data_stage_4__3528_,data_stage_4__3527_,data_stage_4__3526_,
  data_stage_4__3525_,data_stage_4__3524_,data_stage_4__3523_,data_stage_4__3522_,
  data_stage_4__3521_,data_stage_4__3520_,data_stage_4__3519_,data_stage_4__3518_,
  data_stage_4__3517_,data_stage_4__3516_,data_stage_4__3515_,data_stage_4__3514_,
  data_stage_4__3513_,data_stage_4__3512_,data_stage_4__3511_,data_stage_4__3510_,
  data_stage_4__3509_,data_stage_4__3508_,data_stage_4__3507_,data_stage_4__3506_,
  data_stage_4__3505_,data_stage_4__3504_,data_stage_4__3503_,data_stage_4__3502_,
  data_stage_4__3501_,data_stage_4__3500_,data_stage_4__3499_,data_stage_4__3498_,
  data_stage_4__3497_,data_stage_4__3496_,data_stage_4__3495_,data_stage_4__3494_,
  data_stage_4__3493_,data_stage_4__3492_,data_stage_4__3491_,data_stage_4__3490_,
  data_stage_4__3489_,data_stage_4__3488_,data_stage_4__3487_,data_stage_4__3486_,
  data_stage_4__3485_,data_stage_4__3484_,data_stage_4__3483_,data_stage_4__3482_,
  data_stage_4__3481_,data_stage_4__3480_,data_stage_4__3479_,data_stage_4__3478_,
  data_stage_4__3477_,data_stage_4__3476_,data_stage_4__3475_,data_stage_4__3474_,
  data_stage_4__3473_,data_stage_4__3472_,data_stage_4__3471_,data_stage_4__3470_,
  data_stage_4__3469_,data_stage_4__3468_,data_stage_4__3467_,data_stage_4__3466_,
  data_stage_4__3465_,data_stage_4__3464_,data_stage_4__3463_,data_stage_4__3462_,
  data_stage_4__3461_,data_stage_4__3460_,data_stage_4__3459_,data_stage_4__3458_,
  data_stage_4__3457_,data_stage_4__3456_,data_stage_4__3455_,data_stage_4__3454_,
  data_stage_4__3453_,data_stage_4__3452_,data_stage_4__3451_,data_stage_4__3450_,
  data_stage_4__3449_,data_stage_4__3448_,data_stage_4__3447_,data_stage_4__3446_,
  data_stage_4__3445_,data_stage_4__3444_,data_stage_4__3443_,data_stage_4__3442_,
  data_stage_4__3441_,data_stage_4__3440_,data_stage_4__3439_,data_stage_4__3438_,
  data_stage_4__3437_,data_stage_4__3436_,data_stage_4__3435_,data_stage_4__3434_,
  data_stage_4__3433_,data_stage_4__3432_,data_stage_4__3431_,data_stage_4__3430_,
  data_stage_4__3429_,data_stage_4__3428_,data_stage_4__3427_,data_stage_4__3426_,
  data_stage_4__3425_,data_stage_4__3424_,data_stage_4__3423_,data_stage_4__3422_,
  data_stage_4__3421_,data_stage_4__3420_,data_stage_4__3419_,data_stage_4__3418_,
  data_stage_4__3417_,data_stage_4__3416_,data_stage_4__3415_,data_stage_4__3414_,
  data_stage_4__3413_,data_stage_4__3412_,data_stage_4__3411_,data_stage_4__3410_,
  data_stage_4__3409_,data_stage_4__3408_,data_stage_4__3407_,data_stage_4__3406_,
  data_stage_4__3405_,data_stage_4__3404_,data_stage_4__3403_,data_stage_4__3402_,
  data_stage_4__3401_,data_stage_4__3400_,data_stage_4__3399_,data_stage_4__3398_,
  data_stage_4__3397_,data_stage_4__3396_,data_stage_4__3395_,data_stage_4__3394_,
  data_stage_4__3393_,data_stage_4__3392_,data_stage_4__3391_,data_stage_4__3390_,
  data_stage_4__3389_,data_stage_4__3388_,data_stage_4__3387_,data_stage_4__3386_,
  data_stage_4__3385_,data_stage_4__3384_,data_stage_4__3383_,data_stage_4__3382_,
  data_stage_4__3381_,data_stage_4__3380_,data_stage_4__3379_,data_stage_4__3378_,
  data_stage_4__3377_,data_stage_4__3376_,data_stage_4__3375_,data_stage_4__3374_,
  data_stage_4__3373_,data_stage_4__3372_,data_stage_4__3371_,data_stage_4__3370_,
  data_stage_4__3369_,data_stage_4__3368_,data_stage_4__3367_,data_stage_4__3366_,
  data_stage_4__3365_,data_stage_4__3364_,data_stage_4__3363_,data_stage_4__3362_,
  data_stage_4__3361_,data_stage_4__3360_,data_stage_4__3359_,data_stage_4__3358_,
  data_stage_4__3357_,data_stage_4__3356_,data_stage_4__3355_,data_stage_4__3354_,
  data_stage_4__3353_,data_stage_4__3352_,data_stage_4__3351_,data_stage_4__3350_,
  data_stage_4__3349_,data_stage_4__3348_,data_stage_4__3347_,data_stage_4__3346_,
  data_stage_4__3345_,data_stage_4__3344_,data_stage_4__3343_,data_stage_4__3342_,
  data_stage_4__3341_,data_stage_4__3340_,data_stage_4__3339_,data_stage_4__3338_,
  data_stage_4__3337_,data_stage_4__3336_,data_stage_4__3335_,data_stage_4__3334_,
  data_stage_4__3333_,data_stage_4__3332_,data_stage_4__3331_,data_stage_4__3330_,
  data_stage_4__3329_,data_stage_4__3328_,data_stage_4__3327_,data_stage_4__3326_,
  data_stage_4__3325_,data_stage_4__3324_,data_stage_4__3323_,data_stage_4__3322_,
  data_stage_4__3321_,data_stage_4__3320_,data_stage_4__3319_,data_stage_4__3318_,
  data_stage_4__3317_,data_stage_4__3316_,data_stage_4__3315_,data_stage_4__3314_,
  data_stage_4__3313_,data_stage_4__3312_,data_stage_4__3311_,data_stage_4__3310_,
  data_stage_4__3309_,data_stage_4__3308_,data_stage_4__3307_,data_stage_4__3306_,
  data_stage_4__3305_,data_stage_4__3304_,data_stage_4__3303_,data_stage_4__3302_,
  data_stage_4__3301_,data_stage_4__3300_,data_stage_4__3299_,data_stage_4__3298_,
  data_stage_4__3297_,data_stage_4__3296_,data_stage_4__3295_,data_stage_4__3294_,
  data_stage_4__3293_,data_stage_4__3292_,data_stage_4__3291_,data_stage_4__3290_,
  data_stage_4__3289_,data_stage_4__3288_,data_stage_4__3287_,data_stage_4__3286_,
  data_stage_4__3285_,data_stage_4__3284_,data_stage_4__3283_,data_stage_4__3282_,
  data_stage_4__3281_,data_stage_4__3280_,data_stage_4__3279_,data_stage_4__3278_,
  data_stage_4__3277_,data_stage_4__3276_,data_stage_4__3275_,data_stage_4__3274_,
  data_stage_4__3273_,data_stage_4__3272_,data_stage_4__3271_,data_stage_4__3270_,
  data_stage_4__3269_,data_stage_4__3268_,data_stage_4__3267_,data_stage_4__3266_,
  data_stage_4__3265_,data_stage_4__3264_,data_stage_4__3263_,data_stage_4__3262_,
  data_stage_4__3261_,data_stage_4__3260_,data_stage_4__3259_,data_stage_4__3258_,
  data_stage_4__3257_,data_stage_4__3256_,data_stage_4__3255_,data_stage_4__3254_,
  data_stage_4__3253_,data_stage_4__3252_,data_stage_4__3251_,data_stage_4__3250_,
  data_stage_4__3249_,data_stage_4__3248_,data_stage_4__3247_,data_stage_4__3246_,
  data_stage_4__3245_,data_stage_4__3244_,data_stage_4__3243_,data_stage_4__3242_,
  data_stage_4__3241_,data_stage_4__3240_,data_stage_4__3239_,data_stage_4__3238_,
  data_stage_4__3237_,data_stage_4__3236_,data_stage_4__3235_,data_stage_4__3234_,
  data_stage_4__3233_,data_stage_4__3232_,data_stage_4__3231_,data_stage_4__3230_,
  data_stage_4__3229_,data_stage_4__3228_,data_stage_4__3227_,data_stage_4__3226_,
  data_stage_4__3225_,data_stage_4__3224_,data_stage_4__3223_,data_stage_4__3222_,
  data_stage_4__3221_,data_stage_4__3220_,data_stage_4__3219_,data_stage_4__3218_,
  data_stage_4__3217_,data_stage_4__3216_,data_stage_4__3215_,data_stage_4__3214_,
  data_stage_4__3213_,data_stage_4__3212_,data_stage_4__3211_,data_stage_4__3210_,
  data_stage_4__3209_,data_stage_4__3208_,data_stage_4__3207_,data_stage_4__3206_,
  data_stage_4__3205_,data_stage_4__3204_,data_stage_4__3203_,data_stage_4__3202_,
  data_stage_4__3201_,data_stage_4__3200_,data_stage_4__3199_,data_stage_4__3198_,
  data_stage_4__3197_,data_stage_4__3196_,data_stage_4__3195_,data_stage_4__3194_,
  data_stage_4__3193_,data_stage_4__3192_,data_stage_4__3191_,data_stage_4__3190_,
  data_stage_4__3189_,data_stage_4__3188_,data_stage_4__3187_,data_stage_4__3186_,
  data_stage_4__3185_,data_stage_4__3184_,data_stage_4__3183_,data_stage_4__3182_,
  data_stage_4__3181_,data_stage_4__3180_,data_stage_4__3179_,data_stage_4__3178_,
  data_stage_4__3177_,data_stage_4__3176_,data_stage_4__3175_,data_stage_4__3174_,
  data_stage_4__3173_,data_stage_4__3172_,data_stage_4__3171_,data_stage_4__3170_,
  data_stage_4__3169_,data_stage_4__3168_,data_stage_4__3167_,data_stage_4__3166_,
  data_stage_4__3165_,data_stage_4__3164_,data_stage_4__3163_,data_stage_4__3162_,
  data_stage_4__3161_,data_stage_4__3160_,data_stage_4__3159_,data_stage_4__3158_,
  data_stage_4__3157_,data_stage_4__3156_,data_stage_4__3155_,data_stage_4__3154_,
  data_stage_4__3153_,data_stage_4__3152_,data_stage_4__3151_,data_stage_4__3150_,
  data_stage_4__3149_,data_stage_4__3148_,data_stage_4__3147_,data_stage_4__3146_,
  data_stage_4__3145_,data_stage_4__3144_,data_stage_4__3143_,data_stage_4__3142_,
  data_stage_4__3141_,data_stage_4__3140_,data_stage_4__3139_,data_stage_4__3138_,
  data_stage_4__3137_,data_stage_4__3136_,data_stage_4__3135_,data_stage_4__3134_,
  data_stage_4__3133_,data_stage_4__3132_,data_stage_4__3131_,data_stage_4__3130_,
  data_stage_4__3129_,data_stage_4__3128_,data_stage_4__3127_,data_stage_4__3126_,
  data_stage_4__3125_,data_stage_4__3124_,data_stage_4__3123_,data_stage_4__3122_,
  data_stage_4__3121_,data_stage_4__3120_,data_stage_4__3119_,data_stage_4__3118_,
  data_stage_4__3117_,data_stage_4__3116_,data_stage_4__3115_,data_stage_4__3114_,
  data_stage_4__3113_,data_stage_4__3112_,data_stage_4__3111_,data_stage_4__3110_,
  data_stage_4__3109_,data_stage_4__3108_,data_stage_4__3107_,data_stage_4__3106_,
  data_stage_4__3105_,data_stage_4__3104_,data_stage_4__3103_,data_stage_4__3102_,
  data_stage_4__3101_,data_stage_4__3100_,data_stage_4__3099_,data_stage_4__3098_,
  data_stage_4__3097_,data_stage_4__3096_,data_stage_4__3095_,data_stage_4__3094_,
  data_stage_4__3093_,data_stage_4__3092_,data_stage_4__3091_,data_stage_4__3090_,
  data_stage_4__3089_,data_stage_4__3088_,data_stage_4__3087_,data_stage_4__3086_,
  data_stage_4__3085_,data_stage_4__3084_,data_stage_4__3083_,data_stage_4__3082_,
  data_stage_4__3081_,data_stage_4__3080_,data_stage_4__3079_,data_stage_4__3078_,
  data_stage_4__3077_,data_stage_4__3076_,data_stage_4__3075_,data_stage_4__3074_,
  data_stage_4__3073_,data_stage_4__3072_,data_stage_4__3071_,data_stage_4__3070_,
  data_stage_4__3069_,data_stage_4__3068_,data_stage_4__3067_,data_stage_4__3066_,
  data_stage_4__3065_,data_stage_4__3064_,data_stage_4__3063_,data_stage_4__3062_,
  data_stage_4__3061_,data_stage_4__3060_,data_stage_4__3059_,data_stage_4__3058_,
  data_stage_4__3057_,data_stage_4__3056_,data_stage_4__3055_,data_stage_4__3054_,
  data_stage_4__3053_,data_stage_4__3052_,data_stage_4__3051_,data_stage_4__3050_,
  data_stage_4__3049_,data_stage_4__3048_,data_stage_4__3047_,data_stage_4__3046_,
  data_stage_4__3045_,data_stage_4__3044_,data_stage_4__3043_,data_stage_4__3042_,
  data_stage_4__3041_,data_stage_4__3040_,data_stage_4__3039_,data_stage_4__3038_,
  data_stage_4__3037_,data_stage_4__3036_,data_stage_4__3035_,data_stage_4__3034_,
  data_stage_4__3033_,data_stage_4__3032_,data_stage_4__3031_,data_stage_4__3030_,
  data_stage_4__3029_,data_stage_4__3028_,data_stage_4__3027_,data_stage_4__3026_,
  data_stage_4__3025_,data_stage_4__3024_,data_stage_4__3023_,data_stage_4__3022_,
  data_stage_4__3021_,data_stage_4__3020_,data_stage_4__3019_,data_stage_4__3018_,
  data_stage_4__3017_,data_stage_4__3016_,data_stage_4__3015_,data_stage_4__3014_,
  data_stage_4__3013_,data_stage_4__3012_,data_stage_4__3011_,data_stage_4__3010_,
  data_stage_4__3009_,data_stage_4__3008_,data_stage_4__3007_,data_stage_4__3006_,
  data_stage_4__3005_,data_stage_4__3004_,data_stage_4__3003_,data_stage_4__3002_,
  data_stage_4__3001_,data_stage_4__3000_,data_stage_4__2999_,data_stage_4__2998_,
  data_stage_4__2997_,data_stage_4__2996_,data_stage_4__2995_,data_stage_4__2994_,
  data_stage_4__2993_,data_stage_4__2992_,data_stage_4__2991_,data_stage_4__2990_,
  data_stage_4__2989_,data_stage_4__2988_,data_stage_4__2987_,data_stage_4__2986_,
  data_stage_4__2985_,data_stage_4__2984_,data_stage_4__2983_,data_stage_4__2982_,
  data_stage_4__2981_,data_stage_4__2980_,data_stage_4__2979_,data_stage_4__2978_,
  data_stage_4__2977_,data_stage_4__2976_,data_stage_4__2975_,data_stage_4__2974_,
  data_stage_4__2973_,data_stage_4__2972_,data_stage_4__2971_,data_stage_4__2970_,
  data_stage_4__2969_,data_stage_4__2968_,data_stage_4__2967_,data_stage_4__2966_,
  data_stage_4__2965_,data_stage_4__2964_,data_stage_4__2963_,data_stage_4__2962_,
  data_stage_4__2961_,data_stage_4__2960_,data_stage_4__2959_,data_stage_4__2958_,
  data_stage_4__2957_,data_stage_4__2956_,data_stage_4__2955_,data_stage_4__2954_,
  data_stage_4__2953_,data_stage_4__2952_,data_stage_4__2951_,data_stage_4__2950_,
  data_stage_4__2949_,data_stage_4__2948_,data_stage_4__2947_,data_stage_4__2946_,
  data_stage_4__2945_,data_stage_4__2944_,data_stage_4__2943_,data_stage_4__2942_,
  data_stage_4__2941_,data_stage_4__2940_,data_stage_4__2939_,data_stage_4__2938_,
  data_stage_4__2937_,data_stage_4__2936_,data_stage_4__2935_,data_stage_4__2934_,
  data_stage_4__2933_,data_stage_4__2932_,data_stage_4__2931_,data_stage_4__2930_,
  data_stage_4__2929_,data_stage_4__2928_,data_stage_4__2927_,data_stage_4__2926_,
  data_stage_4__2925_,data_stage_4__2924_,data_stage_4__2923_,data_stage_4__2922_,
  data_stage_4__2921_,data_stage_4__2920_,data_stage_4__2919_,data_stage_4__2918_,
  data_stage_4__2917_,data_stage_4__2916_,data_stage_4__2915_,data_stage_4__2914_,
  data_stage_4__2913_,data_stage_4__2912_,data_stage_4__2911_,data_stage_4__2910_,
  data_stage_4__2909_,data_stage_4__2908_,data_stage_4__2907_,data_stage_4__2906_,
  data_stage_4__2905_,data_stage_4__2904_,data_stage_4__2903_,data_stage_4__2902_,
  data_stage_4__2901_,data_stage_4__2900_,data_stage_4__2899_,data_stage_4__2898_,
  data_stage_4__2897_,data_stage_4__2896_,data_stage_4__2895_,data_stage_4__2894_,
  data_stage_4__2893_,data_stage_4__2892_,data_stage_4__2891_,data_stage_4__2890_,
  data_stage_4__2889_,data_stage_4__2888_,data_stage_4__2887_,data_stage_4__2886_,
  data_stage_4__2885_,data_stage_4__2884_,data_stage_4__2883_,data_stage_4__2882_,
  data_stage_4__2881_,data_stage_4__2880_,data_stage_4__2879_,data_stage_4__2878_,
  data_stage_4__2877_,data_stage_4__2876_,data_stage_4__2875_,data_stage_4__2874_,
  data_stage_4__2873_,data_stage_4__2872_,data_stage_4__2871_,data_stage_4__2870_,
  data_stage_4__2869_,data_stage_4__2868_,data_stage_4__2867_,data_stage_4__2866_,
  data_stage_4__2865_,data_stage_4__2864_,data_stage_4__2863_,data_stage_4__2862_,
  data_stage_4__2861_,data_stage_4__2860_,data_stage_4__2859_,data_stage_4__2858_,
  data_stage_4__2857_,data_stage_4__2856_,data_stage_4__2855_,data_stage_4__2854_,
  data_stage_4__2853_,data_stage_4__2852_,data_stage_4__2851_,data_stage_4__2850_,
  data_stage_4__2849_,data_stage_4__2848_,data_stage_4__2847_,data_stage_4__2846_,
  data_stage_4__2845_,data_stage_4__2844_,data_stage_4__2843_,data_stage_4__2842_,
  data_stage_4__2841_,data_stage_4__2840_,data_stage_4__2839_,data_stage_4__2838_,
  data_stage_4__2837_,data_stage_4__2836_,data_stage_4__2835_,data_stage_4__2834_,
  data_stage_4__2833_,data_stage_4__2832_,data_stage_4__2831_,data_stage_4__2830_,
  data_stage_4__2829_,data_stage_4__2828_,data_stage_4__2827_,data_stage_4__2826_,
  data_stage_4__2825_,data_stage_4__2824_,data_stage_4__2823_,data_stage_4__2822_,
  data_stage_4__2821_,data_stage_4__2820_,data_stage_4__2819_,data_stage_4__2818_,
  data_stage_4__2817_,data_stage_4__2816_,data_stage_4__2815_,data_stage_4__2814_,
  data_stage_4__2813_,data_stage_4__2812_,data_stage_4__2811_,data_stage_4__2810_,
  data_stage_4__2809_,data_stage_4__2808_,data_stage_4__2807_,data_stage_4__2806_,
  data_stage_4__2805_,data_stage_4__2804_,data_stage_4__2803_,data_stage_4__2802_,
  data_stage_4__2801_,data_stage_4__2800_,data_stage_4__2799_,data_stage_4__2798_,
  data_stage_4__2797_,data_stage_4__2796_,data_stage_4__2795_,data_stage_4__2794_,
  data_stage_4__2793_,data_stage_4__2792_,data_stage_4__2791_,data_stage_4__2790_,
  data_stage_4__2789_,data_stage_4__2788_,data_stage_4__2787_,data_stage_4__2786_,
  data_stage_4__2785_,data_stage_4__2784_,data_stage_4__2783_,data_stage_4__2782_,
  data_stage_4__2781_,data_stage_4__2780_,data_stage_4__2779_,data_stage_4__2778_,
  data_stage_4__2777_,data_stage_4__2776_,data_stage_4__2775_,data_stage_4__2774_,
  data_stage_4__2773_,data_stage_4__2772_,data_stage_4__2771_,data_stage_4__2770_,
  data_stage_4__2769_,data_stage_4__2768_,data_stage_4__2767_,data_stage_4__2766_,
  data_stage_4__2765_,data_stage_4__2764_,data_stage_4__2763_,data_stage_4__2762_,
  data_stage_4__2761_,data_stage_4__2760_,data_stage_4__2759_,data_stage_4__2758_,
  data_stage_4__2757_,data_stage_4__2756_,data_stage_4__2755_,data_stage_4__2754_,
  data_stage_4__2753_,data_stage_4__2752_,data_stage_4__2751_,data_stage_4__2750_,
  data_stage_4__2749_,data_stage_4__2748_,data_stage_4__2747_,data_stage_4__2746_,
  data_stage_4__2745_,data_stage_4__2744_,data_stage_4__2743_,data_stage_4__2742_,
  data_stage_4__2741_,data_stage_4__2740_,data_stage_4__2739_,data_stage_4__2738_,
  data_stage_4__2737_,data_stage_4__2736_,data_stage_4__2735_,data_stage_4__2734_,
  data_stage_4__2733_,data_stage_4__2732_,data_stage_4__2731_,data_stage_4__2730_,
  data_stage_4__2729_,data_stage_4__2728_,data_stage_4__2727_,data_stage_4__2726_,
  data_stage_4__2725_,data_stage_4__2724_,data_stage_4__2723_,data_stage_4__2722_,
  data_stage_4__2721_,data_stage_4__2720_,data_stage_4__2719_,data_stage_4__2718_,
  data_stage_4__2717_,data_stage_4__2716_,data_stage_4__2715_,data_stage_4__2714_,
  data_stage_4__2713_,data_stage_4__2712_,data_stage_4__2711_,data_stage_4__2710_,
  data_stage_4__2709_,data_stage_4__2708_,data_stage_4__2707_,data_stage_4__2706_,
  data_stage_4__2705_,data_stage_4__2704_,data_stage_4__2703_,data_stage_4__2702_,
  data_stage_4__2701_,data_stage_4__2700_,data_stage_4__2699_,data_stage_4__2698_,
  data_stage_4__2697_,data_stage_4__2696_,data_stage_4__2695_,data_stage_4__2694_,
  data_stage_4__2693_,data_stage_4__2692_,data_stage_4__2691_,data_stage_4__2690_,
  data_stage_4__2689_,data_stage_4__2688_,data_stage_4__2687_,data_stage_4__2686_,
  data_stage_4__2685_,data_stage_4__2684_,data_stage_4__2683_,data_stage_4__2682_,
  data_stage_4__2681_,data_stage_4__2680_,data_stage_4__2679_,data_stage_4__2678_,
  data_stage_4__2677_,data_stage_4__2676_,data_stage_4__2675_,data_stage_4__2674_,
  data_stage_4__2673_,data_stage_4__2672_,data_stage_4__2671_,data_stage_4__2670_,
  data_stage_4__2669_,data_stage_4__2668_,data_stage_4__2667_,data_stage_4__2666_,
  data_stage_4__2665_,data_stage_4__2664_,data_stage_4__2663_,data_stage_4__2662_,
  data_stage_4__2661_,data_stage_4__2660_,data_stage_4__2659_,data_stage_4__2658_,
  data_stage_4__2657_,data_stage_4__2656_,data_stage_4__2655_,data_stage_4__2654_,
  data_stage_4__2653_,data_stage_4__2652_,data_stage_4__2651_,data_stage_4__2650_,
  data_stage_4__2649_,data_stage_4__2648_,data_stage_4__2647_,data_stage_4__2646_,
  data_stage_4__2645_,data_stage_4__2644_,data_stage_4__2643_,data_stage_4__2642_,
  data_stage_4__2641_,data_stage_4__2640_,data_stage_4__2639_,data_stage_4__2638_,
  data_stage_4__2637_,data_stage_4__2636_,data_stage_4__2635_,data_stage_4__2634_,
  data_stage_4__2633_,data_stage_4__2632_,data_stage_4__2631_,data_stage_4__2630_,
  data_stage_4__2629_,data_stage_4__2628_,data_stage_4__2627_,data_stage_4__2626_,
  data_stage_4__2625_,data_stage_4__2624_,data_stage_4__2623_,data_stage_4__2622_,
  data_stage_4__2621_,data_stage_4__2620_,data_stage_4__2619_,data_stage_4__2618_,
  data_stage_4__2617_,data_stage_4__2616_,data_stage_4__2615_,data_stage_4__2614_,
  data_stage_4__2613_,data_stage_4__2612_,data_stage_4__2611_,data_stage_4__2610_,
  data_stage_4__2609_,data_stage_4__2608_,data_stage_4__2607_,data_stage_4__2606_,
  data_stage_4__2605_,data_stage_4__2604_,data_stage_4__2603_,data_stage_4__2602_,
  data_stage_4__2601_,data_stage_4__2600_,data_stage_4__2599_,data_stage_4__2598_,
  data_stage_4__2597_,data_stage_4__2596_,data_stage_4__2595_,data_stage_4__2594_,
  data_stage_4__2593_,data_stage_4__2592_,data_stage_4__2591_,data_stage_4__2590_,
  data_stage_4__2589_,data_stage_4__2588_,data_stage_4__2587_,data_stage_4__2586_,
  data_stage_4__2585_,data_stage_4__2584_,data_stage_4__2583_,data_stage_4__2582_,
  data_stage_4__2581_,data_stage_4__2580_,data_stage_4__2579_,data_stage_4__2578_,
  data_stage_4__2577_,data_stage_4__2576_,data_stage_4__2575_,data_stage_4__2574_,
  data_stage_4__2573_,data_stage_4__2572_,data_stage_4__2571_,data_stage_4__2570_,
  data_stage_4__2569_,data_stage_4__2568_,data_stage_4__2567_,data_stage_4__2566_,
  data_stage_4__2565_,data_stage_4__2564_,data_stage_4__2563_,data_stage_4__2562_,
  data_stage_4__2561_,data_stage_4__2560_,data_stage_4__2559_,data_stage_4__2558_,
  data_stage_4__2557_,data_stage_4__2556_,data_stage_4__2555_,data_stage_4__2554_,
  data_stage_4__2553_,data_stage_4__2552_,data_stage_4__2551_,data_stage_4__2550_,
  data_stage_4__2549_,data_stage_4__2548_,data_stage_4__2547_,data_stage_4__2546_,
  data_stage_4__2545_,data_stage_4__2544_,data_stage_4__2543_,data_stage_4__2542_,
  data_stage_4__2541_,data_stage_4__2540_,data_stage_4__2539_,data_stage_4__2538_,
  data_stage_4__2537_,data_stage_4__2536_,data_stage_4__2535_,data_stage_4__2534_,
  data_stage_4__2533_,data_stage_4__2532_,data_stage_4__2531_,data_stage_4__2530_,
  data_stage_4__2529_,data_stage_4__2528_,data_stage_4__2527_,data_stage_4__2526_,
  data_stage_4__2525_,data_stage_4__2524_,data_stage_4__2523_,data_stage_4__2522_,
  data_stage_4__2521_,data_stage_4__2520_,data_stage_4__2519_,data_stage_4__2518_,
  data_stage_4__2517_,data_stage_4__2516_,data_stage_4__2515_,data_stage_4__2514_,
  data_stage_4__2513_,data_stage_4__2512_,data_stage_4__2511_,data_stage_4__2510_,
  data_stage_4__2509_,data_stage_4__2508_,data_stage_4__2507_,data_stage_4__2506_,
  data_stage_4__2505_,data_stage_4__2504_,data_stage_4__2503_,data_stage_4__2502_,
  data_stage_4__2501_,data_stage_4__2500_,data_stage_4__2499_,data_stage_4__2498_,
  data_stage_4__2497_,data_stage_4__2496_,data_stage_4__2495_,data_stage_4__2494_,
  data_stage_4__2493_,data_stage_4__2492_,data_stage_4__2491_,data_stage_4__2490_,
  data_stage_4__2489_,data_stage_4__2488_,data_stage_4__2487_,data_stage_4__2486_,
  data_stage_4__2485_,data_stage_4__2484_,data_stage_4__2483_,data_stage_4__2482_,
  data_stage_4__2481_,data_stage_4__2480_,data_stage_4__2479_,data_stage_4__2478_,
  data_stage_4__2477_,data_stage_4__2476_,data_stage_4__2475_,data_stage_4__2474_,
  data_stage_4__2473_,data_stage_4__2472_,data_stage_4__2471_,data_stage_4__2470_,
  data_stage_4__2469_,data_stage_4__2468_,data_stage_4__2467_,data_stage_4__2466_,
  data_stage_4__2465_,data_stage_4__2464_,data_stage_4__2463_,data_stage_4__2462_,
  data_stage_4__2461_,data_stage_4__2460_,data_stage_4__2459_,data_stage_4__2458_,
  data_stage_4__2457_,data_stage_4__2456_,data_stage_4__2455_,data_stage_4__2454_,
  data_stage_4__2453_,data_stage_4__2452_,data_stage_4__2451_,data_stage_4__2450_,
  data_stage_4__2449_,data_stage_4__2448_,data_stage_4__2447_,data_stage_4__2446_,
  data_stage_4__2445_,data_stage_4__2444_,data_stage_4__2443_,data_stage_4__2442_,
  data_stage_4__2441_,data_stage_4__2440_,data_stage_4__2439_,data_stage_4__2438_,
  data_stage_4__2437_,data_stage_4__2436_,data_stage_4__2435_,data_stage_4__2434_,
  data_stage_4__2433_,data_stage_4__2432_,data_stage_4__2431_,data_stage_4__2430_,
  data_stage_4__2429_,data_stage_4__2428_,data_stage_4__2427_,data_stage_4__2426_,
  data_stage_4__2425_,data_stage_4__2424_,data_stage_4__2423_,data_stage_4__2422_,
  data_stage_4__2421_,data_stage_4__2420_,data_stage_4__2419_,data_stage_4__2418_,
  data_stage_4__2417_,data_stage_4__2416_,data_stage_4__2415_,data_stage_4__2414_,
  data_stage_4__2413_,data_stage_4__2412_,data_stage_4__2411_,data_stage_4__2410_,
  data_stage_4__2409_,data_stage_4__2408_,data_stage_4__2407_,data_stage_4__2406_,
  data_stage_4__2405_,data_stage_4__2404_,data_stage_4__2403_,data_stage_4__2402_,
  data_stage_4__2401_,data_stage_4__2400_,data_stage_4__2399_,data_stage_4__2398_,
  data_stage_4__2397_,data_stage_4__2396_,data_stage_4__2395_,data_stage_4__2394_,
  data_stage_4__2393_,data_stage_4__2392_,data_stage_4__2391_,data_stage_4__2390_,
  data_stage_4__2389_,data_stage_4__2388_,data_stage_4__2387_,data_stage_4__2386_,
  data_stage_4__2385_,data_stage_4__2384_,data_stage_4__2383_,data_stage_4__2382_,
  data_stage_4__2381_,data_stage_4__2380_,data_stage_4__2379_,data_stage_4__2378_,
  data_stage_4__2377_,data_stage_4__2376_,data_stage_4__2375_,data_stage_4__2374_,
  data_stage_4__2373_,data_stage_4__2372_,data_stage_4__2371_,data_stage_4__2370_,
  data_stage_4__2369_,data_stage_4__2368_,data_stage_4__2367_,data_stage_4__2366_,
  data_stage_4__2365_,data_stage_4__2364_,data_stage_4__2363_,data_stage_4__2362_,
  data_stage_4__2361_,data_stage_4__2360_,data_stage_4__2359_,data_stage_4__2358_,
  data_stage_4__2357_,data_stage_4__2356_,data_stage_4__2355_,data_stage_4__2354_,
  data_stage_4__2353_,data_stage_4__2352_,data_stage_4__2351_,data_stage_4__2350_,
  data_stage_4__2349_,data_stage_4__2348_,data_stage_4__2347_,data_stage_4__2346_,
  data_stage_4__2345_,data_stage_4__2344_,data_stage_4__2343_,data_stage_4__2342_,
  data_stage_4__2341_,data_stage_4__2340_,data_stage_4__2339_,data_stage_4__2338_,
  data_stage_4__2337_,data_stage_4__2336_,data_stage_4__2335_,data_stage_4__2334_,
  data_stage_4__2333_,data_stage_4__2332_,data_stage_4__2331_,data_stage_4__2330_,
  data_stage_4__2329_,data_stage_4__2328_,data_stage_4__2327_,data_stage_4__2326_,
  data_stage_4__2325_,data_stage_4__2324_,data_stage_4__2323_,data_stage_4__2322_,
  data_stage_4__2321_,data_stage_4__2320_,data_stage_4__2319_,data_stage_4__2318_,
  data_stage_4__2317_,data_stage_4__2316_,data_stage_4__2315_,data_stage_4__2314_,
  data_stage_4__2313_,data_stage_4__2312_,data_stage_4__2311_,data_stage_4__2310_,
  data_stage_4__2309_,data_stage_4__2308_,data_stage_4__2307_,data_stage_4__2306_,
  data_stage_4__2305_,data_stage_4__2304_,data_stage_4__2303_,data_stage_4__2302_,
  data_stage_4__2301_,data_stage_4__2300_,data_stage_4__2299_,data_stage_4__2298_,
  data_stage_4__2297_,data_stage_4__2296_,data_stage_4__2295_,data_stage_4__2294_,
  data_stage_4__2293_,data_stage_4__2292_,data_stage_4__2291_,data_stage_4__2290_,
  data_stage_4__2289_,data_stage_4__2288_,data_stage_4__2287_,data_stage_4__2286_,
  data_stage_4__2285_,data_stage_4__2284_,data_stage_4__2283_,data_stage_4__2282_,
  data_stage_4__2281_,data_stage_4__2280_,data_stage_4__2279_,data_stage_4__2278_,
  data_stage_4__2277_,data_stage_4__2276_,data_stage_4__2275_,data_stage_4__2274_,
  data_stage_4__2273_,data_stage_4__2272_,data_stage_4__2271_,data_stage_4__2270_,
  data_stage_4__2269_,data_stage_4__2268_,data_stage_4__2267_,data_stage_4__2266_,
  data_stage_4__2265_,data_stage_4__2264_,data_stage_4__2263_,data_stage_4__2262_,
  data_stage_4__2261_,data_stage_4__2260_,data_stage_4__2259_,data_stage_4__2258_,
  data_stage_4__2257_,data_stage_4__2256_,data_stage_4__2255_,data_stage_4__2254_,
  data_stage_4__2253_,data_stage_4__2252_,data_stage_4__2251_,data_stage_4__2250_,
  data_stage_4__2249_,data_stage_4__2248_,data_stage_4__2247_,data_stage_4__2246_,
  data_stage_4__2245_,data_stage_4__2244_,data_stage_4__2243_,data_stage_4__2242_,
  data_stage_4__2241_,data_stage_4__2240_,data_stage_4__2239_,data_stage_4__2238_,
  data_stage_4__2237_,data_stage_4__2236_,data_stage_4__2235_,data_stage_4__2234_,
  data_stage_4__2233_,data_stage_4__2232_,data_stage_4__2231_,data_stage_4__2230_,
  data_stage_4__2229_,data_stage_4__2228_,data_stage_4__2227_,data_stage_4__2226_,
  data_stage_4__2225_,data_stage_4__2224_,data_stage_4__2223_,data_stage_4__2222_,
  data_stage_4__2221_,data_stage_4__2220_,data_stage_4__2219_,data_stage_4__2218_,
  data_stage_4__2217_,data_stage_4__2216_,data_stage_4__2215_,data_stage_4__2214_,
  data_stage_4__2213_,data_stage_4__2212_,data_stage_4__2211_,data_stage_4__2210_,
  data_stage_4__2209_,data_stage_4__2208_,data_stage_4__2207_,data_stage_4__2206_,
  data_stage_4__2205_,data_stage_4__2204_,data_stage_4__2203_,data_stage_4__2202_,
  data_stage_4__2201_,data_stage_4__2200_,data_stage_4__2199_,data_stage_4__2198_,
  data_stage_4__2197_,data_stage_4__2196_,data_stage_4__2195_,data_stage_4__2194_,
  data_stage_4__2193_,data_stage_4__2192_,data_stage_4__2191_,data_stage_4__2190_,
  data_stage_4__2189_,data_stage_4__2188_,data_stage_4__2187_,data_stage_4__2186_,
  data_stage_4__2185_,data_stage_4__2184_,data_stage_4__2183_,data_stage_4__2182_,
  data_stage_4__2181_,data_stage_4__2180_,data_stage_4__2179_,data_stage_4__2178_,
  data_stage_4__2177_,data_stage_4__2176_,data_stage_4__2175_,data_stage_4__2174_,
  data_stage_4__2173_,data_stage_4__2172_,data_stage_4__2171_,data_stage_4__2170_,
  data_stage_4__2169_,data_stage_4__2168_,data_stage_4__2167_,data_stage_4__2166_,
  data_stage_4__2165_,data_stage_4__2164_,data_stage_4__2163_,data_stage_4__2162_,
  data_stage_4__2161_,data_stage_4__2160_,data_stage_4__2159_,data_stage_4__2158_,
  data_stage_4__2157_,data_stage_4__2156_,data_stage_4__2155_,data_stage_4__2154_,
  data_stage_4__2153_,data_stage_4__2152_,data_stage_4__2151_,data_stage_4__2150_,
  data_stage_4__2149_,data_stage_4__2148_,data_stage_4__2147_,data_stage_4__2146_,
  data_stage_4__2145_,data_stage_4__2144_,data_stage_4__2143_,data_stage_4__2142_,
  data_stage_4__2141_,data_stage_4__2140_,data_stage_4__2139_,data_stage_4__2138_,
  data_stage_4__2137_,data_stage_4__2136_,data_stage_4__2135_,data_stage_4__2134_,
  data_stage_4__2133_,data_stage_4__2132_,data_stage_4__2131_,data_stage_4__2130_,
  data_stage_4__2129_,data_stage_4__2128_,data_stage_4__2127_,data_stage_4__2126_,
  data_stage_4__2125_,data_stage_4__2124_,data_stage_4__2123_,data_stage_4__2122_,
  data_stage_4__2121_,data_stage_4__2120_,data_stage_4__2119_,data_stage_4__2118_,
  data_stage_4__2117_,data_stage_4__2116_,data_stage_4__2115_,data_stage_4__2114_,
  data_stage_4__2113_,data_stage_4__2112_,data_stage_4__2111_,data_stage_4__2110_,
  data_stage_4__2109_,data_stage_4__2108_,data_stage_4__2107_,data_stage_4__2106_,
  data_stage_4__2105_,data_stage_4__2104_,data_stage_4__2103_,data_stage_4__2102_,
  data_stage_4__2101_,data_stage_4__2100_,data_stage_4__2099_,data_stage_4__2098_,
  data_stage_4__2097_,data_stage_4__2096_,data_stage_4__2095_,data_stage_4__2094_,
  data_stage_4__2093_,data_stage_4__2092_,data_stage_4__2091_,data_stage_4__2090_,
  data_stage_4__2089_,data_stage_4__2088_,data_stage_4__2087_,data_stage_4__2086_,
  data_stage_4__2085_,data_stage_4__2084_,data_stage_4__2083_,data_stage_4__2082_,
  data_stage_4__2081_,data_stage_4__2080_,data_stage_4__2079_,data_stage_4__2078_,
  data_stage_4__2077_,data_stage_4__2076_,data_stage_4__2075_,data_stage_4__2074_,
  data_stage_4__2073_,data_stage_4__2072_,data_stage_4__2071_,data_stage_4__2070_,
  data_stage_4__2069_,data_stage_4__2068_,data_stage_4__2067_,data_stage_4__2066_,
  data_stage_4__2065_,data_stage_4__2064_,data_stage_4__2063_,data_stage_4__2062_,
  data_stage_4__2061_,data_stage_4__2060_,data_stage_4__2059_,data_stage_4__2058_,
  data_stage_4__2057_,data_stage_4__2056_,data_stage_4__2055_,data_stage_4__2054_,
  data_stage_4__2053_,data_stage_4__2052_,data_stage_4__2051_,data_stage_4__2050_,
  data_stage_4__2049_,data_stage_4__2048_,data_stage_4__2047_,data_stage_4__2046_,
  data_stage_4__2045_,data_stage_4__2044_,data_stage_4__2043_,data_stage_4__2042_,
  data_stage_4__2041_,data_stage_4__2040_,data_stage_4__2039_,data_stage_4__2038_,
  data_stage_4__2037_,data_stage_4__2036_,data_stage_4__2035_,data_stage_4__2034_,
  data_stage_4__2033_,data_stage_4__2032_,data_stage_4__2031_,data_stage_4__2030_,
  data_stage_4__2029_,data_stage_4__2028_,data_stage_4__2027_,data_stage_4__2026_,
  data_stage_4__2025_,data_stage_4__2024_,data_stage_4__2023_,data_stage_4__2022_,
  data_stage_4__2021_,data_stage_4__2020_,data_stage_4__2019_,data_stage_4__2018_,
  data_stage_4__2017_,data_stage_4__2016_,data_stage_4__2015_,data_stage_4__2014_,
  data_stage_4__2013_,data_stage_4__2012_,data_stage_4__2011_,data_stage_4__2010_,
  data_stage_4__2009_,data_stage_4__2008_,data_stage_4__2007_,data_stage_4__2006_,
  data_stage_4__2005_,data_stage_4__2004_,data_stage_4__2003_,data_stage_4__2002_,
  data_stage_4__2001_,data_stage_4__2000_,data_stage_4__1999_,data_stage_4__1998_,
  data_stage_4__1997_,data_stage_4__1996_,data_stage_4__1995_,data_stage_4__1994_,
  data_stage_4__1993_,data_stage_4__1992_,data_stage_4__1991_,data_stage_4__1990_,
  data_stage_4__1989_,data_stage_4__1988_,data_stage_4__1987_,data_stage_4__1986_,
  data_stage_4__1985_,data_stage_4__1984_,data_stage_4__1983_,data_stage_4__1982_,
  data_stage_4__1981_,data_stage_4__1980_,data_stage_4__1979_,data_stage_4__1978_,
  data_stage_4__1977_,data_stage_4__1976_,data_stage_4__1975_,data_stage_4__1974_,
  data_stage_4__1973_,data_stage_4__1972_,data_stage_4__1971_,data_stage_4__1970_,
  data_stage_4__1969_,data_stage_4__1968_,data_stage_4__1967_,data_stage_4__1966_,
  data_stage_4__1965_,data_stage_4__1964_,data_stage_4__1963_,data_stage_4__1962_,
  data_stage_4__1961_,data_stage_4__1960_,data_stage_4__1959_,data_stage_4__1958_,
  data_stage_4__1957_,data_stage_4__1956_,data_stage_4__1955_,data_stage_4__1954_,
  data_stage_4__1953_,data_stage_4__1952_,data_stage_4__1951_,data_stage_4__1950_,
  data_stage_4__1949_,data_stage_4__1948_,data_stage_4__1947_,data_stage_4__1946_,
  data_stage_4__1945_,data_stage_4__1944_,data_stage_4__1943_,data_stage_4__1942_,
  data_stage_4__1941_,data_stage_4__1940_,data_stage_4__1939_,data_stage_4__1938_,
  data_stage_4__1937_,data_stage_4__1936_,data_stage_4__1935_,data_stage_4__1934_,
  data_stage_4__1933_,data_stage_4__1932_,data_stage_4__1931_,data_stage_4__1930_,
  data_stage_4__1929_,data_stage_4__1928_,data_stage_4__1927_,data_stage_4__1926_,
  data_stage_4__1925_,data_stage_4__1924_,data_stage_4__1923_,data_stage_4__1922_,
  data_stage_4__1921_,data_stage_4__1920_,data_stage_4__1919_,data_stage_4__1918_,
  data_stage_4__1917_,data_stage_4__1916_,data_stage_4__1915_,data_stage_4__1914_,
  data_stage_4__1913_,data_stage_4__1912_,data_stage_4__1911_,data_stage_4__1910_,
  data_stage_4__1909_,data_stage_4__1908_,data_stage_4__1907_,data_stage_4__1906_,
  data_stage_4__1905_,data_stage_4__1904_,data_stage_4__1903_,data_stage_4__1902_,
  data_stage_4__1901_,data_stage_4__1900_,data_stage_4__1899_,data_stage_4__1898_,
  data_stage_4__1897_,data_stage_4__1896_,data_stage_4__1895_,data_stage_4__1894_,
  data_stage_4__1893_,data_stage_4__1892_,data_stage_4__1891_,data_stage_4__1890_,
  data_stage_4__1889_,data_stage_4__1888_,data_stage_4__1887_,data_stage_4__1886_,
  data_stage_4__1885_,data_stage_4__1884_,data_stage_4__1883_,data_stage_4__1882_,
  data_stage_4__1881_,data_stage_4__1880_,data_stage_4__1879_,data_stage_4__1878_,
  data_stage_4__1877_,data_stage_4__1876_,data_stage_4__1875_,data_stage_4__1874_,
  data_stage_4__1873_,data_stage_4__1872_,data_stage_4__1871_,data_stage_4__1870_,
  data_stage_4__1869_,data_stage_4__1868_,data_stage_4__1867_,data_stage_4__1866_,
  data_stage_4__1865_,data_stage_4__1864_,data_stage_4__1863_,data_stage_4__1862_,
  data_stage_4__1861_,data_stage_4__1860_,data_stage_4__1859_,data_stage_4__1858_,
  data_stage_4__1857_,data_stage_4__1856_,data_stage_4__1855_,data_stage_4__1854_,
  data_stage_4__1853_,data_stage_4__1852_,data_stage_4__1851_,data_stage_4__1850_,
  data_stage_4__1849_,data_stage_4__1848_,data_stage_4__1847_,data_stage_4__1846_,
  data_stage_4__1845_,data_stage_4__1844_,data_stage_4__1843_,data_stage_4__1842_,
  data_stage_4__1841_,data_stage_4__1840_,data_stage_4__1839_,data_stage_4__1838_,
  data_stage_4__1837_,data_stage_4__1836_,data_stage_4__1835_,data_stage_4__1834_,
  data_stage_4__1833_,data_stage_4__1832_,data_stage_4__1831_,data_stage_4__1830_,
  data_stage_4__1829_,data_stage_4__1828_,data_stage_4__1827_,data_stage_4__1826_,
  data_stage_4__1825_,data_stage_4__1824_,data_stage_4__1823_,data_stage_4__1822_,
  data_stage_4__1821_,data_stage_4__1820_,data_stage_4__1819_,data_stage_4__1818_,
  data_stage_4__1817_,data_stage_4__1816_,data_stage_4__1815_,data_stage_4__1814_,
  data_stage_4__1813_,data_stage_4__1812_,data_stage_4__1811_,data_stage_4__1810_,
  data_stage_4__1809_,data_stage_4__1808_,data_stage_4__1807_,data_stage_4__1806_,
  data_stage_4__1805_,data_stage_4__1804_,data_stage_4__1803_,data_stage_4__1802_,
  data_stage_4__1801_,data_stage_4__1800_,data_stage_4__1799_,data_stage_4__1798_,
  data_stage_4__1797_,data_stage_4__1796_,data_stage_4__1795_,data_stage_4__1794_,
  data_stage_4__1793_,data_stage_4__1792_,data_stage_4__1791_,data_stage_4__1790_,
  data_stage_4__1789_,data_stage_4__1788_,data_stage_4__1787_,data_stage_4__1786_,
  data_stage_4__1785_,data_stage_4__1784_,data_stage_4__1783_,data_stage_4__1782_,
  data_stage_4__1781_,data_stage_4__1780_,data_stage_4__1779_,data_stage_4__1778_,
  data_stage_4__1777_,data_stage_4__1776_,data_stage_4__1775_,data_stage_4__1774_,
  data_stage_4__1773_,data_stage_4__1772_,data_stage_4__1771_,data_stage_4__1770_,
  data_stage_4__1769_,data_stage_4__1768_,data_stage_4__1767_,data_stage_4__1766_,
  data_stage_4__1765_,data_stage_4__1764_,data_stage_4__1763_,data_stage_4__1762_,
  data_stage_4__1761_,data_stage_4__1760_,data_stage_4__1759_,data_stage_4__1758_,
  data_stage_4__1757_,data_stage_4__1756_,data_stage_4__1755_,data_stage_4__1754_,
  data_stage_4__1753_,data_stage_4__1752_,data_stage_4__1751_,data_stage_4__1750_,
  data_stage_4__1749_,data_stage_4__1748_,data_stage_4__1747_,data_stage_4__1746_,
  data_stage_4__1745_,data_stage_4__1744_,data_stage_4__1743_,data_stage_4__1742_,
  data_stage_4__1741_,data_stage_4__1740_,data_stage_4__1739_,data_stage_4__1738_,
  data_stage_4__1737_,data_stage_4__1736_,data_stage_4__1735_,data_stage_4__1734_,
  data_stage_4__1733_,data_stage_4__1732_,data_stage_4__1731_,data_stage_4__1730_,
  data_stage_4__1729_,data_stage_4__1728_,data_stage_4__1727_,data_stage_4__1726_,
  data_stage_4__1725_,data_stage_4__1724_,data_stage_4__1723_,data_stage_4__1722_,
  data_stage_4__1721_,data_stage_4__1720_,data_stage_4__1719_,data_stage_4__1718_,
  data_stage_4__1717_,data_stage_4__1716_,data_stage_4__1715_,data_stage_4__1714_,
  data_stage_4__1713_,data_stage_4__1712_,data_stage_4__1711_,data_stage_4__1710_,
  data_stage_4__1709_,data_stage_4__1708_,data_stage_4__1707_,data_stage_4__1706_,
  data_stage_4__1705_,data_stage_4__1704_,data_stage_4__1703_,data_stage_4__1702_,
  data_stage_4__1701_,data_stage_4__1700_,data_stage_4__1699_,data_stage_4__1698_,
  data_stage_4__1697_,data_stage_4__1696_,data_stage_4__1695_,data_stage_4__1694_,
  data_stage_4__1693_,data_stage_4__1692_,data_stage_4__1691_,data_stage_4__1690_,
  data_stage_4__1689_,data_stage_4__1688_,data_stage_4__1687_,data_stage_4__1686_,
  data_stage_4__1685_,data_stage_4__1684_,data_stage_4__1683_,data_stage_4__1682_,
  data_stage_4__1681_,data_stage_4__1680_,data_stage_4__1679_,data_stage_4__1678_,
  data_stage_4__1677_,data_stage_4__1676_,data_stage_4__1675_,data_stage_4__1674_,
  data_stage_4__1673_,data_stage_4__1672_,data_stage_4__1671_,data_stage_4__1670_,
  data_stage_4__1669_,data_stage_4__1668_,data_stage_4__1667_,data_stage_4__1666_,
  data_stage_4__1665_,data_stage_4__1664_,data_stage_4__1663_,data_stage_4__1662_,
  data_stage_4__1661_,data_stage_4__1660_,data_stage_4__1659_,data_stage_4__1658_,
  data_stage_4__1657_,data_stage_4__1656_,data_stage_4__1655_,data_stage_4__1654_,
  data_stage_4__1653_,data_stage_4__1652_,data_stage_4__1651_,data_stage_4__1650_,
  data_stage_4__1649_,data_stage_4__1648_,data_stage_4__1647_,data_stage_4__1646_,
  data_stage_4__1645_,data_stage_4__1644_,data_stage_4__1643_,data_stage_4__1642_,
  data_stage_4__1641_,data_stage_4__1640_,data_stage_4__1639_,data_stage_4__1638_,
  data_stage_4__1637_,data_stage_4__1636_,data_stage_4__1635_,data_stage_4__1634_,
  data_stage_4__1633_,data_stage_4__1632_,data_stage_4__1631_,data_stage_4__1630_,
  data_stage_4__1629_,data_stage_4__1628_,data_stage_4__1627_,data_stage_4__1626_,
  data_stage_4__1625_,data_stage_4__1624_,data_stage_4__1623_,data_stage_4__1622_,
  data_stage_4__1621_,data_stage_4__1620_,data_stage_4__1619_,data_stage_4__1618_,
  data_stage_4__1617_,data_stage_4__1616_,data_stage_4__1615_,data_stage_4__1614_,
  data_stage_4__1613_,data_stage_4__1612_,data_stage_4__1611_,data_stage_4__1610_,
  data_stage_4__1609_,data_stage_4__1608_,data_stage_4__1607_,data_stage_4__1606_,
  data_stage_4__1605_,data_stage_4__1604_,data_stage_4__1603_,data_stage_4__1602_,
  data_stage_4__1601_,data_stage_4__1600_,data_stage_4__1599_,data_stage_4__1598_,
  data_stage_4__1597_,data_stage_4__1596_,data_stage_4__1595_,data_stage_4__1594_,
  data_stage_4__1593_,data_stage_4__1592_,data_stage_4__1591_,data_stage_4__1590_,
  data_stage_4__1589_,data_stage_4__1588_,data_stage_4__1587_,data_stage_4__1586_,
  data_stage_4__1585_,data_stage_4__1584_,data_stage_4__1583_,data_stage_4__1582_,
  data_stage_4__1581_,data_stage_4__1580_,data_stage_4__1579_,data_stage_4__1578_,
  data_stage_4__1577_,data_stage_4__1576_,data_stage_4__1575_,data_stage_4__1574_,
  data_stage_4__1573_,data_stage_4__1572_,data_stage_4__1571_,data_stage_4__1570_,
  data_stage_4__1569_,data_stage_4__1568_,data_stage_4__1567_,data_stage_4__1566_,
  data_stage_4__1565_,data_stage_4__1564_,data_stage_4__1563_,data_stage_4__1562_,
  data_stage_4__1561_,data_stage_4__1560_,data_stage_4__1559_,data_stage_4__1558_,
  data_stage_4__1557_,data_stage_4__1556_,data_stage_4__1555_,data_stage_4__1554_,
  data_stage_4__1553_,data_stage_4__1552_,data_stage_4__1551_,data_stage_4__1550_,
  data_stage_4__1549_,data_stage_4__1548_,data_stage_4__1547_,data_stage_4__1546_,
  data_stage_4__1545_,data_stage_4__1544_,data_stage_4__1543_,data_stage_4__1542_,
  data_stage_4__1541_,data_stage_4__1540_,data_stage_4__1539_,data_stage_4__1538_,
  data_stage_4__1537_,data_stage_4__1536_,data_stage_4__1535_,data_stage_4__1534_,
  data_stage_4__1533_,data_stage_4__1532_,data_stage_4__1531_,data_stage_4__1530_,
  data_stage_4__1529_,data_stage_4__1528_,data_stage_4__1527_,data_stage_4__1526_,
  data_stage_4__1525_,data_stage_4__1524_,data_stage_4__1523_,data_stage_4__1522_,
  data_stage_4__1521_,data_stage_4__1520_,data_stage_4__1519_,data_stage_4__1518_,
  data_stage_4__1517_,data_stage_4__1516_,data_stage_4__1515_,data_stage_4__1514_,
  data_stage_4__1513_,data_stage_4__1512_,data_stage_4__1511_,data_stage_4__1510_,
  data_stage_4__1509_,data_stage_4__1508_,data_stage_4__1507_,data_stage_4__1506_,
  data_stage_4__1505_,data_stage_4__1504_,data_stage_4__1503_,data_stage_4__1502_,
  data_stage_4__1501_,data_stage_4__1500_,data_stage_4__1499_,data_stage_4__1498_,
  data_stage_4__1497_,data_stage_4__1496_,data_stage_4__1495_,data_stage_4__1494_,
  data_stage_4__1493_,data_stage_4__1492_,data_stage_4__1491_,data_stage_4__1490_,
  data_stage_4__1489_,data_stage_4__1488_,data_stage_4__1487_,data_stage_4__1486_,
  data_stage_4__1485_,data_stage_4__1484_,data_stage_4__1483_,data_stage_4__1482_,
  data_stage_4__1481_,data_stage_4__1480_,data_stage_4__1479_,data_stage_4__1478_,
  data_stage_4__1477_,data_stage_4__1476_,data_stage_4__1475_,data_stage_4__1474_,
  data_stage_4__1473_,data_stage_4__1472_,data_stage_4__1471_,data_stage_4__1470_,
  data_stage_4__1469_,data_stage_4__1468_,data_stage_4__1467_,data_stage_4__1466_,
  data_stage_4__1465_,data_stage_4__1464_,data_stage_4__1463_,data_stage_4__1462_,
  data_stage_4__1461_,data_stage_4__1460_,data_stage_4__1459_,data_stage_4__1458_,
  data_stage_4__1457_,data_stage_4__1456_,data_stage_4__1455_,data_stage_4__1454_,
  data_stage_4__1453_,data_stage_4__1452_,data_stage_4__1451_,data_stage_4__1450_,
  data_stage_4__1449_,data_stage_4__1448_,data_stage_4__1447_,data_stage_4__1446_,
  data_stage_4__1445_,data_stage_4__1444_,data_stage_4__1443_,data_stage_4__1442_,
  data_stage_4__1441_,data_stage_4__1440_,data_stage_4__1439_,data_stage_4__1438_,
  data_stage_4__1437_,data_stage_4__1436_,data_stage_4__1435_,data_stage_4__1434_,
  data_stage_4__1433_,data_stage_4__1432_,data_stage_4__1431_,data_stage_4__1430_,
  data_stage_4__1429_,data_stage_4__1428_,data_stage_4__1427_,data_stage_4__1426_,
  data_stage_4__1425_,data_stage_4__1424_,data_stage_4__1423_,data_stage_4__1422_,
  data_stage_4__1421_,data_stage_4__1420_,data_stage_4__1419_,data_stage_4__1418_,
  data_stage_4__1417_,data_stage_4__1416_,data_stage_4__1415_,data_stage_4__1414_,
  data_stage_4__1413_,data_stage_4__1412_,data_stage_4__1411_,data_stage_4__1410_,
  data_stage_4__1409_,data_stage_4__1408_,data_stage_4__1407_,data_stage_4__1406_,
  data_stage_4__1405_,data_stage_4__1404_,data_stage_4__1403_,data_stage_4__1402_,
  data_stage_4__1401_,data_stage_4__1400_,data_stage_4__1399_,data_stage_4__1398_,
  data_stage_4__1397_,data_stage_4__1396_,data_stage_4__1395_,data_stage_4__1394_,
  data_stage_4__1393_,data_stage_4__1392_,data_stage_4__1391_,data_stage_4__1390_,
  data_stage_4__1389_,data_stage_4__1388_,data_stage_4__1387_,data_stage_4__1386_,
  data_stage_4__1385_,data_stage_4__1384_,data_stage_4__1383_,data_stage_4__1382_,
  data_stage_4__1381_,data_stage_4__1380_,data_stage_4__1379_,data_stage_4__1378_,
  data_stage_4__1377_,data_stage_4__1376_,data_stage_4__1375_,data_stage_4__1374_,
  data_stage_4__1373_,data_stage_4__1372_,data_stage_4__1371_,data_stage_4__1370_,
  data_stage_4__1369_,data_stage_4__1368_,data_stage_4__1367_,data_stage_4__1366_,
  data_stage_4__1365_,data_stage_4__1364_,data_stage_4__1363_,data_stage_4__1362_,
  data_stage_4__1361_,data_stage_4__1360_,data_stage_4__1359_,data_stage_4__1358_,
  data_stage_4__1357_,data_stage_4__1356_,data_stage_4__1355_,data_stage_4__1354_,
  data_stage_4__1353_,data_stage_4__1352_,data_stage_4__1351_,data_stage_4__1350_,
  data_stage_4__1349_,data_stage_4__1348_,data_stage_4__1347_,data_stage_4__1346_,
  data_stage_4__1345_,data_stage_4__1344_,data_stage_4__1343_,data_stage_4__1342_,
  data_stage_4__1341_,data_stage_4__1340_,data_stage_4__1339_,data_stage_4__1338_,
  data_stage_4__1337_,data_stage_4__1336_,data_stage_4__1335_,data_stage_4__1334_,
  data_stage_4__1333_,data_stage_4__1332_,data_stage_4__1331_,data_stage_4__1330_,
  data_stage_4__1329_,data_stage_4__1328_,data_stage_4__1327_,data_stage_4__1326_,
  data_stage_4__1325_,data_stage_4__1324_,data_stage_4__1323_,data_stage_4__1322_,
  data_stage_4__1321_,data_stage_4__1320_,data_stage_4__1319_,data_stage_4__1318_,
  data_stage_4__1317_,data_stage_4__1316_,data_stage_4__1315_,data_stage_4__1314_,
  data_stage_4__1313_,data_stage_4__1312_,data_stage_4__1311_,data_stage_4__1310_,
  data_stage_4__1309_,data_stage_4__1308_,data_stage_4__1307_,data_stage_4__1306_,
  data_stage_4__1305_,data_stage_4__1304_,data_stage_4__1303_,data_stage_4__1302_,
  data_stage_4__1301_,data_stage_4__1300_,data_stage_4__1299_,data_stage_4__1298_,
  data_stage_4__1297_,data_stage_4__1296_,data_stage_4__1295_,data_stage_4__1294_,
  data_stage_4__1293_,data_stage_4__1292_,data_stage_4__1291_,data_stage_4__1290_,
  data_stage_4__1289_,data_stage_4__1288_,data_stage_4__1287_,data_stage_4__1286_,
  data_stage_4__1285_,data_stage_4__1284_,data_stage_4__1283_,data_stage_4__1282_,
  data_stage_4__1281_,data_stage_4__1280_,data_stage_4__1279_,data_stage_4__1278_,
  data_stage_4__1277_,data_stage_4__1276_,data_stage_4__1275_,data_stage_4__1274_,
  data_stage_4__1273_,data_stage_4__1272_,data_stage_4__1271_,data_stage_4__1270_,
  data_stage_4__1269_,data_stage_4__1268_,data_stage_4__1267_,data_stage_4__1266_,
  data_stage_4__1265_,data_stage_4__1264_,data_stage_4__1263_,data_stage_4__1262_,
  data_stage_4__1261_,data_stage_4__1260_,data_stage_4__1259_,data_stage_4__1258_,
  data_stage_4__1257_,data_stage_4__1256_,data_stage_4__1255_,data_stage_4__1254_,
  data_stage_4__1253_,data_stage_4__1252_,data_stage_4__1251_,data_stage_4__1250_,
  data_stage_4__1249_,data_stage_4__1248_,data_stage_4__1247_,data_stage_4__1246_,
  data_stage_4__1245_,data_stage_4__1244_,data_stage_4__1243_,data_stage_4__1242_,
  data_stage_4__1241_,data_stage_4__1240_,data_stage_4__1239_,data_stage_4__1238_,
  data_stage_4__1237_,data_stage_4__1236_,data_stage_4__1235_,data_stage_4__1234_,
  data_stage_4__1233_,data_stage_4__1232_,data_stage_4__1231_,data_stage_4__1230_,
  data_stage_4__1229_,data_stage_4__1228_,data_stage_4__1227_,data_stage_4__1226_,
  data_stage_4__1225_,data_stage_4__1224_,data_stage_4__1223_,data_stage_4__1222_,
  data_stage_4__1221_,data_stage_4__1220_,data_stage_4__1219_,data_stage_4__1218_,
  data_stage_4__1217_,data_stage_4__1216_,data_stage_4__1215_,data_stage_4__1214_,
  data_stage_4__1213_,data_stage_4__1212_,data_stage_4__1211_,data_stage_4__1210_,
  data_stage_4__1209_,data_stage_4__1208_,data_stage_4__1207_,data_stage_4__1206_,
  data_stage_4__1205_,data_stage_4__1204_,data_stage_4__1203_,data_stage_4__1202_,
  data_stage_4__1201_,data_stage_4__1200_,data_stage_4__1199_,data_stage_4__1198_,
  data_stage_4__1197_,data_stage_4__1196_,data_stage_4__1195_,data_stage_4__1194_,
  data_stage_4__1193_,data_stage_4__1192_,data_stage_4__1191_,data_stage_4__1190_,
  data_stage_4__1189_,data_stage_4__1188_,data_stage_4__1187_,data_stage_4__1186_,
  data_stage_4__1185_,data_stage_4__1184_,data_stage_4__1183_,data_stage_4__1182_,
  data_stage_4__1181_,data_stage_4__1180_,data_stage_4__1179_,data_stage_4__1178_,
  data_stage_4__1177_,data_stage_4__1176_,data_stage_4__1175_,data_stage_4__1174_,
  data_stage_4__1173_,data_stage_4__1172_,data_stage_4__1171_,data_stage_4__1170_,
  data_stage_4__1169_,data_stage_4__1168_,data_stage_4__1167_,data_stage_4__1166_,
  data_stage_4__1165_,data_stage_4__1164_,data_stage_4__1163_,data_stage_4__1162_,
  data_stage_4__1161_,data_stage_4__1160_,data_stage_4__1159_,data_stage_4__1158_,
  data_stage_4__1157_,data_stage_4__1156_,data_stage_4__1155_,data_stage_4__1154_,
  data_stage_4__1153_,data_stage_4__1152_,data_stage_4__1151_,data_stage_4__1150_,
  data_stage_4__1149_,data_stage_4__1148_,data_stage_4__1147_,data_stage_4__1146_,
  data_stage_4__1145_,data_stage_4__1144_,data_stage_4__1143_,data_stage_4__1142_,
  data_stage_4__1141_,data_stage_4__1140_,data_stage_4__1139_,data_stage_4__1138_,
  data_stage_4__1137_,data_stage_4__1136_,data_stage_4__1135_,data_stage_4__1134_,
  data_stage_4__1133_,data_stage_4__1132_,data_stage_4__1131_,data_stage_4__1130_,
  data_stage_4__1129_,data_stage_4__1128_,data_stage_4__1127_,data_stage_4__1126_,
  data_stage_4__1125_,data_stage_4__1124_,data_stage_4__1123_,data_stage_4__1122_,
  data_stage_4__1121_,data_stage_4__1120_,data_stage_4__1119_,data_stage_4__1118_,
  data_stage_4__1117_,data_stage_4__1116_,data_stage_4__1115_,data_stage_4__1114_,
  data_stage_4__1113_,data_stage_4__1112_,data_stage_4__1111_,data_stage_4__1110_,
  data_stage_4__1109_,data_stage_4__1108_,data_stage_4__1107_,data_stage_4__1106_,
  data_stage_4__1105_,data_stage_4__1104_,data_stage_4__1103_,data_stage_4__1102_,
  data_stage_4__1101_,data_stage_4__1100_,data_stage_4__1099_,data_stage_4__1098_,
  data_stage_4__1097_,data_stage_4__1096_,data_stage_4__1095_,data_stage_4__1094_,
  data_stage_4__1093_,data_stage_4__1092_,data_stage_4__1091_,data_stage_4__1090_,
  data_stage_4__1089_,data_stage_4__1088_,data_stage_4__1087_,data_stage_4__1086_,
  data_stage_4__1085_,data_stage_4__1084_,data_stage_4__1083_,data_stage_4__1082_,
  data_stage_4__1081_,data_stage_4__1080_,data_stage_4__1079_,data_stage_4__1078_,
  data_stage_4__1077_,data_stage_4__1076_,data_stage_4__1075_,data_stage_4__1074_,
  data_stage_4__1073_,data_stage_4__1072_,data_stage_4__1071_,data_stage_4__1070_,
  data_stage_4__1069_,data_stage_4__1068_,data_stage_4__1067_,data_stage_4__1066_,
  data_stage_4__1065_,data_stage_4__1064_,data_stage_4__1063_,data_stage_4__1062_,
  data_stage_4__1061_,data_stage_4__1060_,data_stage_4__1059_,data_stage_4__1058_,
  data_stage_4__1057_,data_stage_4__1056_,data_stage_4__1055_,data_stage_4__1054_,
  data_stage_4__1053_,data_stage_4__1052_,data_stage_4__1051_,data_stage_4__1050_,
  data_stage_4__1049_,data_stage_4__1048_,data_stage_4__1047_,data_stage_4__1046_,
  data_stage_4__1045_,data_stage_4__1044_,data_stage_4__1043_,data_stage_4__1042_,
  data_stage_4__1041_,data_stage_4__1040_,data_stage_4__1039_,data_stage_4__1038_,
  data_stage_4__1037_,data_stage_4__1036_,data_stage_4__1035_,data_stage_4__1034_,
  data_stage_4__1033_,data_stage_4__1032_,data_stage_4__1031_,data_stage_4__1030_,
  data_stage_4__1029_,data_stage_4__1028_,data_stage_4__1027_,data_stage_4__1026_,
  data_stage_4__1025_,data_stage_4__1024_,data_stage_4__1023_,data_stage_4__1022_,
  data_stage_4__1021_,data_stage_4__1020_,data_stage_4__1019_,data_stage_4__1018_,
  data_stage_4__1017_,data_stage_4__1016_,data_stage_4__1015_,data_stage_4__1014_,
  data_stage_4__1013_,data_stage_4__1012_,data_stage_4__1011_,data_stage_4__1010_,
  data_stage_4__1009_,data_stage_4__1008_,data_stage_4__1007_,data_stage_4__1006_,
  data_stage_4__1005_,data_stage_4__1004_,data_stage_4__1003_,data_stage_4__1002_,
  data_stage_4__1001_,data_stage_4__1000_,data_stage_4__999_,data_stage_4__998_,
  data_stage_4__997_,data_stage_4__996_,data_stage_4__995_,data_stage_4__994_,
  data_stage_4__993_,data_stage_4__992_,data_stage_4__991_,data_stage_4__990_,data_stage_4__989_,
  data_stage_4__988_,data_stage_4__987_,data_stage_4__986_,data_stage_4__985_,
  data_stage_4__984_,data_stage_4__983_,data_stage_4__982_,data_stage_4__981_,
  data_stage_4__980_,data_stage_4__979_,data_stage_4__978_,data_stage_4__977_,
  data_stage_4__976_,data_stage_4__975_,data_stage_4__974_,data_stage_4__973_,
  data_stage_4__972_,data_stage_4__971_,data_stage_4__970_,data_stage_4__969_,data_stage_4__968_,
  data_stage_4__967_,data_stage_4__966_,data_stage_4__965_,data_stage_4__964_,
  data_stage_4__963_,data_stage_4__962_,data_stage_4__961_,data_stage_4__960_,
  data_stage_4__959_,data_stage_4__958_,data_stage_4__957_,data_stage_4__956_,
  data_stage_4__955_,data_stage_4__954_,data_stage_4__953_,data_stage_4__952_,
  data_stage_4__951_,data_stage_4__950_,data_stage_4__949_,data_stage_4__948_,data_stage_4__947_,
  data_stage_4__946_,data_stage_4__945_,data_stage_4__944_,data_stage_4__943_,
  data_stage_4__942_,data_stage_4__941_,data_stage_4__940_,data_stage_4__939_,
  data_stage_4__938_,data_stage_4__937_,data_stage_4__936_,data_stage_4__935_,
  data_stage_4__934_,data_stage_4__933_,data_stage_4__932_,data_stage_4__931_,data_stage_4__930_,
  data_stage_4__929_,data_stage_4__928_,data_stage_4__927_,data_stage_4__926_,
  data_stage_4__925_,data_stage_4__924_,data_stage_4__923_,data_stage_4__922_,
  data_stage_4__921_,data_stage_4__920_,data_stage_4__919_,data_stage_4__918_,
  data_stage_4__917_,data_stage_4__916_,data_stage_4__915_,data_stage_4__914_,
  data_stage_4__913_,data_stage_4__912_,data_stage_4__911_,data_stage_4__910_,data_stage_4__909_,
  data_stage_4__908_,data_stage_4__907_,data_stage_4__906_,data_stage_4__905_,
  data_stage_4__904_,data_stage_4__903_,data_stage_4__902_,data_stage_4__901_,
  data_stage_4__900_,data_stage_4__899_,data_stage_4__898_,data_stage_4__897_,
  data_stage_4__896_,data_stage_4__895_,data_stage_4__894_,data_stage_4__893_,
  data_stage_4__892_,data_stage_4__891_,data_stage_4__890_,data_stage_4__889_,data_stage_4__888_,
  data_stage_4__887_,data_stage_4__886_,data_stage_4__885_,data_stage_4__884_,
  data_stage_4__883_,data_stage_4__882_,data_stage_4__881_,data_stage_4__880_,
  data_stage_4__879_,data_stage_4__878_,data_stage_4__877_,data_stage_4__876_,
  data_stage_4__875_,data_stage_4__874_,data_stage_4__873_,data_stage_4__872_,
  data_stage_4__871_,data_stage_4__870_,data_stage_4__869_,data_stage_4__868_,data_stage_4__867_,
  data_stage_4__866_,data_stage_4__865_,data_stage_4__864_,data_stage_4__863_,
  data_stage_4__862_,data_stage_4__861_,data_stage_4__860_,data_stage_4__859_,
  data_stage_4__858_,data_stage_4__857_,data_stage_4__856_,data_stage_4__855_,
  data_stage_4__854_,data_stage_4__853_,data_stage_4__852_,data_stage_4__851_,data_stage_4__850_,
  data_stage_4__849_,data_stage_4__848_,data_stage_4__847_,data_stage_4__846_,
  data_stage_4__845_,data_stage_4__844_,data_stage_4__843_,data_stage_4__842_,
  data_stage_4__841_,data_stage_4__840_,data_stage_4__839_,data_stage_4__838_,
  data_stage_4__837_,data_stage_4__836_,data_stage_4__835_,data_stage_4__834_,
  data_stage_4__833_,data_stage_4__832_,data_stage_4__831_,data_stage_4__830_,data_stage_4__829_,
  data_stage_4__828_,data_stage_4__827_,data_stage_4__826_,data_stage_4__825_,
  data_stage_4__824_,data_stage_4__823_,data_stage_4__822_,data_stage_4__821_,
  data_stage_4__820_,data_stage_4__819_,data_stage_4__818_,data_stage_4__817_,
  data_stage_4__816_,data_stage_4__815_,data_stage_4__814_,data_stage_4__813_,
  data_stage_4__812_,data_stage_4__811_,data_stage_4__810_,data_stage_4__809_,data_stage_4__808_,
  data_stage_4__807_,data_stage_4__806_,data_stage_4__805_,data_stage_4__804_,
  data_stage_4__803_,data_stage_4__802_,data_stage_4__801_,data_stage_4__800_,
  data_stage_4__799_,data_stage_4__798_,data_stage_4__797_,data_stage_4__796_,
  data_stage_4__795_,data_stage_4__794_,data_stage_4__793_,data_stage_4__792_,
  data_stage_4__791_,data_stage_4__790_,data_stage_4__789_,data_stage_4__788_,data_stage_4__787_,
  data_stage_4__786_,data_stage_4__785_,data_stage_4__784_,data_stage_4__783_,
  data_stage_4__782_,data_stage_4__781_,data_stage_4__780_,data_stage_4__779_,
  data_stage_4__778_,data_stage_4__777_,data_stage_4__776_,data_stage_4__775_,
  data_stage_4__774_,data_stage_4__773_,data_stage_4__772_,data_stage_4__771_,data_stage_4__770_,
  data_stage_4__769_,data_stage_4__768_,data_stage_4__767_,data_stage_4__766_,
  data_stage_4__765_,data_stage_4__764_,data_stage_4__763_,data_stage_4__762_,
  data_stage_4__761_,data_stage_4__760_,data_stage_4__759_,data_stage_4__758_,
  data_stage_4__757_,data_stage_4__756_,data_stage_4__755_,data_stage_4__754_,
  data_stage_4__753_,data_stage_4__752_,data_stage_4__751_,data_stage_4__750_,data_stage_4__749_,
  data_stage_4__748_,data_stage_4__747_,data_stage_4__746_,data_stage_4__745_,
  data_stage_4__744_,data_stage_4__743_,data_stage_4__742_,data_stage_4__741_,
  data_stage_4__740_,data_stage_4__739_,data_stage_4__738_,data_stage_4__737_,
  data_stage_4__736_,data_stage_4__735_,data_stage_4__734_,data_stage_4__733_,
  data_stage_4__732_,data_stage_4__731_,data_stage_4__730_,data_stage_4__729_,data_stage_4__728_,
  data_stage_4__727_,data_stage_4__726_,data_stage_4__725_,data_stage_4__724_,
  data_stage_4__723_,data_stage_4__722_,data_stage_4__721_,data_stage_4__720_,
  data_stage_4__719_,data_stage_4__718_,data_stage_4__717_,data_stage_4__716_,
  data_stage_4__715_,data_stage_4__714_,data_stage_4__713_,data_stage_4__712_,
  data_stage_4__711_,data_stage_4__710_,data_stage_4__709_,data_stage_4__708_,data_stage_4__707_,
  data_stage_4__706_,data_stage_4__705_,data_stage_4__704_,data_stage_4__703_,
  data_stage_4__702_,data_stage_4__701_,data_stage_4__700_,data_stage_4__699_,
  data_stage_4__698_,data_stage_4__697_,data_stage_4__696_,data_stage_4__695_,
  data_stage_4__694_,data_stage_4__693_,data_stage_4__692_,data_stage_4__691_,data_stage_4__690_,
  data_stage_4__689_,data_stage_4__688_,data_stage_4__687_,data_stage_4__686_,
  data_stage_4__685_,data_stage_4__684_,data_stage_4__683_,data_stage_4__682_,
  data_stage_4__681_,data_stage_4__680_,data_stage_4__679_,data_stage_4__678_,
  data_stage_4__677_,data_stage_4__676_,data_stage_4__675_,data_stage_4__674_,
  data_stage_4__673_,data_stage_4__672_,data_stage_4__671_,data_stage_4__670_,data_stage_4__669_,
  data_stage_4__668_,data_stage_4__667_,data_stage_4__666_,data_stage_4__665_,
  data_stage_4__664_,data_stage_4__663_,data_stage_4__662_,data_stage_4__661_,
  data_stage_4__660_,data_stage_4__659_,data_stage_4__658_,data_stage_4__657_,
  data_stage_4__656_,data_stage_4__655_,data_stage_4__654_,data_stage_4__653_,
  data_stage_4__652_,data_stage_4__651_,data_stage_4__650_,data_stage_4__649_,data_stage_4__648_,
  data_stage_4__647_,data_stage_4__646_,data_stage_4__645_,data_stage_4__644_,
  data_stage_4__643_,data_stage_4__642_,data_stage_4__641_,data_stage_4__640_,
  data_stage_4__639_,data_stage_4__638_,data_stage_4__637_,data_stage_4__636_,
  data_stage_4__635_,data_stage_4__634_,data_stage_4__633_,data_stage_4__632_,
  data_stage_4__631_,data_stage_4__630_,data_stage_4__629_,data_stage_4__628_,data_stage_4__627_,
  data_stage_4__626_,data_stage_4__625_,data_stage_4__624_,data_stage_4__623_,
  data_stage_4__622_,data_stage_4__621_,data_stage_4__620_,data_stage_4__619_,
  data_stage_4__618_,data_stage_4__617_,data_stage_4__616_,data_stage_4__615_,
  data_stage_4__614_,data_stage_4__613_,data_stage_4__612_,data_stage_4__611_,data_stage_4__610_,
  data_stage_4__609_,data_stage_4__608_,data_stage_4__607_,data_stage_4__606_,
  data_stage_4__605_,data_stage_4__604_,data_stage_4__603_,data_stage_4__602_,
  data_stage_4__601_,data_stage_4__600_,data_stage_4__599_,data_stage_4__598_,
  data_stage_4__597_,data_stage_4__596_,data_stage_4__595_,data_stage_4__594_,
  data_stage_4__593_,data_stage_4__592_,data_stage_4__591_,data_stage_4__590_,data_stage_4__589_,
  data_stage_4__588_,data_stage_4__587_,data_stage_4__586_,data_stage_4__585_,
  data_stage_4__584_,data_stage_4__583_,data_stage_4__582_,data_stage_4__581_,
  data_stage_4__580_,data_stage_4__579_,data_stage_4__578_,data_stage_4__577_,
  data_stage_4__576_,data_stage_4__575_,data_stage_4__574_,data_stage_4__573_,
  data_stage_4__572_,data_stage_4__571_,data_stage_4__570_,data_stage_4__569_,data_stage_4__568_,
  data_stage_4__567_,data_stage_4__566_,data_stage_4__565_,data_stage_4__564_,
  data_stage_4__563_,data_stage_4__562_,data_stage_4__561_,data_stage_4__560_,
  data_stage_4__559_,data_stage_4__558_,data_stage_4__557_,data_stage_4__556_,
  data_stage_4__555_,data_stage_4__554_,data_stage_4__553_,data_stage_4__552_,
  data_stage_4__551_,data_stage_4__550_,data_stage_4__549_,data_stage_4__548_,data_stage_4__547_,
  data_stage_4__546_,data_stage_4__545_,data_stage_4__544_,data_stage_4__543_,
  data_stage_4__542_,data_stage_4__541_,data_stage_4__540_,data_stage_4__539_,
  data_stage_4__538_,data_stage_4__537_,data_stage_4__536_,data_stage_4__535_,
  data_stage_4__534_,data_stage_4__533_,data_stage_4__532_,data_stage_4__531_,data_stage_4__530_,
  data_stage_4__529_,data_stage_4__528_,data_stage_4__527_,data_stage_4__526_,
  data_stage_4__525_,data_stage_4__524_,data_stage_4__523_,data_stage_4__522_,
  data_stage_4__521_,data_stage_4__520_,data_stage_4__519_,data_stage_4__518_,
  data_stage_4__517_,data_stage_4__516_,data_stage_4__515_,data_stage_4__514_,
  data_stage_4__513_,data_stage_4__512_,data_stage_4__511_,data_stage_4__510_,data_stage_4__509_,
  data_stage_4__508_,data_stage_4__507_,data_stage_4__506_,data_stage_4__505_,
  data_stage_4__504_,data_stage_4__503_,data_stage_4__502_,data_stage_4__501_,
  data_stage_4__500_,data_stage_4__499_,data_stage_4__498_,data_stage_4__497_,
  data_stage_4__496_,data_stage_4__495_,data_stage_4__494_,data_stage_4__493_,
  data_stage_4__492_,data_stage_4__491_,data_stage_4__490_,data_stage_4__489_,data_stage_4__488_,
  data_stage_4__487_,data_stage_4__486_,data_stage_4__485_,data_stage_4__484_,
  data_stage_4__483_,data_stage_4__482_,data_stage_4__481_,data_stage_4__480_,
  data_stage_4__479_,data_stage_4__478_,data_stage_4__477_,data_stage_4__476_,
  data_stage_4__475_,data_stage_4__474_,data_stage_4__473_,data_stage_4__472_,
  data_stage_4__471_,data_stage_4__470_,data_stage_4__469_,data_stage_4__468_,data_stage_4__467_,
  data_stage_4__466_,data_stage_4__465_,data_stage_4__464_,data_stage_4__463_,
  data_stage_4__462_,data_stage_4__461_,data_stage_4__460_,data_stage_4__459_,
  data_stage_4__458_,data_stage_4__457_,data_stage_4__456_,data_stage_4__455_,
  data_stage_4__454_,data_stage_4__453_,data_stage_4__452_,data_stage_4__451_,data_stage_4__450_,
  data_stage_4__449_,data_stage_4__448_,data_stage_4__447_,data_stage_4__446_,
  data_stage_4__445_,data_stage_4__444_,data_stage_4__443_,data_stage_4__442_,
  data_stage_4__441_,data_stage_4__440_,data_stage_4__439_,data_stage_4__438_,
  data_stage_4__437_,data_stage_4__436_,data_stage_4__435_,data_stage_4__434_,
  data_stage_4__433_,data_stage_4__432_,data_stage_4__431_,data_stage_4__430_,data_stage_4__429_,
  data_stage_4__428_,data_stage_4__427_,data_stage_4__426_,data_stage_4__425_,
  data_stage_4__424_,data_stage_4__423_,data_stage_4__422_,data_stage_4__421_,
  data_stage_4__420_,data_stage_4__419_,data_stage_4__418_,data_stage_4__417_,
  data_stage_4__416_,data_stage_4__415_,data_stage_4__414_,data_stage_4__413_,
  data_stage_4__412_,data_stage_4__411_,data_stage_4__410_,data_stage_4__409_,data_stage_4__408_,
  data_stage_4__407_,data_stage_4__406_,data_stage_4__405_,data_stage_4__404_,
  data_stage_4__403_,data_stage_4__402_,data_stage_4__401_,data_stage_4__400_,
  data_stage_4__399_,data_stage_4__398_,data_stage_4__397_,data_stage_4__396_,
  data_stage_4__395_,data_stage_4__394_,data_stage_4__393_,data_stage_4__392_,
  data_stage_4__391_,data_stage_4__390_,data_stage_4__389_,data_stage_4__388_,data_stage_4__387_,
  data_stage_4__386_,data_stage_4__385_,data_stage_4__384_,data_stage_4__383_,
  data_stage_4__382_,data_stage_4__381_,data_stage_4__380_,data_stage_4__379_,
  data_stage_4__378_,data_stage_4__377_,data_stage_4__376_,data_stage_4__375_,
  data_stage_4__374_,data_stage_4__373_,data_stage_4__372_,data_stage_4__371_,data_stage_4__370_,
  data_stage_4__369_,data_stage_4__368_,data_stage_4__367_,data_stage_4__366_,
  data_stage_4__365_,data_stage_4__364_,data_stage_4__363_,data_stage_4__362_,
  data_stage_4__361_,data_stage_4__360_,data_stage_4__359_,data_stage_4__358_,
  data_stage_4__357_,data_stage_4__356_,data_stage_4__355_,data_stage_4__354_,
  data_stage_4__353_,data_stage_4__352_,data_stage_4__351_,data_stage_4__350_,data_stage_4__349_,
  data_stage_4__348_,data_stage_4__347_,data_stage_4__346_,data_stage_4__345_,
  data_stage_4__344_,data_stage_4__343_,data_stage_4__342_,data_stage_4__341_,
  data_stage_4__340_,data_stage_4__339_,data_stage_4__338_,data_stage_4__337_,
  data_stage_4__336_,data_stage_4__335_,data_stage_4__334_,data_stage_4__333_,
  data_stage_4__332_,data_stage_4__331_,data_stage_4__330_,data_stage_4__329_,data_stage_4__328_,
  data_stage_4__327_,data_stage_4__326_,data_stage_4__325_,data_stage_4__324_,
  data_stage_4__323_,data_stage_4__322_,data_stage_4__321_,data_stage_4__320_,
  data_stage_4__319_,data_stage_4__318_,data_stage_4__317_,data_stage_4__316_,
  data_stage_4__315_,data_stage_4__314_,data_stage_4__313_,data_stage_4__312_,
  data_stage_4__311_,data_stage_4__310_,data_stage_4__309_,data_stage_4__308_,data_stage_4__307_,
  data_stage_4__306_,data_stage_4__305_,data_stage_4__304_,data_stage_4__303_,
  data_stage_4__302_,data_stage_4__301_,data_stage_4__300_,data_stage_4__299_,
  data_stage_4__298_,data_stage_4__297_,data_stage_4__296_,data_stage_4__295_,
  data_stage_4__294_,data_stage_4__293_,data_stage_4__292_,data_stage_4__291_,data_stage_4__290_,
  data_stage_4__289_,data_stage_4__288_,data_stage_4__287_,data_stage_4__286_,
  data_stage_4__285_,data_stage_4__284_,data_stage_4__283_,data_stage_4__282_,
  data_stage_4__281_,data_stage_4__280_,data_stage_4__279_,data_stage_4__278_,
  data_stage_4__277_,data_stage_4__276_,data_stage_4__275_,data_stage_4__274_,
  data_stage_4__273_,data_stage_4__272_,data_stage_4__271_,data_stage_4__270_,data_stage_4__269_,
  data_stage_4__268_,data_stage_4__267_,data_stage_4__266_,data_stage_4__265_,
  data_stage_4__264_,data_stage_4__263_,data_stage_4__262_,data_stage_4__261_,
  data_stage_4__260_,data_stage_4__259_,data_stage_4__258_,data_stage_4__257_,
  data_stage_4__256_,data_stage_4__255_,data_stage_4__254_,data_stage_4__253_,
  data_stage_4__252_,data_stage_4__251_,data_stage_4__250_,data_stage_4__249_,data_stage_4__248_,
  data_stage_4__247_,data_stage_4__246_,data_stage_4__245_,data_stage_4__244_,
  data_stage_4__243_,data_stage_4__242_,data_stage_4__241_,data_stage_4__240_,
  data_stage_4__239_,data_stage_4__238_,data_stage_4__237_,data_stage_4__236_,
  data_stage_4__235_,data_stage_4__234_,data_stage_4__233_,data_stage_4__232_,
  data_stage_4__231_,data_stage_4__230_,data_stage_4__229_,data_stage_4__228_,data_stage_4__227_,
  data_stage_4__226_,data_stage_4__225_,data_stage_4__224_,data_stage_4__223_,
  data_stage_4__222_,data_stage_4__221_,data_stage_4__220_,data_stage_4__219_,
  data_stage_4__218_,data_stage_4__217_,data_stage_4__216_,data_stage_4__215_,
  data_stage_4__214_,data_stage_4__213_,data_stage_4__212_,data_stage_4__211_,data_stage_4__210_,
  data_stage_4__209_,data_stage_4__208_,data_stage_4__207_,data_stage_4__206_,
  data_stage_4__205_,data_stage_4__204_,data_stage_4__203_,data_stage_4__202_,
  data_stage_4__201_,data_stage_4__200_,data_stage_4__199_,data_stage_4__198_,
  data_stage_4__197_,data_stage_4__196_,data_stage_4__195_,data_stage_4__194_,
  data_stage_4__193_,data_stage_4__192_,data_stage_4__191_,data_stage_4__190_,data_stage_4__189_,
  data_stage_4__188_,data_stage_4__187_,data_stage_4__186_,data_stage_4__185_,
  data_stage_4__184_,data_stage_4__183_,data_stage_4__182_,data_stage_4__181_,
  data_stage_4__180_,data_stage_4__179_,data_stage_4__178_,data_stage_4__177_,
  data_stage_4__176_,data_stage_4__175_,data_stage_4__174_,data_stage_4__173_,
  data_stage_4__172_,data_stage_4__171_,data_stage_4__170_,data_stage_4__169_,data_stage_4__168_,
  data_stage_4__167_,data_stage_4__166_,data_stage_4__165_,data_stage_4__164_,
  data_stage_4__163_,data_stage_4__162_,data_stage_4__161_,data_stage_4__160_,
  data_stage_4__159_,data_stage_4__158_,data_stage_4__157_,data_stage_4__156_,
  data_stage_4__155_,data_stage_4__154_,data_stage_4__153_,data_stage_4__152_,
  data_stage_4__151_,data_stage_4__150_,data_stage_4__149_,data_stage_4__148_,data_stage_4__147_,
  data_stage_4__146_,data_stage_4__145_,data_stage_4__144_,data_stage_4__143_,
  data_stage_4__142_,data_stage_4__141_,data_stage_4__140_,data_stage_4__139_,
  data_stage_4__138_,data_stage_4__137_,data_stage_4__136_,data_stage_4__135_,
  data_stage_4__134_,data_stage_4__133_,data_stage_4__132_,data_stage_4__131_,data_stage_4__130_,
  data_stage_4__129_,data_stage_4__128_,data_stage_4__127_,data_stage_4__126_,
  data_stage_4__125_,data_stage_4__124_,data_stage_4__123_,data_stage_4__122_,
  data_stage_4__121_,data_stage_4__120_,data_stage_4__119_,data_stage_4__118_,
  data_stage_4__117_,data_stage_4__116_,data_stage_4__115_,data_stage_4__114_,
  data_stage_4__113_,data_stage_4__112_,data_stage_4__111_,data_stage_4__110_,data_stage_4__109_,
  data_stage_4__108_,data_stage_4__107_,data_stage_4__106_,data_stage_4__105_,
  data_stage_4__104_,data_stage_4__103_,data_stage_4__102_,data_stage_4__101_,
  data_stage_4__100_,data_stage_4__99_,data_stage_4__98_,data_stage_4__97_,
  data_stage_4__96_,data_stage_4__95_,data_stage_4__94_,data_stage_4__93_,data_stage_4__92_,
  data_stage_4__91_,data_stage_4__90_,data_stage_4__89_,data_stage_4__88_,
  data_stage_4__87_,data_stage_4__86_,data_stage_4__85_,data_stage_4__84_,data_stage_4__83_,
  data_stage_4__82_,data_stage_4__81_,data_stage_4__80_,data_stage_4__79_,
  data_stage_4__78_,data_stage_4__77_,data_stage_4__76_,data_stage_4__75_,data_stage_4__74_,
  data_stage_4__73_,data_stage_4__72_,data_stage_4__71_,data_stage_4__70_,
  data_stage_4__69_,data_stage_4__68_,data_stage_4__67_,data_stage_4__66_,data_stage_4__65_,
  data_stage_4__64_,data_stage_4__63_,data_stage_4__62_,data_stage_4__61_,
  data_stage_4__60_,data_stage_4__59_,data_stage_4__58_,data_stage_4__57_,
  data_stage_4__56_,data_stage_4__55_,data_stage_4__54_,data_stage_4__53_,data_stage_4__52_,
  data_stage_4__51_,data_stage_4__50_,data_stage_4__49_,data_stage_4__48_,
  data_stage_4__47_,data_stage_4__46_,data_stage_4__45_,data_stage_4__44_,data_stage_4__43_,
  data_stage_4__42_,data_stage_4__41_,data_stage_4__40_,data_stage_4__39_,
  data_stage_4__38_,data_stage_4__37_,data_stage_4__36_,data_stage_4__35_,data_stage_4__34_,
  data_stage_4__33_,data_stage_4__32_,data_stage_4__31_,data_stage_4__30_,
  data_stage_4__29_,data_stage_4__28_,data_stage_4__27_,data_stage_4__26_,data_stage_4__25_,
  data_stage_4__24_,data_stage_4__23_,data_stage_4__22_,data_stage_4__21_,
  data_stage_4__20_,data_stage_4__19_,data_stage_4__18_,data_stage_4__17_,
  data_stage_4__16_,data_stage_4__15_,data_stage_4__14_,data_stage_4__13_,data_stage_4__12_,
  data_stage_4__11_,data_stage_4__10_,data_stage_4__9_,data_stage_4__8_,
  data_stage_4__7_,data_stage_4__6_,data_stage_4__5_,data_stage_4__4_,data_stage_4__3_,
  data_stage_4__2_,data_stage_4__1_,data_stage_4__0_,data_stage_5__4095_,data_stage_5__4094_,
  data_stage_5__4093_,data_stage_5__4092_,data_stage_5__4091_,data_stage_5__4090_,
  data_stage_5__4089_,data_stage_5__4088_,data_stage_5__4087_,data_stage_5__4086_,
  data_stage_5__4085_,data_stage_5__4084_,data_stage_5__4083_,data_stage_5__4082_,
  data_stage_5__4081_,data_stage_5__4080_,data_stage_5__4079_,data_stage_5__4078_,
  data_stage_5__4077_,data_stage_5__4076_,data_stage_5__4075_,data_stage_5__4074_,
  data_stage_5__4073_,data_stage_5__4072_,data_stage_5__4071_,data_stage_5__4070_,
  data_stage_5__4069_,data_stage_5__4068_,data_stage_5__4067_,data_stage_5__4066_,
  data_stage_5__4065_,data_stage_5__4064_,data_stage_5__4063_,data_stage_5__4062_,
  data_stage_5__4061_,data_stage_5__4060_,data_stage_5__4059_,data_stage_5__4058_,
  data_stage_5__4057_,data_stage_5__4056_,data_stage_5__4055_,data_stage_5__4054_,
  data_stage_5__4053_,data_stage_5__4052_,data_stage_5__4051_,data_stage_5__4050_,
  data_stage_5__4049_,data_stage_5__4048_,data_stage_5__4047_,data_stage_5__4046_,
  data_stage_5__4045_,data_stage_5__4044_,data_stage_5__4043_,data_stage_5__4042_,
  data_stage_5__4041_,data_stage_5__4040_,data_stage_5__4039_,data_stage_5__4038_,
  data_stage_5__4037_,data_stage_5__4036_,data_stage_5__4035_,data_stage_5__4034_,
  data_stage_5__4033_,data_stage_5__4032_,data_stage_5__4031_,data_stage_5__4030_,
  data_stage_5__4029_,data_stage_5__4028_,data_stage_5__4027_,data_stage_5__4026_,
  data_stage_5__4025_,data_stage_5__4024_,data_stage_5__4023_,data_stage_5__4022_,
  data_stage_5__4021_,data_stage_5__4020_,data_stage_5__4019_,data_stage_5__4018_,
  data_stage_5__4017_,data_stage_5__4016_,data_stage_5__4015_,data_stage_5__4014_,
  data_stage_5__4013_,data_stage_5__4012_,data_stage_5__4011_,data_stage_5__4010_,
  data_stage_5__4009_,data_stage_5__4008_,data_stage_5__4007_,data_stage_5__4006_,
  data_stage_5__4005_,data_stage_5__4004_,data_stage_5__4003_,data_stage_5__4002_,
  data_stage_5__4001_,data_stage_5__4000_,data_stage_5__3999_,data_stage_5__3998_,
  data_stage_5__3997_,data_stage_5__3996_,data_stage_5__3995_,data_stage_5__3994_,
  data_stage_5__3993_,data_stage_5__3992_,data_stage_5__3991_,data_stage_5__3990_,
  data_stage_5__3989_,data_stage_5__3988_,data_stage_5__3987_,data_stage_5__3986_,
  data_stage_5__3985_,data_stage_5__3984_,data_stage_5__3983_,data_stage_5__3982_,
  data_stage_5__3981_,data_stage_5__3980_,data_stage_5__3979_,data_stage_5__3978_,
  data_stage_5__3977_,data_stage_5__3976_,data_stage_5__3975_,data_stage_5__3974_,
  data_stage_5__3973_,data_stage_5__3972_,data_stage_5__3971_,data_stage_5__3970_,
  data_stage_5__3969_,data_stage_5__3968_,data_stage_5__3967_,data_stage_5__3966_,
  data_stage_5__3965_,data_stage_5__3964_,data_stage_5__3963_,data_stage_5__3962_,
  data_stage_5__3961_,data_stage_5__3960_,data_stage_5__3959_,data_stage_5__3958_,
  data_stage_5__3957_,data_stage_5__3956_,data_stage_5__3955_,data_stage_5__3954_,
  data_stage_5__3953_,data_stage_5__3952_,data_stage_5__3951_,data_stage_5__3950_,
  data_stage_5__3949_,data_stage_5__3948_,data_stage_5__3947_,data_stage_5__3946_,
  data_stage_5__3945_,data_stage_5__3944_,data_stage_5__3943_,data_stage_5__3942_,
  data_stage_5__3941_,data_stage_5__3940_,data_stage_5__3939_,data_stage_5__3938_,
  data_stage_5__3937_,data_stage_5__3936_,data_stage_5__3935_,data_stage_5__3934_,
  data_stage_5__3933_,data_stage_5__3932_,data_stage_5__3931_,data_stage_5__3930_,
  data_stage_5__3929_,data_stage_5__3928_,data_stage_5__3927_,data_stage_5__3926_,
  data_stage_5__3925_,data_stage_5__3924_,data_stage_5__3923_,data_stage_5__3922_,
  data_stage_5__3921_,data_stage_5__3920_,data_stage_5__3919_,data_stage_5__3918_,
  data_stage_5__3917_,data_stage_5__3916_,data_stage_5__3915_,data_stage_5__3914_,
  data_stage_5__3913_,data_stage_5__3912_,data_stage_5__3911_,data_stage_5__3910_,
  data_stage_5__3909_,data_stage_5__3908_,data_stage_5__3907_,data_stage_5__3906_,
  data_stage_5__3905_,data_stage_5__3904_,data_stage_5__3903_,data_stage_5__3902_,
  data_stage_5__3901_,data_stage_5__3900_,data_stage_5__3899_,data_stage_5__3898_,
  data_stage_5__3897_,data_stage_5__3896_,data_stage_5__3895_,data_stage_5__3894_,
  data_stage_5__3893_,data_stage_5__3892_,data_stage_5__3891_,data_stage_5__3890_,
  data_stage_5__3889_,data_stage_5__3888_,data_stage_5__3887_,data_stage_5__3886_,
  data_stage_5__3885_,data_stage_5__3884_,data_stage_5__3883_,data_stage_5__3882_,
  data_stage_5__3881_,data_stage_5__3880_,data_stage_5__3879_,data_stage_5__3878_,
  data_stage_5__3877_,data_stage_5__3876_,data_stage_5__3875_,data_stage_5__3874_,
  data_stage_5__3873_,data_stage_5__3872_,data_stage_5__3871_,data_stage_5__3870_,
  data_stage_5__3869_,data_stage_5__3868_,data_stage_5__3867_,data_stage_5__3866_,
  data_stage_5__3865_,data_stage_5__3864_,data_stage_5__3863_,data_stage_5__3862_,
  data_stage_5__3861_,data_stage_5__3860_,data_stage_5__3859_,data_stage_5__3858_,
  data_stage_5__3857_,data_stage_5__3856_,data_stage_5__3855_,data_stage_5__3854_,
  data_stage_5__3853_,data_stage_5__3852_,data_stage_5__3851_,data_stage_5__3850_,
  data_stage_5__3849_,data_stage_5__3848_,data_stage_5__3847_,data_stage_5__3846_,
  data_stage_5__3845_,data_stage_5__3844_,data_stage_5__3843_,data_stage_5__3842_,
  data_stage_5__3841_,data_stage_5__3840_,data_stage_5__3839_,data_stage_5__3838_,
  data_stage_5__3837_,data_stage_5__3836_,data_stage_5__3835_,data_stage_5__3834_,
  data_stage_5__3833_,data_stage_5__3832_,data_stage_5__3831_,data_stage_5__3830_,
  data_stage_5__3829_,data_stage_5__3828_,data_stage_5__3827_,data_stage_5__3826_,
  data_stage_5__3825_,data_stage_5__3824_,data_stage_5__3823_,data_stage_5__3822_,
  data_stage_5__3821_,data_stage_5__3820_,data_stage_5__3819_,data_stage_5__3818_,
  data_stage_5__3817_,data_stage_5__3816_,data_stage_5__3815_,data_stage_5__3814_,
  data_stage_5__3813_,data_stage_5__3812_,data_stage_5__3811_,data_stage_5__3810_,
  data_stage_5__3809_,data_stage_5__3808_,data_stage_5__3807_,data_stage_5__3806_,
  data_stage_5__3805_,data_stage_5__3804_,data_stage_5__3803_,data_stage_5__3802_,
  data_stage_5__3801_,data_stage_5__3800_,data_stage_5__3799_,data_stage_5__3798_,
  data_stage_5__3797_,data_stage_5__3796_,data_stage_5__3795_,data_stage_5__3794_,
  data_stage_5__3793_,data_stage_5__3792_,data_stage_5__3791_,data_stage_5__3790_,
  data_stage_5__3789_,data_stage_5__3788_,data_stage_5__3787_,data_stage_5__3786_,
  data_stage_5__3785_,data_stage_5__3784_,data_stage_5__3783_,data_stage_5__3782_,
  data_stage_5__3781_,data_stage_5__3780_,data_stage_5__3779_,data_stage_5__3778_,
  data_stage_5__3777_,data_stage_5__3776_,data_stage_5__3775_,data_stage_5__3774_,
  data_stage_5__3773_,data_stage_5__3772_,data_stage_5__3771_,data_stage_5__3770_,
  data_stage_5__3769_,data_stage_5__3768_,data_stage_5__3767_,data_stage_5__3766_,
  data_stage_5__3765_,data_stage_5__3764_,data_stage_5__3763_,data_stage_5__3762_,
  data_stage_5__3761_,data_stage_5__3760_,data_stage_5__3759_,data_stage_5__3758_,
  data_stage_5__3757_,data_stage_5__3756_,data_stage_5__3755_,data_stage_5__3754_,
  data_stage_5__3753_,data_stage_5__3752_,data_stage_5__3751_,data_stage_5__3750_,
  data_stage_5__3749_,data_stage_5__3748_,data_stage_5__3747_,data_stage_5__3746_,
  data_stage_5__3745_,data_stage_5__3744_,data_stage_5__3743_,data_stage_5__3742_,
  data_stage_5__3741_,data_stage_5__3740_,data_stage_5__3739_,data_stage_5__3738_,
  data_stage_5__3737_,data_stage_5__3736_,data_stage_5__3735_,data_stage_5__3734_,
  data_stage_5__3733_,data_stage_5__3732_,data_stage_5__3731_,data_stage_5__3730_,
  data_stage_5__3729_,data_stage_5__3728_,data_stage_5__3727_,data_stage_5__3726_,
  data_stage_5__3725_,data_stage_5__3724_,data_stage_5__3723_,data_stage_5__3722_,
  data_stage_5__3721_,data_stage_5__3720_,data_stage_5__3719_,data_stage_5__3718_,
  data_stage_5__3717_,data_stage_5__3716_,data_stage_5__3715_,data_stage_5__3714_,
  data_stage_5__3713_,data_stage_5__3712_,data_stage_5__3711_,data_stage_5__3710_,
  data_stage_5__3709_,data_stage_5__3708_,data_stage_5__3707_,data_stage_5__3706_,
  data_stage_5__3705_,data_stage_5__3704_,data_stage_5__3703_,data_stage_5__3702_,
  data_stage_5__3701_,data_stage_5__3700_,data_stage_5__3699_,data_stage_5__3698_,
  data_stage_5__3697_,data_stage_5__3696_,data_stage_5__3695_,data_stage_5__3694_,
  data_stage_5__3693_,data_stage_5__3692_,data_stage_5__3691_,data_stage_5__3690_,
  data_stage_5__3689_,data_stage_5__3688_,data_stage_5__3687_,data_stage_5__3686_,
  data_stage_5__3685_,data_stage_5__3684_,data_stage_5__3683_,data_stage_5__3682_,
  data_stage_5__3681_,data_stage_5__3680_,data_stage_5__3679_,data_stage_5__3678_,
  data_stage_5__3677_,data_stage_5__3676_,data_stage_5__3675_,data_stage_5__3674_,
  data_stage_5__3673_,data_stage_5__3672_,data_stage_5__3671_,data_stage_5__3670_,
  data_stage_5__3669_,data_stage_5__3668_,data_stage_5__3667_,data_stage_5__3666_,
  data_stage_5__3665_,data_stage_5__3664_,data_stage_5__3663_,data_stage_5__3662_,
  data_stage_5__3661_,data_stage_5__3660_,data_stage_5__3659_,data_stage_5__3658_,
  data_stage_5__3657_,data_stage_5__3656_,data_stage_5__3655_,data_stage_5__3654_,
  data_stage_5__3653_,data_stage_5__3652_,data_stage_5__3651_,data_stage_5__3650_,
  data_stage_5__3649_,data_stage_5__3648_,data_stage_5__3647_,data_stage_5__3646_,
  data_stage_5__3645_,data_stage_5__3644_,data_stage_5__3643_,data_stage_5__3642_,
  data_stage_5__3641_,data_stage_5__3640_,data_stage_5__3639_,data_stage_5__3638_,
  data_stage_5__3637_,data_stage_5__3636_,data_stage_5__3635_,data_stage_5__3634_,
  data_stage_5__3633_,data_stage_5__3632_,data_stage_5__3631_,data_stage_5__3630_,
  data_stage_5__3629_,data_stage_5__3628_,data_stage_5__3627_,data_stage_5__3626_,
  data_stage_5__3625_,data_stage_5__3624_,data_stage_5__3623_,data_stage_5__3622_,
  data_stage_5__3621_,data_stage_5__3620_,data_stage_5__3619_,data_stage_5__3618_,
  data_stage_5__3617_,data_stage_5__3616_,data_stage_5__3615_,data_stage_5__3614_,
  data_stage_5__3613_,data_stage_5__3612_,data_stage_5__3611_,data_stage_5__3610_,
  data_stage_5__3609_,data_stage_5__3608_,data_stage_5__3607_,data_stage_5__3606_,
  data_stage_5__3605_,data_stage_5__3604_,data_stage_5__3603_,data_stage_5__3602_,
  data_stage_5__3601_,data_stage_5__3600_,data_stage_5__3599_,data_stage_5__3598_,
  data_stage_5__3597_,data_stage_5__3596_,data_stage_5__3595_,data_stage_5__3594_,
  data_stage_5__3593_,data_stage_5__3592_,data_stage_5__3591_,data_stage_5__3590_,
  data_stage_5__3589_,data_stage_5__3588_,data_stage_5__3587_,data_stage_5__3586_,
  data_stage_5__3585_,data_stage_5__3584_,data_stage_5__3583_,data_stage_5__3582_,
  data_stage_5__3581_,data_stage_5__3580_,data_stage_5__3579_,data_stage_5__3578_,
  data_stage_5__3577_,data_stage_5__3576_,data_stage_5__3575_,data_stage_5__3574_,
  data_stage_5__3573_,data_stage_5__3572_,data_stage_5__3571_,data_stage_5__3570_,
  data_stage_5__3569_,data_stage_5__3568_,data_stage_5__3567_,data_stage_5__3566_,
  data_stage_5__3565_,data_stage_5__3564_,data_stage_5__3563_,data_stage_5__3562_,
  data_stage_5__3561_,data_stage_5__3560_,data_stage_5__3559_,data_stage_5__3558_,
  data_stage_5__3557_,data_stage_5__3556_,data_stage_5__3555_,data_stage_5__3554_,
  data_stage_5__3553_,data_stage_5__3552_,data_stage_5__3551_,data_stage_5__3550_,
  data_stage_5__3549_,data_stage_5__3548_,data_stage_5__3547_,data_stage_5__3546_,
  data_stage_5__3545_,data_stage_5__3544_,data_stage_5__3543_,data_stage_5__3542_,
  data_stage_5__3541_,data_stage_5__3540_,data_stage_5__3539_,data_stage_5__3538_,
  data_stage_5__3537_,data_stage_5__3536_,data_stage_5__3535_,data_stage_5__3534_,
  data_stage_5__3533_,data_stage_5__3532_,data_stage_5__3531_,data_stage_5__3530_,
  data_stage_5__3529_,data_stage_5__3528_,data_stage_5__3527_,data_stage_5__3526_,
  data_stage_5__3525_,data_stage_5__3524_,data_stage_5__3523_,data_stage_5__3522_,
  data_stage_5__3521_,data_stage_5__3520_,data_stage_5__3519_,data_stage_5__3518_,
  data_stage_5__3517_,data_stage_5__3516_,data_stage_5__3515_,data_stage_5__3514_,
  data_stage_5__3513_,data_stage_5__3512_,data_stage_5__3511_,data_stage_5__3510_,
  data_stage_5__3509_,data_stage_5__3508_,data_stage_5__3507_,data_stage_5__3506_,
  data_stage_5__3505_,data_stage_5__3504_,data_stage_5__3503_,data_stage_5__3502_,
  data_stage_5__3501_,data_stage_5__3500_,data_stage_5__3499_,data_stage_5__3498_,
  data_stage_5__3497_,data_stage_5__3496_,data_stage_5__3495_,data_stage_5__3494_,
  data_stage_5__3493_,data_stage_5__3492_,data_stage_5__3491_,data_stage_5__3490_,
  data_stage_5__3489_,data_stage_5__3488_,data_stage_5__3487_,data_stage_5__3486_,
  data_stage_5__3485_,data_stage_5__3484_,data_stage_5__3483_,data_stage_5__3482_,
  data_stage_5__3481_,data_stage_5__3480_,data_stage_5__3479_,data_stage_5__3478_,
  data_stage_5__3477_,data_stage_5__3476_,data_stage_5__3475_,data_stage_5__3474_,
  data_stage_5__3473_,data_stage_5__3472_,data_stage_5__3471_,data_stage_5__3470_,
  data_stage_5__3469_,data_stage_5__3468_,data_stage_5__3467_,data_stage_5__3466_,
  data_stage_5__3465_,data_stage_5__3464_,data_stage_5__3463_,data_stage_5__3462_,
  data_stage_5__3461_,data_stage_5__3460_,data_stage_5__3459_,data_stage_5__3458_,
  data_stage_5__3457_,data_stage_5__3456_,data_stage_5__3455_,data_stage_5__3454_,
  data_stage_5__3453_,data_stage_5__3452_,data_stage_5__3451_,data_stage_5__3450_,
  data_stage_5__3449_,data_stage_5__3448_,data_stage_5__3447_,data_stage_5__3446_,
  data_stage_5__3445_,data_stage_5__3444_,data_stage_5__3443_,data_stage_5__3442_,
  data_stage_5__3441_,data_stage_5__3440_,data_stage_5__3439_,data_stage_5__3438_,
  data_stage_5__3437_,data_stage_5__3436_,data_stage_5__3435_,data_stage_5__3434_,
  data_stage_5__3433_,data_stage_5__3432_,data_stage_5__3431_,data_stage_5__3430_,
  data_stage_5__3429_,data_stage_5__3428_,data_stage_5__3427_,data_stage_5__3426_,
  data_stage_5__3425_,data_stage_5__3424_,data_stage_5__3423_,data_stage_5__3422_,
  data_stage_5__3421_,data_stage_5__3420_,data_stage_5__3419_,data_stage_5__3418_,
  data_stage_5__3417_,data_stage_5__3416_,data_stage_5__3415_,data_stage_5__3414_,
  data_stage_5__3413_,data_stage_5__3412_,data_stage_5__3411_,data_stage_5__3410_,
  data_stage_5__3409_,data_stage_5__3408_,data_stage_5__3407_,data_stage_5__3406_,
  data_stage_5__3405_,data_stage_5__3404_,data_stage_5__3403_,data_stage_5__3402_,
  data_stage_5__3401_,data_stage_5__3400_,data_stage_5__3399_,data_stage_5__3398_,
  data_stage_5__3397_,data_stage_5__3396_,data_stage_5__3395_,data_stage_5__3394_,
  data_stage_5__3393_,data_stage_5__3392_,data_stage_5__3391_,data_stage_5__3390_,
  data_stage_5__3389_,data_stage_5__3388_,data_stage_5__3387_,data_stage_5__3386_,
  data_stage_5__3385_,data_stage_5__3384_,data_stage_5__3383_,data_stage_5__3382_,
  data_stage_5__3381_,data_stage_5__3380_,data_stage_5__3379_,data_stage_5__3378_,
  data_stage_5__3377_,data_stage_5__3376_,data_stage_5__3375_,data_stage_5__3374_,
  data_stage_5__3373_,data_stage_5__3372_,data_stage_5__3371_,data_stage_5__3370_,
  data_stage_5__3369_,data_stage_5__3368_,data_stage_5__3367_,data_stage_5__3366_,
  data_stage_5__3365_,data_stage_5__3364_,data_stage_5__3363_,data_stage_5__3362_,
  data_stage_5__3361_,data_stage_5__3360_,data_stage_5__3359_,data_stage_5__3358_,
  data_stage_5__3357_,data_stage_5__3356_,data_stage_5__3355_,data_stage_5__3354_,
  data_stage_5__3353_,data_stage_5__3352_,data_stage_5__3351_,data_stage_5__3350_,
  data_stage_5__3349_,data_stage_5__3348_,data_stage_5__3347_,data_stage_5__3346_,
  data_stage_5__3345_,data_stage_5__3344_,data_stage_5__3343_,data_stage_5__3342_,
  data_stage_5__3341_,data_stage_5__3340_,data_stage_5__3339_,data_stage_5__3338_,
  data_stage_5__3337_,data_stage_5__3336_,data_stage_5__3335_,data_stage_5__3334_,
  data_stage_5__3333_,data_stage_5__3332_,data_stage_5__3331_,data_stage_5__3330_,
  data_stage_5__3329_,data_stage_5__3328_,data_stage_5__3327_,data_stage_5__3326_,
  data_stage_5__3325_,data_stage_5__3324_,data_stage_5__3323_,data_stage_5__3322_,
  data_stage_5__3321_,data_stage_5__3320_,data_stage_5__3319_,data_stage_5__3318_,
  data_stage_5__3317_,data_stage_5__3316_,data_stage_5__3315_,data_stage_5__3314_,
  data_stage_5__3313_,data_stage_5__3312_,data_stage_5__3311_,data_stage_5__3310_,
  data_stage_5__3309_,data_stage_5__3308_,data_stage_5__3307_,data_stage_5__3306_,
  data_stage_5__3305_,data_stage_5__3304_,data_stage_5__3303_,data_stage_5__3302_,
  data_stage_5__3301_,data_stage_5__3300_,data_stage_5__3299_,data_stage_5__3298_,
  data_stage_5__3297_,data_stage_5__3296_,data_stage_5__3295_,data_stage_5__3294_,
  data_stage_5__3293_,data_stage_5__3292_,data_stage_5__3291_,data_stage_5__3290_,
  data_stage_5__3289_,data_stage_5__3288_,data_stage_5__3287_,data_stage_5__3286_,
  data_stage_5__3285_,data_stage_5__3284_,data_stage_5__3283_,data_stage_5__3282_,
  data_stage_5__3281_,data_stage_5__3280_,data_stage_5__3279_,data_stage_5__3278_,
  data_stage_5__3277_,data_stage_5__3276_,data_stage_5__3275_,data_stage_5__3274_,
  data_stage_5__3273_,data_stage_5__3272_,data_stage_5__3271_,data_stage_5__3270_,
  data_stage_5__3269_,data_stage_5__3268_,data_stage_5__3267_,data_stage_5__3266_,
  data_stage_5__3265_,data_stage_5__3264_,data_stage_5__3263_,data_stage_5__3262_,
  data_stage_5__3261_,data_stage_5__3260_,data_stage_5__3259_,data_stage_5__3258_,
  data_stage_5__3257_,data_stage_5__3256_,data_stage_5__3255_,data_stage_5__3254_,
  data_stage_5__3253_,data_stage_5__3252_,data_stage_5__3251_,data_stage_5__3250_,
  data_stage_5__3249_,data_stage_5__3248_,data_stage_5__3247_,data_stage_5__3246_,
  data_stage_5__3245_,data_stage_5__3244_,data_stage_5__3243_,data_stage_5__3242_,
  data_stage_5__3241_,data_stage_5__3240_,data_stage_5__3239_,data_stage_5__3238_,
  data_stage_5__3237_,data_stage_5__3236_,data_stage_5__3235_,data_stage_5__3234_,
  data_stage_5__3233_,data_stage_5__3232_,data_stage_5__3231_,data_stage_5__3230_,
  data_stage_5__3229_,data_stage_5__3228_,data_stage_5__3227_,data_stage_5__3226_,
  data_stage_5__3225_,data_stage_5__3224_,data_stage_5__3223_,data_stage_5__3222_,
  data_stage_5__3221_,data_stage_5__3220_,data_stage_5__3219_,data_stage_5__3218_,
  data_stage_5__3217_,data_stage_5__3216_,data_stage_5__3215_,data_stage_5__3214_,
  data_stage_5__3213_,data_stage_5__3212_,data_stage_5__3211_,data_stage_5__3210_,
  data_stage_5__3209_,data_stage_5__3208_,data_stage_5__3207_,data_stage_5__3206_,
  data_stage_5__3205_,data_stage_5__3204_,data_stage_5__3203_,data_stage_5__3202_,
  data_stage_5__3201_,data_stage_5__3200_,data_stage_5__3199_,data_stage_5__3198_,
  data_stage_5__3197_,data_stage_5__3196_,data_stage_5__3195_,data_stage_5__3194_,
  data_stage_5__3193_,data_stage_5__3192_,data_stage_5__3191_,data_stage_5__3190_,
  data_stage_5__3189_,data_stage_5__3188_,data_stage_5__3187_,data_stage_5__3186_,
  data_stage_5__3185_,data_stage_5__3184_,data_stage_5__3183_,data_stage_5__3182_,
  data_stage_5__3181_,data_stage_5__3180_,data_stage_5__3179_,data_stage_5__3178_,
  data_stage_5__3177_,data_stage_5__3176_,data_stage_5__3175_,data_stage_5__3174_,
  data_stage_5__3173_,data_stage_5__3172_,data_stage_5__3171_,data_stage_5__3170_,
  data_stage_5__3169_,data_stage_5__3168_,data_stage_5__3167_,data_stage_5__3166_,
  data_stage_5__3165_,data_stage_5__3164_,data_stage_5__3163_,data_stage_5__3162_,
  data_stage_5__3161_,data_stage_5__3160_,data_stage_5__3159_,data_stage_5__3158_,
  data_stage_5__3157_,data_stage_5__3156_,data_stage_5__3155_,data_stage_5__3154_,
  data_stage_5__3153_,data_stage_5__3152_,data_stage_5__3151_,data_stage_5__3150_,
  data_stage_5__3149_,data_stage_5__3148_,data_stage_5__3147_,data_stage_5__3146_,
  data_stage_5__3145_,data_stage_5__3144_,data_stage_5__3143_,data_stage_5__3142_,
  data_stage_5__3141_,data_stage_5__3140_,data_stage_5__3139_,data_stage_5__3138_,
  data_stage_5__3137_,data_stage_5__3136_,data_stage_5__3135_,data_stage_5__3134_,
  data_stage_5__3133_,data_stage_5__3132_,data_stage_5__3131_,data_stage_5__3130_,
  data_stage_5__3129_,data_stage_5__3128_,data_stage_5__3127_,data_stage_5__3126_,
  data_stage_5__3125_,data_stage_5__3124_,data_stage_5__3123_,data_stage_5__3122_,
  data_stage_5__3121_,data_stage_5__3120_,data_stage_5__3119_,data_stage_5__3118_,
  data_stage_5__3117_,data_stage_5__3116_,data_stage_5__3115_,data_stage_5__3114_,
  data_stage_5__3113_,data_stage_5__3112_,data_stage_5__3111_,data_stage_5__3110_,
  data_stage_5__3109_,data_stage_5__3108_,data_stage_5__3107_,data_stage_5__3106_,
  data_stage_5__3105_,data_stage_5__3104_,data_stage_5__3103_,data_stage_5__3102_,
  data_stage_5__3101_,data_stage_5__3100_,data_stage_5__3099_,data_stage_5__3098_,
  data_stage_5__3097_,data_stage_5__3096_,data_stage_5__3095_,data_stage_5__3094_,
  data_stage_5__3093_,data_stage_5__3092_,data_stage_5__3091_,data_stage_5__3090_,
  data_stage_5__3089_,data_stage_5__3088_,data_stage_5__3087_,data_stage_5__3086_,
  data_stage_5__3085_,data_stage_5__3084_,data_stage_5__3083_,data_stage_5__3082_,
  data_stage_5__3081_,data_stage_5__3080_,data_stage_5__3079_,data_stage_5__3078_,
  data_stage_5__3077_,data_stage_5__3076_,data_stage_5__3075_,data_stage_5__3074_,
  data_stage_5__3073_,data_stage_5__3072_,data_stage_5__3071_,data_stage_5__3070_,
  data_stage_5__3069_,data_stage_5__3068_,data_stage_5__3067_,data_stage_5__3066_,
  data_stage_5__3065_,data_stage_5__3064_,data_stage_5__3063_,data_stage_5__3062_,
  data_stage_5__3061_,data_stage_5__3060_,data_stage_5__3059_,data_stage_5__3058_,
  data_stage_5__3057_,data_stage_5__3056_,data_stage_5__3055_,data_stage_5__3054_,
  data_stage_5__3053_,data_stage_5__3052_,data_stage_5__3051_,data_stage_5__3050_,
  data_stage_5__3049_,data_stage_5__3048_,data_stage_5__3047_,data_stage_5__3046_,
  data_stage_5__3045_,data_stage_5__3044_,data_stage_5__3043_,data_stage_5__3042_,
  data_stage_5__3041_,data_stage_5__3040_,data_stage_5__3039_,data_stage_5__3038_,
  data_stage_5__3037_,data_stage_5__3036_,data_stage_5__3035_,data_stage_5__3034_,
  data_stage_5__3033_,data_stage_5__3032_,data_stage_5__3031_,data_stage_5__3030_,
  data_stage_5__3029_,data_stage_5__3028_,data_stage_5__3027_,data_stage_5__3026_,
  data_stage_5__3025_,data_stage_5__3024_,data_stage_5__3023_,data_stage_5__3022_,
  data_stage_5__3021_,data_stage_5__3020_,data_stage_5__3019_,data_stage_5__3018_,
  data_stage_5__3017_,data_stage_5__3016_,data_stage_5__3015_,data_stage_5__3014_,
  data_stage_5__3013_,data_stage_5__3012_,data_stage_5__3011_,data_stage_5__3010_,
  data_stage_5__3009_,data_stage_5__3008_,data_stage_5__3007_,data_stage_5__3006_,
  data_stage_5__3005_,data_stage_5__3004_,data_stage_5__3003_,data_stage_5__3002_,
  data_stage_5__3001_,data_stage_5__3000_,data_stage_5__2999_,data_stage_5__2998_,
  data_stage_5__2997_,data_stage_5__2996_,data_stage_5__2995_,data_stage_5__2994_,
  data_stage_5__2993_,data_stage_5__2992_,data_stage_5__2991_,data_stage_5__2990_,
  data_stage_5__2989_,data_stage_5__2988_,data_stage_5__2987_,data_stage_5__2986_,
  data_stage_5__2985_,data_stage_5__2984_,data_stage_5__2983_,data_stage_5__2982_,
  data_stage_5__2981_,data_stage_5__2980_,data_stage_5__2979_,data_stage_5__2978_,
  data_stage_5__2977_,data_stage_5__2976_,data_stage_5__2975_,data_stage_5__2974_,
  data_stage_5__2973_,data_stage_5__2972_,data_stage_5__2971_,data_stage_5__2970_,
  data_stage_5__2969_,data_stage_5__2968_,data_stage_5__2967_,data_stage_5__2966_,
  data_stage_5__2965_,data_stage_5__2964_,data_stage_5__2963_,data_stage_5__2962_,
  data_stage_5__2961_,data_stage_5__2960_,data_stage_5__2959_,data_stage_5__2958_,
  data_stage_5__2957_,data_stage_5__2956_,data_stage_5__2955_,data_stage_5__2954_,
  data_stage_5__2953_,data_stage_5__2952_,data_stage_5__2951_,data_stage_5__2950_,
  data_stage_5__2949_,data_stage_5__2948_,data_stage_5__2947_,data_stage_5__2946_,
  data_stage_5__2945_,data_stage_5__2944_,data_stage_5__2943_,data_stage_5__2942_,
  data_stage_5__2941_,data_stage_5__2940_,data_stage_5__2939_,data_stage_5__2938_,
  data_stage_5__2937_,data_stage_5__2936_,data_stage_5__2935_,data_stage_5__2934_,
  data_stage_5__2933_,data_stage_5__2932_,data_stage_5__2931_,data_stage_5__2930_,
  data_stage_5__2929_,data_stage_5__2928_,data_stage_5__2927_,data_stage_5__2926_,
  data_stage_5__2925_,data_stage_5__2924_,data_stage_5__2923_,data_stage_5__2922_,
  data_stage_5__2921_,data_stage_5__2920_,data_stage_5__2919_,data_stage_5__2918_,
  data_stage_5__2917_,data_stage_5__2916_,data_stage_5__2915_,data_stage_5__2914_,
  data_stage_5__2913_,data_stage_5__2912_,data_stage_5__2911_,data_stage_5__2910_,
  data_stage_5__2909_,data_stage_5__2908_,data_stage_5__2907_,data_stage_5__2906_,
  data_stage_5__2905_,data_stage_5__2904_,data_stage_5__2903_,data_stage_5__2902_,
  data_stage_5__2901_,data_stage_5__2900_,data_stage_5__2899_,data_stage_5__2898_,
  data_stage_5__2897_,data_stage_5__2896_,data_stage_5__2895_,data_stage_5__2894_,
  data_stage_5__2893_,data_stage_5__2892_,data_stage_5__2891_,data_stage_5__2890_,
  data_stage_5__2889_,data_stage_5__2888_,data_stage_5__2887_,data_stage_5__2886_,
  data_stage_5__2885_,data_stage_5__2884_,data_stage_5__2883_,data_stage_5__2882_,
  data_stage_5__2881_,data_stage_5__2880_,data_stage_5__2879_,data_stage_5__2878_,
  data_stage_5__2877_,data_stage_5__2876_,data_stage_5__2875_,data_stage_5__2874_,
  data_stage_5__2873_,data_stage_5__2872_,data_stage_5__2871_,data_stage_5__2870_,
  data_stage_5__2869_,data_stage_5__2868_,data_stage_5__2867_,data_stage_5__2866_,
  data_stage_5__2865_,data_stage_5__2864_,data_stage_5__2863_,data_stage_5__2862_,
  data_stage_5__2861_,data_stage_5__2860_,data_stage_5__2859_,data_stage_5__2858_,
  data_stage_5__2857_,data_stage_5__2856_,data_stage_5__2855_,data_stage_5__2854_,
  data_stage_5__2853_,data_stage_5__2852_,data_stage_5__2851_,data_stage_5__2850_,
  data_stage_5__2849_,data_stage_5__2848_,data_stage_5__2847_,data_stage_5__2846_,
  data_stage_5__2845_,data_stage_5__2844_,data_stage_5__2843_,data_stage_5__2842_,
  data_stage_5__2841_,data_stage_5__2840_,data_stage_5__2839_,data_stage_5__2838_,
  data_stage_5__2837_,data_stage_5__2836_,data_stage_5__2835_,data_stage_5__2834_,
  data_stage_5__2833_,data_stage_5__2832_,data_stage_5__2831_,data_stage_5__2830_,
  data_stage_5__2829_,data_stage_5__2828_,data_stage_5__2827_,data_stage_5__2826_,
  data_stage_5__2825_,data_stage_5__2824_,data_stage_5__2823_,data_stage_5__2822_,
  data_stage_5__2821_,data_stage_5__2820_,data_stage_5__2819_,data_stage_5__2818_,
  data_stage_5__2817_,data_stage_5__2816_,data_stage_5__2815_,data_stage_5__2814_,
  data_stage_5__2813_,data_stage_5__2812_,data_stage_5__2811_,data_stage_5__2810_,
  data_stage_5__2809_,data_stage_5__2808_,data_stage_5__2807_,data_stage_5__2806_,
  data_stage_5__2805_,data_stage_5__2804_,data_stage_5__2803_,data_stage_5__2802_,
  data_stage_5__2801_,data_stage_5__2800_,data_stage_5__2799_,data_stage_5__2798_,
  data_stage_5__2797_,data_stage_5__2796_,data_stage_5__2795_,data_stage_5__2794_,
  data_stage_5__2793_,data_stage_5__2792_,data_stage_5__2791_,data_stage_5__2790_,
  data_stage_5__2789_,data_stage_5__2788_,data_stage_5__2787_,data_stage_5__2786_,
  data_stage_5__2785_,data_stage_5__2784_,data_stage_5__2783_,data_stage_5__2782_,
  data_stage_5__2781_,data_stage_5__2780_,data_stage_5__2779_,data_stage_5__2778_,
  data_stage_5__2777_,data_stage_5__2776_,data_stage_5__2775_,data_stage_5__2774_,
  data_stage_5__2773_,data_stage_5__2772_,data_stage_5__2771_,data_stage_5__2770_,
  data_stage_5__2769_,data_stage_5__2768_,data_stage_5__2767_,data_stage_5__2766_,
  data_stage_5__2765_,data_stage_5__2764_,data_stage_5__2763_,data_stage_5__2762_,
  data_stage_5__2761_,data_stage_5__2760_,data_stage_5__2759_,data_stage_5__2758_,
  data_stage_5__2757_,data_stage_5__2756_,data_stage_5__2755_,data_stage_5__2754_,
  data_stage_5__2753_,data_stage_5__2752_,data_stage_5__2751_,data_stage_5__2750_,
  data_stage_5__2749_,data_stage_5__2748_,data_stage_5__2747_,data_stage_5__2746_,
  data_stage_5__2745_,data_stage_5__2744_,data_stage_5__2743_,data_stage_5__2742_,
  data_stage_5__2741_,data_stage_5__2740_,data_stage_5__2739_,data_stage_5__2738_,
  data_stage_5__2737_,data_stage_5__2736_,data_stage_5__2735_,data_stage_5__2734_,
  data_stage_5__2733_,data_stage_5__2732_,data_stage_5__2731_,data_stage_5__2730_,
  data_stage_5__2729_,data_stage_5__2728_,data_stage_5__2727_,data_stage_5__2726_,
  data_stage_5__2725_,data_stage_5__2724_,data_stage_5__2723_,data_stage_5__2722_,
  data_stage_5__2721_,data_stage_5__2720_,data_stage_5__2719_,data_stage_5__2718_,
  data_stage_5__2717_,data_stage_5__2716_,data_stage_5__2715_,data_stage_5__2714_,
  data_stage_5__2713_,data_stage_5__2712_,data_stage_5__2711_,data_stage_5__2710_,
  data_stage_5__2709_,data_stage_5__2708_,data_stage_5__2707_,data_stage_5__2706_,
  data_stage_5__2705_,data_stage_5__2704_,data_stage_5__2703_,data_stage_5__2702_,
  data_stage_5__2701_,data_stage_5__2700_,data_stage_5__2699_,data_stage_5__2698_,
  data_stage_5__2697_,data_stage_5__2696_,data_stage_5__2695_,data_stage_5__2694_,
  data_stage_5__2693_,data_stage_5__2692_,data_stage_5__2691_,data_stage_5__2690_,
  data_stage_5__2689_,data_stage_5__2688_,data_stage_5__2687_,data_stage_5__2686_,
  data_stage_5__2685_,data_stage_5__2684_,data_stage_5__2683_,data_stage_5__2682_,
  data_stage_5__2681_,data_stage_5__2680_,data_stage_5__2679_,data_stage_5__2678_,
  data_stage_5__2677_,data_stage_5__2676_,data_stage_5__2675_,data_stage_5__2674_,
  data_stage_5__2673_,data_stage_5__2672_,data_stage_5__2671_,data_stage_5__2670_,
  data_stage_5__2669_,data_stage_5__2668_,data_stage_5__2667_,data_stage_5__2666_,
  data_stage_5__2665_,data_stage_5__2664_,data_stage_5__2663_,data_stage_5__2662_,
  data_stage_5__2661_,data_stage_5__2660_,data_stage_5__2659_,data_stage_5__2658_,
  data_stage_5__2657_,data_stage_5__2656_,data_stage_5__2655_,data_stage_5__2654_,
  data_stage_5__2653_,data_stage_5__2652_,data_stage_5__2651_,data_stage_5__2650_,
  data_stage_5__2649_,data_stage_5__2648_,data_stage_5__2647_,data_stage_5__2646_,
  data_stage_5__2645_,data_stage_5__2644_,data_stage_5__2643_,data_stage_5__2642_,
  data_stage_5__2641_,data_stage_5__2640_,data_stage_5__2639_,data_stage_5__2638_,
  data_stage_5__2637_,data_stage_5__2636_,data_stage_5__2635_,data_stage_5__2634_,
  data_stage_5__2633_,data_stage_5__2632_,data_stage_5__2631_,data_stage_5__2630_,
  data_stage_5__2629_,data_stage_5__2628_,data_stage_5__2627_,data_stage_5__2626_,
  data_stage_5__2625_,data_stage_5__2624_,data_stage_5__2623_,data_stage_5__2622_,
  data_stage_5__2621_,data_stage_5__2620_,data_stage_5__2619_,data_stage_5__2618_,
  data_stage_5__2617_,data_stage_5__2616_,data_stage_5__2615_,data_stage_5__2614_,
  data_stage_5__2613_,data_stage_5__2612_,data_stage_5__2611_,data_stage_5__2610_,
  data_stage_5__2609_,data_stage_5__2608_,data_stage_5__2607_,data_stage_5__2606_,
  data_stage_5__2605_,data_stage_5__2604_,data_stage_5__2603_,data_stage_5__2602_,
  data_stage_5__2601_,data_stage_5__2600_,data_stage_5__2599_,data_stage_5__2598_,
  data_stage_5__2597_,data_stage_5__2596_,data_stage_5__2595_,data_stage_5__2594_,
  data_stage_5__2593_,data_stage_5__2592_,data_stage_5__2591_,data_stage_5__2590_,
  data_stage_5__2589_,data_stage_5__2588_,data_stage_5__2587_,data_stage_5__2586_,
  data_stage_5__2585_,data_stage_5__2584_,data_stage_5__2583_,data_stage_5__2582_,
  data_stage_5__2581_,data_stage_5__2580_,data_stage_5__2579_,data_stage_5__2578_,
  data_stage_5__2577_,data_stage_5__2576_,data_stage_5__2575_,data_stage_5__2574_,
  data_stage_5__2573_,data_stage_5__2572_,data_stage_5__2571_,data_stage_5__2570_,
  data_stage_5__2569_,data_stage_5__2568_,data_stage_5__2567_,data_stage_5__2566_,
  data_stage_5__2565_,data_stage_5__2564_,data_stage_5__2563_,data_stage_5__2562_,
  data_stage_5__2561_,data_stage_5__2560_,data_stage_5__2559_,data_stage_5__2558_,
  data_stage_5__2557_,data_stage_5__2556_,data_stage_5__2555_,data_stage_5__2554_,
  data_stage_5__2553_,data_stage_5__2552_,data_stage_5__2551_,data_stage_5__2550_,
  data_stage_5__2549_,data_stage_5__2548_,data_stage_5__2547_,data_stage_5__2546_,
  data_stage_5__2545_,data_stage_5__2544_,data_stage_5__2543_,data_stage_5__2542_,
  data_stage_5__2541_,data_stage_5__2540_,data_stage_5__2539_,data_stage_5__2538_,
  data_stage_5__2537_,data_stage_5__2536_,data_stage_5__2535_,data_stage_5__2534_,
  data_stage_5__2533_,data_stage_5__2532_,data_stage_5__2531_,data_stage_5__2530_,
  data_stage_5__2529_,data_stage_5__2528_,data_stage_5__2527_,data_stage_5__2526_,
  data_stage_5__2525_,data_stage_5__2524_,data_stage_5__2523_,data_stage_5__2522_,
  data_stage_5__2521_,data_stage_5__2520_,data_stage_5__2519_,data_stage_5__2518_,
  data_stage_5__2517_,data_stage_5__2516_,data_stage_5__2515_,data_stage_5__2514_,
  data_stage_5__2513_,data_stage_5__2512_,data_stage_5__2511_,data_stage_5__2510_,
  data_stage_5__2509_,data_stage_5__2508_,data_stage_5__2507_,data_stage_5__2506_,
  data_stage_5__2505_,data_stage_5__2504_,data_stage_5__2503_,data_stage_5__2502_,
  data_stage_5__2501_,data_stage_5__2500_,data_stage_5__2499_,data_stage_5__2498_,
  data_stage_5__2497_,data_stage_5__2496_,data_stage_5__2495_,data_stage_5__2494_,
  data_stage_5__2493_,data_stage_5__2492_,data_stage_5__2491_,data_stage_5__2490_,
  data_stage_5__2489_,data_stage_5__2488_,data_stage_5__2487_,data_stage_5__2486_,
  data_stage_5__2485_,data_stage_5__2484_,data_stage_5__2483_,data_stage_5__2482_,
  data_stage_5__2481_,data_stage_5__2480_,data_stage_5__2479_,data_stage_5__2478_,
  data_stage_5__2477_,data_stage_5__2476_,data_stage_5__2475_,data_stage_5__2474_,
  data_stage_5__2473_,data_stage_5__2472_,data_stage_5__2471_,data_stage_5__2470_,
  data_stage_5__2469_,data_stage_5__2468_,data_stage_5__2467_,data_stage_5__2466_,
  data_stage_5__2465_,data_stage_5__2464_,data_stage_5__2463_,data_stage_5__2462_,
  data_stage_5__2461_,data_stage_5__2460_,data_stage_5__2459_,data_stage_5__2458_,
  data_stage_5__2457_,data_stage_5__2456_,data_stage_5__2455_,data_stage_5__2454_,
  data_stage_5__2453_,data_stage_5__2452_,data_stage_5__2451_,data_stage_5__2450_,
  data_stage_5__2449_,data_stage_5__2448_,data_stage_5__2447_,data_stage_5__2446_,
  data_stage_5__2445_,data_stage_5__2444_,data_stage_5__2443_,data_stage_5__2442_,
  data_stage_5__2441_,data_stage_5__2440_,data_stage_5__2439_,data_stage_5__2438_,
  data_stage_5__2437_,data_stage_5__2436_,data_stage_5__2435_,data_stage_5__2434_,
  data_stage_5__2433_,data_stage_5__2432_,data_stage_5__2431_,data_stage_5__2430_,
  data_stage_5__2429_,data_stage_5__2428_,data_stage_5__2427_,data_stage_5__2426_,
  data_stage_5__2425_,data_stage_5__2424_,data_stage_5__2423_,data_stage_5__2422_,
  data_stage_5__2421_,data_stage_5__2420_,data_stage_5__2419_,data_stage_5__2418_,
  data_stage_5__2417_,data_stage_5__2416_,data_stage_5__2415_,data_stage_5__2414_,
  data_stage_5__2413_,data_stage_5__2412_,data_stage_5__2411_,data_stage_5__2410_,
  data_stage_5__2409_,data_stage_5__2408_,data_stage_5__2407_,data_stage_5__2406_,
  data_stage_5__2405_,data_stage_5__2404_,data_stage_5__2403_,data_stage_5__2402_,
  data_stage_5__2401_,data_stage_5__2400_,data_stage_5__2399_,data_stage_5__2398_,
  data_stage_5__2397_,data_stage_5__2396_,data_stage_5__2395_,data_stage_5__2394_,
  data_stage_5__2393_,data_stage_5__2392_,data_stage_5__2391_,data_stage_5__2390_,
  data_stage_5__2389_,data_stage_5__2388_,data_stage_5__2387_,data_stage_5__2386_,
  data_stage_5__2385_,data_stage_5__2384_,data_stage_5__2383_,data_stage_5__2382_,
  data_stage_5__2381_,data_stage_5__2380_,data_stage_5__2379_,data_stage_5__2378_,
  data_stage_5__2377_,data_stage_5__2376_,data_stage_5__2375_,data_stage_5__2374_,
  data_stage_5__2373_,data_stage_5__2372_,data_stage_5__2371_,data_stage_5__2370_,
  data_stage_5__2369_,data_stage_5__2368_,data_stage_5__2367_,data_stage_5__2366_,
  data_stage_5__2365_,data_stage_5__2364_,data_stage_5__2363_,data_stage_5__2362_,
  data_stage_5__2361_,data_stage_5__2360_,data_stage_5__2359_,data_stage_5__2358_,
  data_stage_5__2357_,data_stage_5__2356_,data_stage_5__2355_,data_stage_5__2354_,
  data_stage_5__2353_,data_stage_5__2352_,data_stage_5__2351_,data_stage_5__2350_,
  data_stage_5__2349_,data_stage_5__2348_,data_stage_5__2347_,data_stage_5__2346_,
  data_stage_5__2345_,data_stage_5__2344_,data_stage_5__2343_,data_stage_5__2342_,
  data_stage_5__2341_,data_stage_5__2340_,data_stage_5__2339_,data_stage_5__2338_,
  data_stage_5__2337_,data_stage_5__2336_,data_stage_5__2335_,data_stage_5__2334_,
  data_stage_5__2333_,data_stage_5__2332_,data_stage_5__2331_,data_stage_5__2330_,
  data_stage_5__2329_,data_stage_5__2328_,data_stage_5__2327_,data_stage_5__2326_,
  data_stage_5__2325_,data_stage_5__2324_,data_stage_5__2323_,data_stage_5__2322_,
  data_stage_5__2321_,data_stage_5__2320_,data_stage_5__2319_,data_stage_5__2318_,
  data_stage_5__2317_,data_stage_5__2316_,data_stage_5__2315_,data_stage_5__2314_,
  data_stage_5__2313_,data_stage_5__2312_,data_stage_5__2311_,data_stage_5__2310_,
  data_stage_5__2309_,data_stage_5__2308_,data_stage_5__2307_,data_stage_5__2306_,
  data_stage_5__2305_,data_stage_5__2304_,data_stage_5__2303_,data_stage_5__2302_,
  data_stage_5__2301_,data_stage_5__2300_,data_stage_5__2299_,data_stage_5__2298_,
  data_stage_5__2297_,data_stage_5__2296_,data_stage_5__2295_,data_stage_5__2294_,
  data_stage_5__2293_,data_stage_5__2292_,data_stage_5__2291_,data_stage_5__2290_,
  data_stage_5__2289_,data_stage_5__2288_,data_stage_5__2287_,data_stage_5__2286_,
  data_stage_5__2285_,data_stage_5__2284_,data_stage_5__2283_,data_stage_5__2282_,
  data_stage_5__2281_,data_stage_5__2280_,data_stage_5__2279_,data_stage_5__2278_,
  data_stage_5__2277_,data_stage_5__2276_,data_stage_5__2275_,data_stage_5__2274_,
  data_stage_5__2273_,data_stage_5__2272_,data_stage_5__2271_,data_stage_5__2270_,
  data_stage_5__2269_,data_stage_5__2268_,data_stage_5__2267_,data_stage_5__2266_,
  data_stage_5__2265_,data_stage_5__2264_,data_stage_5__2263_,data_stage_5__2262_,
  data_stage_5__2261_,data_stage_5__2260_,data_stage_5__2259_,data_stage_5__2258_,
  data_stage_5__2257_,data_stage_5__2256_,data_stage_5__2255_,data_stage_5__2254_,
  data_stage_5__2253_,data_stage_5__2252_,data_stage_5__2251_,data_stage_5__2250_,
  data_stage_5__2249_,data_stage_5__2248_,data_stage_5__2247_,data_stage_5__2246_,
  data_stage_5__2245_,data_stage_5__2244_,data_stage_5__2243_,data_stage_5__2242_,
  data_stage_5__2241_,data_stage_5__2240_,data_stage_5__2239_,data_stage_5__2238_,
  data_stage_5__2237_,data_stage_5__2236_,data_stage_5__2235_,data_stage_5__2234_,
  data_stage_5__2233_,data_stage_5__2232_,data_stage_5__2231_,data_stage_5__2230_,
  data_stage_5__2229_,data_stage_5__2228_,data_stage_5__2227_,data_stage_5__2226_,
  data_stage_5__2225_,data_stage_5__2224_,data_stage_5__2223_,data_stage_5__2222_,
  data_stage_5__2221_,data_stage_5__2220_,data_stage_5__2219_,data_stage_5__2218_,
  data_stage_5__2217_,data_stage_5__2216_,data_stage_5__2215_,data_stage_5__2214_,
  data_stage_5__2213_,data_stage_5__2212_,data_stage_5__2211_,data_stage_5__2210_,
  data_stage_5__2209_,data_stage_5__2208_,data_stage_5__2207_,data_stage_5__2206_,
  data_stage_5__2205_,data_stage_5__2204_,data_stage_5__2203_,data_stage_5__2202_,
  data_stage_5__2201_,data_stage_5__2200_,data_stage_5__2199_,data_stage_5__2198_,
  data_stage_5__2197_,data_stage_5__2196_,data_stage_5__2195_,data_stage_5__2194_,
  data_stage_5__2193_,data_stage_5__2192_,data_stage_5__2191_,data_stage_5__2190_,
  data_stage_5__2189_,data_stage_5__2188_,data_stage_5__2187_,data_stage_5__2186_,
  data_stage_5__2185_,data_stage_5__2184_,data_stage_5__2183_,data_stage_5__2182_,
  data_stage_5__2181_,data_stage_5__2180_,data_stage_5__2179_,data_stage_5__2178_,
  data_stage_5__2177_,data_stage_5__2176_,data_stage_5__2175_,data_stage_5__2174_,
  data_stage_5__2173_,data_stage_5__2172_,data_stage_5__2171_,data_stage_5__2170_,
  data_stage_5__2169_,data_stage_5__2168_,data_stage_5__2167_,data_stage_5__2166_,
  data_stage_5__2165_,data_stage_5__2164_,data_stage_5__2163_,data_stage_5__2162_,
  data_stage_5__2161_,data_stage_5__2160_,data_stage_5__2159_,data_stage_5__2158_,
  data_stage_5__2157_,data_stage_5__2156_,data_stage_5__2155_,data_stage_5__2154_,
  data_stage_5__2153_,data_stage_5__2152_,data_stage_5__2151_,data_stage_5__2150_,
  data_stage_5__2149_,data_stage_5__2148_,data_stage_5__2147_,data_stage_5__2146_,
  data_stage_5__2145_,data_stage_5__2144_,data_stage_5__2143_,data_stage_5__2142_,
  data_stage_5__2141_,data_stage_5__2140_,data_stage_5__2139_,data_stage_5__2138_,
  data_stage_5__2137_,data_stage_5__2136_,data_stage_5__2135_,data_stage_5__2134_,
  data_stage_5__2133_,data_stage_5__2132_,data_stage_5__2131_,data_stage_5__2130_,
  data_stage_5__2129_,data_stage_5__2128_,data_stage_5__2127_,data_stage_5__2126_,
  data_stage_5__2125_,data_stage_5__2124_,data_stage_5__2123_,data_stage_5__2122_,
  data_stage_5__2121_,data_stage_5__2120_,data_stage_5__2119_,data_stage_5__2118_,
  data_stage_5__2117_,data_stage_5__2116_,data_stage_5__2115_,data_stage_5__2114_,
  data_stage_5__2113_,data_stage_5__2112_,data_stage_5__2111_,data_stage_5__2110_,
  data_stage_5__2109_,data_stage_5__2108_,data_stage_5__2107_,data_stage_5__2106_,
  data_stage_5__2105_,data_stage_5__2104_,data_stage_5__2103_,data_stage_5__2102_,
  data_stage_5__2101_,data_stage_5__2100_,data_stage_5__2099_,data_stage_5__2098_,
  data_stage_5__2097_,data_stage_5__2096_,data_stage_5__2095_,data_stage_5__2094_,
  data_stage_5__2093_,data_stage_5__2092_,data_stage_5__2091_,data_stage_5__2090_,
  data_stage_5__2089_,data_stage_5__2088_,data_stage_5__2087_,data_stage_5__2086_,
  data_stage_5__2085_,data_stage_5__2084_,data_stage_5__2083_,data_stage_5__2082_,
  data_stage_5__2081_,data_stage_5__2080_,data_stage_5__2079_,data_stage_5__2078_,
  data_stage_5__2077_,data_stage_5__2076_,data_stage_5__2075_,data_stage_5__2074_,
  data_stage_5__2073_,data_stage_5__2072_,data_stage_5__2071_,data_stage_5__2070_,
  data_stage_5__2069_,data_stage_5__2068_,data_stage_5__2067_,data_stage_5__2066_,
  data_stage_5__2065_,data_stage_5__2064_,data_stage_5__2063_,data_stage_5__2062_,
  data_stage_5__2061_,data_stage_5__2060_,data_stage_5__2059_,data_stage_5__2058_,
  data_stage_5__2057_,data_stage_5__2056_,data_stage_5__2055_,data_stage_5__2054_,
  data_stage_5__2053_,data_stage_5__2052_,data_stage_5__2051_,data_stage_5__2050_,
  data_stage_5__2049_,data_stage_5__2048_,data_stage_5__2047_,data_stage_5__2046_,
  data_stage_5__2045_,data_stage_5__2044_,data_stage_5__2043_,data_stage_5__2042_,
  data_stage_5__2041_,data_stage_5__2040_,data_stage_5__2039_,data_stage_5__2038_,
  data_stage_5__2037_,data_stage_5__2036_,data_stage_5__2035_,data_stage_5__2034_,
  data_stage_5__2033_,data_stage_5__2032_,data_stage_5__2031_,data_stage_5__2030_,
  data_stage_5__2029_,data_stage_5__2028_,data_stage_5__2027_,data_stage_5__2026_,
  data_stage_5__2025_,data_stage_5__2024_,data_stage_5__2023_,data_stage_5__2022_,
  data_stage_5__2021_,data_stage_5__2020_,data_stage_5__2019_,data_stage_5__2018_,
  data_stage_5__2017_,data_stage_5__2016_,data_stage_5__2015_,data_stage_5__2014_,
  data_stage_5__2013_,data_stage_5__2012_,data_stage_5__2011_,data_stage_5__2010_,
  data_stage_5__2009_,data_stage_5__2008_,data_stage_5__2007_,data_stage_5__2006_,
  data_stage_5__2005_,data_stage_5__2004_,data_stage_5__2003_,data_stage_5__2002_,
  data_stage_5__2001_,data_stage_5__2000_,data_stage_5__1999_,data_stage_5__1998_,
  data_stage_5__1997_,data_stage_5__1996_,data_stage_5__1995_,data_stage_5__1994_,
  data_stage_5__1993_,data_stage_5__1992_,data_stage_5__1991_,data_stage_5__1990_,
  data_stage_5__1989_,data_stage_5__1988_,data_stage_5__1987_,data_stage_5__1986_,
  data_stage_5__1985_,data_stage_5__1984_,data_stage_5__1983_,data_stage_5__1982_,
  data_stage_5__1981_,data_stage_5__1980_,data_stage_5__1979_,data_stage_5__1978_,
  data_stage_5__1977_,data_stage_5__1976_,data_stage_5__1975_,data_stage_5__1974_,
  data_stage_5__1973_,data_stage_5__1972_,data_stage_5__1971_,data_stage_5__1970_,
  data_stage_5__1969_,data_stage_5__1968_,data_stage_5__1967_,data_stage_5__1966_,
  data_stage_5__1965_,data_stage_5__1964_,data_stage_5__1963_,data_stage_5__1962_,
  data_stage_5__1961_,data_stage_5__1960_,data_stage_5__1959_,data_stage_5__1958_,
  data_stage_5__1957_,data_stage_5__1956_,data_stage_5__1955_,data_stage_5__1954_,
  data_stage_5__1953_,data_stage_5__1952_,data_stage_5__1951_,data_stage_5__1950_,
  data_stage_5__1949_,data_stage_5__1948_,data_stage_5__1947_,data_stage_5__1946_,
  data_stage_5__1945_,data_stage_5__1944_,data_stage_5__1943_,data_stage_5__1942_,
  data_stage_5__1941_,data_stage_5__1940_,data_stage_5__1939_,data_stage_5__1938_,
  data_stage_5__1937_,data_stage_5__1936_,data_stage_5__1935_,data_stage_5__1934_,
  data_stage_5__1933_,data_stage_5__1932_,data_stage_5__1931_,data_stage_5__1930_,
  data_stage_5__1929_,data_stage_5__1928_,data_stage_5__1927_,data_stage_5__1926_,
  data_stage_5__1925_,data_stage_5__1924_,data_stage_5__1923_,data_stage_5__1922_,
  data_stage_5__1921_,data_stage_5__1920_,data_stage_5__1919_,data_stage_5__1918_,
  data_stage_5__1917_,data_stage_5__1916_,data_stage_5__1915_,data_stage_5__1914_,
  data_stage_5__1913_,data_stage_5__1912_,data_stage_5__1911_,data_stage_5__1910_,
  data_stage_5__1909_,data_stage_5__1908_,data_stage_5__1907_,data_stage_5__1906_,
  data_stage_5__1905_,data_stage_5__1904_,data_stage_5__1903_,data_stage_5__1902_,
  data_stage_5__1901_,data_stage_5__1900_,data_stage_5__1899_,data_stage_5__1898_,
  data_stage_5__1897_,data_stage_5__1896_,data_stage_5__1895_,data_stage_5__1894_,
  data_stage_5__1893_,data_stage_5__1892_,data_stage_5__1891_,data_stage_5__1890_,
  data_stage_5__1889_,data_stage_5__1888_,data_stage_5__1887_,data_stage_5__1886_,
  data_stage_5__1885_,data_stage_5__1884_,data_stage_5__1883_,data_stage_5__1882_,
  data_stage_5__1881_,data_stage_5__1880_,data_stage_5__1879_,data_stage_5__1878_,
  data_stage_5__1877_,data_stage_5__1876_,data_stage_5__1875_,data_stage_5__1874_,
  data_stage_5__1873_,data_stage_5__1872_,data_stage_5__1871_,data_stage_5__1870_,
  data_stage_5__1869_,data_stage_5__1868_,data_stage_5__1867_,data_stage_5__1866_,
  data_stage_5__1865_,data_stage_5__1864_,data_stage_5__1863_,data_stage_5__1862_,
  data_stage_5__1861_,data_stage_5__1860_,data_stage_5__1859_,data_stage_5__1858_,
  data_stage_5__1857_,data_stage_5__1856_,data_stage_5__1855_,data_stage_5__1854_,
  data_stage_5__1853_,data_stage_5__1852_,data_stage_5__1851_,data_stage_5__1850_,
  data_stage_5__1849_,data_stage_5__1848_,data_stage_5__1847_,data_stage_5__1846_,
  data_stage_5__1845_,data_stage_5__1844_,data_stage_5__1843_,data_stage_5__1842_,
  data_stage_5__1841_,data_stage_5__1840_,data_stage_5__1839_,data_stage_5__1838_,
  data_stage_5__1837_,data_stage_5__1836_,data_stage_5__1835_,data_stage_5__1834_,
  data_stage_5__1833_,data_stage_5__1832_,data_stage_5__1831_,data_stage_5__1830_,
  data_stage_5__1829_,data_stage_5__1828_,data_stage_5__1827_,data_stage_5__1826_,
  data_stage_5__1825_,data_stage_5__1824_,data_stage_5__1823_,data_stage_5__1822_,
  data_stage_5__1821_,data_stage_5__1820_,data_stage_5__1819_,data_stage_5__1818_,
  data_stage_5__1817_,data_stage_5__1816_,data_stage_5__1815_,data_stage_5__1814_,
  data_stage_5__1813_,data_stage_5__1812_,data_stage_5__1811_,data_stage_5__1810_,
  data_stage_5__1809_,data_stage_5__1808_,data_stage_5__1807_,data_stage_5__1806_,
  data_stage_5__1805_,data_stage_5__1804_,data_stage_5__1803_,data_stage_5__1802_,
  data_stage_5__1801_,data_stage_5__1800_,data_stage_5__1799_,data_stage_5__1798_,
  data_stage_5__1797_,data_stage_5__1796_,data_stage_5__1795_,data_stage_5__1794_,
  data_stage_5__1793_,data_stage_5__1792_,data_stage_5__1791_,data_stage_5__1790_,
  data_stage_5__1789_,data_stage_5__1788_,data_stage_5__1787_,data_stage_5__1786_,
  data_stage_5__1785_,data_stage_5__1784_,data_stage_5__1783_,data_stage_5__1782_,
  data_stage_5__1781_,data_stage_5__1780_,data_stage_5__1779_,data_stage_5__1778_,
  data_stage_5__1777_,data_stage_5__1776_,data_stage_5__1775_,data_stage_5__1774_,
  data_stage_5__1773_,data_stage_5__1772_,data_stage_5__1771_,data_stage_5__1770_,
  data_stage_5__1769_,data_stage_5__1768_,data_stage_5__1767_,data_stage_5__1766_,
  data_stage_5__1765_,data_stage_5__1764_,data_stage_5__1763_,data_stage_5__1762_,
  data_stage_5__1761_,data_stage_5__1760_,data_stage_5__1759_,data_stage_5__1758_,
  data_stage_5__1757_,data_stage_5__1756_,data_stage_5__1755_,data_stage_5__1754_,
  data_stage_5__1753_,data_stage_5__1752_,data_stage_5__1751_,data_stage_5__1750_,
  data_stage_5__1749_,data_stage_5__1748_,data_stage_5__1747_,data_stage_5__1746_,
  data_stage_5__1745_,data_stage_5__1744_,data_stage_5__1743_,data_stage_5__1742_,
  data_stage_5__1741_,data_stage_5__1740_,data_stage_5__1739_,data_stage_5__1738_,
  data_stage_5__1737_,data_stage_5__1736_,data_stage_5__1735_,data_stage_5__1734_,
  data_stage_5__1733_,data_stage_5__1732_,data_stage_5__1731_,data_stage_5__1730_,
  data_stage_5__1729_,data_stage_5__1728_,data_stage_5__1727_,data_stage_5__1726_,
  data_stage_5__1725_,data_stage_5__1724_,data_stage_5__1723_,data_stage_5__1722_,
  data_stage_5__1721_,data_stage_5__1720_,data_stage_5__1719_,data_stage_5__1718_,
  data_stage_5__1717_,data_stage_5__1716_,data_stage_5__1715_,data_stage_5__1714_,
  data_stage_5__1713_,data_stage_5__1712_,data_stage_5__1711_,data_stage_5__1710_,
  data_stage_5__1709_,data_stage_5__1708_,data_stage_5__1707_,data_stage_5__1706_,
  data_stage_5__1705_,data_stage_5__1704_,data_stage_5__1703_,data_stage_5__1702_,
  data_stage_5__1701_,data_stage_5__1700_,data_stage_5__1699_,data_stage_5__1698_,
  data_stage_5__1697_,data_stage_5__1696_,data_stage_5__1695_,data_stage_5__1694_,
  data_stage_5__1693_,data_stage_5__1692_,data_stage_5__1691_,data_stage_5__1690_,
  data_stage_5__1689_,data_stage_5__1688_,data_stage_5__1687_,data_stage_5__1686_,
  data_stage_5__1685_,data_stage_5__1684_,data_stage_5__1683_,data_stage_5__1682_,
  data_stage_5__1681_,data_stage_5__1680_,data_stage_5__1679_,data_stage_5__1678_,
  data_stage_5__1677_,data_stage_5__1676_,data_stage_5__1675_,data_stage_5__1674_,
  data_stage_5__1673_,data_stage_5__1672_,data_stage_5__1671_,data_stage_5__1670_,
  data_stage_5__1669_,data_stage_5__1668_,data_stage_5__1667_,data_stage_5__1666_,
  data_stage_5__1665_,data_stage_5__1664_,data_stage_5__1663_,data_stage_5__1662_,
  data_stage_5__1661_,data_stage_5__1660_,data_stage_5__1659_,data_stage_5__1658_,
  data_stage_5__1657_,data_stage_5__1656_,data_stage_5__1655_,data_stage_5__1654_,
  data_stage_5__1653_,data_stage_5__1652_,data_stage_5__1651_,data_stage_5__1650_,
  data_stage_5__1649_,data_stage_5__1648_,data_stage_5__1647_,data_stage_5__1646_,
  data_stage_5__1645_,data_stage_5__1644_,data_stage_5__1643_,data_stage_5__1642_,
  data_stage_5__1641_,data_stage_5__1640_,data_stage_5__1639_,data_stage_5__1638_,
  data_stage_5__1637_,data_stage_5__1636_,data_stage_5__1635_,data_stage_5__1634_,
  data_stage_5__1633_,data_stage_5__1632_,data_stage_5__1631_,data_stage_5__1630_,
  data_stage_5__1629_,data_stage_5__1628_,data_stage_5__1627_,data_stage_5__1626_,
  data_stage_5__1625_,data_stage_5__1624_,data_stage_5__1623_,data_stage_5__1622_,
  data_stage_5__1621_,data_stage_5__1620_,data_stage_5__1619_,data_stage_5__1618_,
  data_stage_5__1617_,data_stage_5__1616_,data_stage_5__1615_,data_stage_5__1614_,
  data_stage_5__1613_,data_stage_5__1612_,data_stage_5__1611_,data_stage_5__1610_,
  data_stage_5__1609_,data_stage_5__1608_,data_stage_5__1607_,data_stage_5__1606_,
  data_stage_5__1605_,data_stage_5__1604_,data_stage_5__1603_,data_stage_5__1602_,
  data_stage_5__1601_,data_stage_5__1600_,data_stage_5__1599_,data_stage_5__1598_,
  data_stage_5__1597_,data_stage_5__1596_,data_stage_5__1595_,data_stage_5__1594_,
  data_stage_5__1593_,data_stage_5__1592_,data_stage_5__1591_,data_stage_5__1590_,
  data_stage_5__1589_,data_stage_5__1588_,data_stage_5__1587_,data_stage_5__1586_,
  data_stage_5__1585_,data_stage_5__1584_,data_stage_5__1583_,data_stage_5__1582_,
  data_stage_5__1581_,data_stage_5__1580_,data_stage_5__1579_,data_stage_5__1578_,
  data_stage_5__1577_,data_stage_5__1576_,data_stage_5__1575_,data_stage_5__1574_,
  data_stage_5__1573_,data_stage_5__1572_,data_stage_5__1571_,data_stage_5__1570_,
  data_stage_5__1569_,data_stage_5__1568_,data_stage_5__1567_,data_stage_5__1566_,
  data_stage_5__1565_,data_stage_5__1564_,data_stage_5__1563_,data_stage_5__1562_,
  data_stage_5__1561_,data_stage_5__1560_,data_stage_5__1559_,data_stage_5__1558_,
  data_stage_5__1557_,data_stage_5__1556_,data_stage_5__1555_,data_stage_5__1554_,
  data_stage_5__1553_,data_stage_5__1552_,data_stage_5__1551_,data_stage_5__1550_,
  data_stage_5__1549_,data_stage_5__1548_,data_stage_5__1547_,data_stage_5__1546_,
  data_stage_5__1545_,data_stage_5__1544_,data_stage_5__1543_,data_stage_5__1542_,
  data_stage_5__1541_,data_stage_5__1540_,data_stage_5__1539_,data_stage_5__1538_,
  data_stage_5__1537_,data_stage_5__1536_,data_stage_5__1535_,data_stage_5__1534_,
  data_stage_5__1533_,data_stage_5__1532_,data_stage_5__1531_,data_stage_5__1530_,
  data_stage_5__1529_,data_stage_5__1528_,data_stage_5__1527_,data_stage_5__1526_,
  data_stage_5__1525_,data_stage_5__1524_,data_stage_5__1523_,data_stage_5__1522_,
  data_stage_5__1521_,data_stage_5__1520_,data_stage_5__1519_,data_stage_5__1518_,
  data_stage_5__1517_,data_stage_5__1516_,data_stage_5__1515_,data_stage_5__1514_,
  data_stage_5__1513_,data_stage_5__1512_,data_stage_5__1511_,data_stage_5__1510_,
  data_stage_5__1509_,data_stage_5__1508_,data_stage_5__1507_,data_stage_5__1506_,
  data_stage_5__1505_,data_stage_5__1504_,data_stage_5__1503_,data_stage_5__1502_,
  data_stage_5__1501_,data_stage_5__1500_,data_stage_5__1499_,data_stage_5__1498_,
  data_stage_5__1497_,data_stage_5__1496_,data_stage_5__1495_,data_stage_5__1494_,
  data_stage_5__1493_,data_stage_5__1492_,data_stage_5__1491_,data_stage_5__1490_,
  data_stage_5__1489_,data_stage_5__1488_,data_stage_5__1487_,data_stage_5__1486_,
  data_stage_5__1485_,data_stage_5__1484_,data_stage_5__1483_,data_stage_5__1482_,
  data_stage_5__1481_,data_stage_5__1480_,data_stage_5__1479_,data_stage_5__1478_,
  data_stage_5__1477_,data_stage_5__1476_,data_stage_5__1475_,data_stage_5__1474_,
  data_stage_5__1473_,data_stage_5__1472_,data_stage_5__1471_,data_stage_5__1470_,
  data_stage_5__1469_,data_stage_5__1468_,data_stage_5__1467_,data_stage_5__1466_,
  data_stage_5__1465_,data_stage_5__1464_,data_stage_5__1463_,data_stage_5__1462_,
  data_stage_5__1461_,data_stage_5__1460_,data_stage_5__1459_,data_stage_5__1458_,
  data_stage_5__1457_,data_stage_5__1456_,data_stage_5__1455_,data_stage_5__1454_,
  data_stage_5__1453_,data_stage_5__1452_,data_stage_5__1451_,data_stage_5__1450_,
  data_stage_5__1449_,data_stage_5__1448_,data_stage_5__1447_,data_stage_5__1446_,
  data_stage_5__1445_,data_stage_5__1444_,data_stage_5__1443_,data_stage_5__1442_,
  data_stage_5__1441_,data_stage_5__1440_,data_stage_5__1439_,data_stage_5__1438_,
  data_stage_5__1437_,data_stage_5__1436_,data_stage_5__1435_,data_stage_5__1434_,
  data_stage_5__1433_,data_stage_5__1432_,data_stage_5__1431_,data_stage_5__1430_,
  data_stage_5__1429_,data_stage_5__1428_,data_stage_5__1427_,data_stage_5__1426_,
  data_stage_5__1425_,data_stage_5__1424_,data_stage_5__1423_,data_stage_5__1422_,
  data_stage_5__1421_,data_stage_5__1420_,data_stage_5__1419_,data_stage_5__1418_,
  data_stage_5__1417_,data_stage_5__1416_,data_stage_5__1415_,data_stage_5__1414_,
  data_stage_5__1413_,data_stage_5__1412_,data_stage_5__1411_,data_stage_5__1410_,
  data_stage_5__1409_,data_stage_5__1408_,data_stage_5__1407_,data_stage_5__1406_,
  data_stage_5__1405_,data_stage_5__1404_,data_stage_5__1403_,data_stage_5__1402_,
  data_stage_5__1401_,data_stage_5__1400_,data_stage_5__1399_,data_stage_5__1398_,
  data_stage_5__1397_,data_stage_5__1396_,data_stage_5__1395_,data_stage_5__1394_,
  data_stage_5__1393_,data_stage_5__1392_,data_stage_5__1391_,data_stage_5__1390_,
  data_stage_5__1389_,data_stage_5__1388_,data_stage_5__1387_,data_stage_5__1386_,
  data_stage_5__1385_,data_stage_5__1384_,data_stage_5__1383_,data_stage_5__1382_,
  data_stage_5__1381_,data_stage_5__1380_,data_stage_5__1379_,data_stage_5__1378_,
  data_stage_5__1377_,data_stage_5__1376_,data_stage_5__1375_,data_stage_5__1374_,
  data_stage_5__1373_,data_stage_5__1372_,data_stage_5__1371_,data_stage_5__1370_,
  data_stage_5__1369_,data_stage_5__1368_,data_stage_5__1367_,data_stage_5__1366_,
  data_stage_5__1365_,data_stage_5__1364_,data_stage_5__1363_,data_stage_5__1362_,
  data_stage_5__1361_,data_stage_5__1360_,data_stage_5__1359_,data_stage_5__1358_,
  data_stage_5__1357_,data_stage_5__1356_,data_stage_5__1355_,data_stage_5__1354_,
  data_stage_5__1353_,data_stage_5__1352_,data_stage_5__1351_,data_stage_5__1350_,
  data_stage_5__1349_,data_stage_5__1348_,data_stage_5__1347_,data_stage_5__1346_,
  data_stage_5__1345_,data_stage_5__1344_,data_stage_5__1343_,data_stage_5__1342_,
  data_stage_5__1341_,data_stage_5__1340_,data_stage_5__1339_,data_stage_5__1338_,
  data_stage_5__1337_,data_stage_5__1336_,data_stage_5__1335_,data_stage_5__1334_,
  data_stage_5__1333_,data_stage_5__1332_,data_stage_5__1331_,data_stage_5__1330_,
  data_stage_5__1329_,data_stage_5__1328_,data_stage_5__1327_,data_stage_5__1326_,
  data_stage_5__1325_,data_stage_5__1324_,data_stage_5__1323_,data_stage_5__1322_,
  data_stage_5__1321_,data_stage_5__1320_,data_stage_5__1319_,data_stage_5__1318_,
  data_stage_5__1317_,data_stage_5__1316_,data_stage_5__1315_,data_stage_5__1314_,
  data_stage_5__1313_,data_stage_5__1312_,data_stage_5__1311_,data_stage_5__1310_,
  data_stage_5__1309_,data_stage_5__1308_,data_stage_5__1307_,data_stage_5__1306_,
  data_stage_5__1305_,data_stage_5__1304_,data_stage_5__1303_,data_stage_5__1302_,
  data_stage_5__1301_,data_stage_5__1300_,data_stage_5__1299_,data_stage_5__1298_,
  data_stage_5__1297_,data_stage_5__1296_,data_stage_5__1295_,data_stage_5__1294_,
  data_stage_5__1293_,data_stage_5__1292_,data_stage_5__1291_,data_stage_5__1290_,
  data_stage_5__1289_,data_stage_5__1288_,data_stage_5__1287_,data_stage_5__1286_,
  data_stage_5__1285_,data_stage_5__1284_,data_stage_5__1283_,data_stage_5__1282_,
  data_stage_5__1281_,data_stage_5__1280_,data_stage_5__1279_,data_stage_5__1278_,
  data_stage_5__1277_,data_stage_5__1276_,data_stage_5__1275_,data_stage_5__1274_,
  data_stage_5__1273_,data_stage_5__1272_,data_stage_5__1271_,data_stage_5__1270_,
  data_stage_5__1269_,data_stage_5__1268_,data_stage_5__1267_,data_stage_5__1266_,
  data_stage_5__1265_,data_stage_5__1264_,data_stage_5__1263_,data_stage_5__1262_,
  data_stage_5__1261_,data_stage_5__1260_,data_stage_5__1259_,data_stage_5__1258_,
  data_stage_5__1257_,data_stage_5__1256_,data_stage_5__1255_,data_stage_5__1254_,
  data_stage_5__1253_,data_stage_5__1252_,data_stage_5__1251_,data_stage_5__1250_,
  data_stage_5__1249_,data_stage_5__1248_,data_stage_5__1247_,data_stage_5__1246_,
  data_stage_5__1245_,data_stage_5__1244_,data_stage_5__1243_,data_stage_5__1242_,
  data_stage_5__1241_,data_stage_5__1240_,data_stage_5__1239_,data_stage_5__1238_,
  data_stage_5__1237_,data_stage_5__1236_,data_stage_5__1235_,data_stage_5__1234_,
  data_stage_5__1233_,data_stage_5__1232_,data_stage_5__1231_,data_stage_5__1230_,
  data_stage_5__1229_,data_stage_5__1228_,data_stage_5__1227_,data_stage_5__1226_,
  data_stage_5__1225_,data_stage_5__1224_,data_stage_5__1223_,data_stage_5__1222_,
  data_stage_5__1221_,data_stage_5__1220_,data_stage_5__1219_,data_stage_5__1218_,
  data_stage_5__1217_,data_stage_5__1216_,data_stage_5__1215_,data_stage_5__1214_,
  data_stage_5__1213_,data_stage_5__1212_,data_stage_5__1211_,data_stage_5__1210_,
  data_stage_5__1209_,data_stage_5__1208_,data_stage_5__1207_,data_stage_5__1206_,
  data_stage_5__1205_,data_stage_5__1204_,data_stage_5__1203_,data_stage_5__1202_,
  data_stage_5__1201_,data_stage_5__1200_,data_stage_5__1199_,data_stage_5__1198_,
  data_stage_5__1197_,data_stage_5__1196_,data_stage_5__1195_,data_stage_5__1194_,
  data_stage_5__1193_,data_stage_5__1192_,data_stage_5__1191_,data_stage_5__1190_,
  data_stage_5__1189_,data_stage_5__1188_,data_stage_5__1187_,data_stage_5__1186_,
  data_stage_5__1185_,data_stage_5__1184_,data_stage_5__1183_,data_stage_5__1182_,
  data_stage_5__1181_,data_stage_5__1180_,data_stage_5__1179_,data_stage_5__1178_,
  data_stage_5__1177_,data_stage_5__1176_,data_stage_5__1175_,data_stage_5__1174_,
  data_stage_5__1173_,data_stage_5__1172_,data_stage_5__1171_,data_stage_5__1170_,
  data_stage_5__1169_,data_stage_5__1168_,data_stage_5__1167_,data_stage_5__1166_,
  data_stage_5__1165_,data_stage_5__1164_,data_stage_5__1163_,data_stage_5__1162_,
  data_stage_5__1161_,data_stage_5__1160_,data_stage_5__1159_,data_stage_5__1158_,
  data_stage_5__1157_,data_stage_5__1156_,data_stage_5__1155_,data_stage_5__1154_,
  data_stage_5__1153_,data_stage_5__1152_,data_stage_5__1151_,data_stage_5__1150_,
  data_stage_5__1149_,data_stage_5__1148_,data_stage_5__1147_,data_stage_5__1146_,
  data_stage_5__1145_,data_stage_5__1144_,data_stage_5__1143_,data_stage_5__1142_,
  data_stage_5__1141_,data_stage_5__1140_,data_stage_5__1139_,data_stage_5__1138_,
  data_stage_5__1137_,data_stage_5__1136_,data_stage_5__1135_,data_stage_5__1134_,
  data_stage_5__1133_,data_stage_5__1132_,data_stage_5__1131_,data_stage_5__1130_,
  data_stage_5__1129_,data_stage_5__1128_,data_stage_5__1127_,data_stage_5__1126_,
  data_stage_5__1125_,data_stage_5__1124_,data_stage_5__1123_,data_stage_5__1122_,
  data_stage_5__1121_,data_stage_5__1120_,data_stage_5__1119_,data_stage_5__1118_,
  data_stage_5__1117_,data_stage_5__1116_,data_stage_5__1115_,data_stage_5__1114_,
  data_stage_5__1113_,data_stage_5__1112_,data_stage_5__1111_,data_stage_5__1110_,
  data_stage_5__1109_,data_stage_5__1108_,data_stage_5__1107_,data_stage_5__1106_,
  data_stage_5__1105_,data_stage_5__1104_,data_stage_5__1103_,data_stage_5__1102_,
  data_stage_5__1101_,data_stage_5__1100_,data_stage_5__1099_,data_stage_5__1098_,
  data_stage_5__1097_,data_stage_5__1096_,data_stage_5__1095_,data_stage_5__1094_,
  data_stage_5__1093_,data_stage_5__1092_,data_stage_5__1091_,data_stage_5__1090_,
  data_stage_5__1089_,data_stage_5__1088_,data_stage_5__1087_,data_stage_5__1086_,
  data_stage_5__1085_,data_stage_5__1084_,data_stage_5__1083_,data_stage_5__1082_,
  data_stage_5__1081_,data_stage_5__1080_,data_stage_5__1079_,data_stage_5__1078_,
  data_stage_5__1077_,data_stage_5__1076_,data_stage_5__1075_,data_stage_5__1074_,
  data_stage_5__1073_,data_stage_5__1072_,data_stage_5__1071_,data_stage_5__1070_,
  data_stage_5__1069_,data_stage_5__1068_,data_stage_5__1067_,data_stage_5__1066_,
  data_stage_5__1065_,data_stage_5__1064_,data_stage_5__1063_,data_stage_5__1062_,
  data_stage_5__1061_,data_stage_5__1060_,data_stage_5__1059_,data_stage_5__1058_,
  data_stage_5__1057_,data_stage_5__1056_,data_stage_5__1055_,data_stage_5__1054_,
  data_stage_5__1053_,data_stage_5__1052_,data_stage_5__1051_,data_stage_5__1050_,
  data_stage_5__1049_,data_stage_5__1048_,data_stage_5__1047_,data_stage_5__1046_,
  data_stage_5__1045_,data_stage_5__1044_,data_stage_5__1043_,data_stage_5__1042_,
  data_stage_5__1041_,data_stage_5__1040_,data_stage_5__1039_,data_stage_5__1038_,
  data_stage_5__1037_,data_stage_5__1036_,data_stage_5__1035_,data_stage_5__1034_,
  data_stage_5__1033_,data_stage_5__1032_,data_stage_5__1031_,data_stage_5__1030_,
  data_stage_5__1029_,data_stage_5__1028_,data_stage_5__1027_,data_stage_5__1026_,
  data_stage_5__1025_,data_stage_5__1024_,data_stage_5__1023_,data_stage_5__1022_,
  data_stage_5__1021_,data_stage_5__1020_,data_stage_5__1019_,data_stage_5__1018_,
  data_stage_5__1017_,data_stage_5__1016_,data_stage_5__1015_,data_stage_5__1014_,
  data_stage_5__1013_,data_stage_5__1012_,data_stage_5__1011_,data_stage_5__1010_,
  data_stage_5__1009_,data_stage_5__1008_,data_stage_5__1007_,data_stage_5__1006_,
  data_stage_5__1005_,data_stage_5__1004_,data_stage_5__1003_,data_stage_5__1002_,
  data_stage_5__1001_,data_stage_5__1000_,data_stage_5__999_,data_stage_5__998_,
  data_stage_5__997_,data_stage_5__996_,data_stage_5__995_,data_stage_5__994_,
  data_stage_5__993_,data_stage_5__992_,data_stage_5__991_,data_stage_5__990_,
  data_stage_5__989_,data_stage_5__988_,data_stage_5__987_,data_stage_5__986_,
  data_stage_5__985_,data_stage_5__984_,data_stage_5__983_,data_stage_5__982_,
  data_stage_5__981_,data_stage_5__980_,data_stage_5__979_,data_stage_5__978_,data_stage_5__977_,
  data_stage_5__976_,data_stage_5__975_,data_stage_5__974_,data_stage_5__973_,
  data_stage_5__972_,data_stage_5__971_,data_stage_5__970_,data_stage_5__969_,
  data_stage_5__968_,data_stage_5__967_,data_stage_5__966_,data_stage_5__965_,
  data_stage_5__964_,data_stage_5__963_,data_stage_5__962_,data_stage_5__961_,data_stage_5__960_,
  data_stage_5__959_,data_stage_5__958_,data_stage_5__957_,data_stage_5__956_,
  data_stage_5__955_,data_stage_5__954_,data_stage_5__953_,data_stage_5__952_,
  data_stage_5__951_,data_stage_5__950_,data_stage_5__949_,data_stage_5__948_,
  data_stage_5__947_,data_stage_5__946_,data_stage_5__945_,data_stage_5__944_,
  data_stage_5__943_,data_stage_5__942_,data_stage_5__941_,data_stage_5__940_,data_stage_5__939_,
  data_stage_5__938_,data_stage_5__937_,data_stage_5__936_,data_stage_5__935_,
  data_stage_5__934_,data_stage_5__933_,data_stage_5__932_,data_stage_5__931_,
  data_stage_5__930_,data_stage_5__929_,data_stage_5__928_,data_stage_5__927_,
  data_stage_5__926_,data_stage_5__925_,data_stage_5__924_,data_stage_5__923_,
  data_stage_5__922_,data_stage_5__921_,data_stage_5__920_,data_stage_5__919_,data_stage_5__918_,
  data_stage_5__917_,data_stage_5__916_,data_stage_5__915_,data_stage_5__914_,
  data_stage_5__913_,data_stage_5__912_,data_stage_5__911_,data_stage_5__910_,
  data_stage_5__909_,data_stage_5__908_,data_stage_5__907_,data_stage_5__906_,
  data_stage_5__905_,data_stage_5__904_,data_stage_5__903_,data_stage_5__902_,
  data_stage_5__901_,data_stage_5__900_,data_stage_5__899_,data_stage_5__898_,data_stage_5__897_,
  data_stage_5__896_,data_stage_5__895_,data_stage_5__894_,data_stage_5__893_,
  data_stage_5__892_,data_stage_5__891_,data_stage_5__890_,data_stage_5__889_,
  data_stage_5__888_,data_stage_5__887_,data_stage_5__886_,data_stage_5__885_,
  data_stage_5__884_,data_stage_5__883_,data_stage_5__882_,data_stage_5__881_,data_stage_5__880_,
  data_stage_5__879_,data_stage_5__878_,data_stage_5__877_,data_stage_5__876_,
  data_stage_5__875_,data_stage_5__874_,data_stage_5__873_,data_stage_5__872_,
  data_stage_5__871_,data_stage_5__870_,data_stage_5__869_,data_stage_5__868_,
  data_stage_5__867_,data_stage_5__866_,data_stage_5__865_,data_stage_5__864_,
  data_stage_5__863_,data_stage_5__862_,data_stage_5__861_,data_stage_5__860_,data_stage_5__859_,
  data_stage_5__858_,data_stage_5__857_,data_stage_5__856_,data_stage_5__855_,
  data_stage_5__854_,data_stage_5__853_,data_stage_5__852_,data_stage_5__851_,
  data_stage_5__850_,data_stage_5__849_,data_stage_5__848_,data_stage_5__847_,
  data_stage_5__846_,data_stage_5__845_,data_stage_5__844_,data_stage_5__843_,
  data_stage_5__842_,data_stage_5__841_,data_stage_5__840_,data_stage_5__839_,data_stage_5__838_,
  data_stage_5__837_,data_stage_5__836_,data_stage_5__835_,data_stage_5__834_,
  data_stage_5__833_,data_stage_5__832_,data_stage_5__831_,data_stage_5__830_,
  data_stage_5__829_,data_stage_5__828_,data_stage_5__827_,data_stage_5__826_,
  data_stage_5__825_,data_stage_5__824_,data_stage_5__823_,data_stage_5__822_,
  data_stage_5__821_,data_stage_5__820_,data_stage_5__819_,data_stage_5__818_,data_stage_5__817_,
  data_stage_5__816_,data_stage_5__815_,data_stage_5__814_,data_stage_5__813_,
  data_stage_5__812_,data_stage_5__811_,data_stage_5__810_,data_stage_5__809_,
  data_stage_5__808_,data_stage_5__807_,data_stage_5__806_,data_stage_5__805_,
  data_stage_5__804_,data_stage_5__803_,data_stage_5__802_,data_stage_5__801_,data_stage_5__800_,
  data_stage_5__799_,data_stage_5__798_,data_stage_5__797_,data_stage_5__796_,
  data_stage_5__795_,data_stage_5__794_,data_stage_5__793_,data_stage_5__792_,
  data_stage_5__791_,data_stage_5__790_,data_stage_5__789_,data_stage_5__788_,
  data_stage_5__787_,data_stage_5__786_,data_stage_5__785_,data_stage_5__784_,
  data_stage_5__783_,data_stage_5__782_,data_stage_5__781_,data_stage_5__780_,data_stage_5__779_,
  data_stage_5__778_,data_stage_5__777_,data_stage_5__776_,data_stage_5__775_,
  data_stage_5__774_,data_stage_5__773_,data_stage_5__772_,data_stage_5__771_,
  data_stage_5__770_,data_stage_5__769_,data_stage_5__768_,data_stage_5__767_,
  data_stage_5__766_,data_stage_5__765_,data_stage_5__764_,data_stage_5__763_,
  data_stage_5__762_,data_stage_5__761_,data_stage_5__760_,data_stage_5__759_,data_stage_5__758_,
  data_stage_5__757_,data_stage_5__756_,data_stage_5__755_,data_stage_5__754_,
  data_stage_5__753_,data_stage_5__752_,data_stage_5__751_,data_stage_5__750_,
  data_stage_5__749_,data_stage_5__748_,data_stage_5__747_,data_stage_5__746_,
  data_stage_5__745_,data_stage_5__744_,data_stage_5__743_,data_stage_5__742_,
  data_stage_5__741_,data_stage_5__740_,data_stage_5__739_,data_stage_5__738_,data_stage_5__737_,
  data_stage_5__736_,data_stage_5__735_,data_stage_5__734_,data_stage_5__733_,
  data_stage_5__732_,data_stage_5__731_,data_stage_5__730_,data_stage_5__729_,
  data_stage_5__728_,data_stage_5__727_,data_stage_5__726_,data_stage_5__725_,
  data_stage_5__724_,data_stage_5__723_,data_stage_5__722_,data_stage_5__721_,data_stage_5__720_,
  data_stage_5__719_,data_stage_5__718_,data_stage_5__717_,data_stage_5__716_,
  data_stage_5__715_,data_stage_5__714_,data_stage_5__713_,data_stage_5__712_,
  data_stage_5__711_,data_stage_5__710_,data_stage_5__709_,data_stage_5__708_,
  data_stage_5__707_,data_stage_5__706_,data_stage_5__705_,data_stage_5__704_,
  data_stage_5__703_,data_stage_5__702_,data_stage_5__701_,data_stage_5__700_,data_stage_5__699_,
  data_stage_5__698_,data_stage_5__697_,data_stage_5__696_,data_stage_5__695_,
  data_stage_5__694_,data_stage_5__693_,data_stage_5__692_,data_stage_5__691_,
  data_stage_5__690_,data_stage_5__689_,data_stage_5__688_,data_stage_5__687_,
  data_stage_5__686_,data_stage_5__685_,data_stage_5__684_,data_stage_5__683_,
  data_stage_5__682_,data_stage_5__681_,data_stage_5__680_,data_stage_5__679_,data_stage_5__678_,
  data_stage_5__677_,data_stage_5__676_,data_stage_5__675_,data_stage_5__674_,
  data_stage_5__673_,data_stage_5__672_,data_stage_5__671_,data_stage_5__670_,
  data_stage_5__669_,data_stage_5__668_,data_stage_5__667_,data_stage_5__666_,
  data_stage_5__665_,data_stage_5__664_,data_stage_5__663_,data_stage_5__662_,
  data_stage_5__661_,data_stage_5__660_,data_stage_5__659_,data_stage_5__658_,data_stage_5__657_,
  data_stage_5__656_,data_stage_5__655_,data_stage_5__654_,data_stage_5__653_,
  data_stage_5__652_,data_stage_5__651_,data_stage_5__650_,data_stage_5__649_,
  data_stage_5__648_,data_stage_5__647_,data_stage_5__646_,data_stage_5__645_,
  data_stage_5__644_,data_stage_5__643_,data_stage_5__642_,data_stage_5__641_,data_stage_5__640_,
  data_stage_5__639_,data_stage_5__638_,data_stage_5__637_,data_stage_5__636_,
  data_stage_5__635_,data_stage_5__634_,data_stage_5__633_,data_stage_5__632_,
  data_stage_5__631_,data_stage_5__630_,data_stage_5__629_,data_stage_5__628_,
  data_stage_5__627_,data_stage_5__626_,data_stage_5__625_,data_stage_5__624_,
  data_stage_5__623_,data_stage_5__622_,data_stage_5__621_,data_stage_5__620_,data_stage_5__619_,
  data_stage_5__618_,data_stage_5__617_,data_stage_5__616_,data_stage_5__615_,
  data_stage_5__614_,data_stage_5__613_,data_stage_5__612_,data_stage_5__611_,
  data_stage_5__610_,data_stage_5__609_,data_stage_5__608_,data_stage_5__607_,
  data_stage_5__606_,data_stage_5__605_,data_stage_5__604_,data_stage_5__603_,
  data_stage_5__602_,data_stage_5__601_,data_stage_5__600_,data_stage_5__599_,data_stage_5__598_,
  data_stage_5__597_,data_stage_5__596_,data_stage_5__595_,data_stage_5__594_,
  data_stage_5__593_,data_stage_5__592_,data_stage_5__591_,data_stage_5__590_,
  data_stage_5__589_,data_stage_5__588_,data_stage_5__587_,data_stage_5__586_,
  data_stage_5__585_,data_stage_5__584_,data_stage_5__583_,data_stage_5__582_,
  data_stage_5__581_,data_stage_5__580_,data_stage_5__579_,data_stage_5__578_,data_stage_5__577_,
  data_stage_5__576_,data_stage_5__575_,data_stage_5__574_,data_stage_5__573_,
  data_stage_5__572_,data_stage_5__571_,data_stage_5__570_,data_stage_5__569_,
  data_stage_5__568_,data_stage_5__567_,data_stage_5__566_,data_stage_5__565_,
  data_stage_5__564_,data_stage_5__563_,data_stage_5__562_,data_stage_5__561_,data_stage_5__560_,
  data_stage_5__559_,data_stage_5__558_,data_stage_5__557_,data_stage_5__556_,
  data_stage_5__555_,data_stage_5__554_,data_stage_5__553_,data_stage_5__552_,
  data_stage_5__551_,data_stage_5__550_,data_stage_5__549_,data_stage_5__548_,
  data_stage_5__547_,data_stage_5__546_,data_stage_5__545_,data_stage_5__544_,
  data_stage_5__543_,data_stage_5__542_,data_stage_5__541_,data_stage_5__540_,data_stage_5__539_,
  data_stage_5__538_,data_stage_5__537_,data_stage_5__536_,data_stage_5__535_,
  data_stage_5__534_,data_stage_5__533_,data_stage_5__532_,data_stage_5__531_,
  data_stage_5__530_,data_stage_5__529_,data_stage_5__528_,data_stage_5__527_,
  data_stage_5__526_,data_stage_5__525_,data_stage_5__524_,data_stage_5__523_,
  data_stage_5__522_,data_stage_5__521_,data_stage_5__520_,data_stage_5__519_,data_stage_5__518_,
  data_stage_5__517_,data_stage_5__516_,data_stage_5__515_,data_stage_5__514_,
  data_stage_5__513_,data_stage_5__512_,data_stage_5__511_,data_stage_5__510_,
  data_stage_5__509_,data_stage_5__508_,data_stage_5__507_,data_stage_5__506_,
  data_stage_5__505_,data_stage_5__504_,data_stage_5__503_,data_stage_5__502_,
  data_stage_5__501_,data_stage_5__500_,data_stage_5__499_,data_stage_5__498_,data_stage_5__497_,
  data_stage_5__496_,data_stage_5__495_,data_stage_5__494_,data_stage_5__493_,
  data_stage_5__492_,data_stage_5__491_,data_stage_5__490_,data_stage_5__489_,
  data_stage_5__488_,data_stage_5__487_,data_stage_5__486_,data_stage_5__485_,
  data_stage_5__484_,data_stage_5__483_,data_stage_5__482_,data_stage_5__481_,data_stage_5__480_,
  data_stage_5__479_,data_stage_5__478_,data_stage_5__477_,data_stage_5__476_,
  data_stage_5__475_,data_stage_5__474_,data_stage_5__473_,data_stage_5__472_,
  data_stage_5__471_,data_stage_5__470_,data_stage_5__469_,data_stage_5__468_,
  data_stage_5__467_,data_stage_5__466_,data_stage_5__465_,data_stage_5__464_,
  data_stage_5__463_,data_stage_5__462_,data_stage_5__461_,data_stage_5__460_,data_stage_5__459_,
  data_stage_5__458_,data_stage_5__457_,data_stage_5__456_,data_stage_5__455_,
  data_stage_5__454_,data_stage_5__453_,data_stage_5__452_,data_stage_5__451_,
  data_stage_5__450_,data_stage_5__449_,data_stage_5__448_,data_stage_5__447_,
  data_stage_5__446_,data_stage_5__445_,data_stage_5__444_,data_stage_5__443_,
  data_stage_5__442_,data_stage_5__441_,data_stage_5__440_,data_stage_5__439_,data_stage_5__438_,
  data_stage_5__437_,data_stage_5__436_,data_stage_5__435_,data_stage_5__434_,
  data_stage_5__433_,data_stage_5__432_,data_stage_5__431_,data_stage_5__430_,
  data_stage_5__429_,data_stage_5__428_,data_stage_5__427_,data_stage_5__426_,
  data_stage_5__425_,data_stage_5__424_,data_stage_5__423_,data_stage_5__422_,
  data_stage_5__421_,data_stage_5__420_,data_stage_5__419_,data_stage_5__418_,data_stage_5__417_,
  data_stage_5__416_,data_stage_5__415_,data_stage_5__414_,data_stage_5__413_,
  data_stage_5__412_,data_stage_5__411_,data_stage_5__410_,data_stage_5__409_,
  data_stage_5__408_,data_stage_5__407_,data_stage_5__406_,data_stage_5__405_,
  data_stage_5__404_,data_stage_5__403_,data_stage_5__402_,data_stage_5__401_,data_stage_5__400_,
  data_stage_5__399_,data_stage_5__398_,data_stage_5__397_,data_stage_5__396_,
  data_stage_5__395_,data_stage_5__394_,data_stage_5__393_,data_stage_5__392_,
  data_stage_5__391_,data_stage_5__390_,data_stage_5__389_,data_stage_5__388_,
  data_stage_5__387_,data_stage_5__386_,data_stage_5__385_,data_stage_5__384_,
  data_stage_5__383_,data_stage_5__382_,data_stage_5__381_,data_stage_5__380_,data_stage_5__379_,
  data_stage_5__378_,data_stage_5__377_,data_stage_5__376_,data_stage_5__375_,
  data_stage_5__374_,data_stage_5__373_,data_stage_5__372_,data_stage_5__371_,
  data_stage_5__370_,data_stage_5__369_,data_stage_5__368_,data_stage_5__367_,
  data_stage_5__366_,data_stage_5__365_,data_stage_5__364_,data_stage_5__363_,
  data_stage_5__362_,data_stage_5__361_,data_stage_5__360_,data_stage_5__359_,data_stage_5__358_,
  data_stage_5__357_,data_stage_5__356_,data_stage_5__355_,data_stage_5__354_,
  data_stage_5__353_,data_stage_5__352_,data_stage_5__351_,data_stage_5__350_,
  data_stage_5__349_,data_stage_5__348_,data_stage_5__347_,data_stage_5__346_,
  data_stage_5__345_,data_stage_5__344_,data_stage_5__343_,data_stage_5__342_,
  data_stage_5__341_,data_stage_5__340_,data_stage_5__339_,data_stage_5__338_,data_stage_5__337_,
  data_stage_5__336_,data_stage_5__335_,data_stage_5__334_,data_stage_5__333_,
  data_stage_5__332_,data_stage_5__331_,data_stage_5__330_,data_stage_5__329_,
  data_stage_5__328_,data_stage_5__327_,data_stage_5__326_,data_stage_5__325_,
  data_stage_5__324_,data_stage_5__323_,data_stage_5__322_,data_stage_5__321_,data_stage_5__320_,
  data_stage_5__319_,data_stage_5__318_,data_stage_5__317_,data_stage_5__316_,
  data_stage_5__315_,data_stage_5__314_,data_stage_5__313_,data_stage_5__312_,
  data_stage_5__311_,data_stage_5__310_,data_stage_5__309_,data_stage_5__308_,
  data_stage_5__307_,data_stage_5__306_,data_stage_5__305_,data_stage_5__304_,
  data_stage_5__303_,data_stage_5__302_,data_stage_5__301_,data_stage_5__300_,data_stage_5__299_,
  data_stage_5__298_,data_stage_5__297_,data_stage_5__296_,data_stage_5__295_,
  data_stage_5__294_,data_stage_5__293_,data_stage_5__292_,data_stage_5__291_,
  data_stage_5__290_,data_stage_5__289_,data_stage_5__288_,data_stage_5__287_,
  data_stage_5__286_,data_stage_5__285_,data_stage_5__284_,data_stage_5__283_,
  data_stage_5__282_,data_stage_5__281_,data_stage_5__280_,data_stage_5__279_,data_stage_5__278_,
  data_stage_5__277_,data_stage_5__276_,data_stage_5__275_,data_stage_5__274_,
  data_stage_5__273_,data_stage_5__272_,data_stage_5__271_,data_stage_5__270_,
  data_stage_5__269_,data_stage_5__268_,data_stage_5__267_,data_stage_5__266_,
  data_stage_5__265_,data_stage_5__264_,data_stage_5__263_,data_stage_5__262_,
  data_stage_5__261_,data_stage_5__260_,data_stage_5__259_,data_stage_5__258_,data_stage_5__257_,
  data_stage_5__256_,data_stage_5__255_,data_stage_5__254_,data_stage_5__253_,
  data_stage_5__252_,data_stage_5__251_,data_stage_5__250_,data_stage_5__249_,
  data_stage_5__248_,data_stage_5__247_,data_stage_5__246_,data_stage_5__245_,
  data_stage_5__244_,data_stage_5__243_,data_stage_5__242_,data_stage_5__241_,data_stage_5__240_,
  data_stage_5__239_,data_stage_5__238_,data_stage_5__237_,data_stage_5__236_,
  data_stage_5__235_,data_stage_5__234_,data_stage_5__233_,data_stage_5__232_,
  data_stage_5__231_,data_stage_5__230_,data_stage_5__229_,data_stage_5__228_,
  data_stage_5__227_,data_stage_5__226_,data_stage_5__225_,data_stage_5__224_,
  data_stage_5__223_,data_stage_5__222_,data_stage_5__221_,data_stage_5__220_,data_stage_5__219_,
  data_stage_5__218_,data_stage_5__217_,data_stage_5__216_,data_stage_5__215_,
  data_stage_5__214_,data_stage_5__213_,data_stage_5__212_,data_stage_5__211_,
  data_stage_5__210_,data_stage_5__209_,data_stage_5__208_,data_stage_5__207_,
  data_stage_5__206_,data_stage_5__205_,data_stage_5__204_,data_stage_5__203_,
  data_stage_5__202_,data_stage_5__201_,data_stage_5__200_,data_stage_5__199_,data_stage_5__198_,
  data_stage_5__197_,data_stage_5__196_,data_stage_5__195_,data_stage_5__194_,
  data_stage_5__193_,data_stage_5__192_,data_stage_5__191_,data_stage_5__190_,
  data_stage_5__189_,data_stage_5__188_,data_stage_5__187_,data_stage_5__186_,
  data_stage_5__185_,data_stage_5__184_,data_stage_5__183_,data_stage_5__182_,
  data_stage_5__181_,data_stage_5__180_,data_stage_5__179_,data_stage_5__178_,data_stage_5__177_,
  data_stage_5__176_,data_stage_5__175_,data_stage_5__174_,data_stage_5__173_,
  data_stage_5__172_,data_stage_5__171_,data_stage_5__170_,data_stage_5__169_,
  data_stage_5__168_,data_stage_5__167_,data_stage_5__166_,data_stage_5__165_,
  data_stage_5__164_,data_stage_5__163_,data_stage_5__162_,data_stage_5__161_,data_stage_5__160_,
  data_stage_5__159_,data_stage_5__158_,data_stage_5__157_,data_stage_5__156_,
  data_stage_5__155_,data_stage_5__154_,data_stage_5__153_,data_stage_5__152_,
  data_stage_5__151_,data_stage_5__150_,data_stage_5__149_,data_stage_5__148_,
  data_stage_5__147_,data_stage_5__146_,data_stage_5__145_,data_stage_5__144_,
  data_stage_5__143_,data_stage_5__142_,data_stage_5__141_,data_stage_5__140_,data_stage_5__139_,
  data_stage_5__138_,data_stage_5__137_,data_stage_5__136_,data_stage_5__135_,
  data_stage_5__134_,data_stage_5__133_,data_stage_5__132_,data_stage_5__131_,
  data_stage_5__130_,data_stage_5__129_,data_stage_5__128_,data_stage_5__127_,
  data_stage_5__126_,data_stage_5__125_,data_stage_5__124_,data_stage_5__123_,
  data_stage_5__122_,data_stage_5__121_,data_stage_5__120_,data_stage_5__119_,data_stage_5__118_,
  data_stage_5__117_,data_stage_5__116_,data_stage_5__115_,data_stage_5__114_,
  data_stage_5__113_,data_stage_5__112_,data_stage_5__111_,data_stage_5__110_,
  data_stage_5__109_,data_stage_5__108_,data_stage_5__107_,data_stage_5__106_,
  data_stage_5__105_,data_stage_5__104_,data_stage_5__103_,data_stage_5__102_,
  data_stage_5__101_,data_stage_5__100_,data_stage_5__99_,data_stage_5__98_,data_stage_5__97_,
  data_stage_5__96_,data_stage_5__95_,data_stage_5__94_,data_stage_5__93_,
  data_stage_5__92_,data_stage_5__91_,data_stage_5__90_,data_stage_5__89_,data_stage_5__88_,
  data_stage_5__87_,data_stage_5__86_,data_stage_5__85_,data_stage_5__84_,
  data_stage_5__83_,data_stage_5__82_,data_stage_5__81_,data_stage_5__80_,data_stage_5__79_,
  data_stage_5__78_,data_stage_5__77_,data_stage_5__76_,data_stage_5__75_,
  data_stage_5__74_,data_stage_5__73_,data_stage_5__72_,data_stage_5__71_,data_stage_5__70_,
  data_stage_5__69_,data_stage_5__68_,data_stage_5__67_,data_stage_5__66_,
  data_stage_5__65_,data_stage_5__64_,data_stage_5__63_,data_stage_5__62_,
  data_stage_5__61_,data_stage_5__60_,data_stage_5__59_,data_stage_5__58_,data_stage_5__57_,
  data_stage_5__56_,data_stage_5__55_,data_stage_5__54_,data_stage_5__53_,
  data_stage_5__52_,data_stage_5__51_,data_stage_5__50_,data_stage_5__49_,data_stage_5__48_,
  data_stage_5__47_,data_stage_5__46_,data_stage_5__45_,data_stage_5__44_,
  data_stage_5__43_,data_stage_5__42_,data_stage_5__41_,data_stage_5__40_,data_stage_5__39_,
  data_stage_5__38_,data_stage_5__37_,data_stage_5__36_,data_stage_5__35_,
  data_stage_5__34_,data_stage_5__33_,data_stage_5__32_,data_stage_5__31_,data_stage_5__30_,
  data_stage_5__29_,data_stage_5__28_,data_stage_5__27_,data_stage_5__26_,
  data_stage_5__25_,data_stage_5__24_,data_stage_5__23_,data_stage_5__22_,
  data_stage_5__21_,data_stage_5__20_,data_stage_5__19_,data_stage_5__18_,data_stage_5__17_,
  data_stage_5__16_,data_stage_5__15_,data_stage_5__14_,data_stage_5__13_,
  data_stage_5__12_,data_stage_5__11_,data_stage_5__10_,data_stage_5__9_,data_stage_5__8_,
  data_stage_5__7_,data_stage_5__6_,data_stage_5__5_,data_stage_5__4_,data_stage_5__3_,
  data_stage_5__2_,data_stage_5__1_,data_stage_5__0_;

  bsg_swap_width_p64
  mux_stage_0__mux_swap_0__swap_inst
  (
    .data_i(data_i[127:0]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__127_, data_stage_1__126_, data_stage_1__125_, data_stage_1__124_, data_stage_1__123_, data_stage_1__122_, data_stage_1__121_, data_stage_1__120_, data_stage_1__119_, data_stage_1__118_, data_stage_1__117_, data_stage_1__116_, data_stage_1__115_, data_stage_1__114_, data_stage_1__113_, data_stage_1__112_, data_stage_1__111_, data_stage_1__110_, data_stage_1__109_, data_stage_1__108_, data_stage_1__107_, data_stage_1__106_, data_stage_1__105_, data_stage_1__104_, data_stage_1__103_, data_stage_1__102_, data_stage_1__101_, data_stage_1__100_, data_stage_1__99_, data_stage_1__98_, data_stage_1__97_, data_stage_1__96_, data_stage_1__95_, data_stage_1__94_, data_stage_1__93_, data_stage_1__92_, data_stage_1__91_, data_stage_1__90_, data_stage_1__89_, data_stage_1__88_, data_stage_1__87_, data_stage_1__86_, data_stage_1__85_, data_stage_1__84_, data_stage_1__83_, data_stage_1__82_, data_stage_1__81_, data_stage_1__80_, data_stage_1__79_, data_stage_1__78_, data_stage_1__77_, data_stage_1__76_, data_stage_1__75_, data_stage_1__74_, data_stage_1__73_, data_stage_1__72_, data_stage_1__71_, data_stage_1__70_, data_stage_1__69_, data_stage_1__68_, data_stage_1__67_, data_stage_1__66_, data_stage_1__65_, data_stage_1__64_, data_stage_1__63_, data_stage_1__62_, data_stage_1__61_, data_stage_1__60_, data_stage_1__59_, data_stage_1__58_, data_stage_1__57_, data_stage_1__56_, data_stage_1__55_, data_stage_1__54_, data_stage_1__53_, data_stage_1__52_, data_stage_1__51_, data_stage_1__50_, data_stage_1__49_, data_stage_1__48_, data_stage_1__47_, data_stage_1__46_, data_stage_1__45_, data_stage_1__44_, data_stage_1__43_, data_stage_1__42_, data_stage_1__41_, data_stage_1__40_, data_stage_1__39_, data_stage_1__38_, data_stage_1__37_, data_stage_1__36_, data_stage_1__35_, data_stage_1__34_, data_stage_1__33_, data_stage_1__32_, data_stage_1__31_, data_stage_1__30_, data_stage_1__29_, data_stage_1__28_, data_stage_1__27_, data_stage_1__26_, data_stage_1__25_, data_stage_1__24_, data_stage_1__23_, data_stage_1__22_, data_stage_1__21_, data_stage_1__20_, data_stage_1__19_, data_stage_1__18_, data_stage_1__17_, data_stage_1__16_, data_stage_1__15_, data_stage_1__14_, data_stage_1__13_, data_stage_1__12_, data_stage_1__11_, data_stage_1__10_, data_stage_1__9_, data_stage_1__8_, data_stage_1__7_, data_stage_1__6_, data_stage_1__5_, data_stage_1__4_, data_stage_1__3_, data_stage_1__2_, data_stage_1__1_, data_stage_1__0_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_1__swap_inst
  (
    .data_i(data_i[255:128]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__255_, data_stage_1__254_, data_stage_1__253_, data_stage_1__252_, data_stage_1__251_, data_stage_1__250_, data_stage_1__249_, data_stage_1__248_, data_stage_1__247_, data_stage_1__246_, data_stage_1__245_, data_stage_1__244_, data_stage_1__243_, data_stage_1__242_, data_stage_1__241_, data_stage_1__240_, data_stage_1__239_, data_stage_1__238_, data_stage_1__237_, data_stage_1__236_, data_stage_1__235_, data_stage_1__234_, data_stage_1__233_, data_stage_1__232_, data_stage_1__231_, data_stage_1__230_, data_stage_1__229_, data_stage_1__228_, data_stage_1__227_, data_stage_1__226_, data_stage_1__225_, data_stage_1__224_, data_stage_1__223_, data_stage_1__222_, data_stage_1__221_, data_stage_1__220_, data_stage_1__219_, data_stage_1__218_, data_stage_1__217_, data_stage_1__216_, data_stage_1__215_, data_stage_1__214_, data_stage_1__213_, data_stage_1__212_, data_stage_1__211_, data_stage_1__210_, data_stage_1__209_, data_stage_1__208_, data_stage_1__207_, data_stage_1__206_, data_stage_1__205_, data_stage_1__204_, data_stage_1__203_, data_stage_1__202_, data_stage_1__201_, data_stage_1__200_, data_stage_1__199_, data_stage_1__198_, data_stage_1__197_, data_stage_1__196_, data_stage_1__195_, data_stage_1__194_, data_stage_1__193_, data_stage_1__192_, data_stage_1__191_, data_stage_1__190_, data_stage_1__189_, data_stage_1__188_, data_stage_1__187_, data_stage_1__186_, data_stage_1__185_, data_stage_1__184_, data_stage_1__183_, data_stage_1__182_, data_stage_1__181_, data_stage_1__180_, data_stage_1__179_, data_stage_1__178_, data_stage_1__177_, data_stage_1__176_, data_stage_1__175_, data_stage_1__174_, data_stage_1__173_, data_stage_1__172_, data_stage_1__171_, data_stage_1__170_, data_stage_1__169_, data_stage_1__168_, data_stage_1__167_, data_stage_1__166_, data_stage_1__165_, data_stage_1__164_, data_stage_1__163_, data_stage_1__162_, data_stage_1__161_, data_stage_1__160_, data_stage_1__159_, data_stage_1__158_, data_stage_1__157_, data_stage_1__156_, data_stage_1__155_, data_stage_1__154_, data_stage_1__153_, data_stage_1__152_, data_stage_1__151_, data_stage_1__150_, data_stage_1__149_, data_stage_1__148_, data_stage_1__147_, data_stage_1__146_, data_stage_1__145_, data_stage_1__144_, data_stage_1__143_, data_stage_1__142_, data_stage_1__141_, data_stage_1__140_, data_stage_1__139_, data_stage_1__138_, data_stage_1__137_, data_stage_1__136_, data_stage_1__135_, data_stage_1__134_, data_stage_1__133_, data_stage_1__132_, data_stage_1__131_, data_stage_1__130_, data_stage_1__129_, data_stage_1__128_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_2__swap_inst
  (
    .data_i(data_i[383:256]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__383_, data_stage_1__382_, data_stage_1__381_, data_stage_1__380_, data_stage_1__379_, data_stage_1__378_, data_stage_1__377_, data_stage_1__376_, data_stage_1__375_, data_stage_1__374_, data_stage_1__373_, data_stage_1__372_, data_stage_1__371_, data_stage_1__370_, data_stage_1__369_, data_stage_1__368_, data_stage_1__367_, data_stage_1__366_, data_stage_1__365_, data_stage_1__364_, data_stage_1__363_, data_stage_1__362_, data_stage_1__361_, data_stage_1__360_, data_stage_1__359_, data_stage_1__358_, data_stage_1__357_, data_stage_1__356_, data_stage_1__355_, data_stage_1__354_, data_stage_1__353_, data_stage_1__352_, data_stage_1__351_, data_stage_1__350_, data_stage_1__349_, data_stage_1__348_, data_stage_1__347_, data_stage_1__346_, data_stage_1__345_, data_stage_1__344_, data_stage_1__343_, data_stage_1__342_, data_stage_1__341_, data_stage_1__340_, data_stage_1__339_, data_stage_1__338_, data_stage_1__337_, data_stage_1__336_, data_stage_1__335_, data_stage_1__334_, data_stage_1__333_, data_stage_1__332_, data_stage_1__331_, data_stage_1__330_, data_stage_1__329_, data_stage_1__328_, data_stage_1__327_, data_stage_1__326_, data_stage_1__325_, data_stage_1__324_, data_stage_1__323_, data_stage_1__322_, data_stage_1__321_, data_stage_1__320_, data_stage_1__319_, data_stage_1__318_, data_stage_1__317_, data_stage_1__316_, data_stage_1__315_, data_stage_1__314_, data_stage_1__313_, data_stage_1__312_, data_stage_1__311_, data_stage_1__310_, data_stage_1__309_, data_stage_1__308_, data_stage_1__307_, data_stage_1__306_, data_stage_1__305_, data_stage_1__304_, data_stage_1__303_, data_stage_1__302_, data_stage_1__301_, data_stage_1__300_, data_stage_1__299_, data_stage_1__298_, data_stage_1__297_, data_stage_1__296_, data_stage_1__295_, data_stage_1__294_, data_stage_1__293_, data_stage_1__292_, data_stage_1__291_, data_stage_1__290_, data_stage_1__289_, data_stage_1__288_, data_stage_1__287_, data_stage_1__286_, data_stage_1__285_, data_stage_1__284_, data_stage_1__283_, data_stage_1__282_, data_stage_1__281_, data_stage_1__280_, data_stage_1__279_, data_stage_1__278_, data_stage_1__277_, data_stage_1__276_, data_stage_1__275_, data_stage_1__274_, data_stage_1__273_, data_stage_1__272_, data_stage_1__271_, data_stage_1__270_, data_stage_1__269_, data_stage_1__268_, data_stage_1__267_, data_stage_1__266_, data_stage_1__265_, data_stage_1__264_, data_stage_1__263_, data_stage_1__262_, data_stage_1__261_, data_stage_1__260_, data_stage_1__259_, data_stage_1__258_, data_stage_1__257_, data_stage_1__256_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_3__swap_inst
  (
    .data_i(data_i[511:384]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__511_, data_stage_1__510_, data_stage_1__509_, data_stage_1__508_, data_stage_1__507_, data_stage_1__506_, data_stage_1__505_, data_stage_1__504_, data_stage_1__503_, data_stage_1__502_, data_stage_1__501_, data_stage_1__500_, data_stage_1__499_, data_stage_1__498_, data_stage_1__497_, data_stage_1__496_, data_stage_1__495_, data_stage_1__494_, data_stage_1__493_, data_stage_1__492_, data_stage_1__491_, data_stage_1__490_, data_stage_1__489_, data_stage_1__488_, data_stage_1__487_, data_stage_1__486_, data_stage_1__485_, data_stage_1__484_, data_stage_1__483_, data_stage_1__482_, data_stage_1__481_, data_stage_1__480_, data_stage_1__479_, data_stage_1__478_, data_stage_1__477_, data_stage_1__476_, data_stage_1__475_, data_stage_1__474_, data_stage_1__473_, data_stage_1__472_, data_stage_1__471_, data_stage_1__470_, data_stage_1__469_, data_stage_1__468_, data_stage_1__467_, data_stage_1__466_, data_stage_1__465_, data_stage_1__464_, data_stage_1__463_, data_stage_1__462_, data_stage_1__461_, data_stage_1__460_, data_stage_1__459_, data_stage_1__458_, data_stage_1__457_, data_stage_1__456_, data_stage_1__455_, data_stage_1__454_, data_stage_1__453_, data_stage_1__452_, data_stage_1__451_, data_stage_1__450_, data_stage_1__449_, data_stage_1__448_, data_stage_1__447_, data_stage_1__446_, data_stage_1__445_, data_stage_1__444_, data_stage_1__443_, data_stage_1__442_, data_stage_1__441_, data_stage_1__440_, data_stage_1__439_, data_stage_1__438_, data_stage_1__437_, data_stage_1__436_, data_stage_1__435_, data_stage_1__434_, data_stage_1__433_, data_stage_1__432_, data_stage_1__431_, data_stage_1__430_, data_stage_1__429_, data_stage_1__428_, data_stage_1__427_, data_stage_1__426_, data_stage_1__425_, data_stage_1__424_, data_stage_1__423_, data_stage_1__422_, data_stage_1__421_, data_stage_1__420_, data_stage_1__419_, data_stage_1__418_, data_stage_1__417_, data_stage_1__416_, data_stage_1__415_, data_stage_1__414_, data_stage_1__413_, data_stage_1__412_, data_stage_1__411_, data_stage_1__410_, data_stage_1__409_, data_stage_1__408_, data_stage_1__407_, data_stage_1__406_, data_stage_1__405_, data_stage_1__404_, data_stage_1__403_, data_stage_1__402_, data_stage_1__401_, data_stage_1__400_, data_stage_1__399_, data_stage_1__398_, data_stage_1__397_, data_stage_1__396_, data_stage_1__395_, data_stage_1__394_, data_stage_1__393_, data_stage_1__392_, data_stage_1__391_, data_stage_1__390_, data_stage_1__389_, data_stage_1__388_, data_stage_1__387_, data_stage_1__386_, data_stage_1__385_, data_stage_1__384_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_4__swap_inst
  (
    .data_i(data_i[639:512]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__639_, data_stage_1__638_, data_stage_1__637_, data_stage_1__636_, data_stage_1__635_, data_stage_1__634_, data_stage_1__633_, data_stage_1__632_, data_stage_1__631_, data_stage_1__630_, data_stage_1__629_, data_stage_1__628_, data_stage_1__627_, data_stage_1__626_, data_stage_1__625_, data_stage_1__624_, data_stage_1__623_, data_stage_1__622_, data_stage_1__621_, data_stage_1__620_, data_stage_1__619_, data_stage_1__618_, data_stage_1__617_, data_stage_1__616_, data_stage_1__615_, data_stage_1__614_, data_stage_1__613_, data_stage_1__612_, data_stage_1__611_, data_stage_1__610_, data_stage_1__609_, data_stage_1__608_, data_stage_1__607_, data_stage_1__606_, data_stage_1__605_, data_stage_1__604_, data_stage_1__603_, data_stage_1__602_, data_stage_1__601_, data_stage_1__600_, data_stage_1__599_, data_stage_1__598_, data_stage_1__597_, data_stage_1__596_, data_stage_1__595_, data_stage_1__594_, data_stage_1__593_, data_stage_1__592_, data_stage_1__591_, data_stage_1__590_, data_stage_1__589_, data_stage_1__588_, data_stage_1__587_, data_stage_1__586_, data_stage_1__585_, data_stage_1__584_, data_stage_1__583_, data_stage_1__582_, data_stage_1__581_, data_stage_1__580_, data_stage_1__579_, data_stage_1__578_, data_stage_1__577_, data_stage_1__576_, data_stage_1__575_, data_stage_1__574_, data_stage_1__573_, data_stage_1__572_, data_stage_1__571_, data_stage_1__570_, data_stage_1__569_, data_stage_1__568_, data_stage_1__567_, data_stage_1__566_, data_stage_1__565_, data_stage_1__564_, data_stage_1__563_, data_stage_1__562_, data_stage_1__561_, data_stage_1__560_, data_stage_1__559_, data_stage_1__558_, data_stage_1__557_, data_stage_1__556_, data_stage_1__555_, data_stage_1__554_, data_stage_1__553_, data_stage_1__552_, data_stage_1__551_, data_stage_1__550_, data_stage_1__549_, data_stage_1__548_, data_stage_1__547_, data_stage_1__546_, data_stage_1__545_, data_stage_1__544_, data_stage_1__543_, data_stage_1__542_, data_stage_1__541_, data_stage_1__540_, data_stage_1__539_, data_stage_1__538_, data_stage_1__537_, data_stage_1__536_, data_stage_1__535_, data_stage_1__534_, data_stage_1__533_, data_stage_1__532_, data_stage_1__531_, data_stage_1__530_, data_stage_1__529_, data_stage_1__528_, data_stage_1__527_, data_stage_1__526_, data_stage_1__525_, data_stage_1__524_, data_stage_1__523_, data_stage_1__522_, data_stage_1__521_, data_stage_1__520_, data_stage_1__519_, data_stage_1__518_, data_stage_1__517_, data_stage_1__516_, data_stage_1__515_, data_stage_1__514_, data_stage_1__513_, data_stage_1__512_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_5__swap_inst
  (
    .data_i(data_i[767:640]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__767_, data_stage_1__766_, data_stage_1__765_, data_stage_1__764_, data_stage_1__763_, data_stage_1__762_, data_stage_1__761_, data_stage_1__760_, data_stage_1__759_, data_stage_1__758_, data_stage_1__757_, data_stage_1__756_, data_stage_1__755_, data_stage_1__754_, data_stage_1__753_, data_stage_1__752_, data_stage_1__751_, data_stage_1__750_, data_stage_1__749_, data_stage_1__748_, data_stage_1__747_, data_stage_1__746_, data_stage_1__745_, data_stage_1__744_, data_stage_1__743_, data_stage_1__742_, data_stage_1__741_, data_stage_1__740_, data_stage_1__739_, data_stage_1__738_, data_stage_1__737_, data_stage_1__736_, data_stage_1__735_, data_stage_1__734_, data_stage_1__733_, data_stage_1__732_, data_stage_1__731_, data_stage_1__730_, data_stage_1__729_, data_stage_1__728_, data_stage_1__727_, data_stage_1__726_, data_stage_1__725_, data_stage_1__724_, data_stage_1__723_, data_stage_1__722_, data_stage_1__721_, data_stage_1__720_, data_stage_1__719_, data_stage_1__718_, data_stage_1__717_, data_stage_1__716_, data_stage_1__715_, data_stage_1__714_, data_stage_1__713_, data_stage_1__712_, data_stage_1__711_, data_stage_1__710_, data_stage_1__709_, data_stage_1__708_, data_stage_1__707_, data_stage_1__706_, data_stage_1__705_, data_stage_1__704_, data_stage_1__703_, data_stage_1__702_, data_stage_1__701_, data_stage_1__700_, data_stage_1__699_, data_stage_1__698_, data_stage_1__697_, data_stage_1__696_, data_stage_1__695_, data_stage_1__694_, data_stage_1__693_, data_stage_1__692_, data_stage_1__691_, data_stage_1__690_, data_stage_1__689_, data_stage_1__688_, data_stage_1__687_, data_stage_1__686_, data_stage_1__685_, data_stage_1__684_, data_stage_1__683_, data_stage_1__682_, data_stage_1__681_, data_stage_1__680_, data_stage_1__679_, data_stage_1__678_, data_stage_1__677_, data_stage_1__676_, data_stage_1__675_, data_stage_1__674_, data_stage_1__673_, data_stage_1__672_, data_stage_1__671_, data_stage_1__670_, data_stage_1__669_, data_stage_1__668_, data_stage_1__667_, data_stage_1__666_, data_stage_1__665_, data_stage_1__664_, data_stage_1__663_, data_stage_1__662_, data_stage_1__661_, data_stage_1__660_, data_stage_1__659_, data_stage_1__658_, data_stage_1__657_, data_stage_1__656_, data_stage_1__655_, data_stage_1__654_, data_stage_1__653_, data_stage_1__652_, data_stage_1__651_, data_stage_1__650_, data_stage_1__649_, data_stage_1__648_, data_stage_1__647_, data_stage_1__646_, data_stage_1__645_, data_stage_1__644_, data_stage_1__643_, data_stage_1__642_, data_stage_1__641_, data_stage_1__640_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_6__swap_inst
  (
    .data_i(data_i[895:768]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__895_, data_stage_1__894_, data_stage_1__893_, data_stage_1__892_, data_stage_1__891_, data_stage_1__890_, data_stage_1__889_, data_stage_1__888_, data_stage_1__887_, data_stage_1__886_, data_stage_1__885_, data_stage_1__884_, data_stage_1__883_, data_stage_1__882_, data_stage_1__881_, data_stage_1__880_, data_stage_1__879_, data_stage_1__878_, data_stage_1__877_, data_stage_1__876_, data_stage_1__875_, data_stage_1__874_, data_stage_1__873_, data_stage_1__872_, data_stage_1__871_, data_stage_1__870_, data_stage_1__869_, data_stage_1__868_, data_stage_1__867_, data_stage_1__866_, data_stage_1__865_, data_stage_1__864_, data_stage_1__863_, data_stage_1__862_, data_stage_1__861_, data_stage_1__860_, data_stage_1__859_, data_stage_1__858_, data_stage_1__857_, data_stage_1__856_, data_stage_1__855_, data_stage_1__854_, data_stage_1__853_, data_stage_1__852_, data_stage_1__851_, data_stage_1__850_, data_stage_1__849_, data_stage_1__848_, data_stage_1__847_, data_stage_1__846_, data_stage_1__845_, data_stage_1__844_, data_stage_1__843_, data_stage_1__842_, data_stage_1__841_, data_stage_1__840_, data_stage_1__839_, data_stage_1__838_, data_stage_1__837_, data_stage_1__836_, data_stage_1__835_, data_stage_1__834_, data_stage_1__833_, data_stage_1__832_, data_stage_1__831_, data_stage_1__830_, data_stage_1__829_, data_stage_1__828_, data_stage_1__827_, data_stage_1__826_, data_stage_1__825_, data_stage_1__824_, data_stage_1__823_, data_stage_1__822_, data_stage_1__821_, data_stage_1__820_, data_stage_1__819_, data_stage_1__818_, data_stage_1__817_, data_stage_1__816_, data_stage_1__815_, data_stage_1__814_, data_stage_1__813_, data_stage_1__812_, data_stage_1__811_, data_stage_1__810_, data_stage_1__809_, data_stage_1__808_, data_stage_1__807_, data_stage_1__806_, data_stage_1__805_, data_stage_1__804_, data_stage_1__803_, data_stage_1__802_, data_stage_1__801_, data_stage_1__800_, data_stage_1__799_, data_stage_1__798_, data_stage_1__797_, data_stage_1__796_, data_stage_1__795_, data_stage_1__794_, data_stage_1__793_, data_stage_1__792_, data_stage_1__791_, data_stage_1__790_, data_stage_1__789_, data_stage_1__788_, data_stage_1__787_, data_stage_1__786_, data_stage_1__785_, data_stage_1__784_, data_stage_1__783_, data_stage_1__782_, data_stage_1__781_, data_stage_1__780_, data_stage_1__779_, data_stage_1__778_, data_stage_1__777_, data_stage_1__776_, data_stage_1__775_, data_stage_1__774_, data_stage_1__773_, data_stage_1__772_, data_stage_1__771_, data_stage_1__770_, data_stage_1__769_, data_stage_1__768_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_7__swap_inst
  (
    .data_i(data_i[1023:896]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__1023_, data_stage_1__1022_, data_stage_1__1021_, data_stage_1__1020_, data_stage_1__1019_, data_stage_1__1018_, data_stage_1__1017_, data_stage_1__1016_, data_stage_1__1015_, data_stage_1__1014_, data_stage_1__1013_, data_stage_1__1012_, data_stage_1__1011_, data_stage_1__1010_, data_stage_1__1009_, data_stage_1__1008_, data_stage_1__1007_, data_stage_1__1006_, data_stage_1__1005_, data_stage_1__1004_, data_stage_1__1003_, data_stage_1__1002_, data_stage_1__1001_, data_stage_1__1000_, data_stage_1__999_, data_stage_1__998_, data_stage_1__997_, data_stage_1__996_, data_stage_1__995_, data_stage_1__994_, data_stage_1__993_, data_stage_1__992_, data_stage_1__991_, data_stage_1__990_, data_stage_1__989_, data_stage_1__988_, data_stage_1__987_, data_stage_1__986_, data_stage_1__985_, data_stage_1__984_, data_stage_1__983_, data_stage_1__982_, data_stage_1__981_, data_stage_1__980_, data_stage_1__979_, data_stage_1__978_, data_stage_1__977_, data_stage_1__976_, data_stage_1__975_, data_stage_1__974_, data_stage_1__973_, data_stage_1__972_, data_stage_1__971_, data_stage_1__970_, data_stage_1__969_, data_stage_1__968_, data_stage_1__967_, data_stage_1__966_, data_stage_1__965_, data_stage_1__964_, data_stage_1__963_, data_stage_1__962_, data_stage_1__961_, data_stage_1__960_, data_stage_1__959_, data_stage_1__958_, data_stage_1__957_, data_stage_1__956_, data_stage_1__955_, data_stage_1__954_, data_stage_1__953_, data_stage_1__952_, data_stage_1__951_, data_stage_1__950_, data_stage_1__949_, data_stage_1__948_, data_stage_1__947_, data_stage_1__946_, data_stage_1__945_, data_stage_1__944_, data_stage_1__943_, data_stage_1__942_, data_stage_1__941_, data_stage_1__940_, data_stage_1__939_, data_stage_1__938_, data_stage_1__937_, data_stage_1__936_, data_stage_1__935_, data_stage_1__934_, data_stage_1__933_, data_stage_1__932_, data_stage_1__931_, data_stage_1__930_, data_stage_1__929_, data_stage_1__928_, data_stage_1__927_, data_stage_1__926_, data_stage_1__925_, data_stage_1__924_, data_stage_1__923_, data_stage_1__922_, data_stage_1__921_, data_stage_1__920_, data_stage_1__919_, data_stage_1__918_, data_stage_1__917_, data_stage_1__916_, data_stage_1__915_, data_stage_1__914_, data_stage_1__913_, data_stage_1__912_, data_stage_1__911_, data_stage_1__910_, data_stage_1__909_, data_stage_1__908_, data_stage_1__907_, data_stage_1__906_, data_stage_1__905_, data_stage_1__904_, data_stage_1__903_, data_stage_1__902_, data_stage_1__901_, data_stage_1__900_, data_stage_1__899_, data_stage_1__898_, data_stage_1__897_, data_stage_1__896_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_8__swap_inst
  (
    .data_i(data_i[1151:1024]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__1151_, data_stage_1__1150_, data_stage_1__1149_, data_stage_1__1148_, data_stage_1__1147_, data_stage_1__1146_, data_stage_1__1145_, data_stage_1__1144_, data_stage_1__1143_, data_stage_1__1142_, data_stage_1__1141_, data_stage_1__1140_, data_stage_1__1139_, data_stage_1__1138_, data_stage_1__1137_, data_stage_1__1136_, data_stage_1__1135_, data_stage_1__1134_, data_stage_1__1133_, data_stage_1__1132_, data_stage_1__1131_, data_stage_1__1130_, data_stage_1__1129_, data_stage_1__1128_, data_stage_1__1127_, data_stage_1__1126_, data_stage_1__1125_, data_stage_1__1124_, data_stage_1__1123_, data_stage_1__1122_, data_stage_1__1121_, data_stage_1__1120_, data_stage_1__1119_, data_stage_1__1118_, data_stage_1__1117_, data_stage_1__1116_, data_stage_1__1115_, data_stage_1__1114_, data_stage_1__1113_, data_stage_1__1112_, data_stage_1__1111_, data_stage_1__1110_, data_stage_1__1109_, data_stage_1__1108_, data_stage_1__1107_, data_stage_1__1106_, data_stage_1__1105_, data_stage_1__1104_, data_stage_1__1103_, data_stage_1__1102_, data_stage_1__1101_, data_stage_1__1100_, data_stage_1__1099_, data_stage_1__1098_, data_stage_1__1097_, data_stage_1__1096_, data_stage_1__1095_, data_stage_1__1094_, data_stage_1__1093_, data_stage_1__1092_, data_stage_1__1091_, data_stage_1__1090_, data_stage_1__1089_, data_stage_1__1088_, data_stage_1__1087_, data_stage_1__1086_, data_stage_1__1085_, data_stage_1__1084_, data_stage_1__1083_, data_stage_1__1082_, data_stage_1__1081_, data_stage_1__1080_, data_stage_1__1079_, data_stage_1__1078_, data_stage_1__1077_, data_stage_1__1076_, data_stage_1__1075_, data_stage_1__1074_, data_stage_1__1073_, data_stage_1__1072_, data_stage_1__1071_, data_stage_1__1070_, data_stage_1__1069_, data_stage_1__1068_, data_stage_1__1067_, data_stage_1__1066_, data_stage_1__1065_, data_stage_1__1064_, data_stage_1__1063_, data_stage_1__1062_, data_stage_1__1061_, data_stage_1__1060_, data_stage_1__1059_, data_stage_1__1058_, data_stage_1__1057_, data_stage_1__1056_, data_stage_1__1055_, data_stage_1__1054_, data_stage_1__1053_, data_stage_1__1052_, data_stage_1__1051_, data_stage_1__1050_, data_stage_1__1049_, data_stage_1__1048_, data_stage_1__1047_, data_stage_1__1046_, data_stage_1__1045_, data_stage_1__1044_, data_stage_1__1043_, data_stage_1__1042_, data_stage_1__1041_, data_stage_1__1040_, data_stage_1__1039_, data_stage_1__1038_, data_stage_1__1037_, data_stage_1__1036_, data_stage_1__1035_, data_stage_1__1034_, data_stage_1__1033_, data_stage_1__1032_, data_stage_1__1031_, data_stage_1__1030_, data_stage_1__1029_, data_stage_1__1028_, data_stage_1__1027_, data_stage_1__1026_, data_stage_1__1025_, data_stage_1__1024_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_9__swap_inst
  (
    .data_i(data_i[1279:1152]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__1279_, data_stage_1__1278_, data_stage_1__1277_, data_stage_1__1276_, data_stage_1__1275_, data_stage_1__1274_, data_stage_1__1273_, data_stage_1__1272_, data_stage_1__1271_, data_stage_1__1270_, data_stage_1__1269_, data_stage_1__1268_, data_stage_1__1267_, data_stage_1__1266_, data_stage_1__1265_, data_stage_1__1264_, data_stage_1__1263_, data_stage_1__1262_, data_stage_1__1261_, data_stage_1__1260_, data_stage_1__1259_, data_stage_1__1258_, data_stage_1__1257_, data_stage_1__1256_, data_stage_1__1255_, data_stage_1__1254_, data_stage_1__1253_, data_stage_1__1252_, data_stage_1__1251_, data_stage_1__1250_, data_stage_1__1249_, data_stage_1__1248_, data_stage_1__1247_, data_stage_1__1246_, data_stage_1__1245_, data_stage_1__1244_, data_stage_1__1243_, data_stage_1__1242_, data_stage_1__1241_, data_stage_1__1240_, data_stage_1__1239_, data_stage_1__1238_, data_stage_1__1237_, data_stage_1__1236_, data_stage_1__1235_, data_stage_1__1234_, data_stage_1__1233_, data_stage_1__1232_, data_stage_1__1231_, data_stage_1__1230_, data_stage_1__1229_, data_stage_1__1228_, data_stage_1__1227_, data_stage_1__1226_, data_stage_1__1225_, data_stage_1__1224_, data_stage_1__1223_, data_stage_1__1222_, data_stage_1__1221_, data_stage_1__1220_, data_stage_1__1219_, data_stage_1__1218_, data_stage_1__1217_, data_stage_1__1216_, data_stage_1__1215_, data_stage_1__1214_, data_stage_1__1213_, data_stage_1__1212_, data_stage_1__1211_, data_stage_1__1210_, data_stage_1__1209_, data_stage_1__1208_, data_stage_1__1207_, data_stage_1__1206_, data_stage_1__1205_, data_stage_1__1204_, data_stage_1__1203_, data_stage_1__1202_, data_stage_1__1201_, data_stage_1__1200_, data_stage_1__1199_, data_stage_1__1198_, data_stage_1__1197_, data_stage_1__1196_, data_stage_1__1195_, data_stage_1__1194_, data_stage_1__1193_, data_stage_1__1192_, data_stage_1__1191_, data_stage_1__1190_, data_stage_1__1189_, data_stage_1__1188_, data_stage_1__1187_, data_stage_1__1186_, data_stage_1__1185_, data_stage_1__1184_, data_stage_1__1183_, data_stage_1__1182_, data_stage_1__1181_, data_stage_1__1180_, data_stage_1__1179_, data_stage_1__1178_, data_stage_1__1177_, data_stage_1__1176_, data_stage_1__1175_, data_stage_1__1174_, data_stage_1__1173_, data_stage_1__1172_, data_stage_1__1171_, data_stage_1__1170_, data_stage_1__1169_, data_stage_1__1168_, data_stage_1__1167_, data_stage_1__1166_, data_stage_1__1165_, data_stage_1__1164_, data_stage_1__1163_, data_stage_1__1162_, data_stage_1__1161_, data_stage_1__1160_, data_stage_1__1159_, data_stage_1__1158_, data_stage_1__1157_, data_stage_1__1156_, data_stage_1__1155_, data_stage_1__1154_, data_stage_1__1153_, data_stage_1__1152_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_10__swap_inst
  (
    .data_i(data_i[1407:1280]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__1407_, data_stage_1__1406_, data_stage_1__1405_, data_stage_1__1404_, data_stage_1__1403_, data_stage_1__1402_, data_stage_1__1401_, data_stage_1__1400_, data_stage_1__1399_, data_stage_1__1398_, data_stage_1__1397_, data_stage_1__1396_, data_stage_1__1395_, data_stage_1__1394_, data_stage_1__1393_, data_stage_1__1392_, data_stage_1__1391_, data_stage_1__1390_, data_stage_1__1389_, data_stage_1__1388_, data_stage_1__1387_, data_stage_1__1386_, data_stage_1__1385_, data_stage_1__1384_, data_stage_1__1383_, data_stage_1__1382_, data_stage_1__1381_, data_stage_1__1380_, data_stage_1__1379_, data_stage_1__1378_, data_stage_1__1377_, data_stage_1__1376_, data_stage_1__1375_, data_stage_1__1374_, data_stage_1__1373_, data_stage_1__1372_, data_stage_1__1371_, data_stage_1__1370_, data_stage_1__1369_, data_stage_1__1368_, data_stage_1__1367_, data_stage_1__1366_, data_stage_1__1365_, data_stage_1__1364_, data_stage_1__1363_, data_stage_1__1362_, data_stage_1__1361_, data_stage_1__1360_, data_stage_1__1359_, data_stage_1__1358_, data_stage_1__1357_, data_stage_1__1356_, data_stage_1__1355_, data_stage_1__1354_, data_stage_1__1353_, data_stage_1__1352_, data_stage_1__1351_, data_stage_1__1350_, data_stage_1__1349_, data_stage_1__1348_, data_stage_1__1347_, data_stage_1__1346_, data_stage_1__1345_, data_stage_1__1344_, data_stage_1__1343_, data_stage_1__1342_, data_stage_1__1341_, data_stage_1__1340_, data_stage_1__1339_, data_stage_1__1338_, data_stage_1__1337_, data_stage_1__1336_, data_stage_1__1335_, data_stage_1__1334_, data_stage_1__1333_, data_stage_1__1332_, data_stage_1__1331_, data_stage_1__1330_, data_stage_1__1329_, data_stage_1__1328_, data_stage_1__1327_, data_stage_1__1326_, data_stage_1__1325_, data_stage_1__1324_, data_stage_1__1323_, data_stage_1__1322_, data_stage_1__1321_, data_stage_1__1320_, data_stage_1__1319_, data_stage_1__1318_, data_stage_1__1317_, data_stage_1__1316_, data_stage_1__1315_, data_stage_1__1314_, data_stage_1__1313_, data_stage_1__1312_, data_stage_1__1311_, data_stage_1__1310_, data_stage_1__1309_, data_stage_1__1308_, data_stage_1__1307_, data_stage_1__1306_, data_stage_1__1305_, data_stage_1__1304_, data_stage_1__1303_, data_stage_1__1302_, data_stage_1__1301_, data_stage_1__1300_, data_stage_1__1299_, data_stage_1__1298_, data_stage_1__1297_, data_stage_1__1296_, data_stage_1__1295_, data_stage_1__1294_, data_stage_1__1293_, data_stage_1__1292_, data_stage_1__1291_, data_stage_1__1290_, data_stage_1__1289_, data_stage_1__1288_, data_stage_1__1287_, data_stage_1__1286_, data_stage_1__1285_, data_stage_1__1284_, data_stage_1__1283_, data_stage_1__1282_, data_stage_1__1281_, data_stage_1__1280_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_11__swap_inst
  (
    .data_i(data_i[1535:1408]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__1535_, data_stage_1__1534_, data_stage_1__1533_, data_stage_1__1532_, data_stage_1__1531_, data_stage_1__1530_, data_stage_1__1529_, data_stage_1__1528_, data_stage_1__1527_, data_stage_1__1526_, data_stage_1__1525_, data_stage_1__1524_, data_stage_1__1523_, data_stage_1__1522_, data_stage_1__1521_, data_stage_1__1520_, data_stage_1__1519_, data_stage_1__1518_, data_stage_1__1517_, data_stage_1__1516_, data_stage_1__1515_, data_stage_1__1514_, data_stage_1__1513_, data_stage_1__1512_, data_stage_1__1511_, data_stage_1__1510_, data_stage_1__1509_, data_stage_1__1508_, data_stage_1__1507_, data_stage_1__1506_, data_stage_1__1505_, data_stage_1__1504_, data_stage_1__1503_, data_stage_1__1502_, data_stage_1__1501_, data_stage_1__1500_, data_stage_1__1499_, data_stage_1__1498_, data_stage_1__1497_, data_stage_1__1496_, data_stage_1__1495_, data_stage_1__1494_, data_stage_1__1493_, data_stage_1__1492_, data_stage_1__1491_, data_stage_1__1490_, data_stage_1__1489_, data_stage_1__1488_, data_stage_1__1487_, data_stage_1__1486_, data_stage_1__1485_, data_stage_1__1484_, data_stage_1__1483_, data_stage_1__1482_, data_stage_1__1481_, data_stage_1__1480_, data_stage_1__1479_, data_stage_1__1478_, data_stage_1__1477_, data_stage_1__1476_, data_stage_1__1475_, data_stage_1__1474_, data_stage_1__1473_, data_stage_1__1472_, data_stage_1__1471_, data_stage_1__1470_, data_stage_1__1469_, data_stage_1__1468_, data_stage_1__1467_, data_stage_1__1466_, data_stage_1__1465_, data_stage_1__1464_, data_stage_1__1463_, data_stage_1__1462_, data_stage_1__1461_, data_stage_1__1460_, data_stage_1__1459_, data_stage_1__1458_, data_stage_1__1457_, data_stage_1__1456_, data_stage_1__1455_, data_stage_1__1454_, data_stage_1__1453_, data_stage_1__1452_, data_stage_1__1451_, data_stage_1__1450_, data_stage_1__1449_, data_stage_1__1448_, data_stage_1__1447_, data_stage_1__1446_, data_stage_1__1445_, data_stage_1__1444_, data_stage_1__1443_, data_stage_1__1442_, data_stage_1__1441_, data_stage_1__1440_, data_stage_1__1439_, data_stage_1__1438_, data_stage_1__1437_, data_stage_1__1436_, data_stage_1__1435_, data_stage_1__1434_, data_stage_1__1433_, data_stage_1__1432_, data_stage_1__1431_, data_stage_1__1430_, data_stage_1__1429_, data_stage_1__1428_, data_stage_1__1427_, data_stage_1__1426_, data_stage_1__1425_, data_stage_1__1424_, data_stage_1__1423_, data_stage_1__1422_, data_stage_1__1421_, data_stage_1__1420_, data_stage_1__1419_, data_stage_1__1418_, data_stage_1__1417_, data_stage_1__1416_, data_stage_1__1415_, data_stage_1__1414_, data_stage_1__1413_, data_stage_1__1412_, data_stage_1__1411_, data_stage_1__1410_, data_stage_1__1409_, data_stage_1__1408_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_12__swap_inst
  (
    .data_i(data_i[1663:1536]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__1663_, data_stage_1__1662_, data_stage_1__1661_, data_stage_1__1660_, data_stage_1__1659_, data_stage_1__1658_, data_stage_1__1657_, data_stage_1__1656_, data_stage_1__1655_, data_stage_1__1654_, data_stage_1__1653_, data_stage_1__1652_, data_stage_1__1651_, data_stage_1__1650_, data_stage_1__1649_, data_stage_1__1648_, data_stage_1__1647_, data_stage_1__1646_, data_stage_1__1645_, data_stage_1__1644_, data_stage_1__1643_, data_stage_1__1642_, data_stage_1__1641_, data_stage_1__1640_, data_stage_1__1639_, data_stage_1__1638_, data_stage_1__1637_, data_stage_1__1636_, data_stage_1__1635_, data_stage_1__1634_, data_stage_1__1633_, data_stage_1__1632_, data_stage_1__1631_, data_stage_1__1630_, data_stage_1__1629_, data_stage_1__1628_, data_stage_1__1627_, data_stage_1__1626_, data_stage_1__1625_, data_stage_1__1624_, data_stage_1__1623_, data_stage_1__1622_, data_stage_1__1621_, data_stage_1__1620_, data_stage_1__1619_, data_stage_1__1618_, data_stage_1__1617_, data_stage_1__1616_, data_stage_1__1615_, data_stage_1__1614_, data_stage_1__1613_, data_stage_1__1612_, data_stage_1__1611_, data_stage_1__1610_, data_stage_1__1609_, data_stage_1__1608_, data_stage_1__1607_, data_stage_1__1606_, data_stage_1__1605_, data_stage_1__1604_, data_stage_1__1603_, data_stage_1__1602_, data_stage_1__1601_, data_stage_1__1600_, data_stage_1__1599_, data_stage_1__1598_, data_stage_1__1597_, data_stage_1__1596_, data_stage_1__1595_, data_stage_1__1594_, data_stage_1__1593_, data_stage_1__1592_, data_stage_1__1591_, data_stage_1__1590_, data_stage_1__1589_, data_stage_1__1588_, data_stage_1__1587_, data_stage_1__1586_, data_stage_1__1585_, data_stage_1__1584_, data_stage_1__1583_, data_stage_1__1582_, data_stage_1__1581_, data_stage_1__1580_, data_stage_1__1579_, data_stage_1__1578_, data_stage_1__1577_, data_stage_1__1576_, data_stage_1__1575_, data_stage_1__1574_, data_stage_1__1573_, data_stage_1__1572_, data_stage_1__1571_, data_stage_1__1570_, data_stage_1__1569_, data_stage_1__1568_, data_stage_1__1567_, data_stage_1__1566_, data_stage_1__1565_, data_stage_1__1564_, data_stage_1__1563_, data_stage_1__1562_, data_stage_1__1561_, data_stage_1__1560_, data_stage_1__1559_, data_stage_1__1558_, data_stage_1__1557_, data_stage_1__1556_, data_stage_1__1555_, data_stage_1__1554_, data_stage_1__1553_, data_stage_1__1552_, data_stage_1__1551_, data_stage_1__1550_, data_stage_1__1549_, data_stage_1__1548_, data_stage_1__1547_, data_stage_1__1546_, data_stage_1__1545_, data_stage_1__1544_, data_stage_1__1543_, data_stage_1__1542_, data_stage_1__1541_, data_stage_1__1540_, data_stage_1__1539_, data_stage_1__1538_, data_stage_1__1537_, data_stage_1__1536_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_13__swap_inst
  (
    .data_i(data_i[1791:1664]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__1791_, data_stage_1__1790_, data_stage_1__1789_, data_stage_1__1788_, data_stage_1__1787_, data_stage_1__1786_, data_stage_1__1785_, data_stage_1__1784_, data_stage_1__1783_, data_stage_1__1782_, data_stage_1__1781_, data_stage_1__1780_, data_stage_1__1779_, data_stage_1__1778_, data_stage_1__1777_, data_stage_1__1776_, data_stage_1__1775_, data_stage_1__1774_, data_stage_1__1773_, data_stage_1__1772_, data_stage_1__1771_, data_stage_1__1770_, data_stage_1__1769_, data_stage_1__1768_, data_stage_1__1767_, data_stage_1__1766_, data_stage_1__1765_, data_stage_1__1764_, data_stage_1__1763_, data_stage_1__1762_, data_stage_1__1761_, data_stage_1__1760_, data_stage_1__1759_, data_stage_1__1758_, data_stage_1__1757_, data_stage_1__1756_, data_stage_1__1755_, data_stage_1__1754_, data_stage_1__1753_, data_stage_1__1752_, data_stage_1__1751_, data_stage_1__1750_, data_stage_1__1749_, data_stage_1__1748_, data_stage_1__1747_, data_stage_1__1746_, data_stage_1__1745_, data_stage_1__1744_, data_stage_1__1743_, data_stage_1__1742_, data_stage_1__1741_, data_stage_1__1740_, data_stage_1__1739_, data_stage_1__1738_, data_stage_1__1737_, data_stage_1__1736_, data_stage_1__1735_, data_stage_1__1734_, data_stage_1__1733_, data_stage_1__1732_, data_stage_1__1731_, data_stage_1__1730_, data_stage_1__1729_, data_stage_1__1728_, data_stage_1__1727_, data_stage_1__1726_, data_stage_1__1725_, data_stage_1__1724_, data_stage_1__1723_, data_stage_1__1722_, data_stage_1__1721_, data_stage_1__1720_, data_stage_1__1719_, data_stage_1__1718_, data_stage_1__1717_, data_stage_1__1716_, data_stage_1__1715_, data_stage_1__1714_, data_stage_1__1713_, data_stage_1__1712_, data_stage_1__1711_, data_stage_1__1710_, data_stage_1__1709_, data_stage_1__1708_, data_stage_1__1707_, data_stage_1__1706_, data_stage_1__1705_, data_stage_1__1704_, data_stage_1__1703_, data_stage_1__1702_, data_stage_1__1701_, data_stage_1__1700_, data_stage_1__1699_, data_stage_1__1698_, data_stage_1__1697_, data_stage_1__1696_, data_stage_1__1695_, data_stage_1__1694_, data_stage_1__1693_, data_stage_1__1692_, data_stage_1__1691_, data_stage_1__1690_, data_stage_1__1689_, data_stage_1__1688_, data_stage_1__1687_, data_stage_1__1686_, data_stage_1__1685_, data_stage_1__1684_, data_stage_1__1683_, data_stage_1__1682_, data_stage_1__1681_, data_stage_1__1680_, data_stage_1__1679_, data_stage_1__1678_, data_stage_1__1677_, data_stage_1__1676_, data_stage_1__1675_, data_stage_1__1674_, data_stage_1__1673_, data_stage_1__1672_, data_stage_1__1671_, data_stage_1__1670_, data_stage_1__1669_, data_stage_1__1668_, data_stage_1__1667_, data_stage_1__1666_, data_stage_1__1665_, data_stage_1__1664_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_14__swap_inst
  (
    .data_i(data_i[1919:1792]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__1919_, data_stage_1__1918_, data_stage_1__1917_, data_stage_1__1916_, data_stage_1__1915_, data_stage_1__1914_, data_stage_1__1913_, data_stage_1__1912_, data_stage_1__1911_, data_stage_1__1910_, data_stage_1__1909_, data_stage_1__1908_, data_stage_1__1907_, data_stage_1__1906_, data_stage_1__1905_, data_stage_1__1904_, data_stage_1__1903_, data_stage_1__1902_, data_stage_1__1901_, data_stage_1__1900_, data_stage_1__1899_, data_stage_1__1898_, data_stage_1__1897_, data_stage_1__1896_, data_stage_1__1895_, data_stage_1__1894_, data_stage_1__1893_, data_stage_1__1892_, data_stage_1__1891_, data_stage_1__1890_, data_stage_1__1889_, data_stage_1__1888_, data_stage_1__1887_, data_stage_1__1886_, data_stage_1__1885_, data_stage_1__1884_, data_stage_1__1883_, data_stage_1__1882_, data_stage_1__1881_, data_stage_1__1880_, data_stage_1__1879_, data_stage_1__1878_, data_stage_1__1877_, data_stage_1__1876_, data_stage_1__1875_, data_stage_1__1874_, data_stage_1__1873_, data_stage_1__1872_, data_stage_1__1871_, data_stage_1__1870_, data_stage_1__1869_, data_stage_1__1868_, data_stage_1__1867_, data_stage_1__1866_, data_stage_1__1865_, data_stage_1__1864_, data_stage_1__1863_, data_stage_1__1862_, data_stage_1__1861_, data_stage_1__1860_, data_stage_1__1859_, data_stage_1__1858_, data_stage_1__1857_, data_stage_1__1856_, data_stage_1__1855_, data_stage_1__1854_, data_stage_1__1853_, data_stage_1__1852_, data_stage_1__1851_, data_stage_1__1850_, data_stage_1__1849_, data_stage_1__1848_, data_stage_1__1847_, data_stage_1__1846_, data_stage_1__1845_, data_stage_1__1844_, data_stage_1__1843_, data_stage_1__1842_, data_stage_1__1841_, data_stage_1__1840_, data_stage_1__1839_, data_stage_1__1838_, data_stage_1__1837_, data_stage_1__1836_, data_stage_1__1835_, data_stage_1__1834_, data_stage_1__1833_, data_stage_1__1832_, data_stage_1__1831_, data_stage_1__1830_, data_stage_1__1829_, data_stage_1__1828_, data_stage_1__1827_, data_stage_1__1826_, data_stage_1__1825_, data_stage_1__1824_, data_stage_1__1823_, data_stage_1__1822_, data_stage_1__1821_, data_stage_1__1820_, data_stage_1__1819_, data_stage_1__1818_, data_stage_1__1817_, data_stage_1__1816_, data_stage_1__1815_, data_stage_1__1814_, data_stage_1__1813_, data_stage_1__1812_, data_stage_1__1811_, data_stage_1__1810_, data_stage_1__1809_, data_stage_1__1808_, data_stage_1__1807_, data_stage_1__1806_, data_stage_1__1805_, data_stage_1__1804_, data_stage_1__1803_, data_stage_1__1802_, data_stage_1__1801_, data_stage_1__1800_, data_stage_1__1799_, data_stage_1__1798_, data_stage_1__1797_, data_stage_1__1796_, data_stage_1__1795_, data_stage_1__1794_, data_stage_1__1793_, data_stage_1__1792_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_15__swap_inst
  (
    .data_i(data_i[2047:1920]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__2047_, data_stage_1__2046_, data_stage_1__2045_, data_stage_1__2044_, data_stage_1__2043_, data_stage_1__2042_, data_stage_1__2041_, data_stage_1__2040_, data_stage_1__2039_, data_stage_1__2038_, data_stage_1__2037_, data_stage_1__2036_, data_stage_1__2035_, data_stage_1__2034_, data_stage_1__2033_, data_stage_1__2032_, data_stage_1__2031_, data_stage_1__2030_, data_stage_1__2029_, data_stage_1__2028_, data_stage_1__2027_, data_stage_1__2026_, data_stage_1__2025_, data_stage_1__2024_, data_stage_1__2023_, data_stage_1__2022_, data_stage_1__2021_, data_stage_1__2020_, data_stage_1__2019_, data_stage_1__2018_, data_stage_1__2017_, data_stage_1__2016_, data_stage_1__2015_, data_stage_1__2014_, data_stage_1__2013_, data_stage_1__2012_, data_stage_1__2011_, data_stage_1__2010_, data_stage_1__2009_, data_stage_1__2008_, data_stage_1__2007_, data_stage_1__2006_, data_stage_1__2005_, data_stage_1__2004_, data_stage_1__2003_, data_stage_1__2002_, data_stage_1__2001_, data_stage_1__2000_, data_stage_1__1999_, data_stage_1__1998_, data_stage_1__1997_, data_stage_1__1996_, data_stage_1__1995_, data_stage_1__1994_, data_stage_1__1993_, data_stage_1__1992_, data_stage_1__1991_, data_stage_1__1990_, data_stage_1__1989_, data_stage_1__1988_, data_stage_1__1987_, data_stage_1__1986_, data_stage_1__1985_, data_stage_1__1984_, data_stage_1__1983_, data_stage_1__1982_, data_stage_1__1981_, data_stage_1__1980_, data_stage_1__1979_, data_stage_1__1978_, data_stage_1__1977_, data_stage_1__1976_, data_stage_1__1975_, data_stage_1__1974_, data_stage_1__1973_, data_stage_1__1972_, data_stage_1__1971_, data_stage_1__1970_, data_stage_1__1969_, data_stage_1__1968_, data_stage_1__1967_, data_stage_1__1966_, data_stage_1__1965_, data_stage_1__1964_, data_stage_1__1963_, data_stage_1__1962_, data_stage_1__1961_, data_stage_1__1960_, data_stage_1__1959_, data_stage_1__1958_, data_stage_1__1957_, data_stage_1__1956_, data_stage_1__1955_, data_stage_1__1954_, data_stage_1__1953_, data_stage_1__1952_, data_stage_1__1951_, data_stage_1__1950_, data_stage_1__1949_, data_stage_1__1948_, data_stage_1__1947_, data_stage_1__1946_, data_stage_1__1945_, data_stage_1__1944_, data_stage_1__1943_, data_stage_1__1942_, data_stage_1__1941_, data_stage_1__1940_, data_stage_1__1939_, data_stage_1__1938_, data_stage_1__1937_, data_stage_1__1936_, data_stage_1__1935_, data_stage_1__1934_, data_stage_1__1933_, data_stage_1__1932_, data_stage_1__1931_, data_stage_1__1930_, data_stage_1__1929_, data_stage_1__1928_, data_stage_1__1927_, data_stage_1__1926_, data_stage_1__1925_, data_stage_1__1924_, data_stage_1__1923_, data_stage_1__1922_, data_stage_1__1921_, data_stage_1__1920_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_16__swap_inst
  (
    .data_i(data_i[2175:2048]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__2175_, data_stage_1__2174_, data_stage_1__2173_, data_stage_1__2172_, data_stage_1__2171_, data_stage_1__2170_, data_stage_1__2169_, data_stage_1__2168_, data_stage_1__2167_, data_stage_1__2166_, data_stage_1__2165_, data_stage_1__2164_, data_stage_1__2163_, data_stage_1__2162_, data_stage_1__2161_, data_stage_1__2160_, data_stage_1__2159_, data_stage_1__2158_, data_stage_1__2157_, data_stage_1__2156_, data_stage_1__2155_, data_stage_1__2154_, data_stage_1__2153_, data_stage_1__2152_, data_stage_1__2151_, data_stage_1__2150_, data_stage_1__2149_, data_stage_1__2148_, data_stage_1__2147_, data_stage_1__2146_, data_stage_1__2145_, data_stage_1__2144_, data_stage_1__2143_, data_stage_1__2142_, data_stage_1__2141_, data_stage_1__2140_, data_stage_1__2139_, data_stage_1__2138_, data_stage_1__2137_, data_stage_1__2136_, data_stage_1__2135_, data_stage_1__2134_, data_stage_1__2133_, data_stage_1__2132_, data_stage_1__2131_, data_stage_1__2130_, data_stage_1__2129_, data_stage_1__2128_, data_stage_1__2127_, data_stage_1__2126_, data_stage_1__2125_, data_stage_1__2124_, data_stage_1__2123_, data_stage_1__2122_, data_stage_1__2121_, data_stage_1__2120_, data_stage_1__2119_, data_stage_1__2118_, data_stage_1__2117_, data_stage_1__2116_, data_stage_1__2115_, data_stage_1__2114_, data_stage_1__2113_, data_stage_1__2112_, data_stage_1__2111_, data_stage_1__2110_, data_stage_1__2109_, data_stage_1__2108_, data_stage_1__2107_, data_stage_1__2106_, data_stage_1__2105_, data_stage_1__2104_, data_stage_1__2103_, data_stage_1__2102_, data_stage_1__2101_, data_stage_1__2100_, data_stage_1__2099_, data_stage_1__2098_, data_stage_1__2097_, data_stage_1__2096_, data_stage_1__2095_, data_stage_1__2094_, data_stage_1__2093_, data_stage_1__2092_, data_stage_1__2091_, data_stage_1__2090_, data_stage_1__2089_, data_stage_1__2088_, data_stage_1__2087_, data_stage_1__2086_, data_stage_1__2085_, data_stage_1__2084_, data_stage_1__2083_, data_stage_1__2082_, data_stage_1__2081_, data_stage_1__2080_, data_stage_1__2079_, data_stage_1__2078_, data_stage_1__2077_, data_stage_1__2076_, data_stage_1__2075_, data_stage_1__2074_, data_stage_1__2073_, data_stage_1__2072_, data_stage_1__2071_, data_stage_1__2070_, data_stage_1__2069_, data_stage_1__2068_, data_stage_1__2067_, data_stage_1__2066_, data_stage_1__2065_, data_stage_1__2064_, data_stage_1__2063_, data_stage_1__2062_, data_stage_1__2061_, data_stage_1__2060_, data_stage_1__2059_, data_stage_1__2058_, data_stage_1__2057_, data_stage_1__2056_, data_stage_1__2055_, data_stage_1__2054_, data_stage_1__2053_, data_stage_1__2052_, data_stage_1__2051_, data_stage_1__2050_, data_stage_1__2049_, data_stage_1__2048_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_17__swap_inst
  (
    .data_i(data_i[2303:2176]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__2303_, data_stage_1__2302_, data_stage_1__2301_, data_stage_1__2300_, data_stage_1__2299_, data_stage_1__2298_, data_stage_1__2297_, data_stage_1__2296_, data_stage_1__2295_, data_stage_1__2294_, data_stage_1__2293_, data_stage_1__2292_, data_stage_1__2291_, data_stage_1__2290_, data_stage_1__2289_, data_stage_1__2288_, data_stage_1__2287_, data_stage_1__2286_, data_stage_1__2285_, data_stage_1__2284_, data_stage_1__2283_, data_stage_1__2282_, data_stage_1__2281_, data_stage_1__2280_, data_stage_1__2279_, data_stage_1__2278_, data_stage_1__2277_, data_stage_1__2276_, data_stage_1__2275_, data_stage_1__2274_, data_stage_1__2273_, data_stage_1__2272_, data_stage_1__2271_, data_stage_1__2270_, data_stage_1__2269_, data_stage_1__2268_, data_stage_1__2267_, data_stage_1__2266_, data_stage_1__2265_, data_stage_1__2264_, data_stage_1__2263_, data_stage_1__2262_, data_stage_1__2261_, data_stage_1__2260_, data_stage_1__2259_, data_stage_1__2258_, data_stage_1__2257_, data_stage_1__2256_, data_stage_1__2255_, data_stage_1__2254_, data_stage_1__2253_, data_stage_1__2252_, data_stage_1__2251_, data_stage_1__2250_, data_stage_1__2249_, data_stage_1__2248_, data_stage_1__2247_, data_stage_1__2246_, data_stage_1__2245_, data_stage_1__2244_, data_stage_1__2243_, data_stage_1__2242_, data_stage_1__2241_, data_stage_1__2240_, data_stage_1__2239_, data_stage_1__2238_, data_stage_1__2237_, data_stage_1__2236_, data_stage_1__2235_, data_stage_1__2234_, data_stage_1__2233_, data_stage_1__2232_, data_stage_1__2231_, data_stage_1__2230_, data_stage_1__2229_, data_stage_1__2228_, data_stage_1__2227_, data_stage_1__2226_, data_stage_1__2225_, data_stage_1__2224_, data_stage_1__2223_, data_stage_1__2222_, data_stage_1__2221_, data_stage_1__2220_, data_stage_1__2219_, data_stage_1__2218_, data_stage_1__2217_, data_stage_1__2216_, data_stage_1__2215_, data_stage_1__2214_, data_stage_1__2213_, data_stage_1__2212_, data_stage_1__2211_, data_stage_1__2210_, data_stage_1__2209_, data_stage_1__2208_, data_stage_1__2207_, data_stage_1__2206_, data_stage_1__2205_, data_stage_1__2204_, data_stage_1__2203_, data_stage_1__2202_, data_stage_1__2201_, data_stage_1__2200_, data_stage_1__2199_, data_stage_1__2198_, data_stage_1__2197_, data_stage_1__2196_, data_stage_1__2195_, data_stage_1__2194_, data_stage_1__2193_, data_stage_1__2192_, data_stage_1__2191_, data_stage_1__2190_, data_stage_1__2189_, data_stage_1__2188_, data_stage_1__2187_, data_stage_1__2186_, data_stage_1__2185_, data_stage_1__2184_, data_stage_1__2183_, data_stage_1__2182_, data_stage_1__2181_, data_stage_1__2180_, data_stage_1__2179_, data_stage_1__2178_, data_stage_1__2177_, data_stage_1__2176_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_18__swap_inst
  (
    .data_i(data_i[2431:2304]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__2431_, data_stage_1__2430_, data_stage_1__2429_, data_stage_1__2428_, data_stage_1__2427_, data_stage_1__2426_, data_stage_1__2425_, data_stage_1__2424_, data_stage_1__2423_, data_stage_1__2422_, data_stage_1__2421_, data_stage_1__2420_, data_stage_1__2419_, data_stage_1__2418_, data_stage_1__2417_, data_stage_1__2416_, data_stage_1__2415_, data_stage_1__2414_, data_stage_1__2413_, data_stage_1__2412_, data_stage_1__2411_, data_stage_1__2410_, data_stage_1__2409_, data_stage_1__2408_, data_stage_1__2407_, data_stage_1__2406_, data_stage_1__2405_, data_stage_1__2404_, data_stage_1__2403_, data_stage_1__2402_, data_stage_1__2401_, data_stage_1__2400_, data_stage_1__2399_, data_stage_1__2398_, data_stage_1__2397_, data_stage_1__2396_, data_stage_1__2395_, data_stage_1__2394_, data_stage_1__2393_, data_stage_1__2392_, data_stage_1__2391_, data_stage_1__2390_, data_stage_1__2389_, data_stage_1__2388_, data_stage_1__2387_, data_stage_1__2386_, data_stage_1__2385_, data_stage_1__2384_, data_stage_1__2383_, data_stage_1__2382_, data_stage_1__2381_, data_stage_1__2380_, data_stage_1__2379_, data_stage_1__2378_, data_stage_1__2377_, data_stage_1__2376_, data_stage_1__2375_, data_stage_1__2374_, data_stage_1__2373_, data_stage_1__2372_, data_stage_1__2371_, data_stage_1__2370_, data_stage_1__2369_, data_stage_1__2368_, data_stage_1__2367_, data_stage_1__2366_, data_stage_1__2365_, data_stage_1__2364_, data_stage_1__2363_, data_stage_1__2362_, data_stage_1__2361_, data_stage_1__2360_, data_stage_1__2359_, data_stage_1__2358_, data_stage_1__2357_, data_stage_1__2356_, data_stage_1__2355_, data_stage_1__2354_, data_stage_1__2353_, data_stage_1__2352_, data_stage_1__2351_, data_stage_1__2350_, data_stage_1__2349_, data_stage_1__2348_, data_stage_1__2347_, data_stage_1__2346_, data_stage_1__2345_, data_stage_1__2344_, data_stage_1__2343_, data_stage_1__2342_, data_stage_1__2341_, data_stage_1__2340_, data_stage_1__2339_, data_stage_1__2338_, data_stage_1__2337_, data_stage_1__2336_, data_stage_1__2335_, data_stage_1__2334_, data_stage_1__2333_, data_stage_1__2332_, data_stage_1__2331_, data_stage_1__2330_, data_stage_1__2329_, data_stage_1__2328_, data_stage_1__2327_, data_stage_1__2326_, data_stage_1__2325_, data_stage_1__2324_, data_stage_1__2323_, data_stage_1__2322_, data_stage_1__2321_, data_stage_1__2320_, data_stage_1__2319_, data_stage_1__2318_, data_stage_1__2317_, data_stage_1__2316_, data_stage_1__2315_, data_stage_1__2314_, data_stage_1__2313_, data_stage_1__2312_, data_stage_1__2311_, data_stage_1__2310_, data_stage_1__2309_, data_stage_1__2308_, data_stage_1__2307_, data_stage_1__2306_, data_stage_1__2305_, data_stage_1__2304_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_19__swap_inst
  (
    .data_i(data_i[2559:2432]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__2559_, data_stage_1__2558_, data_stage_1__2557_, data_stage_1__2556_, data_stage_1__2555_, data_stage_1__2554_, data_stage_1__2553_, data_stage_1__2552_, data_stage_1__2551_, data_stage_1__2550_, data_stage_1__2549_, data_stage_1__2548_, data_stage_1__2547_, data_stage_1__2546_, data_stage_1__2545_, data_stage_1__2544_, data_stage_1__2543_, data_stage_1__2542_, data_stage_1__2541_, data_stage_1__2540_, data_stage_1__2539_, data_stage_1__2538_, data_stage_1__2537_, data_stage_1__2536_, data_stage_1__2535_, data_stage_1__2534_, data_stage_1__2533_, data_stage_1__2532_, data_stage_1__2531_, data_stage_1__2530_, data_stage_1__2529_, data_stage_1__2528_, data_stage_1__2527_, data_stage_1__2526_, data_stage_1__2525_, data_stage_1__2524_, data_stage_1__2523_, data_stage_1__2522_, data_stage_1__2521_, data_stage_1__2520_, data_stage_1__2519_, data_stage_1__2518_, data_stage_1__2517_, data_stage_1__2516_, data_stage_1__2515_, data_stage_1__2514_, data_stage_1__2513_, data_stage_1__2512_, data_stage_1__2511_, data_stage_1__2510_, data_stage_1__2509_, data_stage_1__2508_, data_stage_1__2507_, data_stage_1__2506_, data_stage_1__2505_, data_stage_1__2504_, data_stage_1__2503_, data_stage_1__2502_, data_stage_1__2501_, data_stage_1__2500_, data_stage_1__2499_, data_stage_1__2498_, data_stage_1__2497_, data_stage_1__2496_, data_stage_1__2495_, data_stage_1__2494_, data_stage_1__2493_, data_stage_1__2492_, data_stage_1__2491_, data_stage_1__2490_, data_stage_1__2489_, data_stage_1__2488_, data_stage_1__2487_, data_stage_1__2486_, data_stage_1__2485_, data_stage_1__2484_, data_stage_1__2483_, data_stage_1__2482_, data_stage_1__2481_, data_stage_1__2480_, data_stage_1__2479_, data_stage_1__2478_, data_stage_1__2477_, data_stage_1__2476_, data_stage_1__2475_, data_stage_1__2474_, data_stage_1__2473_, data_stage_1__2472_, data_stage_1__2471_, data_stage_1__2470_, data_stage_1__2469_, data_stage_1__2468_, data_stage_1__2467_, data_stage_1__2466_, data_stage_1__2465_, data_stage_1__2464_, data_stage_1__2463_, data_stage_1__2462_, data_stage_1__2461_, data_stage_1__2460_, data_stage_1__2459_, data_stage_1__2458_, data_stage_1__2457_, data_stage_1__2456_, data_stage_1__2455_, data_stage_1__2454_, data_stage_1__2453_, data_stage_1__2452_, data_stage_1__2451_, data_stage_1__2450_, data_stage_1__2449_, data_stage_1__2448_, data_stage_1__2447_, data_stage_1__2446_, data_stage_1__2445_, data_stage_1__2444_, data_stage_1__2443_, data_stage_1__2442_, data_stage_1__2441_, data_stage_1__2440_, data_stage_1__2439_, data_stage_1__2438_, data_stage_1__2437_, data_stage_1__2436_, data_stage_1__2435_, data_stage_1__2434_, data_stage_1__2433_, data_stage_1__2432_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_20__swap_inst
  (
    .data_i(data_i[2687:2560]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__2687_, data_stage_1__2686_, data_stage_1__2685_, data_stage_1__2684_, data_stage_1__2683_, data_stage_1__2682_, data_stage_1__2681_, data_stage_1__2680_, data_stage_1__2679_, data_stage_1__2678_, data_stage_1__2677_, data_stage_1__2676_, data_stage_1__2675_, data_stage_1__2674_, data_stage_1__2673_, data_stage_1__2672_, data_stage_1__2671_, data_stage_1__2670_, data_stage_1__2669_, data_stage_1__2668_, data_stage_1__2667_, data_stage_1__2666_, data_stage_1__2665_, data_stage_1__2664_, data_stage_1__2663_, data_stage_1__2662_, data_stage_1__2661_, data_stage_1__2660_, data_stage_1__2659_, data_stage_1__2658_, data_stage_1__2657_, data_stage_1__2656_, data_stage_1__2655_, data_stage_1__2654_, data_stage_1__2653_, data_stage_1__2652_, data_stage_1__2651_, data_stage_1__2650_, data_stage_1__2649_, data_stage_1__2648_, data_stage_1__2647_, data_stage_1__2646_, data_stage_1__2645_, data_stage_1__2644_, data_stage_1__2643_, data_stage_1__2642_, data_stage_1__2641_, data_stage_1__2640_, data_stage_1__2639_, data_stage_1__2638_, data_stage_1__2637_, data_stage_1__2636_, data_stage_1__2635_, data_stage_1__2634_, data_stage_1__2633_, data_stage_1__2632_, data_stage_1__2631_, data_stage_1__2630_, data_stage_1__2629_, data_stage_1__2628_, data_stage_1__2627_, data_stage_1__2626_, data_stage_1__2625_, data_stage_1__2624_, data_stage_1__2623_, data_stage_1__2622_, data_stage_1__2621_, data_stage_1__2620_, data_stage_1__2619_, data_stage_1__2618_, data_stage_1__2617_, data_stage_1__2616_, data_stage_1__2615_, data_stage_1__2614_, data_stage_1__2613_, data_stage_1__2612_, data_stage_1__2611_, data_stage_1__2610_, data_stage_1__2609_, data_stage_1__2608_, data_stage_1__2607_, data_stage_1__2606_, data_stage_1__2605_, data_stage_1__2604_, data_stage_1__2603_, data_stage_1__2602_, data_stage_1__2601_, data_stage_1__2600_, data_stage_1__2599_, data_stage_1__2598_, data_stage_1__2597_, data_stage_1__2596_, data_stage_1__2595_, data_stage_1__2594_, data_stage_1__2593_, data_stage_1__2592_, data_stage_1__2591_, data_stage_1__2590_, data_stage_1__2589_, data_stage_1__2588_, data_stage_1__2587_, data_stage_1__2586_, data_stage_1__2585_, data_stage_1__2584_, data_stage_1__2583_, data_stage_1__2582_, data_stage_1__2581_, data_stage_1__2580_, data_stage_1__2579_, data_stage_1__2578_, data_stage_1__2577_, data_stage_1__2576_, data_stage_1__2575_, data_stage_1__2574_, data_stage_1__2573_, data_stage_1__2572_, data_stage_1__2571_, data_stage_1__2570_, data_stage_1__2569_, data_stage_1__2568_, data_stage_1__2567_, data_stage_1__2566_, data_stage_1__2565_, data_stage_1__2564_, data_stage_1__2563_, data_stage_1__2562_, data_stage_1__2561_, data_stage_1__2560_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_21__swap_inst
  (
    .data_i(data_i[2815:2688]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__2815_, data_stage_1__2814_, data_stage_1__2813_, data_stage_1__2812_, data_stage_1__2811_, data_stage_1__2810_, data_stage_1__2809_, data_stage_1__2808_, data_stage_1__2807_, data_stage_1__2806_, data_stage_1__2805_, data_stage_1__2804_, data_stage_1__2803_, data_stage_1__2802_, data_stage_1__2801_, data_stage_1__2800_, data_stage_1__2799_, data_stage_1__2798_, data_stage_1__2797_, data_stage_1__2796_, data_stage_1__2795_, data_stage_1__2794_, data_stage_1__2793_, data_stage_1__2792_, data_stage_1__2791_, data_stage_1__2790_, data_stage_1__2789_, data_stage_1__2788_, data_stage_1__2787_, data_stage_1__2786_, data_stage_1__2785_, data_stage_1__2784_, data_stage_1__2783_, data_stage_1__2782_, data_stage_1__2781_, data_stage_1__2780_, data_stage_1__2779_, data_stage_1__2778_, data_stage_1__2777_, data_stage_1__2776_, data_stage_1__2775_, data_stage_1__2774_, data_stage_1__2773_, data_stage_1__2772_, data_stage_1__2771_, data_stage_1__2770_, data_stage_1__2769_, data_stage_1__2768_, data_stage_1__2767_, data_stage_1__2766_, data_stage_1__2765_, data_stage_1__2764_, data_stage_1__2763_, data_stage_1__2762_, data_stage_1__2761_, data_stage_1__2760_, data_stage_1__2759_, data_stage_1__2758_, data_stage_1__2757_, data_stage_1__2756_, data_stage_1__2755_, data_stage_1__2754_, data_stage_1__2753_, data_stage_1__2752_, data_stage_1__2751_, data_stage_1__2750_, data_stage_1__2749_, data_stage_1__2748_, data_stage_1__2747_, data_stage_1__2746_, data_stage_1__2745_, data_stage_1__2744_, data_stage_1__2743_, data_stage_1__2742_, data_stage_1__2741_, data_stage_1__2740_, data_stage_1__2739_, data_stage_1__2738_, data_stage_1__2737_, data_stage_1__2736_, data_stage_1__2735_, data_stage_1__2734_, data_stage_1__2733_, data_stage_1__2732_, data_stage_1__2731_, data_stage_1__2730_, data_stage_1__2729_, data_stage_1__2728_, data_stage_1__2727_, data_stage_1__2726_, data_stage_1__2725_, data_stage_1__2724_, data_stage_1__2723_, data_stage_1__2722_, data_stage_1__2721_, data_stage_1__2720_, data_stage_1__2719_, data_stage_1__2718_, data_stage_1__2717_, data_stage_1__2716_, data_stage_1__2715_, data_stage_1__2714_, data_stage_1__2713_, data_stage_1__2712_, data_stage_1__2711_, data_stage_1__2710_, data_stage_1__2709_, data_stage_1__2708_, data_stage_1__2707_, data_stage_1__2706_, data_stage_1__2705_, data_stage_1__2704_, data_stage_1__2703_, data_stage_1__2702_, data_stage_1__2701_, data_stage_1__2700_, data_stage_1__2699_, data_stage_1__2698_, data_stage_1__2697_, data_stage_1__2696_, data_stage_1__2695_, data_stage_1__2694_, data_stage_1__2693_, data_stage_1__2692_, data_stage_1__2691_, data_stage_1__2690_, data_stage_1__2689_, data_stage_1__2688_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_22__swap_inst
  (
    .data_i(data_i[2943:2816]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__2943_, data_stage_1__2942_, data_stage_1__2941_, data_stage_1__2940_, data_stage_1__2939_, data_stage_1__2938_, data_stage_1__2937_, data_stage_1__2936_, data_stage_1__2935_, data_stage_1__2934_, data_stage_1__2933_, data_stage_1__2932_, data_stage_1__2931_, data_stage_1__2930_, data_stage_1__2929_, data_stage_1__2928_, data_stage_1__2927_, data_stage_1__2926_, data_stage_1__2925_, data_stage_1__2924_, data_stage_1__2923_, data_stage_1__2922_, data_stage_1__2921_, data_stage_1__2920_, data_stage_1__2919_, data_stage_1__2918_, data_stage_1__2917_, data_stage_1__2916_, data_stage_1__2915_, data_stage_1__2914_, data_stage_1__2913_, data_stage_1__2912_, data_stage_1__2911_, data_stage_1__2910_, data_stage_1__2909_, data_stage_1__2908_, data_stage_1__2907_, data_stage_1__2906_, data_stage_1__2905_, data_stage_1__2904_, data_stage_1__2903_, data_stage_1__2902_, data_stage_1__2901_, data_stage_1__2900_, data_stage_1__2899_, data_stage_1__2898_, data_stage_1__2897_, data_stage_1__2896_, data_stage_1__2895_, data_stage_1__2894_, data_stage_1__2893_, data_stage_1__2892_, data_stage_1__2891_, data_stage_1__2890_, data_stage_1__2889_, data_stage_1__2888_, data_stage_1__2887_, data_stage_1__2886_, data_stage_1__2885_, data_stage_1__2884_, data_stage_1__2883_, data_stage_1__2882_, data_stage_1__2881_, data_stage_1__2880_, data_stage_1__2879_, data_stage_1__2878_, data_stage_1__2877_, data_stage_1__2876_, data_stage_1__2875_, data_stage_1__2874_, data_stage_1__2873_, data_stage_1__2872_, data_stage_1__2871_, data_stage_1__2870_, data_stage_1__2869_, data_stage_1__2868_, data_stage_1__2867_, data_stage_1__2866_, data_stage_1__2865_, data_stage_1__2864_, data_stage_1__2863_, data_stage_1__2862_, data_stage_1__2861_, data_stage_1__2860_, data_stage_1__2859_, data_stage_1__2858_, data_stage_1__2857_, data_stage_1__2856_, data_stage_1__2855_, data_stage_1__2854_, data_stage_1__2853_, data_stage_1__2852_, data_stage_1__2851_, data_stage_1__2850_, data_stage_1__2849_, data_stage_1__2848_, data_stage_1__2847_, data_stage_1__2846_, data_stage_1__2845_, data_stage_1__2844_, data_stage_1__2843_, data_stage_1__2842_, data_stage_1__2841_, data_stage_1__2840_, data_stage_1__2839_, data_stage_1__2838_, data_stage_1__2837_, data_stage_1__2836_, data_stage_1__2835_, data_stage_1__2834_, data_stage_1__2833_, data_stage_1__2832_, data_stage_1__2831_, data_stage_1__2830_, data_stage_1__2829_, data_stage_1__2828_, data_stage_1__2827_, data_stage_1__2826_, data_stage_1__2825_, data_stage_1__2824_, data_stage_1__2823_, data_stage_1__2822_, data_stage_1__2821_, data_stage_1__2820_, data_stage_1__2819_, data_stage_1__2818_, data_stage_1__2817_, data_stage_1__2816_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_23__swap_inst
  (
    .data_i(data_i[3071:2944]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__3071_, data_stage_1__3070_, data_stage_1__3069_, data_stage_1__3068_, data_stage_1__3067_, data_stage_1__3066_, data_stage_1__3065_, data_stage_1__3064_, data_stage_1__3063_, data_stage_1__3062_, data_stage_1__3061_, data_stage_1__3060_, data_stage_1__3059_, data_stage_1__3058_, data_stage_1__3057_, data_stage_1__3056_, data_stage_1__3055_, data_stage_1__3054_, data_stage_1__3053_, data_stage_1__3052_, data_stage_1__3051_, data_stage_1__3050_, data_stage_1__3049_, data_stage_1__3048_, data_stage_1__3047_, data_stage_1__3046_, data_stage_1__3045_, data_stage_1__3044_, data_stage_1__3043_, data_stage_1__3042_, data_stage_1__3041_, data_stage_1__3040_, data_stage_1__3039_, data_stage_1__3038_, data_stage_1__3037_, data_stage_1__3036_, data_stage_1__3035_, data_stage_1__3034_, data_stage_1__3033_, data_stage_1__3032_, data_stage_1__3031_, data_stage_1__3030_, data_stage_1__3029_, data_stage_1__3028_, data_stage_1__3027_, data_stage_1__3026_, data_stage_1__3025_, data_stage_1__3024_, data_stage_1__3023_, data_stage_1__3022_, data_stage_1__3021_, data_stage_1__3020_, data_stage_1__3019_, data_stage_1__3018_, data_stage_1__3017_, data_stage_1__3016_, data_stage_1__3015_, data_stage_1__3014_, data_stage_1__3013_, data_stage_1__3012_, data_stage_1__3011_, data_stage_1__3010_, data_stage_1__3009_, data_stage_1__3008_, data_stage_1__3007_, data_stage_1__3006_, data_stage_1__3005_, data_stage_1__3004_, data_stage_1__3003_, data_stage_1__3002_, data_stage_1__3001_, data_stage_1__3000_, data_stage_1__2999_, data_stage_1__2998_, data_stage_1__2997_, data_stage_1__2996_, data_stage_1__2995_, data_stage_1__2994_, data_stage_1__2993_, data_stage_1__2992_, data_stage_1__2991_, data_stage_1__2990_, data_stage_1__2989_, data_stage_1__2988_, data_stage_1__2987_, data_stage_1__2986_, data_stage_1__2985_, data_stage_1__2984_, data_stage_1__2983_, data_stage_1__2982_, data_stage_1__2981_, data_stage_1__2980_, data_stage_1__2979_, data_stage_1__2978_, data_stage_1__2977_, data_stage_1__2976_, data_stage_1__2975_, data_stage_1__2974_, data_stage_1__2973_, data_stage_1__2972_, data_stage_1__2971_, data_stage_1__2970_, data_stage_1__2969_, data_stage_1__2968_, data_stage_1__2967_, data_stage_1__2966_, data_stage_1__2965_, data_stage_1__2964_, data_stage_1__2963_, data_stage_1__2962_, data_stage_1__2961_, data_stage_1__2960_, data_stage_1__2959_, data_stage_1__2958_, data_stage_1__2957_, data_stage_1__2956_, data_stage_1__2955_, data_stage_1__2954_, data_stage_1__2953_, data_stage_1__2952_, data_stage_1__2951_, data_stage_1__2950_, data_stage_1__2949_, data_stage_1__2948_, data_stage_1__2947_, data_stage_1__2946_, data_stage_1__2945_, data_stage_1__2944_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_24__swap_inst
  (
    .data_i(data_i[3199:3072]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__3199_, data_stage_1__3198_, data_stage_1__3197_, data_stage_1__3196_, data_stage_1__3195_, data_stage_1__3194_, data_stage_1__3193_, data_stage_1__3192_, data_stage_1__3191_, data_stage_1__3190_, data_stage_1__3189_, data_stage_1__3188_, data_stage_1__3187_, data_stage_1__3186_, data_stage_1__3185_, data_stage_1__3184_, data_stage_1__3183_, data_stage_1__3182_, data_stage_1__3181_, data_stage_1__3180_, data_stage_1__3179_, data_stage_1__3178_, data_stage_1__3177_, data_stage_1__3176_, data_stage_1__3175_, data_stage_1__3174_, data_stage_1__3173_, data_stage_1__3172_, data_stage_1__3171_, data_stage_1__3170_, data_stage_1__3169_, data_stage_1__3168_, data_stage_1__3167_, data_stage_1__3166_, data_stage_1__3165_, data_stage_1__3164_, data_stage_1__3163_, data_stage_1__3162_, data_stage_1__3161_, data_stage_1__3160_, data_stage_1__3159_, data_stage_1__3158_, data_stage_1__3157_, data_stage_1__3156_, data_stage_1__3155_, data_stage_1__3154_, data_stage_1__3153_, data_stage_1__3152_, data_stage_1__3151_, data_stage_1__3150_, data_stage_1__3149_, data_stage_1__3148_, data_stage_1__3147_, data_stage_1__3146_, data_stage_1__3145_, data_stage_1__3144_, data_stage_1__3143_, data_stage_1__3142_, data_stage_1__3141_, data_stage_1__3140_, data_stage_1__3139_, data_stage_1__3138_, data_stage_1__3137_, data_stage_1__3136_, data_stage_1__3135_, data_stage_1__3134_, data_stage_1__3133_, data_stage_1__3132_, data_stage_1__3131_, data_stage_1__3130_, data_stage_1__3129_, data_stage_1__3128_, data_stage_1__3127_, data_stage_1__3126_, data_stage_1__3125_, data_stage_1__3124_, data_stage_1__3123_, data_stage_1__3122_, data_stage_1__3121_, data_stage_1__3120_, data_stage_1__3119_, data_stage_1__3118_, data_stage_1__3117_, data_stage_1__3116_, data_stage_1__3115_, data_stage_1__3114_, data_stage_1__3113_, data_stage_1__3112_, data_stage_1__3111_, data_stage_1__3110_, data_stage_1__3109_, data_stage_1__3108_, data_stage_1__3107_, data_stage_1__3106_, data_stage_1__3105_, data_stage_1__3104_, data_stage_1__3103_, data_stage_1__3102_, data_stage_1__3101_, data_stage_1__3100_, data_stage_1__3099_, data_stage_1__3098_, data_stage_1__3097_, data_stage_1__3096_, data_stage_1__3095_, data_stage_1__3094_, data_stage_1__3093_, data_stage_1__3092_, data_stage_1__3091_, data_stage_1__3090_, data_stage_1__3089_, data_stage_1__3088_, data_stage_1__3087_, data_stage_1__3086_, data_stage_1__3085_, data_stage_1__3084_, data_stage_1__3083_, data_stage_1__3082_, data_stage_1__3081_, data_stage_1__3080_, data_stage_1__3079_, data_stage_1__3078_, data_stage_1__3077_, data_stage_1__3076_, data_stage_1__3075_, data_stage_1__3074_, data_stage_1__3073_, data_stage_1__3072_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_25__swap_inst
  (
    .data_i(data_i[3327:3200]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__3327_, data_stage_1__3326_, data_stage_1__3325_, data_stage_1__3324_, data_stage_1__3323_, data_stage_1__3322_, data_stage_1__3321_, data_stage_1__3320_, data_stage_1__3319_, data_stage_1__3318_, data_stage_1__3317_, data_stage_1__3316_, data_stage_1__3315_, data_stage_1__3314_, data_stage_1__3313_, data_stage_1__3312_, data_stage_1__3311_, data_stage_1__3310_, data_stage_1__3309_, data_stage_1__3308_, data_stage_1__3307_, data_stage_1__3306_, data_stage_1__3305_, data_stage_1__3304_, data_stage_1__3303_, data_stage_1__3302_, data_stage_1__3301_, data_stage_1__3300_, data_stage_1__3299_, data_stage_1__3298_, data_stage_1__3297_, data_stage_1__3296_, data_stage_1__3295_, data_stage_1__3294_, data_stage_1__3293_, data_stage_1__3292_, data_stage_1__3291_, data_stage_1__3290_, data_stage_1__3289_, data_stage_1__3288_, data_stage_1__3287_, data_stage_1__3286_, data_stage_1__3285_, data_stage_1__3284_, data_stage_1__3283_, data_stage_1__3282_, data_stage_1__3281_, data_stage_1__3280_, data_stage_1__3279_, data_stage_1__3278_, data_stage_1__3277_, data_stage_1__3276_, data_stage_1__3275_, data_stage_1__3274_, data_stage_1__3273_, data_stage_1__3272_, data_stage_1__3271_, data_stage_1__3270_, data_stage_1__3269_, data_stage_1__3268_, data_stage_1__3267_, data_stage_1__3266_, data_stage_1__3265_, data_stage_1__3264_, data_stage_1__3263_, data_stage_1__3262_, data_stage_1__3261_, data_stage_1__3260_, data_stage_1__3259_, data_stage_1__3258_, data_stage_1__3257_, data_stage_1__3256_, data_stage_1__3255_, data_stage_1__3254_, data_stage_1__3253_, data_stage_1__3252_, data_stage_1__3251_, data_stage_1__3250_, data_stage_1__3249_, data_stage_1__3248_, data_stage_1__3247_, data_stage_1__3246_, data_stage_1__3245_, data_stage_1__3244_, data_stage_1__3243_, data_stage_1__3242_, data_stage_1__3241_, data_stage_1__3240_, data_stage_1__3239_, data_stage_1__3238_, data_stage_1__3237_, data_stage_1__3236_, data_stage_1__3235_, data_stage_1__3234_, data_stage_1__3233_, data_stage_1__3232_, data_stage_1__3231_, data_stage_1__3230_, data_stage_1__3229_, data_stage_1__3228_, data_stage_1__3227_, data_stage_1__3226_, data_stage_1__3225_, data_stage_1__3224_, data_stage_1__3223_, data_stage_1__3222_, data_stage_1__3221_, data_stage_1__3220_, data_stage_1__3219_, data_stage_1__3218_, data_stage_1__3217_, data_stage_1__3216_, data_stage_1__3215_, data_stage_1__3214_, data_stage_1__3213_, data_stage_1__3212_, data_stage_1__3211_, data_stage_1__3210_, data_stage_1__3209_, data_stage_1__3208_, data_stage_1__3207_, data_stage_1__3206_, data_stage_1__3205_, data_stage_1__3204_, data_stage_1__3203_, data_stage_1__3202_, data_stage_1__3201_, data_stage_1__3200_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_26__swap_inst
  (
    .data_i(data_i[3455:3328]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__3455_, data_stage_1__3454_, data_stage_1__3453_, data_stage_1__3452_, data_stage_1__3451_, data_stage_1__3450_, data_stage_1__3449_, data_stage_1__3448_, data_stage_1__3447_, data_stage_1__3446_, data_stage_1__3445_, data_stage_1__3444_, data_stage_1__3443_, data_stage_1__3442_, data_stage_1__3441_, data_stage_1__3440_, data_stage_1__3439_, data_stage_1__3438_, data_stage_1__3437_, data_stage_1__3436_, data_stage_1__3435_, data_stage_1__3434_, data_stage_1__3433_, data_stage_1__3432_, data_stage_1__3431_, data_stage_1__3430_, data_stage_1__3429_, data_stage_1__3428_, data_stage_1__3427_, data_stage_1__3426_, data_stage_1__3425_, data_stage_1__3424_, data_stage_1__3423_, data_stage_1__3422_, data_stage_1__3421_, data_stage_1__3420_, data_stage_1__3419_, data_stage_1__3418_, data_stage_1__3417_, data_stage_1__3416_, data_stage_1__3415_, data_stage_1__3414_, data_stage_1__3413_, data_stage_1__3412_, data_stage_1__3411_, data_stage_1__3410_, data_stage_1__3409_, data_stage_1__3408_, data_stage_1__3407_, data_stage_1__3406_, data_stage_1__3405_, data_stage_1__3404_, data_stage_1__3403_, data_stage_1__3402_, data_stage_1__3401_, data_stage_1__3400_, data_stage_1__3399_, data_stage_1__3398_, data_stage_1__3397_, data_stage_1__3396_, data_stage_1__3395_, data_stage_1__3394_, data_stage_1__3393_, data_stage_1__3392_, data_stage_1__3391_, data_stage_1__3390_, data_stage_1__3389_, data_stage_1__3388_, data_stage_1__3387_, data_stage_1__3386_, data_stage_1__3385_, data_stage_1__3384_, data_stage_1__3383_, data_stage_1__3382_, data_stage_1__3381_, data_stage_1__3380_, data_stage_1__3379_, data_stage_1__3378_, data_stage_1__3377_, data_stage_1__3376_, data_stage_1__3375_, data_stage_1__3374_, data_stage_1__3373_, data_stage_1__3372_, data_stage_1__3371_, data_stage_1__3370_, data_stage_1__3369_, data_stage_1__3368_, data_stage_1__3367_, data_stage_1__3366_, data_stage_1__3365_, data_stage_1__3364_, data_stage_1__3363_, data_stage_1__3362_, data_stage_1__3361_, data_stage_1__3360_, data_stage_1__3359_, data_stage_1__3358_, data_stage_1__3357_, data_stage_1__3356_, data_stage_1__3355_, data_stage_1__3354_, data_stage_1__3353_, data_stage_1__3352_, data_stage_1__3351_, data_stage_1__3350_, data_stage_1__3349_, data_stage_1__3348_, data_stage_1__3347_, data_stage_1__3346_, data_stage_1__3345_, data_stage_1__3344_, data_stage_1__3343_, data_stage_1__3342_, data_stage_1__3341_, data_stage_1__3340_, data_stage_1__3339_, data_stage_1__3338_, data_stage_1__3337_, data_stage_1__3336_, data_stage_1__3335_, data_stage_1__3334_, data_stage_1__3333_, data_stage_1__3332_, data_stage_1__3331_, data_stage_1__3330_, data_stage_1__3329_, data_stage_1__3328_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_27__swap_inst
  (
    .data_i(data_i[3583:3456]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__3583_, data_stage_1__3582_, data_stage_1__3581_, data_stage_1__3580_, data_stage_1__3579_, data_stage_1__3578_, data_stage_1__3577_, data_stage_1__3576_, data_stage_1__3575_, data_stage_1__3574_, data_stage_1__3573_, data_stage_1__3572_, data_stage_1__3571_, data_stage_1__3570_, data_stage_1__3569_, data_stage_1__3568_, data_stage_1__3567_, data_stage_1__3566_, data_stage_1__3565_, data_stage_1__3564_, data_stage_1__3563_, data_stage_1__3562_, data_stage_1__3561_, data_stage_1__3560_, data_stage_1__3559_, data_stage_1__3558_, data_stage_1__3557_, data_stage_1__3556_, data_stage_1__3555_, data_stage_1__3554_, data_stage_1__3553_, data_stage_1__3552_, data_stage_1__3551_, data_stage_1__3550_, data_stage_1__3549_, data_stage_1__3548_, data_stage_1__3547_, data_stage_1__3546_, data_stage_1__3545_, data_stage_1__3544_, data_stage_1__3543_, data_stage_1__3542_, data_stage_1__3541_, data_stage_1__3540_, data_stage_1__3539_, data_stage_1__3538_, data_stage_1__3537_, data_stage_1__3536_, data_stage_1__3535_, data_stage_1__3534_, data_stage_1__3533_, data_stage_1__3532_, data_stage_1__3531_, data_stage_1__3530_, data_stage_1__3529_, data_stage_1__3528_, data_stage_1__3527_, data_stage_1__3526_, data_stage_1__3525_, data_stage_1__3524_, data_stage_1__3523_, data_stage_1__3522_, data_stage_1__3521_, data_stage_1__3520_, data_stage_1__3519_, data_stage_1__3518_, data_stage_1__3517_, data_stage_1__3516_, data_stage_1__3515_, data_stage_1__3514_, data_stage_1__3513_, data_stage_1__3512_, data_stage_1__3511_, data_stage_1__3510_, data_stage_1__3509_, data_stage_1__3508_, data_stage_1__3507_, data_stage_1__3506_, data_stage_1__3505_, data_stage_1__3504_, data_stage_1__3503_, data_stage_1__3502_, data_stage_1__3501_, data_stage_1__3500_, data_stage_1__3499_, data_stage_1__3498_, data_stage_1__3497_, data_stage_1__3496_, data_stage_1__3495_, data_stage_1__3494_, data_stage_1__3493_, data_stage_1__3492_, data_stage_1__3491_, data_stage_1__3490_, data_stage_1__3489_, data_stage_1__3488_, data_stage_1__3487_, data_stage_1__3486_, data_stage_1__3485_, data_stage_1__3484_, data_stage_1__3483_, data_stage_1__3482_, data_stage_1__3481_, data_stage_1__3480_, data_stage_1__3479_, data_stage_1__3478_, data_stage_1__3477_, data_stage_1__3476_, data_stage_1__3475_, data_stage_1__3474_, data_stage_1__3473_, data_stage_1__3472_, data_stage_1__3471_, data_stage_1__3470_, data_stage_1__3469_, data_stage_1__3468_, data_stage_1__3467_, data_stage_1__3466_, data_stage_1__3465_, data_stage_1__3464_, data_stage_1__3463_, data_stage_1__3462_, data_stage_1__3461_, data_stage_1__3460_, data_stage_1__3459_, data_stage_1__3458_, data_stage_1__3457_, data_stage_1__3456_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_28__swap_inst
  (
    .data_i(data_i[3711:3584]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__3711_, data_stage_1__3710_, data_stage_1__3709_, data_stage_1__3708_, data_stage_1__3707_, data_stage_1__3706_, data_stage_1__3705_, data_stage_1__3704_, data_stage_1__3703_, data_stage_1__3702_, data_stage_1__3701_, data_stage_1__3700_, data_stage_1__3699_, data_stage_1__3698_, data_stage_1__3697_, data_stage_1__3696_, data_stage_1__3695_, data_stage_1__3694_, data_stage_1__3693_, data_stage_1__3692_, data_stage_1__3691_, data_stage_1__3690_, data_stage_1__3689_, data_stage_1__3688_, data_stage_1__3687_, data_stage_1__3686_, data_stage_1__3685_, data_stage_1__3684_, data_stage_1__3683_, data_stage_1__3682_, data_stage_1__3681_, data_stage_1__3680_, data_stage_1__3679_, data_stage_1__3678_, data_stage_1__3677_, data_stage_1__3676_, data_stage_1__3675_, data_stage_1__3674_, data_stage_1__3673_, data_stage_1__3672_, data_stage_1__3671_, data_stage_1__3670_, data_stage_1__3669_, data_stage_1__3668_, data_stage_1__3667_, data_stage_1__3666_, data_stage_1__3665_, data_stage_1__3664_, data_stage_1__3663_, data_stage_1__3662_, data_stage_1__3661_, data_stage_1__3660_, data_stage_1__3659_, data_stage_1__3658_, data_stage_1__3657_, data_stage_1__3656_, data_stage_1__3655_, data_stage_1__3654_, data_stage_1__3653_, data_stage_1__3652_, data_stage_1__3651_, data_stage_1__3650_, data_stage_1__3649_, data_stage_1__3648_, data_stage_1__3647_, data_stage_1__3646_, data_stage_1__3645_, data_stage_1__3644_, data_stage_1__3643_, data_stage_1__3642_, data_stage_1__3641_, data_stage_1__3640_, data_stage_1__3639_, data_stage_1__3638_, data_stage_1__3637_, data_stage_1__3636_, data_stage_1__3635_, data_stage_1__3634_, data_stage_1__3633_, data_stage_1__3632_, data_stage_1__3631_, data_stage_1__3630_, data_stage_1__3629_, data_stage_1__3628_, data_stage_1__3627_, data_stage_1__3626_, data_stage_1__3625_, data_stage_1__3624_, data_stage_1__3623_, data_stage_1__3622_, data_stage_1__3621_, data_stage_1__3620_, data_stage_1__3619_, data_stage_1__3618_, data_stage_1__3617_, data_stage_1__3616_, data_stage_1__3615_, data_stage_1__3614_, data_stage_1__3613_, data_stage_1__3612_, data_stage_1__3611_, data_stage_1__3610_, data_stage_1__3609_, data_stage_1__3608_, data_stage_1__3607_, data_stage_1__3606_, data_stage_1__3605_, data_stage_1__3604_, data_stage_1__3603_, data_stage_1__3602_, data_stage_1__3601_, data_stage_1__3600_, data_stage_1__3599_, data_stage_1__3598_, data_stage_1__3597_, data_stage_1__3596_, data_stage_1__3595_, data_stage_1__3594_, data_stage_1__3593_, data_stage_1__3592_, data_stage_1__3591_, data_stage_1__3590_, data_stage_1__3589_, data_stage_1__3588_, data_stage_1__3587_, data_stage_1__3586_, data_stage_1__3585_, data_stage_1__3584_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_29__swap_inst
  (
    .data_i(data_i[3839:3712]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__3839_, data_stage_1__3838_, data_stage_1__3837_, data_stage_1__3836_, data_stage_1__3835_, data_stage_1__3834_, data_stage_1__3833_, data_stage_1__3832_, data_stage_1__3831_, data_stage_1__3830_, data_stage_1__3829_, data_stage_1__3828_, data_stage_1__3827_, data_stage_1__3826_, data_stage_1__3825_, data_stage_1__3824_, data_stage_1__3823_, data_stage_1__3822_, data_stage_1__3821_, data_stage_1__3820_, data_stage_1__3819_, data_stage_1__3818_, data_stage_1__3817_, data_stage_1__3816_, data_stage_1__3815_, data_stage_1__3814_, data_stage_1__3813_, data_stage_1__3812_, data_stage_1__3811_, data_stage_1__3810_, data_stage_1__3809_, data_stage_1__3808_, data_stage_1__3807_, data_stage_1__3806_, data_stage_1__3805_, data_stage_1__3804_, data_stage_1__3803_, data_stage_1__3802_, data_stage_1__3801_, data_stage_1__3800_, data_stage_1__3799_, data_stage_1__3798_, data_stage_1__3797_, data_stage_1__3796_, data_stage_1__3795_, data_stage_1__3794_, data_stage_1__3793_, data_stage_1__3792_, data_stage_1__3791_, data_stage_1__3790_, data_stage_1__3789_, data_stage_1__3788_, data_stage_1__3787_, data_stage_1__3786_, data_stage_1__3785_, data_stage_1__3784_, data_stage_1__3783_, data_stage_1__3782_, data_stage_1__3781_, data_stage_1__3780_, data_stage_1__3779_, data_stage_1__3778_, data_stage_1__3777_, data_stage_1__3776_, data_stage_1__3775_, data_stage_1__3774_, data_stage_1__3773_, data_stage_1__3772_, data_stage_1__3771_, data_stage_1__3770_, data_stage_1__3769_, data_stage_1__3768_, data_stage_1__3767_, data_stage_1__3766_, data_stage_1__3765_, data_stage_1__3764_, data_stage_1__3763_, data_stage_1__3762_, data_stage_1__3761_, data_stage_1__3760_, data_stage_1__3759_, data_stage_1__3758_, data_stage_1__3757_, data_stage_1__3756_, data_stage_1__3755_, data_stage_1__3754_, data_stage_1__3753_, data_stage_1__3752_, data_stage_1__3751_, data_stage_1__3750_, data_stage_1__3749_, data_stage_1__3748_, data_stage_1__3747_, data_stage_1__3746_, data_stage_1__3745_, data_stage_1__3744_, data_stage_1__3743_, data_stage_1__3742_, data_stage_1__3741_, data_stage_1__3740_, data_stage_1__3739_, data_stage_1__3738_, data_stage_1__3737_, data_stage_1__3736_, data_stage_1__3735_, data_stage_1__3734_, data_stage_1__3733_, data_stage_1__3732_, data_stage_1__3731_, data_stage_1__3730_, data_stage_1__3729_, data_stage_1__3728_, data_stage_1__3727_, data_stage_1__3726_, data_stage_1__3725_, data_stage_1__3724_, data_stage_1__3723_, data_stage_1__3722_, data_stage_1__3721_, data_stage_1__3720_, data_stage_1__3719_, data_stage_1__3718_, data_stage_1__3717_, data_stage_1__3716_, data_stage_1__3715_, data_stage_1__3714_, data_stage_1__3713_, data_stage_1__3712_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_30__swap_inst
  (
    .data_i(data_i[3967:3840]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__3967_, data_stage_1__3966_, data_stage_1__3965_, data_stage_1__3964_, data_stage_1__3963_, data_stage_1__3962_, data_stage_1__3961_, data_stage_1__3960_, data_stage_1__3959_, data_stage_1__3958_, data_stage_1__3957_, data_stage_1__3956_, data_stage_1__3955_, data_stage_1__3954_, data_stage_1__3953_, data_stage_1__3952_, data_stage_1__3951_, data_stage_1__3950_, data_stage_1__3949_, data_stage_1__3948_, data_stage_1__3947_, data_stage_1__3946_, data_stage_1__3945_, data_stage_1__3944_, data_stage_1__3943_, data_stage_1__3942_, data_stage_1__3941_, data_stage_1__3940_, data_stage_1__3939_, data_stage_1__3938_, data_stage_1__3937_, data_stage_1__3936_, data_stage_1__3935_, data_stage_1__3934_, data_stage_1__3933_, data_stage_1__3932_, data_stage_1__3931_, data_stage_1__3930_, data_stage_1__3929_, data_stage_1__3928_, data_stage_1__3927_, data_stage_1__3926_, data_stage_1__3925_, data_stage_1__3924_, data_stage_1__3923_, data_stage_1__3922_, data_stage_1__3921_, data_stage_1__3920_, data_stage_1__3919_, data_stage_1__3918_, data_stage_1__3917_, data_stage_1__3916_, data_stage_1__3915_, data_stage_1__3914_, data_stage_1__3913_, data_stage_1__3912_, data_stage_1__3911_, data_stage_1__3910_, data_stage_1__3909_, data_stage_1__3908_, data_stage_1__3907_, data_stage_1__3906_, data_stage_1__3905_, data_stage_1__3904_, data_stage_1__3903_, data_stage_1__3902_, data_stage_1__3901_, data_stage_1__3900_, data_stage_1__3899_, data_stage_1__3898_, data_stage_1__3897_, data_stage_1__3896_, data_stage_1__3895_, data_stage_1__3894_, data_stage_1__3893_, data_stage_1__3892_, data_stage_1__3891_, data_stage_1__3890_, data_stage_1__3889_, data_stage_1__3888_, data_stage_1__3887_, data_stage_1__3886_, data_stage_1__3885_, data_stage_1__3884_, data_stage_1__3883_, data_stage_1__3882_, data_stage_1__3881_, data_stage_1__3880_, data_stage_1__3879_, data_stage_1__3878_, data_stage_1__3877_, data_stage_1__3876_, data_stage_1__3875_, data_stage_1__3874_, data_stage_1__3873_, data_stage_1__3872_, data_stage_1__3871_, data_stage_1__3870_, data_stage_1__3869_, data_stage_1__3868_, data_stage_1__3867_, data_stage_1__3866_, data_stage_1__3865_, data_stage_1__3864_, data_stage_1__3863_, data_stage_1__3862_, data_stage_1__3861_, data_stage_1__3860_, data_stage_1__3859_, data_stage_1__3858_, data_stage_1__3857_, data_stage_1__3856_, data_stage_1__3855_, data_stage_1__3854_, data_stage_1__3853_, data_stage_1__3852_, data_stage_1__3851_, data_stage_1__3850_, data_stage_1__3849_, data_stage_1__3848_, data_stage_1__3847_, data_stage_1__3846_, data_stage_1__3845_, data_stage_1__3844_, data_stage_1__3843_, data_stage_1__3842_, data_stage_1__3841_, data_stage_1__3840_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_31__swap_inst
  (
    .data_i(data_i[4095:3968]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__4095_, data_stage_1__4094_, data_stage_1__4093_, data_stage_1__4092_, data_stage_1__4091_, data_stage_1__4090_, data_stage_1__4089_, data_stage_1__4088_, data_stage_1__4087_, data_stage_1__4086_, data_stage_1__4085_, data_stage_1__4084_, data_stage_1__4083_, data_stage_1__4082_, data_stage_1__4081_, data_stage_1__4080_, data_stage_1__4079_, data_stage_1__4078_, data_stage_1__4077_, data_stage_1__4076_, data_stage_1__4075_, data_stage_1__4074_, data_stage_1__4073_, data_stage_1__4072_, data_stage_1__4071_, data_stage_1__4070_, data_stage_1__4069_, data_stage_1__4068_, data_stage_1__4067_, data_stage_1__4066_, data_stage_1__4065_, data_stage_1__4064_, data_stage_1__4063_, data_stage_1__4062_, data_stage_1__4061_, data_stage_1__4060_, data_stage_1__4059_, data_stage_1__4058_, data_stage_1__4057_, data_stage_1__4056_, data_stage_1__4055_, data_stage_1__4054_, data_stage_1__4053_, data_stage_1__4052_, data_stage_1__4051_, data_stage_1__4050_, data_stage_1__4049_, data_stage_1__4048_, data_stage_1__4047_, data_stage_1__4046_, data_stage_1__4045_, data_stage_1__4044_, data_stage_1__4043_, data_stage_1__4042_, data_stage_1__4041_, data_stage_1__4040_, data_stage_1__4039_, data_stage_1__4038_, data_stage_1__4037_, data_stage_1__4036_, data_stage_1__4035_, data_stage_1__4034_, data_stage_1__4033_, data_stage_1__4032_, data_stage_1__4031_, data_stage_1__4030_, data_stage_1__4029_, data_stage_1__4028_, data_stage_1__4027_, data_stage_1__4026_, data_stage_1__4025_, data_stage_1__4024_, data_stage_1__4023_, data_stage_1__4022_, data_stage_1__4021_, data_stage_1__4020_, data_stage_1__4019_, data_stage_1__4018_, data_stage_1__4017_, data_stage_1__4016_, data_stage_1__4015_, data_stage_1__4014_, data_stage_1__4013_, data_stage_1__4012_, data_stage_1__4011_, data_stage_1__4010_, data_stage_1__4009_, data_stage_1__4008_, data_stage_1__4007_, data_stage_1__4006_, data_stage_1__4005_, data_stage_1__4004_, data_stage_1__4003_, data_stage_1__4002_, data_stage_1__4001_, data_stage_1__4000_, data_stage_1__3999_, data_stage_1__3998_, data_stage_1__3997_, data_stage_1__3996_, data_stage_1__3995_, data_stage_1__3994_, data_stage_1__3993_, data_stage_1__3992_, data_stage_1__3991_, data_stage_1__3990_, data_stage_1__3989_, data_stage_1__3988_, data_stage_1__3987_, data_stage_1__3986_, data_stage_1__3985_, data_stage_1__3984_, data_stage_1__3983_, data_stage_1__3982_, data_stage_1__3981_, data_stage_1__3980_, data_stage_1__3979_, data_stage_1__3978_, data_stage_1__3977_, data_stage_1__3976_, data_stage_1__3975_, data_stage_1__3974_, data_stage_1__3973_, data_stage_1__3972_, data_stage_1__3971_, data_stage_1__3970_, data_stage_1__3969_, data_stage_1__3968_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_0__swap_inst
  (
    .data_i({ data_stage_1__255_, data_stage_1__254_, data_stage_1__253_, data_stage_1__252_, data_stage_1__251_, data_stage_1__250_, data_stage_1__249_, data_stage_1__248_, data_stage_1__247_, data_stage_1__246_, data_stage_1__245_, data_stage_1__244_, data_stage_1__243_, data_stage_1__242_, data_stage_1__241_, data_stage_1__240_, data_stage_1__239_, data_stage_1__238_, data_stage_1__237_, data_stage_1__236_, data_stage_1__235_, data_stage_1__234_, data_stage_1__233_, data_stage_1__232_, data_stage_1__231_, data_stage_1__230_, data_stage_1__229_, data_stage_1__228_, data_stage_1__227_, data_stage_1__226_, data_stage_1__225_, data_stage_1__224_, data_stage_1__223_, data_stage_1__222_, data_stage_1__221_, data_stage_1__220_, data_stage_1__219_, data_stage_1__218_, data_stage_1__217_, data_stage_1__216_, data_stage_1__215_, data_stage_1__214_, data_stage_1__213_, data_stage_1__212_, data_stage_1__211_, data_stage_1__210_, data_stage_1__209_, data_stage_1__208_, data_stage_1__207_, data_stage_1__206_, data_stage_1__205_, data_stage_1__204_, data_stage_1__203_, data_stage_1__202_, data_stage_1__201_, data_stage_1__200_, data_stage_1__199_, data_stage_1__198_, data_stage_1__197_, data_stage_1__196_, data_stage_1__195_, data_stage_1__194_, data_stage_1__193_, data_stage_1__192_, data_stage_1__191_, data_stage_1__190_, data_stage_1__189_, data_stage_1__188_, data_stage_1__187_, data_stage_1__186_, data_stage_1__185_, data_stage_1__184_, data_stage_1__183_, data_stage_1__182_, data_stage_1__181_, data_stage_1__180_, data_stage_1__179_, data_stage_1__178_, data_stage_1__177_, data_stage_1__176_, data_stage_1__175_, data_stage_1__174_, data_stage_1__173_, data_stage_1__172_, data_stage_1__171_, data_stage_1__170_, data_stage_1__169_, data_stage_1__168_, data_stage_1__167_, data_stage_1__166_, data_stage_1__165_, data_stage_1__164_, data_stage_1__163_, data_stage_1__162_, data_stage_1__161_, data_stage_1__160_, data_stage_1__159_, data_stage_1__158_, data_stage_1__157_, data_stage_1__156_, data_stage_1__155_, data_stage_1__154_, data_stage_1__153_, data_stage_1__152_, data_stage_1__151_, data_stage_1__150_, data_stage_1__149_, data_stage_1__148_, data_stage_1__147_, data_stage_1__146_, data_stage_1__145_, data_stage_1__144_, data_stage_1__143_, data_stage_1__142_, data_stage_1__141_, data_stage_1__140_, data_stage_1__139_, data_stage_1__138_, data_stage_1__137_, data_stage_1__136_, data_stage_1__135_, data_stage_1__134_, data_stage_1__133_, data_stage_1__132_, data_stage_1__131_, data_stage_1__130_, data_stage_1__129_, data_stage_1__128_, data_stage_1__127_, data_stage_1__126_, data_stage_1__125_, data_stage_1__124_, data_stage_1__123_, data_stage_1__122_, data_stage_1__121_, data_stage_1__120_, data_stage_1__119_, data_stage_1__118_, data_stage_1__117_, data_stage_1__116_, data_stage_1__115_, data_stage_1__114_, data_stage_1__113_, data_stage_1__112_, data_stage_1__111_, data_stage_1__110_, data_stage_1__109_, data_stage_1__108_, data_stage_1__107_, data_stage_1__106_, data_stage_1__105_, data_stage_1__104_, data_stage_1__103_, data_stage_1__102_, data_stage_1__101_, data_stage_1__100_, data_stage_1__99_, data_stage_1__98_, data_stage_1__97_, data_stage_1__96_, data_stage_1__95_, data_stage_1__94_, data_stage_1__93_, data_stage_1__92_, data_stage_1__91_, data_stage_1__90_, data_stage_1__89_, data_stage_1__88_, data_stage_1__87_, data_stage_1__86_, data_stage_1__85_, data_stage_1__84_, data_stage_1__83_, data_stage_1__82_, data_stage_1__81_, data_stage_1__80_, data_stage_1__79_, data_stage_1__78_, data_stage_1__77_, data_stage_1__76_, data_stage_1__75_, data_stage_1__74_, data_stage_1__73_, data_stage_1__72_, data_stage_1__71_, data_stage_1__70_, data_stage_1__69_, data_stage_1__68_, data_stage_1__67_, data_stage_1__66_, data_stage_1__65_, data_stage_1__64_, data_stage_1__63_, data_stage_1__62_, data_stage_1__61_, data_stage_1__60_, data_stage_1__59_, data_stage_1__58_, data_stage_1__57_, data_stage_1__56_, data_stage_1__55_, data_stage_1__54_, data_stage_1__53_, data_stage_1__52_, data_stage_1__51_, data_stage_1__50_, data_stage_1__49_, data_stage_1__48_, data_stage_1__47_, data_stage_1__46_, data_stage_1__45_, data_stage_1__44_, data_stage_1__43_, data_stage_1__42_, data_stage_1__41_, data_stage_1__40_, data_stage_1__39_, data_stage_1__38_, data_stage_1__37_, data_stage_1__36_, data_stage_1__35_, data_stage_1__34_, data_stage_1__33_, data_stage_1__32_, data_stage_1__31_, data_stage_1__30_, data_stage_1__29_, data_stage_1__28_, data_stage_1__27_, data_stage_1__26_, data_stage_1__25_, data_stage_1__24_, data_stage_1__23_, data_stage_1__22_, data_stage_1__21_, data_stage_1__20_, data_stage_1__19_, data_stage_1__18_, data_stage_1__17_, data_stage_1__16_, data_stage_1__15_, data_stage_1__14_, data_stage_1__13_, data_stage_1__12_, data_stage_1__11_, data_stage_1__10_, data_stage_1__9_, data_stage_1__8_, data_stage_1__7_, data_stage_1__6_, data_stage_1__5_, data_stage_1__4_, data_stage_1__3_, data_stage_1__2_, data_stage_1__1_, data_stage_1__0_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__255_, data_stage_2__254_, data_stage_2__253_, data_stage_2__252_, data_stage_2__251_, data_stage_2__250_, data_stage_2__249_, data_stage_2__248_, data_stage_2__247_, data_stage_2__246_, data_stage_2__245_, data_stage_2__244_, data_stage_2__243_, data_stage_2__242_, data_stage_2__241_, data_stage_2__240_, data_stage_2__239_, data_stage_2__238_, data_stage_2__237_, data_stage_2__236_, data_stage_2__235_, data_stage_2__234_, data_stage_2__233_, data_stage_2__232_, data_stage_2__231_, data_stage_2__230_, data_stage_2__229_, data_stage_2__228_, data_stage_2__227_, data_stage_2__226_, data_stage_2__225_, data_stage_2__224_, data_stage_2__223_, data_stage_2__222_, data_stage_2__221_, data_stage_2__220_, data_stage_2__219_, data_stage_2__218_, data_stage_2__217_, data_stage_2__216_, data_stage_2__215_, data_stage_2__214_, data_stage_2__213_, data_stage_2__212_, data_stage_2__211_, data_stage_2__210_, data_stage_2__209_, data_stage_2__208_, data_stage_2__207_, data_stage_2__206_, data_stage_2__205_, data_stage_2__204_, data_stage_2__203_, data_stage_2__202_, data_stage_2__201_, data_stage_2__200_, data_stage_2__199_, data_stage_2__198_, data_stage_2__197_, data_stage_2__196_, data_stage_2__195_, data_stage_2__194_, data_stage_2__193_, data_stage_2__192_, data_stage_2__191_, data_stage_2__190_, data_stage_2__189_, data_stage_2__188_, data_stage_2__187_, data_stage_2__186_, data_stage_2__185_, data_stage_2__184_, data_stage_2__183_, data_stage_2__182_, data_stage_2__181_, data_stage_2__180_, data_stage_2__179_, data_stage_2__178_, data_stage_2__177_, data_stage_2__176_, data_stage_2__175_, data_stage_2__174_, data_stage_2__173_, data_stage_2__172_, data_stage_2__171_, data_stage_2__170_, data_stage_2__169_, data_stage_2__168_, data_stage_2__167_, data_stage_2__166_, data_stage_2__165_, data_stage_2__164_, data_stage_2__163_, data_stage_2__162_, data_stage_2__161_, data_stage_2__160_, data_stage_2__159_, data_stage_2__158_, data_stage_2__157_, data_stage_2__156_, data_stage_2__155_, data_stage_2__154_, data_stage_2__153_, data_stage_2__152_, data_stage_2__151_, data_stage_2__150_, data_stage_2__149_, data_stage_2__148_, data_stage_2__147_, data_stage_2__146_, data_stage_2__145_, data_stage_2__144_, data_stage_2__143_, data_stage_2__142_, data_stage_2__141_, data_stage_2__140_, data_stage_2__139_, data_stage_2__138_, data_stage_2__137_, data_stage_2__136_, data_stage_2__135_, data_stage_2__134_, data_stage_2__133_, data_stage_2__132_, data_stage_2__131_, data_stage_2__130_, data_stage_2__129_, data_stage_2__128_, data_stage_2__127_, data_stage_2__126_, data_stage_2__125_, data_stage_2__124_, data_stage_2__123_, data_stage_2__122_, data_stage_2__121_, data_stage_2__120_, data_stage_2__119_, data_stage_2__118_, data_stage_2__117_, data_stage_2__116_, data_stage_2__115_, data_stage_2__114_, data_stage_2__113_, data_stage_2__112_, data_stage_2__111_, data_stage_2__110_, data_stage_2__109_, data_stage_2__108_, data_stage_2__107_, data_stage_2__106_, data_stage_2__105_, data_stage_2__104_, data_stage_2__103_, data_stage_2__102_, data_stage_2__101_, data_stage_2__100_, data_stage_2__99_, data_stage_2__98_, data_stage_2__97_, data_stage_2__96_, data_stage_2__95_, data_stage_2__94_, data_stage_2__93_, data_stage_2__92_, data_stage_2__91_, data_stage_2__90_, data_stage_2__89_, data_stage_2__88_, data_stage_2__87_, data_stage_2__86_, data_stage_2__85_, data_stage_2__84_, data_stage_2__83_, data_stage_2__82_, data_stage_2__81_, data_stage_2__80_, data_stage_2__79_, data_stage_2__78_, data_stage_2__77_, data_stage_2__76_, data_stage_2__75_, data_stage_2__74_, data_stage_2__73_, data_stage_2__72_, data_stage_2__71_, data_stage_2__70_, data_stage_2__69_, data_stage_2__68_, data_stage_2__67_, data_stage_2__66_, data_stage_2__65_, data_stage_2__64_, data_stage_2__63_, data_stage_2__62_, data_stage_2__61_, data_stage_2__60_, data_stage_2__59_, data_stage_2__58_, data_stage_2__57_, data_stage_2__56_, data_stage_2__55_, data_stage_2__54_, data_stage_2__53_, data_stage_2__52_, data_stage_2__51_, data_stage_2__50_, data_stage_2__49_, data_stage_2__48_, data_stage_2__47_, data_stage_2__46_, data_stage_2__45_, data_stage_2__44_, data_stage_2__43_, data_stage_2__42_, data_stage_2__41_, data_stage_2__40_, data_stage_2__39_, data_stage_2__38_, data_stage_2__37_, data_stage_2__36_, data_stage_2__35_, data_stage_2__34_, data_stage_2__33_, data_stage_2__32_, data_stage_2__31_, data_stage_2__30_, data_stage_2__29_, data_stage_2__28_, data_stage_2__27_, data_stage_2__26_, data_stage_2__25_, data_stage_2__24_, data_stage_2__23_, data_stage_2__22_, data_stage_2__21_, data_stage_2__20_, data_stage_2__19_, data_stage_2__18_, data_stage_2__17_, data_stage_2__16_, data_stage_2__15_, data_stage_2__14_, data_stage_2__13_, data_stage_2__12_, data_stage_2__11_, data_stage_2__10_, data_stage_2__9_, data_stage_2__8_, data_stage_2__7_, data_stage_2__6_, data_stage_2__5_, data_stage_2__4_, data_stage_2__3_, data_stage_2__2_, data_stage_2__1_, data_stage_2__0_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_1__swap_inst
  (
    .data_i({ data_stage_1__511_, data_stage_1__510_, data_stage_1__509_, data_stage_1__508_, data_stage_1__507_, data_stage_1__506_, data_stage_1__505_, data_stage_1__504_, data_stage_1__503_, data_stage_1__502_, data_stage_1__501_, data_stage_1__500_, data_stage_1__499_, data_stage_1__498_, data_stage_1__497_, data_stage_1__496_, data_stage_1__495_, data_stage_1__494_, data_stage_1__493_, data_stage_1__492_, data_stage_1__491_, data_stage_1__490_, data_stage_1__489_, data_stage_1__488_, data_stage_1__487_, data_stage_1__486_, data_stage_1__485_, data_stage_1__484_, data_stage_1__483_, data_stage_1__482_, data_stage_1__481_, data_stage_1__480_, data_stage_1__479_, data_stage_1__478_, data_stage_1__477_, data_stage_1__476_, data_stage_1__475_, data_stage_1__474_, data_stage_1__473_, data_stage_1__472_, data_stage_1__471_, data_stage_1__470_, data_stage_1__469_, data_stage_1__468_, data_stage_1__467_, data_stage_1__466_, data_stage_1__465_, data_stage_1__464_, data_stage_1__463_, data_stage_1__462_, data_stage_1__461_, data_stage_1__460_, data_stage_1__459_, data_stage_1__458_, data_stage_1__457_, data_stage_1__456_, data_stage_1__455_, data_stage_1__454_, data_stage_1__453_, data_stage_1__452_, data_stage_1__451_, data_stage_1__450_, data_stage_1__449_, data_stage_1__448_, data_stage_1__447_, data_stage_1__446_, data_stage_1__445_, data_stage_1__444_, data_stage_1__443_, data_stage_1__442_, data_stage_1__441_, data_stage_1__440_, data_stage_1__439_, data_stage_1__438_, data_stage_1__437_, data_stage_1__436_, data_stage_1__435_, data_stage_1__434_, data_stage_1__433_, data_stage_1__432_, data_stage_1__431_, data_stage_1__430_, data_stage_1__429_, data_stage_1__428_, data_stage_1__427_, data_stage_1__426_, data_stage_1__425_, data_stage_1__424_, data_stage_1__423_, data_stage_1__422_, data_stage_1__421_, data_stage_1__420_, data_stage_1__419_, data_stage_1__418_, data_stage_1__417_, data_stage_1__416_, data_stage_1__415_, data_stage_1__414_, data_stage_1__413_, data_stage_1__412_, data_stage_1__411_, data_stage_1__410_, data_stage_1__409_, data_stage_1__408_, data_stage_1__407_, data_stage_1__406_, data_stage_1__405_, data_stage_1__404_, data_stage_1__403_, data_stage_1__402_, data_stage_1__401_, data_stage_1__400_, data_stage_1__399_, data_stage_1__398_, data_stage_1__397_, data_stage_1__396_, data_stage_1__395_, data_stage_1__394_, data_stage_1__393_, data_stage_1__392_, data_stage_1__391_, data_stage_1__390_, data_stage_1__389_, data_stage_1__388_, data_stage_1__387_, data_stage_1__386_, data_stage_1__385_, data_stage_1__384_, data_stage_1__383_, data_stage_1__382_, data_stage_1__381_, data_stage_1__380_, data_stage_1__379_, data_stage_1__378_, data_stage_1__377_, data_stage_1__376_, data_stage_1__375_, data_stage_1__374_, data_stage_1__373_, data_stage_1__372_, data_stage_1__371_, data_stage_1__370_, data_stage_1__369_, data_stage_1__368_, data_stage_1__367_, data_stage_1__366_, data_stage_1__365_, data_stage_1__364_, data_stage_1__363_, data_stage_1__362_, data_stage_1__361_, data_stage_1__360_, data_stage_1__359_, data_stage_1__358_, data_stage_1__357_, data_stage_1__356_, data_stage_1__355_, data_stage_1__354_, data_stage_1__353_, data_stage_1__352_, data_stage_1__351_, data_stage_1__350_, data_stage_1__349_, data_stage_1__348_, data_stage_1__347_, data_stage_1__346_, data_stage_1__345_, data_stage_1__344_, data_stage_1__343_, data_stage_1__342_, data_stage_1__341_, data_stage_1__340_, data_stage_1__339_, data_stage_1__338_, data_stage_1__337_, data_stage_1__336_, data_stage_1__335_, data_stage_1__334_, data_stage_1__333_, data_stage_1__332_, data_stage_1__331_, data_stage_1__330_, data_stage_1__329_, data_stage_1__328_, data_stage_1__327_, data_stage_1__326_, data_stage_1__325_, data_stage_1__324_, data_stage_1__323_, data_stage_1__322_, data_stage_1__321_, data_stage_1__320_, data_stage_1__319_, data_stage_1__318_, data_stage_1__317_, data_stage_1__316_, data_stage_1__315_, data_stage_1__314_, data_stage_1__313_, data_stage_1__312_, data_stage_1__311_, data_stage_1__310_, data_stage_1__309_, data_stage_1__308_, data_stage_1__307_, data_stage_1__306_, data_stage_1__305_, data_stage_1__304_, data_stage_1__303_, data_stage_1__302_, data_stage_1__301_, data_stage_1__300_, data_stage_1__299_, data_stage_1__298_, data_stage_1__297_, data_stage_1__296_, data_stage_1__295_, data_stage_1__294_, data_stage_1__293_, data_stage_1__292_, data_stage_1__291_, data_stage_1__290_, data_stage_1__289_, data_stage_1__288_, data_stage_1__287_, data_stage_1__286_, data_stage_1__285_, data_stage_1__284_, data_stage_1__283_, data_stage_1__282_, data_stage_1__281_, data_stage_1__280_, data_stage_1__279_, data_stage_1__278_, data_stage_1__277_, data_stage_1__276_, data_stage_1__275_, data_stage_1__274_, data_stage_1__273_, data_stage_1__272_, data_stage_1__271_, data_stage_1__270_, data_stage_1__269_, data_stage_1__268_, data_stage_1__267_, data_stage_1__266_, data_stage_1__265_, data_stage_1__264_, data_stage_1__263_, data_stage_1__262_, data_stage_1__261_, data_stage_1__260_, data_stage_1__259_, data_stage_1__258_, data_stage_1__257_, data_stage_1__256_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__511_, data_stage_2__510_, data_stage_2__509_, data_stage_2__508_, data_stage_2__507_, data_stage_2__506_, data_stage_2__505_, data_stage_2__504_, data_stage_2__503_, data_stage_2__502_, data_stage_2__501_, data_stage_2__500_, data_stage_2__499_, data_stage_2__498_, data_stage_2__497_, data_stage_2__496_, data_stage_2__495_, data_stage_2__494_, data_stage_2__493_, data_stage_2__492_, data_stage_2__491_, data_stage_2__490_, data_stage_2__489_, data_stage_2__488_, data_stage_2__487_, data_stage_2__486_, data_stage_2__485_, data_stage_2__484_, data_stage_2__483_, data_stage_2__482_, data_stage_2__481_, data_stage_2__480_, data_stage_2__479_, data_stage_2__478_, data_stage_2__477_, data_stage_2__476_, data_stage_2__475_, data_stage_2__474_, data_stage_2__473_, data_stage_2__472_, data_stage_2__471_, data_stage_2__470_, data_stage_2__469_, data_stage_2__468_, data_stage_2__467_, data_stage_2__466_, data_stage_2__465_, data_stage_2__464_, data_stage_2__463_, data_stage_2__462_, data_stage_2__461_, data_stage_2__460_, data_stage_2__459_, data_stage_2__458_, data_stage_2__457_, data_stage_2__456_, data_stage_2__455_, data_stage_2__454_, data_stage_2__453_, data_stage_2__452_, data_stage_2__451_, data_stage_2__450_, data_stage_2__449_, data_stage_2__448_, data_stage_2__447_, data_stage_2__446_, data_stage_2__445_, data_stage_2__444_, data_stage_2__443_, data_stage_2__442_, data_stage_2__441_, data_stage_2__440_, data_stage_2__439_, data_stage_2__438_, data_stage_2__437_, data_stage_2__436_, data_stage_2__435_, data_stage_2__434_, data_stage_2__433_, data_stage_2__432_, data_stage_2__431_, data_stage_2__430_, data_stage_2__429_, data_stage_2__428_, data_stage_2__427_, data_stage_2__426_, data_stage_2__425_, data_stage_2__424_, data_stage_2__423_, data_stage_2__422_, data_stage_2__421_, data_stage_2__420_, data_stage_2__419_, data_stage_2__418_, data_stage_2__417_, data_stage_2__416_, data_stage_2__415_, data_stage_2__414_, data_stage_2__413_, data_stage_2__412_, data_stage_2__411_, data_stage_2__410_, data_stage_2__409_, data_stage_2__408_, data_stage_2__407_, data_stage_2__406_, data_stage_2__405_, data_stage_2__404_, data_stage_2__403_, data_stage_2__402_, data_stage_2__401_, data_stage_2__400_, data_stage_2__399_, data_stage_2__398_, data_stage_2__397_, data_stage_2__396_, data_stage_2__395_, data_stage_2__394_, data_stage_2__393_, data_stage_2__392_, data_stage_2__391_, data_stage_2__390_, data_stage_2__389_, data_stage_2__388_, data_stage_2__387_, data_stage_2__386_, data_stage_2__385_, data_stage_2__384_, data_stage_2__383_, data_stage_2__382_, data_stage_2__381_, data_stage_2__380_, data_stage_2__379_, data_stage_2__378_, data_stage_2__377_, data_stage_2__376_, data_stage_2__375_, data_stage_2__374_, data_stage_2__373_, data_stage_2__372_, data_stage_2__371_, data_stage_2__370_, data_stage_2__369_, data_stage_2__368_, data_stage_2__367_, data_stage_2__366_, data_stage_2__365_, data_stage_2__364_, data_stage_2__363_, data_stage_2__362_, data_stage_2__361_, data_stage_2__360_, data_stage_2__359_, data_stage_2__358_, data_stage_2__357_, data_stage_2__356_, data_stage_2__355_, data_stage_2__354_, data_stage_2__353_, data_stage_2__352_, data_stage_2__351_, data_stage_2__350_, data_stage_2__349_, data_stage_2__348_, data_stage_2__347_, data_stage_2__346_, data_stage_2__345_, data_stage_2__344_, data_stage_2__343_, data_stage_2__342_, data_stage_2__341_, data_stage_2__340_, data_stage_2__339_, data_stage_2__338_, data_stage_2__337_, data_stage_2__336_, data_stage_2__335_, data_stage_2__334_, data_stage_2__333_, data_stage_2__332_, data_stage_2__331_, data_stage_2__330_, data_stage_2__329_, data_stage_2__328_, data_stage_2__327_, data_stage_2__326_, data_stage_2__325_, data_stage_2__324_, data_stage_2__323_, data_stage_2__322_, data_stage_2__321_, data_stage_2__320_, data_stage_2__319_, data_stage_2__318_, data_stage_2__317_, data_stage_2__316_, data_stage_2__315_, data_stage_2__314_, data_stage_2__313_, data_stage_2__312_, data_stage_2__311_, data_stage_2__310_, data_stage_2__309_, data_stage_2__308_, data_stage_2__307_, data_stage_2__306_, data_stage_2__305_, data_stage_2__304_, data_stage_2__303_, data_stage_2__302_, data_stage_2__301_, data_stage_2__300_, data_stage_2__299_, data_stage_2__298_, data_stage_2__297_, data_stage_2__296_, data_stage_2__295_, data_stage_2__294_, data_stage_2__293_, data_stage_2__292_, data_stage_2__291_, data_stage_2__290_, data_stage_2__289_, data_stage_2__288_, data_stage_2__287_, data_stage_2__286_, data_stage_2__285_, data_stage_2__284_, data_stage_2__283_, data_stage_2__282_, data_stage_2__281_, data_stage_2__280_, data_stage_2__279_, data_stage_2__278_, data_stage_2__277_, data_stage_2__276_, data_stage_2__275_, data_stage_2__274_, data_stage_2__273_, data_stage_2__272_, data_stage_2__271_, data_stage_2__270_, data_stage_2__269_, data_stage_2__268_, data_stage_2__267_, data_stage_2__266_, data_stage_2__265_, data_stage_2__264_, data_stage_2__263_, data_stage_2__262_, data_stage_2__261_, data_stage_2__260_, data_stage_2__259_, data_stage_2__258_, data_stage_2__257_, data_stage_2__256_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_2__swap_inst
  (
    .data_i({ data_stage_1__767_, data_stage_1__766_, data_stage_1__765_, data_stage_1__764_, data_stage_1__763_, data_stage_1__762_, data_stage_1__761_, data_stage_1__760_, data_stage_1__759_, data_stage_1__758_, data_stage_1__757_, data_stage_1__756_, data_stage_1__755_, data_stage_1__754_, data_stage_1__753_, data_stage_1__752_, data_stage_1__751_, data_stage_1__750_, data_stage_1__749_, data_stage_1__748_, data_stage_1__747_, data_stage_1__746_, data_stage_1__745_, data_stage_1__744_, data_stage_1__743_, data_stage_1__742_, data_stage_1__741_, data_stage_1__740_, data_stage_1__739_, data_stage_1__738_, data_stage_1__737_, data_stage_1__736_, data_stage_1__735_, data_stage_1__734_, data_stage_1__733_, data_stage_1__732_, data_stage_1__731_, data_stage_1__730_, data_stage_1__729_, data_stage_1__728_, data_stage_1__727_, data_stage_1__726_, data_stage_1__725_, data_stage_1__724_, data_stage_1__723_, data_stage_1__722_, data_stage_1__721_, data_stage_1__720_, data_stage_1__719_, data_stage_1__718_, data_stage_1__717_, data_stage_1__716_, data_stage_1__715_, data_stage_1__714_, data_stage_1__713_, data_stage_1__712_, data_stage_1__711_, data_stage_1__710_, data_stage_1__709_, data_stage_1__708_, data_stage_1__707_, data_stage_1__706_, data_stage_1__705_, data_stage_1__704_, data_stage_1__703_, data_stage_1__702_, data_stage_1__701_, data_stage_1__700_, data_stage_1__699_, data_stage_1__698_, data_stage_1__697_, data_stage_1__696_, data_stage_1__695_, data_stage_1__694_, data_stage_1__693_, data_stage_1__692_, data_stage_1__691_, data_stage_1__690_, data_stage_1__689_, data_stage_1__688_, data_stage_1__687_, data_stage_1__686_, data_stage_1__685_, data_stage_1__684_, data_stage_1__683_, data_stage_1__682_, data_stage_1__681_, data_stage_1__680_, data_stage_1__679_, data_stage_1__678_, data_stage_1__677_, data_stage_1__676_, data_stage_1__675_, data_stage_1__674_, data_stage_1__673_, data_stage_1__672_, data_stage_1__671_, data_stage_1__670_, data_stage_1__669_, data_stage_1__668_, data_stage_1__667_, data_stage_1__666_, data_stage_1__665_, data_stage_1__664_, data_stage_1__663_, data_stage_1__662_, data_stage_1__661_, data_stage_1__660_, data_stage_1__659_, data_stage_1__658_, data_stage_1__657_, data_stage_1__656_, data_stage_1__655_, data_stage_1__654_, data_stage_1__653_, data_stage_1__652_, data_stage_1__651_, data_stage_1__650_, data_stage_1__649_, data_stage_1__648_, data_stage_1__647_, data_stage_1__646_, data_stage_1__645_, data_stage_1__644_, data_stage_1__643_, data_stage_1__642_, data_stage_1__641_, data_stage_1__640_, data_stage_1__639_, data_stage_1__638_, data_stage_1__637_, data_stage_1__636_, data_stage_1__635_, data_stage_1__634_, data_stage_1__633_, data_stage_1__632_, data_stage_1__631_, data_stage_1__630_, data_stage_1__629_, data_stage_1__628_, data_stage_1__627_, data_stage_1__626_, data_stage_1__625_, data_stage_1__624_, data_stage_1__623_, data_stage_1__622_, data_stage_1__621_, data_stage_1__620_, data_stage_1__619_, data_stage_1__618_, data_stage_1__617_, data_stage_1__616_, data_stage_1__615_, data_stage_1__614_, data_stage_1__613_, data_stage_1__612_, data_stage_1__611_, data_stage_1__610_, data_stage_1__609_, data_stage_1__608_, data_stage_1__607_, data_stage_1__606_, data_stage_1__605_, data_stage_1__604_, data_stage_1__603_, data_stage_1__602_, data_stage_1__601_, data_stage_1__600_, data_stage_1__599_, data_stage_1__598_, data_stage_1__597_, data_stage_1__596_, data_stage_1__595_, data_stage_1__594_, data_stage_1__593_, data_stage_1__592_, data_stage_1__591_, data_stage_1__590_, data_stage_1__589_, data_stage_1__588_, data_stage_1__587_, data_stage_1__586_, data_stage_1__585_, data_stage_1__584_, data_stage_1__583_, data_stage_1__582_, data_stage_1__581_, data_stage_1__580_, data_stage_1__579_, data_stage_1__578_, data_stage_1__577_, data_stage_1__576_, data_stage_1__575_, data_stage_1__574_, data_stage_1__573_, data_stage_1__572_, data_stage_1__571_, data_stage_1__570_, data_stage_1__569_, data_stage_1__568_, data_stage_1__567_, data_stage_1__566_, data_stage_1__565_, data_stage_1__564_, data_stage_1__563_, data_stage_1__562_, data_stage_1__561_, data_stage_1__560_, data_stage_1__559_, data_stage_1__558_, data_stage_1__557_, data_stage_1__556_, data_stage_1__555_, data_stage_1__554_, data_stage_1__553_, data_stage_1__552_, data_stage_1__551_, data_stage_1__550_, data_stage_1__549_, data_stage_1__548_, data_stage_1__547_, data_stage_1__546_, data_stage_1__545_, data_stage_1__544_, data_stage_1__543_, data_stage_1__542_, data_stage_1__541_, data_stage_1__540_, data_stage_1__539_, data_stage_1__538_, data_stage_1__537_, data_stage_1__536_, data_stage_1__535_, data_stage_1__534_, data_stage_1__533_, data_stage_1__532_, data_stage_1__531_, data_stage_1__530_, data_stage_1__529_, data_stage_1__528_, data_stage_1__527_, data_stage_1__526_, data_stage_1__525_, data_stage_1__524_, data_stage_1__523_, data_stage_1__522_, data_stage_1__521_, data_stage_1__520_, data_stage_1__519_, data_stage_1__518_, data_stage_1__517_, data_stage_1__516_, data_stage_1__515_, data_stage_1__514_, data_stage_1__513_, data_stage_1__512_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__767_, data_stage_2__766_, data_stage_2__765_, data_stage_2__764_, data_stage_2__763_, data_stage_2__762_, data_stage_2__761_, data_stage_2__760_, data_stage_2__759_, data_stage_2__758_, data_stage_2__757_, data_stage_2__756_, data_stage_2__755_, data_stage_2__754_, data_stage_2__753_, data_stage_2__752_, data_stage_2__751_, data_stage_2__750_, data_stage_2__749_, data_stage_2__748_, data_stage_2__747_, data_stage_2__746_, data_stage_2__745_, data_stage_2__744_, data_stage_2__743_, data_stage_2__742_, data_stage_2__741_, data_stage_2__740_, data_stage_2__739_, data_stage_2__738_, data_stage_2__737_, data_stage_2__736_, data_stage_2__735_, data_stage_2__734_, data_stage_2__733_, data_stage_2__732_, data_stage_2__731_, data_stage_2__730_, data_stage_2__729_, data_stage_2__728_, data_stage_2__727_, data_stage_2__726_, data_stage_2__725_, data_stage_2__724_, data_stage_2__723_, data_stage_2__722_, data_stage_2__721_, data_stage_2__720_, data_stage_2__719_, data_stage_2__718_, data_stage_2__717_, data_stage_2__716_, data_stage_2__715_, data_stage_2__714_, data_stage_2__713_, data_stage_2__712_, data_stage_2__711_, data_stage_2__710_, data_stage_2__709_, data_stage_2__708_, data_stage_2__707_, data_stage_2__706_, data_stage_2__705_, data_stage_2__704_, data_stage_2__703_, data_stage_2__702_, data_stage_2__701_, data_stage_2__700_, data_stage_2__699_, data_stage_2__698_, data_stage_2__697_, data_stage_2__696_, data_stage_2__695_, data_stage_2__694_, data_stage_2__693_, data_stage_2__692_, data_stage_2__691_, data_stage_2__690_, data_stage_2__689_, data_stage_2__688_, data_stage_2__687_, data_stage_2__686_, data_stage_2__685_, data_stage_2__684_, data_stage_2__683_, data_stage_2__682_, data_stage_2__681_, data_stage_2__680_, data_stage_2__679_, data_stage_2__678_, data_stage_2__677_, data_stage_2__676_, data_stage_2__675_, data_stage_2__674_, data_stage_2__673_, data_stage_2__672_, data_stage_2__671_, data_stage_2__670_, data_stage_2__669_, data_stage_2__668_, data_stage_2__667_, data_stage_2__666_, data_stage_2__665_, data_stage_2__664_, data_stage_2__663_, data_stage_2__662_, data_stage_2__661_, data_stage_2__660_, data_stage_2__659_, data_stage_2__658_, data_stage_2__657_, data_stage_2__656_, data_stage_2__655_, data_stage_2__654_, data_stage_2__653_, data_stage_2__652_, data_stage_2__651_, data_stage_2__650_, data_stage_2__649_, data_stage_2__648_, data_stage_2__647_, data_stage_2__646_, data_stage_2__645_, data_stage_2__644_, data_stage_2__643_, data_stage_2__642_, data_stage_2__641_, data_stage_2__640_, data_stage_2__639_, data_stage_2__638_, data_stage_2__637_, data_stage_2__636_, data_stage_2__635_, data_stage_2__634_, data_stage_2__633_, data_stage_2__632_, data_stage_2__631_, data_stage_2__630_, data_stage_2__629_, data_stage_2__628_, data_stage_2__627_, data_stage_2__626_, data_stage_2__625_, data_stage_2__624_, data_stage_2__623_, data_stage_2__622_, data_stage_2__621_, data_stage_2__620_, data_stage_2__619_, data_stage_2__618_, data_stage_2__617_, data_stage_2__616_, data_stage_2__615_, data_stage_2__614_, data_stage_2__613_, data_stage_2__612_, data_stage_2__611_, data_stage_2__610_, data_stage_2__609_, data_stage_2__608_, data_stage_2__607_, data_stage_2__606_, data_stage_2__605_, data_stage_2__604_, data_stage_2__603_, data_stage_2__602_, data_stage_2__601_, data_stage_2__600_, data_stage_2__599_, data_stage_2__598_, data_stage_2__597_, data_stage_2__596_, data_stage_2__595_, data_stage_2__594_, data_stage_2__593_, data_stage_2__592_, data_stage_2__591_, data_stage_2__590_, data_stage_2__589_, data_stage_2__588_, data_stage_2__587_, data_stage_2__586_, data_stage_2__585_, data_stage_2__584_, data_stage_2__583_, data_stage_2__582_, data_stage_2__581_, data_stage_2__580_, data_stage_2__579_, data_stage_2__578_, data_stage_2__577_, data_stage_2__576_, data_stage_2__575_, data_stage_2__574_, data_stage_2__573_, data_stage_2__572_, data_stage_2__571_, data_stage_2__570_, data_stage_2__569_, data_stage_2__568_, data_stage_2__567_, data_stage_2__566_, data_stage_2__565_, data_stage_2__564_, data_stage_2__563_, data_stage_2__562_, data_stage_2__561_, data_stage_2__560_, data_stage_2__559_, data_stage_2__558_, data_stage_2__557_, data_stage_2__556_, data_stage_2__555_, data_stage_2__554_, data_stage_2__553_, data_stage_2__552_, data_stage_2__551_, data_stage_2__550_, data_stage_2__549_, data_stage_2__548_, data_stage_2__547_, data_stage_2__546_, data_stage_2__545_, data_stage_2__544_, data_stage_2__543_, data_stage_2__542_, data_stage_2__541_, data_stage_2__540_, data_stage_2__539_, data_stage_2__538_, data_stage_2__537_, data_stage_2__536_, data_stage_2__535_, data_stage_2__534_, data_stage_2__533_, data_stage_2__532_, data_stage_2__531_, data_stage_2__530_, data_stage_2__529_, data_stage_2__528_, data_stage_2__527_, data_stage_2__526_, data_stage_2__525_, data_stage_2__524_, data_stage_2__523_, data_stage_2__522_, data_stage_2__521_, data_stage_2__520_, data_stage_2__519_, data_stage_2__518_, data_stage_2__517_, data_stage_2__516_, data_stage_2__515_, data_stage_2__514_, data_stage_2__513_, data_stage_2__512_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_3__swap_inst
  (
    .data_i({ data_stage_1__1023_, data_stage_1__1022_, data_stage_1__1021_, data_stage_1__1020_, data_stage_1__1019_, data_stage_1__1018_, data_stage_1__1017_, data_stage_1__1016_, data_stage_1__1015_, data_stage_1__1014_, data_stage_1__1013_, data_stage_1__1012_, data_stage_1__1011_, data_stage_1__1010_, data_stage_1__1009_, data_stage_1__1008_, data_stage_1__1007_, data_stage_1__1006_, data_stage_1__1005_, data_stage_1__1004_, data_stage_1__1003_, data_stage_1__1002_, data_stage_1__1001_, data_stage_1__1000_, data_stage_1__999_, data_stage_1__998_, data_stage_1__997_, data_stage_1__996_, data_stage_1__995_, data_stage_1__994_, data_stage_1__993_, data_stage_1__992_, data_stage_1__991_, data_stage_1__990_, data_stage_1__989_, data_stage_1__988_, data_stage_1__987_, data_stage_1__986_, data_stage_1__985_, data_stage_1__984_, data_stage_1__983_, data_stage_1__982_, data_stage_1__981_, data_stage_1__980_, data_stage_1__979_, data_stage_1__978_, data_stage_1__977_, data_stage_1__976_, data_stage_1__975_, data_stage_1__974_, data_stage_1__973_, data_stage_1__972_, data_stage_1__971_, data_stage_1__970_, data_stage_1__969_, data_stage_1__968_, data_stage_1__967_, data_stage_1__966_, data_stage_1__965_, data_stage_1__964_, data_stage_1__963_, data_stage_1__962_, data_stage_1__961_, data_stage_1__960_, data_stage_1__959_, data_stage_1__958_, data_stage_1__957_, data_stage_1__956_, data_stage_1__955_, data_stage_1__954_, data_stage_1__953_, data_stage_1__952_, data_stage_1__951_, data_stage_1__950_, data_stage_1__949_, data_stage_1__948_, data_stage_1__947_, data_stage_1__946_, data_stage_1__945_, data_stage_1__944_, data_stage_1__943_, data_stage_1__942_, data_stage_1__941_, data_stage_1__940_, data_stage_1__939_, data_stage_1__938_, data_stage_1__937_, data_stage_1__936_, data_stage_1__935_, data_stage_1__934_, data_stage_1__933_, data_stage_1__932_, data_stage_1__931_, data_stage_1__930_, data_stage_1__929_, data_stage_1__928_, data_stage_1__927_, data_stage_1__926_, data_stage_1__925_, data_stage_1__924_, data_stage_1__923_, data_stage_1__922_, data_stage_1__921_, data_stage_1__920_, data_stage_1__919_, data_stage_1__918_, data_stage_1__917_, data_stage_1__916_, data_stage_1__915_, data_stage_1__914_, data_stage_1__913_, data_stage_1__912_, data_stage_1__911_, data_stage_1__910_, data_stage_1__909_, data_stage_1__908_, data_stage_1__907_, data_stage_1__906_, data_stage_1__905_, data_stage_1__904_, data_stage_1__903_, data_stage_1__902_, data_stage_1__901_, data_stage_1__900_, data_stage_1__899_, data_stage_1__898_, data_stage_1__897_, data_stage_1__896_, data_stage_1__895_, data_stage_1__894_, data_stage_1__893_, data_stage_1__892_, data_stage_1__891_, data_stage_1__890_, data_stage_1__889_, data_stage_1__888_, data_stage_1__887_, data_stage_1__886_, data_stage_1__885_, data_stage_1__884_, data_stage_1__883_, data_stage_1__882_, data_stage_1__881_, data_stage_1__880_, data_stage_1__879_, data_stage_1__878_, data_stage_1__877_, data_stage_1__876_, data_stage_1__875_, data_stage_1__874_, data_stage_1__873_, data_stage_1__872_, data_stage_1__871_, data_stage_1__870_, data_stage_1__869_, data_stage_1__868_, data_stage_1__867_, data_stage_1__866_, data_stage_1__865_, data_stage_1__864_, data_stage_1__863_, data_stage_1__862_, data_stage_1__861_, data_stage_1__860_, data_stage_1__859_, data_stage_1__858_, data_stage_1__857_, data_stage_1__856_, data_stage_1__855_, data_stage_1__854_, data_stage_1__853_, data_stage_1__852_, data_stage_1__851_, data_stage_1__850_, data_stage_1__849_, data_stage_1__848_, data_stage_1__847_, data_stage_1__846_, data_stage_1__845_, data_stage_1__844_, data_stage_1__843_, data_stage_1__842_, data_stage_1__841_, data_stage_1__840_, data_stage_1__839_, data_stage_1__838_, data_stage_1__837_, data_stage_1__836_, data_stage_1__835_, data_stage_1__834_, data_stage_1__833_, data_stage_1__832_, data_stage_1__831_, data_stage_1__830_, data_stage_1__829_, data_stage_1__828_, data_stage_1__827_, data_stage_1__826_, data_stage_1__825_, data_stage_1__824_, data_stage_1__823_, data_stage_1__822_, data_stage_1__821_, data_stage_1__820_, data_stage_1__819_, data_stage_1__818_, data_stage_1__817_, data_stage_1__816_, data_stage_1__815_, data_stage_1__814_, data_stage_1__813_, data_stage_1__812_, data_stage_1__811_, data_stage_1__810_, data_stage_1__809_, data_stage_1__808_, data_stage_1__807_, data_stage_1__806_, data_stage_1__805_, data_stage_1__804_, data_stage_1__803_, data_stage_1__802_, data_stage_1__801_, data_stage_1__800_, data_stage_1__799_, data_stage_1__798_, data_stage_1__797_, data_stage_1__796_, data_stage_1__795_, data_stage_1__794_, data_stage_1__793_, data_stage_1__792_, data_stage_1__791_, data_stage_1__790_, data_stage_1__789_, data_stage_1__788_, data_stage_1__787_, data_stage_1__786_, data_stage_1__785_, data_stage_1__784_, data_stage_1__783_, data_stage_1__782_, data_stage_1__781_, data_stage_1__780_, data_stage_1__779_, data_stage_1__778_, data_stage_1__777_, data_stage_1__776_, data_stage_1__775_, data_stage_1__774_, data_stage_1__773_, data_stage_1__772_, data_stage_1__771_, data_stage_1__770_, data_stage_1__769_, data_stage_1__768_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__1023_, data_stage_2__1022_, data_stage_2__1021_, data_stage_2__1020_, data_stage_2__1019_, data_stage_2__1018_, data_stage_2__1017_, data_stage_2__1016_, data_stage_2__1015_, data_stage_2__1014_, data_stage_2__1013_, data_stage_2__1012_, data_stage_2__1011_, data_stage_2__1010_, data_stage_2__1009_, data_stage_2__1008_, data_stage_2__1007_, data_stage_2__1006_, data_stage_2__1005_, data_stage_2__1004_, data_stage_2__1003_, data_stage_2__1002_, data_stage_2__1001_, data_stage_2__1000_, data_stage_2__999_, data_stage_2__998_, data_stage_2__997_, data_stage_2__996_, data_stage_2__995_, data_stage_2__994_, data_stage_2__993_, data_stage_2__992_, data_stage_2__991_, data_stage_2__990_, data_stage_2__989_, data_stage_2__988_, data_stage_2__987_, data_stage_2__986_, data_stage_2__985_, data_stage_2__984_, data_stage_2__983_, data_stage_2__982_, data_stage_2__981_, data_stage_2__980_, data_stage_2__979_, data_stage_2__978_, data_stage_2__977_, data_stage_2__976_, data_stage_2__975_, data_stage_2__974_, data_stage_2__973_, data_stage_2__972_, data_stage_2__971_, data_stage_2__970_, data_stage_2__969_, data_stage_2__968_, data_stage_2__967_, data_stage_2__966_, data_stage_2__965_, data_stage_2__964_, data_stage_2__963_, data_stage_2__962_, data_stage_2__961_, data_stage_2__960_, data_stage_2__959_, data_stage_2__958_, data_stage_2__957_, data_stage_2__956_, data_stage_2__955_, data_stage_2__954_, data_stage_2__953_, data_stage_2__952_, data_stage_2__951_, data_stage_2__950_, data_stage_2__949_, data_stage_2__948_, data_stage_2__947_, data_stage_2__946_, data_stage_2__945_, data_stage_2__944_, data_stage_2__943_, data_stage_2__942_, data_stage_2__941_, data_stage_2__940_, data_stage_2__939_, data_stage_2__938_, data_stage_2__937_, data_stage_2__936_, data_stage_2__935_, data_stage_2__934_, data_stage_2__933_, data_stage_2__932_, data_stage_2__931_, data_stage_2__930_, data_stage_2__929_, data_stage_2__928_, data_stage_2__927_, data_stage_2__926_, data_stage_2__925_, data_stage_2__924_, data_stage_2__923_, data_stage_2__922_, data_stage_2__921_, data_stage_2__920_, data_stage_2__919_, data_stage_2__918_, data_stage_2__917_, data_stage_2__916_, data_stage_2__915_, data_stage_2__914_, data_stage_2__913_, data_stage_2__912_, data_stage_2__911_, data_stage_2__910_, data_stage_2__909_, data_stage_2__908_, data_stage_2__907_, data_stage_2__906_, data_stage_2__905_, data_stage_2__904_, data_stage_2__903_, data_stage_2__902_, data_stage_2__901_, data_stage_2__900_, data_stage_2__899_, data_stage_2__898_, data_stage_2__897_, data_stage_2__896_, data_stage_2__895_, data_stage_2__894_, data_stage_2__893_, data_stage_2__892_, data_stage_2__891_, data_stage_2__890_, data_stage_2__889_, data_stage_2__888_, data_stage_2__887_, data_stage_2__886_, data_stage_2__885_, data_stage_2__884_, data_stage_2__883_, data_stage_2__882_, data_stage_2__881_, data_stage_2__880_, data_stage_2__879_, data_stage_2__878_, data_stage_2__877_, data_stage_2__876_, data_stage_2__875_, data_stage_2__874_, data_stage_2__873_, data_stage_2__872_, data_stage_2__871_, data_stage_2__870_, data_stage_2__869_, data_stage_2__868_, data_stage_2__867_, data_stage_2__866_, data_stage_2__865_, data_stage_2__864_, data_stage_2__863_, data_stage_2__862_, data_stage_2__861_, data_stage_2__860_, data_stage_2__859_, data_stage_2__858_, data_stage_2__857_, data_stage_2__856_, data_stage_2__855_, data_stage_2__854_, data_stage_2__853_, data_stage_2__852_, data_stage_2__851_, data_stage_2__850_, data_stage_2__849_, data_stage_2__848_, data_stage_2__847_, data_stage_2__846_, data_stage_2__845_, data_stage_2__844_, data_stage_2__843_, data_stage_2__842_, data_stage_2__841_, data_stage_2__840_, data_stage_2__839_, data_stage_2__838_, data_stage_2__837_, data_stage_2__836_, data_stage_2__835_, data_stage_2__834_, data_stage_2__833_, data_stage_2__832_, data_stage_2__831_, data_stage_2__830_, data_stage_2__829_, data_stage_2__828_, data_stage_2__827_, data_stage_2__826_, data_stage_2__825_, data_stage_2__824_, data_stage_2__823_, data_stage_2__822_, data_stage_2__821_, data_stage_2__820_, data_stage_2__819_, data_stage_2__818_, data_stage_2__817_, data_stage_2__816_, data_stage_2__815_, data_stage_2__814_, data_stage_2__813_, data_stage_2__812_, data_stage_2__811_, data_stage_2__810_, data_stage_2__809_, data_stage_2__808_, data_stage_2__807_, data_stage_2__806_, data_stage_2__805_, data_stage_2__804_, data_stage_2__803_, data_stage_2__802_, data_stage_2__801_, data_stage_2__800_, data_stage_2__799_, data_stage_2__798_, data_stage_2__797_, data_stage_2__796_, data_stage_2__795_, data_stage_2__794_, data_stage_2__793_, data_stage_2__792_, data_stage_2__791_, data_stage_2__790_, data_stage_2__789_, data_stage_2__788_, data_stage_2__787_, data_stage_2__786_, data_stage_2__785_, data_stage_2__784_, data_stage_2__783_, data_stage_2__782_, data_stage_2__781_, data_stage_2__780_, data_stage_2__779_, data_stage_2__778_, data_stage_2__777_, data_stage_2__776_, data_stage_2__775_, data_stage_2__774_, data_stage_2__773_, data_stage_2__772_, data_stage_2__771_, data_stage_2__770_, data_stage_2__769_, data_stage_2__768_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_4__swap_inst
  (
    .data_i({ data_stage_1__1279_, data_stage_1__1278_, data_stage_1__1277_, data_stage_1__1276_, data_stage_1__1275_, data_stage_1__1274_, data_stage_1__1273_, data_stage_1__1272_, data_stage_1__1271_, data_stage_1__1270_, data_stage_1__1269_, data_stage_1__1268_, data_stage_1__1267_, data_stage_1__1266_, data_stage_1__1265_, data_stage_1__1264_, data_stage_1__1263_, data_stage_1__1262_, data_stage_1__1261_, data_stage_1__1260_, data_stage_1__1259_, data_stage_1__1258_, data_stage_1__1257_, data_stage_1__1256_, data_stage_1__1255_, data_stage_1__1254_, data_stage_1__1253_, data_stage_1__1252_, data_stage_1__1251_, data_stage_1__1250_, data_stage_1__1249_, data_stage_1__1248_, data_stage_1__1247_, data_stage_1__1246_, data_stage_1__1245_, data_stage_1__1244_, data_stage_1__1243_, data_stage_1__1242_, data_stage_1__1241_, data_stage_1__1240_, data_stage_1__1239_, data_stage_1__1238_, data_stage_1__1237_, data_stage_1__1236_, data_stage_1__1235_, data_stage_1__1234_, data_stage_1__1233_, data_stage_1__1232_, data_stage_1__1231_, data_stage_1__1230_, data_stage_1__1229_, data_stage_1__1228_, data_stage_1__1227_, data_stage_1__1226_, data_stage_1__1225_, data_stage_1__1224_, data_stage_1__1223_, data_stage_1__1222_, data_stage_1__1221_, data_stage_1__1220_, data_stage_1__1219_, data_stage_1__1218_, data_stage_1__1217_, data_stage_1__1216_, data_stage_1__1215_, data_stage_1__1214_, data_stage_1__1213_, data_stage_1__1212_, data_stage_1__1211_, data_stage_1__1210_, data_stage_1__1209_, data_stage_1__1208_, data_stage_1__1207_, data_stage_1__1206_, data_stage_1__1205_, data_stage_1__1204_, data_stage_1__1203_, data_stage_1__1202_, data_stage_1__1201_, data_stage_1__1200_, data_stage_1__1199_, data_stage_1__1198_, data_stage_1__1197_, data_stage_1__1196_, data_stage_1__1195_, data_stage_1__1194_, data_stage_1__1193_, data_stage_1__1192_, data_stage_1__1191_, data_stage_1__1190_, data_stage_1__1189_, data_stage_1__1188_, data_stage_1__1187_, data_stage_1__1186_, data_stage_1__1185_, data_stage_1__1184_, data_stage_1__1183_, data_stage_1__1182_, data_stage_1__1181_, data_stage_1__1180_, data_stage_1__1179_, data_stage_1__1178_, data_stage_1__1177_, data_stage_1__1176_, data_stage_1__1175_, data_stage_1__1174_, data_stage_1__1173_, data_stage_1__1172_, data_stage_1__1171_, data_stage_1__1170_, data_stage_1__1169_, data_stage_1__1168_, data_stage_1__1167_, data_stage_1__1166_, data_stage_1__1165_, data_stage_1__1164_, data_stage_1__1163_, data_stage_1__1162_, data_stage_1__1161_, data_stage_1__1160_, data_stage_1__1159_, data_stage_1__1158_, data_stage_1__1157_, data_stage_1__1156_, data_stage_1__1155_, data_stage_1__1154_, data_stage_1__1153_, data_stage_1__1152_, data_stage_1__1151_, data_stage_1__1150_, data_stage_1__1149_, data_stage_1__1148_, data_stage_1__1147_, data_stage_1__1146_, data_stage_1__1145_, data_stage_1__1144_, data_stage_1__1143_, data_stage_1__1142_, data_stage_1__1141_, data_stage_1__1140_, data_stage_1__1139_, data_stage_1__1138_, data_stage_1__1137_, data_stage_1__1136_, data_stage_1__1135_, data_stage_1__1134_, data_stage_1__1133_, data_stage_1__1132_, data_stage_1__1131_, data_stage_1__1130_, data_stage_1__1129_, data_stage_1__1128_, data_stage_1__1127_, data_stage_1__1126_, data_stage_1__1125_, data_stage_1__1124_, data_stage_1__1123_, data_stage_1__1122_, data_stage_1__1121_, data_stage_1__1120_, data_stage_1__1119_, data_stage_1__1118_, data_stage_1__1117_, data_stage_1__1116_, data_stage_1__1115_, data_stage_1__1114_, data_stage_1__1113_, data_stage_1__1112_, data_stage_1__1111_, data_stage_1__1110_, data_stage_1__1109_, data_stage_1__1108_, data_stage_1__1107_, data_stage_1__1106_, data_stage_1__1105_, data_stage_1__1104_, data_stage_1__1103_, data_stage_1__1102_, data_stage_1__1101_, data_stage_1__1100_, data_stage_1__1099_, data_stage_1__1098_, data_stage_1__1097_, data_stage_1__1096_, data_stage_1__1095_, data_stage_1__1094_, data_stage_1__1093_, data_stage_1__1092_, data_stage_1__1091_, data_stage_1__1090_, data_stage_1__1089_, data_stage_1__1088_, data_stage_1__1087_, data_stage_1__1086_, data_stage_1__1085_, data_stage_1__1084_, data_stage_1__1083_, data_stage_1__1082_, data_stage_1__1081_, data_stage_1__1080_, data_stage_1__1079_, data_stage_1__1078_, data_stage_1__1077_, data_stage_1__1076_, data_stage_1__1075_, data_stage_1__1074_, data_stage_1__1073_, data_stage_1__1072_, data_stage_1__1071_, data_stage_1__1070_, data_stage_1__1069_, data_stage_1__1068_, data_stage_1__1067_, data_stage_1__1066_, data_stage_1__1065_, data_stage_1__1064_, data_stage_1__1063_, data_stage_1__1062_, data_stage_1__1061_, data_stage_1__1060_, data_stage_1__1059_, data_stage_1__1058_, data_stage_1__1057_, data_stage_1__1056_, data_stage_1__1055_, data_stage_1__1054_, data_stage_1__1053_, data_stage_1__1052_, data_stage_1__1051_, data_stage_1__1050_, data_stage_1__1049_, data_stage_1__1048_, data_stage_1__1047_, data_stage_1__1046_, data_stage_1__1045_, data_stage_1__1044_, data_stage_1__1043_, data_stage_1__1042_, data_stage_1__1041_, data_stage_1__1040_, data_stage_1__1039_, data_stage_1__1038_, data_stage_1__1037_, data_stage_1__1036_, data_stage_1__1035_, data_stage_1__1034_, data_stage_1__1033_, data_stage_1__1032_, data_stage_1__1031_, data_stage_1__1030_, data_stage_1__1029_, data_stage_1__1028_, data_stage_1__1027_, data_stage_1__1026_, data_stage_1__1025_, data_stage_1__1024_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__1279_, data_stage_2__1278_, data_stage_2__1277_, data_stage_2__1276_, data_stage_2__1275_, data_stage_2__1274_, data_stage_2__1273_, data_stage_2__1272_, data_stage_2__1271_, data_stage_2__1270_, data_stage_2__1269_, data_stage_2__1268_, data_stage_2__1267_, data_stage_2__1266_, data_stage_2__1265_, data_stage_2__1264_, data_stage_2__1263_, data_stage_2__1262_, data_stage_2__1261_, data_stage_2__1260_, data_stage_2__1259_, data_stage_2__1258_, data_stage_2__1257_, data_stage_2__1256_, data_stage_2__1255_, data_stage_2__1254_, data_stage_2__1253_, data_stage_2__1252_, data_stage_2__1251_, data_stage_2__1250_, data_stage_2__1249_, data_stage_2__1248_, data_stage_2__1247_, data_stage_2__1246_, data_stage_2__1245_, data_stage_2__1244_, data_stage_2__1243_, data_stage_2__1242_, data_stage_2__1241_, data_stage_2__1240_, data_stage_2__1239_, data_stage_2__1238_, data_stage_2__1237_, data_stage_2__1236_, data_stage_2__1235_, data_stage_2__1234_, data_stage_2__1233_, data_stage_2__1232_, data_stage_2__1231_, data_stage_2__1230_, data_stage_2__1229_, data_stage_2__1228_, data_stage_2__1227_, data_stage_2__1226_, data_stage_2__1225_, data_stage_2__1224_, data_stage_2__1223_, data_stage_2__1222_, data_stage_2__1221_, data_stage_2__1220_, data_stage_2__1219_, data_stage_2__1218_, data_stage_2__1217_, data_stage_2__1216_, data_stage_2__1215_, data_stage_2__1214_, data_stage_2__1213_, data_stage_2__1212_, data_stage_2__1211_, data_stage_2__1210_, data_stage_2__1209_, data_stage_2__1208_, data_stage_2__1207_, data_stage_2__1206_, data_stage_2__1205_, data_stage_2__1204_, data_stage_2__1203_, data_stage_2__1202_, data_stage_2__1201_, data_stage_2__1200_, data_stage_2__1199_, data_stage_2__1198_, data_stage_2__1197_, data_stage_2__1196_, data_stage_2__1195_, data_stage_2__1194_, data_stage_2__1193_, data_stage_2__1192_, data_stage_2__1191_, data_stage_2__1190_, data_stage_2__1189_, data_stage_2__1188_, data_stage_2__1187_, data_stage_2__1186_, data_stage_2__1185_, data_stage_2__1184_, data_stage_2__1183_, data_stage_2__1182_, data_stage_2__1181_, data_stage_2__1180_, data_stage_2__1179_, data_stage_2__1178_, data_stage_2__1177_, data_stage_2__1176_, data_stage_2__1175_, data_stage_2__1174_, data_stage_2__1173_, data_stage_2__1172_, data_stage_2__1171_, data_stage_2__1170_, data_stage_2__1169_, data_stage_2__1168_, data_stage_2__1167_, data_stage_2__1166_, data_stage_2__1165_, data_stage_2__1164_, data_stage_2__1163_, data_stage_2__1162_, data_stage_2__1161_, data_stage_2__1160_, data_stage_2__1159_, data_stage_2__1158_, data_stage_2__1157_, data_stage_2__1156_, data_stage_2__1155_, data_stage_2__1154_, data_stage_2__1153_, data_stage_2__1152_, data_stage_2__1151_, data_stage_2__1150_, data_stage_2__1149_, data_stage_2__1148_, data_stage_2__1147_, data_stage_2__1146_, data_stage_2__1145_, data_stage_2__1144_, data_stage_2__1143_, data_stage_2__1142_, data_stage_2__1141_, data_stage_2__1140_, data_stage_2__1139_, data_stage_2__1138_, data_stage_2__1137_, data_stage_2__1136_, data_stage_2__1135_, data_stage_2__1134_, data_stage_2__1133_, data_stage_2__1132_, data_stage_2__1131_, data_stage_2__1130_, data_stage_2__1129_, data_stage_2__1128_, data_stage_2__1127_, data_stage_2__1126_, data_stage_2__1125_, data_stage_2__1124_, data_stage_2__1123_, data_stage_2__1122_, data_stage_2__1121_, data_stage_2__1120_, data_stage_2__1119_, data_stage_2__1118_, data_stage_2__1117_, data_stage_2__1116_, data_stage_2__1115_, data_stage_2__1114_, data_stage_2__1113_, data_stage_2__1112_, data_stage_2__1111_, data_stage_2__1110_, data_stage_2__1109_, data_stage_2__1108_, data_stage_2__1107_, data_stage_2__1106_, data_stage_2__1105_, data_stage_2__1104_, data_stage_2__1103_, data_stage_2__1102_, data_stage_2__1101_, data_stage_2__1100_, data_stage_2__1099_, data_stage_2__1098_, data_stage_2__1097_, data_stage_2__1096_, data_stage_2__1095_, data_stage_2__1094_, data_stage_2__1093_, data_stage_2__1092_, data_stage_2__1091_, data_stage_2__1090_, data_stage_2__1089_, data_stage_2__1088_, data_stage_2__1087_, data_stage_2__1086_, data_stage_2__1085_, data_stage_2__1084_, data_stage_2__1083_, data_stage_2__1082_, data_stage_2__1081_, data_stage_2__1080_, data_stage_2__1079_, data_stage_2__1078_, data_stage_2__1077_, data_stage_2__1076_, data_stage_2__1075_, data_stage_2__1074_, data_stage_2__1073_, data_stage_2__1072_, data_stage_2__1071_, data_stage_2__1070_, data_stage_2__1069_, data_stage_2__1068_, data_stage_2__1067_, data_stage_2__1066_, data_stage_2__1065_, data_stage_2__1064_, data_stage_2__1063_, data_stage_2__1062_, data_stage_2__1061_, data_stage_2__1060_, data_stage_2__1059_, data_stage_2__1058_, data_stage_2__1057_, data_stage_2__1056_, data_stage_2__1055_, data_stage_2__1054_, data_stage_2__1053_, data_stage_2__1052_, data_stage_2__1051_, data_stage_2__1050_, data_stage_2__1049_, data_stage_2__1048_, data_stage_2__1047_, data_stage_2__1046_, data_stage_2__1045_, data_stage_2__1044_, data_stage_2__1043_, data_stage_2__1042_, data_stage_2__1041_, data_stage_2__1040_, data_stage_2__1039_, data_stage_2__1038_, data_stage_2__1037_, data_stage_2__1036_, data_stage_2__1035_, data_stage_2__1034_, data_stage_2__1033_, data_stage_2__1032_, data_stage_2__1031_, data_stage_2__1030_, data_stage_2__1029_, data_stage_2__1028_, data_stage_2__1027_, data_stage_2__1026_, data_stage_2__1025_, data_stage_2__1024_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_5__swap_inst
  (
    .data_i({ data_stage_1__1535_, data_stage_1__1534_, data_stage_1__1533_, data_stage_1__1532_, data_stage_1__1531_, data_stage_1__1530_, data_stage_1__1529_, data_stage_1__1528_, data_stage_1__1527_, data_stage_1__1526_, data_stage_1__1525_, data_stage_1__1524_, data_stage_1__1523_, data_stage_1__1522_, data_stage_1__1521_, data_stage_1__1520_, data_stage_1__1519_, data_stage_1__1518_, data_stage_1__1517_, data_stage_1__1516_, data_stage_1__1515_, data_stage_1__1514_, data_stage_1__1513_, data_stage_1__1512_, data_stage_1__1511_, data_stage_1__1510_, data_stage_1__1509_, data_stage_1__1508_, data_stage_1__1507_, data_stage_1__1506_, data_stage_1__1505_, data_stage_1__1504_, data_stage_1__1503_, data_stage_1__1502_, data_stage_1__1501_, data_stage_1__1500_, data_stage_1__1499_, data_stage_1__1498_, data_stage_1__1497_, data_stage_1__1496_, data_stage_1__1495_, data_stage_1__1494_, data_stage_1__1493_, data_stage_1__1492_, data_stage_1__1491_, data_stage_1__1490_, data_stage_1__1489_, data_stage_1__1488_, data_stage_1__1487_, data_stage_1__1486_, data_stage_1__1485_, data_stage_1__1484_, data_stage_1__1483_, data_stage_1__1482_, data_stage_1__1481_, data_stage_1__1480_, data_stage_1__1479_, data_stage_1__1478_, data_stage_1__1477_, data_stage_1__1476_, data_stage_1__1475_, data_stage_1__1474_, data_stage_1__1473_, data_stage_1__1472_, data_stage_1__1471_, data_stage_1__1470_, data_stage_1__1469_, data_stage_1__1468_, data_stage_1__1467_, data_stage_1__1466_, data_stage_1__1465_, data_stage_1__1464_, data_stage_1__1463_, data_stage_1__1462_, data_stage_1__1461_, data_stage_1__1460_, data_stage_1__1459_, data_stage_1__1458_, data_stage_1__1457_, data_stage_1__1456_, data_stage_1__1455_, data_stage_1__1454_, data_stage_1__1453_, data_stage_1__1452_, data_stage_1__1451_, data_stage_1__1450_, data_stage_1__1449_, data_stage_1__1448_, data_stage_1__1447_, data_stage_1__1446_, data_stage_1__1445_, data_stage_1__1444_, data_stage_1__1443_, data_stage_1__1442_, data_stage_1__1441_, data_stage_1__1440_, data_stage_1__1439_, data_stage_1__1438_, data_stage_1__1437_, data_stage_1__1436_, data_stage_1__1435_, data_stage_1__1434_, data_stage_1__1433_, data_stage_1__1432_, data_stage_1__1431_, data_stage_1__1430_, data_stage_1__1429_, data_stage_1__1428_, data_stage_1__1427_, data_stage_1__1426_, data_stage_1__1425_, data_stage_1__1424_, data_stage_1__1423_, data_stage_1__1422_, data_stage_1__1421_, data_stage_1__1420_, data_stage_1__1419_, data_stage_1__1418_, data_stage_1__1417_, data_stage_1__1416_, data_stage_1__1415_, data_stage_1__1414_, data_stage_1__1413_, data_stage_1__1412_, data_stage_1__1411_, data_stage_1__1410_, data_stage_1__1409_, data_stage_1__1408_, data_stage_1__1407_, data_stage_1__1406_, data_stage_1__1405_, data_stage_1__1404_, data_stage_1__1403_, data_stage_1__1402_, data_stage_1__1401_, data_stage_1__1400_, data_stage_1__1399_, data_stage_1__1398_, data_stage_1__1397_, data_stage_1__1396_, data_stage_1__1395_, data_stage_1__1394_, data_stage_1__1393_, data_stage_1__1392_, data_stage_1__1391_, data_stage_1__1390_, data_stage_1__1389_, data_stage_1__1388_, data_stage_1__1387_, data_stage_1__1386_, data_stage_1__1385_, data_stage_1__1384_, data_stage_1__1383_, data_stage_1__1382_, data_stage_1__1381_, data_stage_1__1380_, data_stage_1__1379_, data_stage_1__1378_, data_stage_1__1377_, data_stage_1__1376_, data_stage_1__1375_, data_stage_1__1374_, data_stage_1__1373_, data_stage_1__1372_, data_stage_1__1371_, data_stage_1__1370_, data_stage_1__1369_, data_stage_1__1368_, data_stage_1__1367_, data_stage_1__1366_, data_stage_1__1365_, data_stage_1__1364_, data_stage_1__1363_, data_stage_1__1362_, data_stage_1__1361_, data_stage_1__1360_, data_stage_1__1359_, data_stage_1__1358_, data_stage_1__1357_, data_stage_1__1356_, data_stage_1__1355_, data_stage_1__1354_, data_stage_1__1353_, data_stage_1__1352_, data_stage_1__1351_, data_stage_1__1350_, data_stage_1__1349_, data_stage_1__1348_, data_stage_1__1347_, data_stage_1__1346_, data_stage_1__1345_, data_stage_1__1344_, data_stage_1__1343_, data_stage_1__1342_, data_stage_1__1341_, data_stage_1__1340_, data_stage_1__1339_, data_stage_1__1338_, data_stage_1__1337_, data_stage_1__1336_, data_stage_1__1335_, data_stage_1__1334_, data_stage_1__1333_, data_stage_1__1332_, data_stage_1__1331_, data_stage_1__1330_, data_stage_1__1329_, data_stage_1__1328_, data_stage_1__1327_, data_stage_1__1326_, data_stage_1__1325_, data_stage_1__1324_, data_stage_1__1323_, data_stage_1__1322_, data_stage_1__1321_, data_stage_1__1320_, data_stage_1__1319_, data_stage_1__1318_, data_stage_1__1317_, data_stage_1__1316_, data_stage_1__1315_, data_stage_1__1314_, data_stage_1__1313_, data_stage_1__1312_, data_stage_1__1311_, data_stage_1__1310_, data_stage_1__1309_, data_stage_1__1308_, data_stage_1__1307_, data_stage_1__1306_, data_stage_1__1305_, data_stage_1__1304_, data_stage_1__1303_, data_stage_1__1302_, data_stage_1__1301_, data_stage_1__1300_, data_stage_1__1299_, data_stage_1__1298_, data_stage_1__1297_, data_stage_1__1296_, data_stage_1__1295_, data_stage_1__1294_, data_stage_1__1293_, data_stage_1__1292_, data_stage_1__1291_, data_stage_1__1290_, data_stage_1__1289_, data_stage_1__1288_, data_stage_1__1287_, data_stage_1__1286_, data_stage_1__1285_, data_stage_1__1284_, data_stage_1__1283_, data_stage_1__1282_, data_stage_1__1281_, data_stage_1__1280_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__1535_, data_stage_2__1534_, data_stage_2__1533_, data_stage_2__1532_, data_stage_2__1531_, data_stage_2__1530_, data_stage_2__1529_, data_stage_2__1528_, data_stage_2__1527_, data_stage_2__1526_, data_stage_2__1525_, data_stage_2__1524_, data_stage_2__1523_, data_stage_2__1522_, data_stage_2__1521_, data_stage_2__1520_, data_stage_2__1519_, data_stage_2__1518_, data_stage_2__1517_, data_stage_2__1516_, data_stage_2__1515_, data_stage_2__1514_, data_stage_2__1513_, data_stage_2__1512_, data_stage_2__1511_, data_stage_2__1510_, data_stage_2__1509_, data_stage_2__1508_, data_stage_2__1507_, data_stage_2__1506_, data_stage_2__1505_, data_stage_2__1504_, data_stage_2__1503_, data_stage_2__1502_, data_stage_2__1501_, data_stage_2__1500_, data_stage_2__1499_, data_stage_2__1498_, data_stage_2__1497_, data_stage_2__1496_, data_stage_2__1495_, data_stage_2__1494_, data_stage_2__1493_, data_stage_2__1492_, data_stage_2__1491_, data_stage_2__1490_, data_stage_2__1489_, data_stage_2__1488_, data_stage_2__1487_, data_stage_2__1486_, data_stage_2__1485_, data_stage_2__1484_, data_stage_2__1483_, data_stage_2__1482_, data_stage_2__1481_, data_stage_2__1480_, data_stage_2__1479_, data_stage_2__1478_, data_stage_2__1477_, data_stage_2__1476_, data_stage_2__1475_, data_stage_2__1474_, data_stage_2__1473_, data_stage_2__1472_, data_stage_2__1471_, data_stage_2__1470_, data_stage_2__1469_, data_stage_2__1468_, data_stage_2__1467_, data_stage_2__1466_, data_stage_2__1465_, data_stage_2__1464_, data_stage_2__1463_, data_stage_2__1462_, data_stage_2__1461_, data_stage_2__1460_, data_stage_2__1459_, data_stage_2__1458_, data_stage_2__1457_, data_stage_2__1456_, data_stage_2__1455_, data_stage_2__1454_, data_stage_2__1453_, data_stage_2__1452_, data_stage_2__1451_, data_stage_2__1450_, data_stage_2__1449_, data_stage_2__1448_, data_stage_2__1447_, data_stage_2__1446_, data_stage_2__1445_, data_stage_2__1444_, data_stage_2__1443_, data_stage_2__1442_, data_stage_2__1441_, data_stage_2__1440_, data_stage_2__1439_, data_stage_2__1438_, data_stage_2__1437_, data_stage_2__1436_, data_stage_2__1435_, data_stage_2__1434_, data_stage_2__1433_, data_stage_2__1432_, data_stage_2__1431_, data_stage_2__1430_, data_stage_2__1429_, data_stage_2__1428_, data_stage_2__1427_, data_stage_2__1426_, data_stage_2__1425_, data_stage_2__1424_, data_stage_2__1423_, data_stage_2__1422_, data_stage_2__1421_, data_stage_2__1420_, data_stage_2__1419_, data_stage_2__1418_, data_stage_2__1417_, data_stage_2__1416_, data_stage_2__1415_, data_stage_2__1414_, data_stage_2__1413_, data_stage_2__1412_, data_stage_2__1411_, data_stage_2__1410_, data_stage_2__1409_, data_stage_2__1408_, data_stage_2__1407_, data_stage_2__1406_, data_stage_2__1405_, data_stage_2__1404_, data_stage_2__1403_, data_stage_2__1402_, data_stage_2__1401_, data_stage_2__1400_, data_stage_2__1399_, data_stage_2__1398_, data_stage_2__1397_, data_stage_2__1396_, data_stage_2__1395_, data_stage_2__1394_, data_stage_2__1393_, data_stage_2__1392_, data_stage_2__1391_, data_stage_2__1390_, data_stage_2__1389_, data_stage_2__1388_, data_stage_2__1387_, data_stage_2__1386_, data_stage_2__1385_, data_stage_2__1384_, data_stage_2__1383_, data_stage_2__1382_, data_stage_2__1381_, data_stage_2__1380_, data_stage_2__1379_, data_stage_2__1378_, data_stage_2__1377_, data_stage_2__1376_, data_stage_2__1375_, data_stage_2__1374_, data_stage_2__1373_, data_stage_2__1372_, data_stage_2__1371_, data_stage_2__1370_, data_stage_2__1369_, data_stage_2__1368_, data_stage_2__1367_, data_stage_2__1366_, data_stage_2__1365_, data_stage_2__1364_, data_stage_2__1363_, data_stage_2__1362_, data_stage_2__1361_, data_stage_2__1360_, data_stage_2__1359_, data_stage_2__1358_, data_stage_2__1357_, data_stage_2__1356_, data_stage_2__1355_, data_stage_2__1354_, data_stage_2__1353_, data_stage_2__1352_, data_stage_2__1351_, data_stage_2__1350_, data_stage_2__1349_, data_stage_2__1348_, data_stage_2__1347_, data_stage_2__1346_, data_stage_2__1345_, data_stage_2__1344_, data_stage_2__1343_, data_stage_2__1342_, data_stage_2__1341_, data_stage_2__1340_, data_stage_2__1339_, data_stage_2__1338_, data_stage_2__1337_, data_stage_2__1336_, data_stage_2__1335_, data_stage_2__1334_, data_stage_2__1333_, data_stage_2__1332_, data_stage_2__1331_, data_stage_2__1330_, data_stage_2__1329_, data_stage_2__1328_, data_stage_2__1327_, data_stage_2__1326_, data_stage_2__1325_, data_stage_2__1324_, data_stage_2__1323_, data_stage_2__1322_, data_stage_2__1321_, data_stage_2__1320_, data_stage_2__1319_, data_stage_2__1318_, data_stage_2__1317_, data_stage_2__1316_, data_stage_2__1315_, data_stage_2__1314_, data_stage_2__1313_, data_stage_2__1312_, data_stage_2__1311_, data_stage_2__1310_, data_stage_2__1309_, data_stage_2__1308_, data_stage_2__1307_, data_stage_2__1306_, data_stage_2__1305_, data_stage_2__1304_, data_stage_2__1303_, data_stage_2__1302_, data_stage_2__1301_, data_stage_2__1300_, data_stage_2__1299_, data_stage_2__1298_, data_stage_2__1297_, data_stage_2__1296_, data_stage_2__1295_, data_stage_2__1294_, data_stage_2__1293_, data_stage_2__1292_, data_stage_2__1291_, data_stage_2__1290_, data_stage_2__1289_, data_stage_2__1288_, data_stage_2__1287_, data_stage_2__1286_, data_stage_2__1285_, data_stage_2__1284_, data_stage_2__1283_, data_stage_2__1282_, data_stage_2__1281_, data_stage_2__1280_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_6__swap_inst
  (
    .data_i({ data_stage_1__1791_, data_stage_1__1790_, data_stage_1__1789_, data_stage_1__1788_, data_stage_1__1787_, data_stage_1__1786_, data_stage_1__1785_, data_stage_1__1784_, data_stage_1__1783_, data_stage_1__1782_, data_stage_1__1781_, data_stage_1__1780_, data_stage_1__1779_, data_stage_1__1778_, data_stage_1__1777_, data_stage_1__1776_, data_stage_1__1775_, data_stage_1__1774_, data_stage_1__1773_, data_stage_1__1772_, data_stage_1__1771_, data_stage_1__1770_, data_stage_1__1769_, data_stage_1__1768_, data_stage_1__1767_, data_stage_1__1766_, data_stage_1__1765_, data_stage_1__1764_, data_stage_1__1763_, data_stage_1__1762_, data_stage_1__1761_, data_stage_1__1760_, data_stage_1__1759_, data_stage_1__1758_, data_stage_1__1757_, data_stage_1__1756_, data_stage_1__1755_, data_stage_1__1754_, data_stage_1__1753_, data_stage_1__1752_, data_stage_1__1751_, data_stage_1__1750_, data_stage_1__1749_, data_stage_1__1748_, data_stage_1__1747_, data_stage_1__1746_, data_stage_1__1745_, data_stage_1__1744_, data_stage_1__1743_, data_stage_1__1742_, data_stage_1__1741_, data_stage_1__1740_, data_stage_1__1739_, data_stage_1__1738_, data_stage_1__1737_, data_stage_1__1736_, data_stage_1__1735_, data_stage_1__1734_, data_stage_1__1733_, data_stage_1__1732_, data_stage_1__1731_, data_stage_1__1730_, data_stage_1__1729_, data_stage_1__1728_, data_stage_1__1727_, data_stage_1__1726_, data_stage_1__1725_, data_stage_1__1724_, data_stage_1__1723_, data_stage_1__1722_, data_stage_1__1721_, data_stage_1__1720_, data_stage_1__1719_, data_stage_1__1718_, data_stage_1__1717_, data_stage_1__1716_, data_stage_1__1715_, data_stage_1__1714_, data_stage_1__1713_, data_stage_1__1712_, data_stage_1__1711_, data_stage_1__1710_, data_stage_1__1709_, data_stage_1__1708_, data_stage_1__1707_, data_stage_1__1706_, data_stage_1__1705_, data_stage_1__1704_, data_stage_1__1703_, data_stage_1__1702_, data_stage_1__1701_, data_stage_1__1700_, data_stage_1__1699_, data_stage_1__1698_, data_stage_1__1697_, data_stage_1__1696_, data_stage_1__1695_, data_stage_1__1694_, data_stage_1__1693_, data_stage_1__1692_, data_stage_1__1691_, data_stage_1__1690_, data_stage_1__1689_, data_stage_1__1688_, data_stage_1__1687_, data_stage_1__1686_, data_stage_1__1685_, data_stage_1__1684_, data_stage_1__1683_, data_stage_1__1682_, data_stage_1__1681_, data_stage_1__1680_, data_stage_1__1679_, data_stage_1__1678_, data_stage_1__1677_, data_stage_1__1676_, data_stage_1__1675_, data_stage_1__1674_, data_stage_1__1673_, data_stage_1__1672_, data_stage_1__1671_, data_stage_1__1670_, data_stage_1__1669_, data_stage_1__1668_, data_stage_1__1667_, data_stage_1__1666_, data_stage_1__1665_, data_stage_1__1664_, data_stage_1__1663_, data_stage_1__1662_, data_stage_1__1661_, data_stage_1__1660_, data_stage_1__1659_, data_stage_1__1658_, data_stage_1__1657_, data_stage_1__1656_, data_stage_1__1655_, data_stage_1__1654_, data_stage_1__1653_, data_stage_1__1652_, data_stage_1__1651_, data_stage_1__1650_, data_stage_1__1649_, data_stage_1__1648_, data_stage_1__1647_, data_stage_1__1646_, data_stage_1__1645_, data_stage_1__1644_, data_stage_1__1643_, data_stage_1__1642_, data_stage_1__1641_, data_stage_1__1640_, data_stage_1__1639_, data_stage_1__1638_, data_stage_1__1637_, data_stage_1__1636_, data_stage_1__1635_, data_stage_1__1634_, data_stage_1__1633_, data_stage_1__1632_, data_stage_1__1631_, data_stage_1__1630_, data_stage_1__1629_, data_stage_1__1628_, data_stage_1__1627_, data_stage_1__1626_, data_stage_1__1625_, data_stage_1__1624_, data_stage_1__1623_, data_stage_1__1622_, data_stage_1__1621_, data_stage_1__1620_, data_stage_1__1619_, data_stage_1__1618_, data_stage_1__1617_, data_stage_1__1616_, data_stage_1__1615_, data_stage_1__1614_, data_stage_1__1613_, data_stage_1__1612_, data_stage_1__1611_, data_stage_1__1610_, data_stage_1__1609_, data_stage_1__1608_, data_stage_1__1607_, data_stage_1__1606_, data_stage_1__1605_, data_stage_1__1604_, data_stage_1__1603_, data_stage_1__1602_, data_stage_1__1601_, data_stage_1__1600_, data_stage_1__1599_, data_stage_1__1598_, data_stage_1__1597_, data_stage_1__1596_, data_stage_1__1595_, data_stage_1__1594_, data_stage_1__1593_, data_stage_1__1592_, data_stage_1__1591_, data_stage_1__1590_, data_stage_1__1589_, data_stage_1__1588_, data_stage_1__1587_, data_stage_1__1586_, data_stage_1__1585_, data_stage_1__1584_, data_stage_1__1583_, data_stage_1__1582_, data_stage_1__1581_, data_stage_1__1580_, data_stage_1__1579_, data_stage_1__1578_, data_stage_1__1577_, data_stage_1__1576_, data_stage_1__1575_, data_stage_1__1574_, data_stage_1__1573_, data_stage_1__1572_, data_stage_1__1571_, data_stage_1__1570_, data_stage_1__1569_, data_stage_1__1568_, data_stage_1__1567_, data_stage_1__1566_, data_stage_1__1565_, data_stage_1__1564_, data_stage_1__1563_, data_stage_1__1562_, data_stage_1__1561_, data_stage_1__1560_, data_stage_1__1559_, data_stage_1__1558_, data_stage_1__1557_, data_stage_1__1556_, data_stage_1__1555_, data_stage_1__1554_, data_stage_1__1553_, data_stage_1__1552_, data_stage_1__1551_, data_stage_1__1550_, data_stage_1__1549_, data_stage_1__1548_, data_stage_1__1547_, data_stage_1__1546_, data_stage_1__1545_, data_stage_1__1544_, data_stage_1__1543_, data_stage_1__1542_, data_stage_1__1541_, data_stage_1__1540_, data_stage_1__1539_, data_stage_1__1538_, data_stage_1__1537_, data_stage_1__1536_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__1791_, data_stage_2__1790_, data_stage_2__1789_, data_stage_2__1788_, data_stage_2__1787_, data_stage_2__1786_, data_stage_2__1785_, data_stage_2__1784_, data_stage_2__1783_, data_stage_2__1782_, data_stage_2__1781_, data_stage_2__1780_, data_stage_2__1779_, data_stage_2__1778_, data_stage_2__1777_, data_stage_2__1776_, data_stage_2__1775_, data_stage_2__1774_, data_stage_2__1773_, data_stage_2__1772_, data_stage_2__1771_, data_stage_2__1770_, data_stage_2__1769_, data_stage_2__1768_, data_stage_2__1767_, data_stage_2__1766_, data_stage_2__1765_, data_stage_2__1764_, data_stage_2__1763_, data_stage_2__1762_, data_stage_2__1761_, data_stage_2__1760_, data_stage_2__1759_, data_stage_2__1758_, data_stage_2__1757_, data_stage_2__1756_, data_stage_2__1755_, data_stage_2__1754_, data_stage_2__1753_, data_stage_2__1752_, data_stage_2__1751_, data_stage_2__1750_, data_stage_2__1749_, data_stage_2__1748_, data_stage_2__1747_, data_stage_2__1746_, data_stage_2__1745_, data_stage_2__1744_, data_stage_2__1743_, data_stage_2__1742_, data_stage_2__1741_, data_stage_2__1740_, data_stage_2__1739_, data_stage_2__1738_, data_stage_2__1737_, data_stage_2__1736_, data_stage_2__1735_, data_stage_2__1734_, data_stage_2__1733_, data_stage_2__1732_, data_stage_2__1731_, data_stage_2__1730_, data_stage_2__1729_, data_stage_2__1728_, data_stage_2__1727_, data_stage_2__1726_, data_stage_2__1725_, data_stage_2__1724_, data_stage_2__1723_, data_stage_2__1722_, data_stage_2__1721_, data_stage_2__1720_, data_stage_2__1719_, data_stage_2__1718_, data_stage_2__1717_, data_stage_2__1716_, data_stage_2__1715_, data_stage_2__1714_, data_stage_2__1713_, data_stage_2__1712_, data_stage_2__1711_, data_stage_2__1710_, data_stage_2__1709_, data_stage_2__1708_, data_stage_2__1707_, data_stage_2__1706_, data_stage_2__1705_, data_stage_2__1704_, data_stage_2__1703_, data_stage_2__1702_, data_stage_2__1701_, data_stage_2__1700_, data_stage_2__1699_, data_stage_2__1698_, data_stage_2__1697_, data_stage_2__1696_, data_stage_2__1695_, data_stage_2__1694_, data_stage_2__1693_, data_stage_2__1692_, data_stage_2__1691_, data_stage_2__1690_, data_stage_2__1689_, data_stage_2__1688_, data_stage_2__1687_, data_stage_2__1686_, data_stage_2__1685_, data_stage_2__1684_, data_stage_2__1683_, data_stage_2__1682_, data_stage_2__1681_, data_stage_2__1680_, data_stage_2__1679_, data_stage_2__1678_, data_stage_2__1677_, data_stage_2__1676_, data_stage_2__1675_, data_stage_2__1674_, data_stage_2__1673_, data_stage_2__1672_, data_stage_2__1671_, data_stage_2__1670_, data_stage_2__1669_, data_stage_2__1668_, data_stage_2__1667_, data_stage_2__1666_, data_stage_2__1665_, data_stage_2__1664_, data_stage_2__1663_, data_stage_2__1662_, data_stage_2__1661_, data_stage_2__1660_, data_stage_2__1659_, data_stage_2__1658_, data_stage_2__1657_, data_stage_2__1656_, data_stage_2__1655_, data_stage_2__1654_, data_stage_2__1653_, data_stage_2__1652_, data_stage_2__1651_, data_stage_2__1650_, data_stage_2__1649_, data_stage_2__1648_, data_stage_2__1647_, data_stage_2__1646_, data_stage_2__1645_, data_stage_2__1644_, data_stage_2__1643_, data_stage_2__1642_, data_stage_2__1641_, data_stage_2__1640_, data_stage_2__1639_, data_stage_2__1638_, data_stage_2__1637_, data_stage_2__1636_, data_stage_2__1635_, data_stage_2__1634_, data_stage_2__1633_, data_stage_2__1632_, data_stage_2__1631_, data_stage_2__1630_, data_stage_2__1629_, data_stage_2__1628_, data_stage_2__1627_, data_stage_2__1626_, data_stage_2__1625_, data_stage_2__1624_, data_stage_2__1623_, data_stage_2__1622_, data_stage_2__1621_, data_stage_2__1620_, data_stage_2__1619_, data_stage_2__1618_, data_stage_2__1617_, data_stage_2__1616_, data_stage_2__1615_, data_stage_2__1614_, data_stage_2__1613_, data_stage_2__1612_, data_stage_2__1611_, data_stage_2__1610_, data_stage_2__1609_, data_stage_2__1608_, data_stage_2__1607_, data_stage_2__1606_, data_stage_2__1605_, data_stage_2__1604_, data_stage_2__1603_, data_stage_2__1602_, data_stage_2__1601_, data_stage_2__1600_, data_stage_2__1599_, data_stage_2__1598_, data_stage_2__1597_, data_stage_2__1596_, data_stage_2__1595_, data_stage_2__1594_, data_stage_2__1593_, data_stage_2__1592_, data_stage_2__1591_, data_stage_2__1590_, data_stage_2__1589_, data_stage_2__1588_, data_stage_2__1587_, data_stage_2__1586_, data_stage_2__1585_, data_stage_2__1584_, data_stage_2__1583_, data_stage_2__1582_, data_stage_2__1581_, data_stage_2__1580_, data_stage_2__1579_, data_stage_2__1578_, data_stage_2__1577_, data_stage_2__1576_, data_stage_2__1575_, data_stage_2__1574_, data_stage_2__1573_, data_stage_2__1572_, data_stage_2__1571_, data_stage_2__1570_, data_stage_2__1569_, data_stage_2__1568_, data_stage_2__1567_, data_stage_2__1566_, data_stage_2__1565_, data_stage_2__1564_, data_stage_2__1563_, data_stage_2__1562_, data_stage_2__1561_, data_stage_2__1560_, data_stage_2__1559_, data_stage_2__1558_, data_stage_2__1557_, data_stage_2__1556_, data_stage_2__1555_, data_stage_2__1554_, data_stage_2__1553_, data_stage_2__1552_, data_stage_2__1551_, data_stage_2__1550_, data_stage_2__1549_, data_stage_2__1548_, data_stage_2__1547_, data_stage_2__1546_, data_stage_2__1545_, data_stage_2__1544_, data_stage_2__1543_, data_stage_2__1542_, data_stage_2__1541_, data_stage_2__1540_, data_stage_2__1539_, data_stage_2__1538_, data_stage_2__1537_, data_stage_2__1536_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_7__swap_inst
  (
    .data_i({ data_stage_1__2047_, data_stage_1__2046_, data_stage_1__2045_, data_stage_1__2044_, data_stage_1__2043_, data_stage_1__2042_, data_stage_1__2041_, data_stage_1__2040_, data_stage_1__2039_, data_stage_1__2038_, data_stage_1__2037_, data_stage_1__2036_, data_stage_1__2035_, data_stage_1__2034_, data_stage_1__2033_, data_stage_1__2032_, data_stage_1__2031_, data_stage_1__2030_, data_stage_1__2029_, data_stage_1__2028_, data_stage_1__2027_, data_stage_1__2026_, data_stage_1__2025_, data_stage_1__2024_, data_stage_1__2023_, data_stage_1__2022_, data_stage_1__2021_, data_stage_1__2020_, data_stage_1__2019_, data_stage_1__2018_, data_stage_1__2017_, data_stage_1__2016_, data_stage_1__2015_, data_stage_1__2014_, data_stage_1__2013_, data_stage_1__2012_, data_stage_1__2011_, data_stage_1__2010_, data_stage_1__2009_, data_stage_1__2008_, data_stage_1__2007_, data_stage_1__2006_, data_stage_1__2005_, data_stage_1__2004_, data_stage_1__2003_, data_stage_1__2002_, data_stage_1__2001_, data_stage_1__2000_, data_stage_1__1999_, data_stage_1__1998_, data_stage_1__1997_, data_stage_1__1996_, data_stage_1__1995_, data_stage_1__1994_, data_stage_1__1993_, data_stage_1__1992_, data_stage_1__1991_, data_stage_1__1990_, data_stage_1__1989_, data_stage_1__1988_, data_stage_1__1987_, data_stage_1__1986_, data_stage_1__1985_, data_stage_1__1984_, data_stage_1__1983_, data_stage_1__1982_, data_stage_1__1981_, data_stage_1__1980_, data_stage_1__1979_, data_stage_1__1978_, data_stage_1__1977_, data_stage_1__1976_, data_stage_1__1975_, data_stage_1__1974_, data_stage_1__1973_, data_stage_1__1972_, data_stage_1__1971_, data_stage_1__1970_, data_stage_1__1969_, data_stage_1__1968_, data_stage_1__1967_, data_stage_1__1966_, data_stage_1__1965_, data_stage_1__1964_, data_stage_1__1963_, data_stage_1__1962_, data_stage_1__1961_, data_stage_1__1960_, data_stage_1__1959_, data_stage_1__1958_, data_stage_1__1957_, data_stage_1__1956_, data_stage_1__1955_, data_stage_1__1954_, data_stage_1__1953_, data_stage_1__1952_, data_stage_1__1951_, data_stage_1__1950_, data_stage_1__1949_, data_stage_1__1948_, data_stage_1__1947_, data_stage_1__1946_, data_stage_1__1945_, data_stage_1__1944_, data_stage_1__1943_, data_stage_1__1942_, data_stage_1__1941_, data_stage_1__1940_, data_stage_1__1939_, data_stage_1__1938_, data_stage_1__1937_, data_stage_1__1936_, data_stage_1__1935_, data_stage_1__1934_, data_stage_1__1933_, data_stage_1__1932_, data_stage_1__1931_, data_stage_1__1930_, data_stage_1__1929_, data_stage_1__1928_, data_stage_1__1927_, data_stage_1__1926_, data_stage_1__1925_, data_stage_1__1924_, data_stage_1__1923_, data_stage_1__1922_, data_stage_1__1921_, data_stage_1__1920_, data_stage_1__1919_, data_stage_1__1918_, data_stage_1__1917_, data_stage_1__1916_, data_stage_1__1915_, data_stage_1__1914_, data_stage_1__1913_, data_stage_1__1912_, data_stage_1__1911_, data_stage_1__1910_, data_stage_1__1909_, data_stage_1__1908_, data_stage_1__1907_, data_stage_1__1906_, data_stage_1__1905_, data_stage_1__1904_, data_stage_1__1903_, data_stage_1__1902_, data_stage_1__1901_, data_stage_1__1900_, data_stage_1__1899_, data_stage_1__1898_, data_stage_1__1897_, data_stage_1__1896_, data_stage_1__1895_, data_stage_1__1894_, data_stage_1__1893_, data_stage_1__1892_, data_stage_1__1891_, data_stage_1__1890_, data_stage_1__1889_, data_stage_1__1888_, data_stage_1__1887_, data_stage_1__1886_, data_stage_1__1885_, data_stage_1__1884_, data_stage_1__1883_, data_stage_1__1882_, data_stage_1__1881_, data_stage_1__1880_, data_stage_1__1879_, data_stage_1__1878_, data_stage_1__1877_, data_stage_1__1876_, data_stage_1__1875_, data_stage_1__1874_, data_stage_1__1873_, data_stage_1__1872_, data_stage_1__1871_, data_stage_1__1870_, data_stage_1__1869_, data_stage_1__1868_, data_stage_1__1867_, data_stage_1__1866_, data_stage_1__1865_, data_stage_1__1864_, data_stage_1__1863_, data_stage_1__1862_, data_stage_1__1861_, data_stage_1__1860_, data_stage_1__1859_, data_stage_1__1858_, data_stage_1__1857_, data_stage_1__1856_, data_stage_1__1855_, data_stage_1__1854_, data_stage_1__1853_, data_stage_1__1852_, data_stage_1__1851_, data_stage_1__1850_, data_stage_1__1849_, data_stage_1__1848_, data_stage_1__1847_, data_stage_1__1846_, data_stage_1__1845_, data_stage_1__1844_, data_stage_1__1843_, data_stage_1__1842_, data_stage_1__1841_, data_stage_1__1840_, data_stage_1__1839_, data_stage_1__1838_, data_stage_1__1837_, data_stage_1__1836_, data_stage_1__1835_, data_stage_1__1834_, data_stage_1__1833_, data_stage_1__1832_, data_stage_1__1831_, data_stage_1__1830_, data_stage_1__1829_, data_stage_1__1828_, data_stage_1__1827_, data_stage_1__1826_, data_stage_1__1825_, data_stage_1__1824_, data_stage_1__1823_, data_stage_1__1822_, data_stage_1__1821_, data_stage_1__1820_, data_stage_1__1819_, data_stage_1__1818_, data_stage_1__1817_, data_stage_1__1816_, data_stage_1__1815_, data_stage_1__1814_, data_stage_1__1813_, data_stage_1__1812_, data_stage_1__1811_, data_stage_1__1810_, data_stage_1__1809_, data_stage_1__1808_, data_stage_1__1807_, data_stage_1__1806_, data_stage_1__1805_, data_stage_1__1804_, data_stage_1__1803_, data_stage_1__1802_, data_stage_1__1801_, data_stage_1__1800_, data_stage_1__1799_, data_stage_1__1798_, data_stage_1__1797_, data_stage_1__1796_, data_stage_1__1795_, data_stage_1__1794_, data_stage_1__1793_, data_stage_1__1792_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__2047_, data_stage_2__2046_, data_stage_2__2045_, data_stage_2__2044_, data_stage_2__2043_, data_stage_2__2042_, data_stage_2__2041_, data_stage_2__2040_, data_stage_2__2039_, data_stage_2__2038_, data_stage_2__2037_, data_stage_2__2036_, data_stage_2__2035_, data_stage_2__2034_, data_stage_2__2033_, data_stage_2__2032_, data_stage_2__2031_, data_stage_2__2030_, data_stage_2__2029_, data_stage_2__2028_, data_stage_2__2027_, data_stage_2__2026_, data_stage_2__2025_, data_stage_2__2024_, data_stage_2__2023_, data_stage_2__2022_, data_stage_2__2021_, data_stage_2__2020_, data_stage_2__2019_, data_stage_2__2018_, data_stage_2__2017_, data_stage_2__2016_, data_stage_2__2015_, data_stage_2__2014_, data_stage_2__2013_, data_stage_2__2012_, data_stage_2__2011_, data_stage_2__2010_, data_stage_2__2009_, data_stage_2__2008_, data_stage_2__2007_, data_stage_2__2006_, data_stage_2__2005_, data_stage_2__2004_, data_stage_2__2003_, data_stage_2__2002_, data_stage_2__2001_, data_stage_2__2000_, data_stage_2__1999_, data_stage_2__1998_, data_stage_2__1997_, data_stage_2__1996_, data_stage_2__1995_, data_stage_2__1994_, data_stage_2__1993_, data_stage_2__1992_, data_stage_2__1991_, data_stage_2__1990_, data_stage_2__1989_, data_stage_2__1988_, data_stage_2__1987_, data_stage_2__1986_, data_stage_2__1985_, data_stage_2__1984_, data_stage_2__1983_, data_stage_2__1982_, data_stage_2__1981_, data_stage_2__1980_, data_stage_2__1979_, data_stage_2__1978_, data_stage_2__1977_, data_stage_2__1976_, data_stage_2__1975_, data_stage_2__1974_, data_stage_2__1973_, data_stage_2__1972_, data_stage_2__1971_, data_stage_2__1970_, data_stage_2__1969_, data_stage_2__1968_, data_stage_2__1967_, data_stage_2__1966_, data_stage_2__1965_, data_stage_2__1964_, data_stage_2__1963_, data_stage_2__1962_, data_stage_2__1961_, data_stage_2__1960_, data_stage_2__1959_, data_stage_2__1958_, data_stage_2__1957_, data_stage_2__1956_, data_stage_2__1955_, data_stage_2__1954_, data_stage_2__1953_, data_stage_2__1952_, data_stage_2__1951_, data_stage_2__1950_, data_stage_2__1949_, data_stage_2__1948_, data_stage_2__1947_, data_stage_2__1946_, data_stage_2__1945_, data_stage_2__1944_, data_stage_2__1943_, data_stage_2__1942_, data_stage_2__1941_, data_stage_2__1940_, data_stage_2__1939_, data_stage_2__1938_, data_stage_2__1937_, data_stage_2__1936_, data_stage_2__1935_, data_stage_2__1934_, data_stage_2__1933_, data_stage_2__1932_, data_stage_2__1931_, data_stage_2__1930_, data_stage_2__1929_, data_stage_2__1928_, data_stage_2__1927_, data_stage_2__1926_, data_stage_2__1925_, data_stage_2__1924_, data_stage_2__1923_, data_stage_2__1922_, data_stage_2__1921_, data_stage_2__1920_, data_stage_2__1919_, data_stage_2__1918_, data_stage_2__1917_, data_stage_2__1916_, data_stage_2__1915_, data_stage_2__1914_, data_stage_2__1913_, data_stage_2__1912_, data_stage_2__1911_, data_stage_2__1910_, data_stage_2__1909_, data_stage_2__1908_, data_stage_2__1907_, data_stage_2__1906_, data_stage_2__1905_, data_stage_2__1904_, data_stage_2__1903_, data_stage_2__1902_, data_stage_2__1901_, data_stage_2__1900_, data_stage_2__1899_, data_stage_2__1898_, data_stage_2__1897_, data_stage_2__1896_, data_stage_2__1895_, data_stage_2__1894_, data_stage_2__1893_, data_stage_2__1892_, data_stage_2__1891_, data_stage_2__1890_, data_stage_2__1889_, data_stage_2__1888_, data_stage_2__1887_, data_stage_2__1886_, data_stage_2__1885_, data_stage_2__1884_, data_stage_2__1883_, data_stage_2__1882_, data_stage_2__1881_, data_stage_2__1880_, data_stage_2__1879_, data_stage_2__1878_, data_stage_2__1877_, data_stage_2__1876_, data_stage_2__1875_, data_stage_2__1874_, data_stage_2__1873_, data_stage_2__1872_, data_stage_2__1871_, data_stage_2__1870_, data_stage_2__1869_, data_stage_2__1868_, data_stage_2__1867_, data_stage_2__1866_, data_stage_2__1865_, data_stage_2__1864_, data_stage_2__1863_, data_stage_2__1862_, data_stage_2__1861_, data_stage_2__1860_, data_stage_2__1859_, data_stage_2__1858_, data_stage_2__1857_, data_stage_2__1856_, data_stage_2__1855_, data_stage_2__1854_, data_stage_2__1853_, data_stage_2__1852_, data_stage_2__1851_, data_stage_2__1850_, data_stage_2__1849_, data_stage_2__1848_, data_stage_2__1847_, data_stage_2__1846_, data_stage_2__1845_, data_stage_2__1844_, data_stage_2__1843_, data_stage_2__1842_, data_stage_2__1841_, data_stage_2__1840_, data_stage_2__1839_, data_stage_2__1838_, data_stage_2__1837_, data_stage_2__1836_, data_stage_2__1835_, data_stage_2__1834_, data_stage_2__1833_, data_stage_2__1832_, data_stage_2__1831_, data_stage_2__1830_, data_stage_2__1829_, data_stage_2__1828_, data_stage_2__1827_, data_stage_2__1826_, data_stage_2__1825_, data_stage_2__1824_, data_stage_2__1823_, data_stage_2__1822_, data_stage_2__1821_, data_stage_2__1820_, data_stage_2__1819_, data_stage_2__1818_, data_stage_2__1817_, data_stage_2__1816_, data_stage_2__1815_, data_stage_2__1814_, data_stage_2__1813_, data_stage_2__1812_, data_stage_2__1811_, data_stage_2__1810_, data_stage_2__1809_, data_stage_2__1808_, data_stage_2__1807_, data_stage_2__1806_, data_stage_2__1805_, data_stage_2__1804_, data_stage_2__1803_, data_stage_2__1802_, data_stage_2__1801_, data_stage_2__1800_, data_stage_2__1799_, data_stage_2__1798_, data_stage_2__1797_, data_stage_2__1796_, data_stage_2__1795_, data_stage_2__1794_, data_stage_2__1793_, data_stage_2__1792_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_8__swap_inst
  (
    .data_i({ data_stage_1__2303_, data_stage_1__2302_, data_stage_1__2301_, data_stage_1__2300_, data_stage_1__2299_, data_stage_1__2298_, data_stage_1__2297_, data_stage_1__2296_, data_stage_1__2295_, data_stage_1__2294_, data_stage_1__2293_, data_stage_1__2292_, data_stage_1__2291_, data_stage_1__2290_, data_stage_1__2289_, data_stage_1__2288_, data_stage_1__2287_, data_stage_1__2286_, data_stage_1__2285_, data_stage_1__2284_, data_stage_1__2283_, data_stage_1__2282_, data_stage_1__2281_, data_stage_1__2280_, data_stage_1__2279_, data_stage_1__2278_, data_stage_1__2277_, data_stage_1__2276_, data_stage_1__2275_, data_stage_1__2274_, data_stage_1__2273_, data_stage_1__2272_, data_stage_1__2271_, data_stage_1__2270_, data_stage_1__2269_, data_stage_1__2268_, data_stage_1__2267_, data_stage_1__2266_, data_stage_1__2265_, data_stage_1__2264_, data_stage_1__2263_, data_stage_1__2262_, data_stage_1__2261_, data_stage_1__2260_, data_stage_1__2259_, data_stage_1__2258_, data_stage_1__2257_, data_stage_1__2256_, data_stage_1__2255_, data_stage_1__2254_, data_stage_1__2253_, data_stage_1__2252_, data_stage_1__2251_, data_stage_1__2250_, data_stage_1__2249_, data_stage_1__2248_, data_stage_1__2247_, data_stage_1__2246_, data_stage_1__2245_, data_stage_1__2244_, data_stage_1__2243_, data_stage_1__2242_, data_stage_1__2241_, data_stage_1__2240_, data_stage_1__2239_, data_stage_1__2238_, data_stage_1__2237_, data_stage_1__2236_, data_stage_1__2235_, data_stage_1__2234_, data_stage_1__2233_, data_stage_1__2232_, data_stage_1__2231_, data_stage_1__2230_, data_stage_1__2229_, data_stage_1__2228_, data_stage_1__2227_, data_stage_1__2226_, data_stage_1__2225_, data_stage_1__2224_, data_stage_1__2223_, data_stage_1__2222_, data_stage_1__2221_, data_stage_1__2220_, data_stage_1__2219_, data_stage_1__2218_, data_stage_1__2217_, data_stage_1__2216_, data_stage_1__2215_, data_stage_1__2214_, data_stage_1__2213_, data_stage_1__2212_, data_stage_1__2211_, data_stage_1__2210_, data_stage_1__2209_, data_stage_1__2208_, data_stage_1__2207_, data_stage_1__2206_, data_stage_1__2205_, data_stage_1__2204_, data_stage_1__2203_, data_stage_1__2202_, data_stage_1__2201_, data_stage_1__2200_, data_stage_1__2199_, data_stage_1__2198_, data_stage_1__2197_, data_stage_1__2196_, data_stage_1__2195_, data_stage_1__2194_, data_stage_1__2193_, data_stage_1__2192_, data_stage_1__2191_, data_stage_1__2190_, data_stage_1__2189_, data_stage_1__2188_, data_stage_1__2187_, data_stage_1__2186_, data_stage_1__2185_, data_stage_1__2184_, data_stage_1__2183_, data_stage_1__2182_, data_stage_1__2181_, data_stage_1__2180_, data_stage_1__2179_, data_stage_1__2178_, data_stage_1__2177_, data_stage_1__2176_, data_stage_1__2175_, data_stage_1__2174_, data_stage_1__2173_, data_stage_1__2172_, data_stage_1__2171_, data_stage_1__2170_, data_stage_1__2169_, data_stage_1__2168_, data_stage_1__2167_, data_stage_1__2166_, data_stage_1__2165_, data_stage_1__2164_, data_stage_1__2163_, data_stage_1__2162_, data_stage_1__2161_, data_stage_1__2160_, data_stage_1__2159_, data_stage_1__2158_, data_stage_1__2157_, data_stage_1__2156_, data_stage_1__2155_, data_stage_1__2154_, data_stage_1__2153_, data_stage_1__2152_, data_stage_1__2151_, data_stage_1__2150_, data_stage_1__2149_, data_stage_1__2148_, data_stage_1__2147_, data_stage_1__2146_, data_stage_1__2145_, data_stage_1__2144_, data_stage_1__2143_, data_stage_1__2142_, data_stage_1__2141_, data_stage_1__2140_, data_stage_1__2139_, data_stage_1__2138_, data_stage_1__2137_, data_stage_1__2136_, data_stage_1__2135_, data_stage_1__2134_, data_stage_1__2133_, data_stage_1__2132_, data_stage_1__2131_, data_stage_1__2130_, data_stage_1__2129_, data_stage_1__2128_, data_stage_1__2127_, data_stage_1__2126_, data_stage_1__2125_, data_stage_1__2124_, data_stage_1__2123_, data_stage_1__2122_, data_stage_1__2121_, data_stage_1__2120_, data_stage_1__2119_, data_stage_1__2118_, data_stage_1__2117_, data_stage_1__2116_, data_stage_1__2115_, data_stage_1__2114_, data_stage_1__2113_, data_stage_1__2112_, data_stage_1__2111_, data_stage_1__2110_, data_stage_1__2109_, data_stage_1__2108_, data_stage_1__2107_, data_stage_1__2106_, data_stage_1__2105_, data_stage_1__2104_, data_stage_1__2103_, data_stage_1__2102_, data_stage_1__2101_, data_stage_1__2100_, data_stage_1__2099_, data_stage_1__2098_, data_stage_1__2097_, data_stage_1__2096_, data_stage_1__2095_, data_stage_1__2094_, data_stage_1__2093_, data_stage_1__2092_, data_stage_1__2091_, data_stage_1__2090_, data_stage_1__2089_, data_stage_1__2088_, data_stage_1__2087_, data_stage_1__2086_, data_stage_1__2085_, data_stage_1__2084_, data_stage_1__2083_, data_stage_1__2082_, data_stage_1__2081_, data_stage_1__2080_, data_stage_1__2079_, data_stage_1__2078_, data_stage_1__2077_, data_stage_1__2076_, data_stage_1__2075_, data_stage_1__2074_, data_stage_1__2073_, data_stage_1__2072_, data_stage_1__2071_, data_stage_1__2070_, data_stage_1__2069_, data_stage_1__2068_, data_stage_1__2067_, data_stage_1__2066_, data_stage_1__2065_, data_stage_1__2064_, data_stage_1__2063_, data_stage_1__2062_, data_stage_1__2061_, data_stage_1__2060_, data_stage_1__2059_, data_stage_1__2058_, data_stage_1__2057_, data_stage_1__2056_, data_stage_1__2055_, data_stage_1__2054_, data_stage_1__2053_, data_stage_1__2052_, data_stage_1__2051_, data_stage_1__2050_, data_stage_1__2049_, data_stage_1__2048_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__2303_, data_stage_2__2302_, data_stage_2__2301_, data_stage_2__2300_, data_stage_2__2299_, data_stage_2__2298_, data_stage_2__2297_, data_stage_2__2296_, data_stage_2__2295_, data_stage_2__2294_, data_stage_2__2293_, data_stage_2__2292_, data_stage_2__2291_, data_stage_2__2290_, data_stage_2__2289_, data_stage_2__2288_, data_stage_2__2287_, data_stage_2__2286_, data_stage_2__2285_, data_stage_2__2284_, data_stage_2__2283_, data_stage_2__2282_, data_stage_2__2281_, data_stage_2__2280_, data_stage_2__2279_, data_stage_2__2278_, data_stage_2__2277_, data_stage_2__2276_, data_stage_2__2275_, data_stage_2__2274_, data_stage_2__2273_, data_stage_2__2272_, data_stage_2__2271_, data_stage_2__2270_, data_stage_2__2269_, data_stage_2__2268_, data_stage_2__2267_, data_stage_2__2266_, data_stage_2__2265_, data_stage_2__2264_, data_stage_2__2263_, data_stage_2__2262_, data_stage_2__2261_, data_stage_2__2260_, data_stage_2__2259_, data_stage_2__2258_, data_stage_2__2257_, data_stage_2__2256_, data_stage_2__2255_, data_stage_2__2254_, data_stage_2__2253_, data_stage_2__2252_, data_stage_2__2251_, data_stage_2__2250_, data_stage_2__2249_, data_stage_2__2248_, data_stage_2__2247_, data_stage_2__2246_, data_stage_2__2245_, data_stage_2__2244_, data_stage_2__2243_, data_stage_2__2242_, data_stage_2__2241_, data_stage_2__2240_, data_stage_2__2239_, data_stage_2__2238_, data_stage_2__2237_, data_stage_2__2236_, data_stage_2__2235_, data_stage_2__2234_, data_stage_2__2233_, data_stage_2__2232_, data_stage_2__2231_, data_stage_2__2230_, data_stage_2__2229_, data_stage_2__2228_, data_stage_2__2227_, data_stage_2__2226_, data_stage_2__2225_, data_stage_2__2224_, data_stage_2__2223_, data_stage_2__2222_, data_stage_2__2221_, data_stage_2__2220_, data_stage_2__2219_, data_stage_2__2218_, data_stage_2__2217_, data_stage_2__2216_, data_stage_2__2215_, data_stage_2__2214_, data_stage_2__2213_, data_stage_2__2212_, data_stage_2__2211_, data_stage_2__2210_, data_stage_2__2209_, data_stage_2__2208_, data_stage_2__2207_, data_stage_2__2206_, data_stage_2__2205_, data_stage_2__2204_, data_stage_2__2203_, data_stage_2__2202_, data_stage_2__2201_, data_stage_2__2200_, data_stage_2__2199_, data_stage_2__2198_, data_stage_2__2197_, data_stage_2__2196_, data_stage_2__2195_, data_stage_2__2194_, data_stage_2__2193_, data_stage_2__2192_, data_stage_2__2191_, data_stage_2__2190_, data_stage_2__2189_, data_stage_2__2188_, data_stage_2__2187_, data_stage_2__2186_, data_stage_2__2185_, data_stage_2__2184_, data_stage_2__2183_, data_stage_2__2182_, data_stage_2__2181_, data_stage_2__2180_, data_stage_2__2179_, data_stage_2__2178_, data_stage_2__2177_, data_stage_2__2176_, data_stage_2__2175_, data_stage_2__2174_, data_stage_2__2173_, data_stage_2__2172_, data_stage_2__2171_, data_stage_2__2170_, data_stage_2__2169_, data_stage_2__2168_, data_stage_2__2167_, data_stage_2__2166_, data_stage_2__2165_, data_stage_2__2164_, data_stage_2__2163_, data_stage_2__2162_, data_stage_2__2161_, data_stage_2__2160_, data_stage_2__2159_, data_stage_2__2158_, data_stage_2__2157_, data_stage_2__2156_, data_stage_2__2155_, data_stage_2__2154_, data_stage_2__2153_, data_stage_2__2152_, data_stage_2__2151_, data_stage_2__2150_, data_stage_2__2149_, data_stage_2__2148_, data_stage_2__2147_, data_stage_2__2146_, data_stage_2__2145_, data_stage_2__2144_, data_stage_2__2143_, data_stage_2__2142_, data_stage_2__2141_, data_stage_2__2140_, data_stage_2__2139_, data_stage_2__2138_, data_stage_2__2137_, data_stage_2__2136_, data_stage_2__2135_, data_stage_2__2134_, data_stage_2__2133_, data_stage_2__2132_, data_stage_2__2131_, data_stage_2__2130_, data_stage_2__2129_, data_stage_2__2128_, data_stage_2__2127_, data_stage_2__2126_, data_stage_2__2125_, data_stage_2__2124_, data_stage_2__2123_, data_stage_2__2122_, data_stage_2__2121_, data_stage_2__2120_, data_stage_2__2119_, data_stage_2__2118_, data_stage_2__2117_, data_stage_2__2116_, data_stage_2__2115_, data_stage_2__2114_, data_stage_2__2113_, data_stage_2__2112_, data_stage_2__2111_, data_stage_2__2110_, data_stage_2__2109_, data_stage_2__2108_, data_stage_2__2107_, data_stage_2__2106_, data_stage_2__2105_, data_stage_2__2104_, data_stage_2__2103_, data_stage_2__2102_, data_stage_2__2101_, data_stage_2__2100_, data_stage_2__2099_, data_stage_2__2098_, data_stage_2__2097_, data_stage_2__2096_, data_stage_2__2095_, data_stage_2__2094_, data_stage_2__2093_, data_stage_2__2092_, data_stage_2__2091_, data_stage_2__2090_, data_stage_2__2089_, data_stage_2__2088_, data_stage_2__2087_, data_stage_2__2086_, data_stage_2__2085_, data_stage_2__2084_, data_stage_2__2083_, data_stage_2__2082_, data_stage_2__2081_, data_stage_2__2080_, data_stage_2__2079_, data_stage_2__2078_, data_stage_2__2077_, data_stage_2__2076_, data_stage_2__2075_, data_stage_2__2074_, data_stage_2__2073_, data_stage_2__2072_, data_stage_2__2071_, data_stage_2__2070_, data_stage_2__2069_, data_stage_2__2068_, data_stage_2__2067_, data_stage_2__2066_, data_stage_2__2065_, data_stage_2__2064_, data_stage_2__2063_, data_stage_2__2062_, data_stage_2__2061_, data_stage_2__2060_, data_stage_2__2059_, data_stage_2__2058_, data_stage_2__2057_, data_stage_2__2056_, data_stage_2__2055_, data_stage_2__2054_, data_stage_2__2053_, data_stage_2__2052_, data_stage_2__2051_, data_stage_2__2050_, data_stage_2__2049_, data_stage_2__2048_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_9__swap_inst
  (
    .data_i({ data_stage_1__2559_, data_stage_1__2558_, data_stage_1__2557_, data_stage_1__2556_, data_stage_1__2555_, data_stage_1__2554_, data_stage_1__2553_, data_stage_1__2552_, data_stage_1__2551_, data_stage_1__2550_, data_stage_1__2549_, data_stage_1__2548_, data_stage_1__2547_, data_stage_1__2546_, data_stage_1__2545_, data_stage_1__2544_, data_stage_1__2543_, data_stage_1__2542_, data_stage_1__2541_, data_stage_1__2540_, data_stage_1__2539_, data_stage_1__2538_, data_stage_1__2537_, data_stage_1__2536_, data_stage_1__2535_, data_stage_1__2534_, data_stage_1__2533_, data_stage_1__2532_, data_stage_1__2531_, data_stage_1__2530_, data_stage_1__2529_, data_stage_1__2528_, data_stage_1__2527_, data_stage_1__2526_, data_stage_1__2525_, data_stage_1__2524_, data_stage_1__2523_, data_stage_1__2522_, data_stage_1__2521_, data_stage_1__2520_, data_stage_1__2519_, data_stage_1__2518_, data_stage_1__2517_, data_stage_1__2516_, data_stage_1__2515_, data_stage_1__2514_, data_stage_1__2513_, data_stage_1__2512_, data_stage_1__2511_, data_stage_1__2510_, data_stage_1__2509_, data_stage_1__2508_, data_stage_1__2507_, data_stage_1__2506_, data_stage_1__2505_, data_stage_1__2504_, data_stage_1__2503_, data_stage_1__2502_, data_stage_1__2501_, data_stage_1__2500_, data_stage_1__2499_, data_stage_1__2498_, data_stage_1__2497_, data_stage_1__2496_, data_stage_1__2495_, data_stage_1__2494_, data_stage_1__2493_, data_stage_1__2492_, data_stage_1__2491_, data_stage_1__2490_, data_stage_1__2489_, data_stage_1__2488_, data_stage_1__2487_, data_stage_1__2486_, data_stage_1__2485_, data_stage_1__2484_, data_stage_1__2483_, data_stage_1__2482_, data_stage_1__2481_, data_stage_1__2480_, data_stage_1__2479_, data_stage_1__2478_, data_stage_1__2477_, data_stage_1__2476_, data_stage_1__2475_, data_stage_1__2474_, data_stage_1__2473_, data_stage_1__2472_, data_stage_1__2471_, data_stage_1__2470_, data_stage_1__2469_, data_stage_1__2468_, data_stage_1__2467_, data_stage_1__2466_, data_stage_1__2465_, data_stage_1__2464_, data_stage_1__2463_, data_stage_1__2462_, data_stage_1__2461_, data_stage_1__2460_, data_stage_1__2459_, data_stage_1__2458_, data_stage_1__2457_, data_stage_1__2456_, data_stage_1__2455_, data_stage_1__2454_, data_stage_1__2453_, data_stage_1__2452_, data_stage_1__2451_, data_stage_1__2450_, data_stage_1__2449_, data_stage_1__2448_, data_stage_1__2447_, data_stage_1__2446_, data_stage_1__2445_, data_stage_1__2444_, data_stage_1__2443_, data_stage_1__2442_, data_stage_1__2441_, data_stage_1__2440_, data_stage_1__2439_, data_stage_1__2438_, data_stage_1__2437_, data_stage_1__2436_, data_stage_1__2435_, data_stage_1__2434_, data_stage_1__2433_, data_stage_1__2432_, data_stage_1__2431_, data_stage_1__2430_, data_stage_1__2429_, data_stage_1__2428_, data_stage_1__2427_, data_stage_1__2426_, data_stage_1__2425_, data_stage_1__2424_, data_stage_1__2423_, data_stage_1__2422_, data_stage_1__2421_, data_stage_1__2420_, data_stage_1__2419_, data_stage_1__2418_, data_stage_1__2417_, data_stage_1__2416_, data_stage_1__2415_, data_stage_1__2414_, data_stage_1__2413_, data_stage_1__2412_, data_stage_1__2411_, data_stage_1__2410_, data_stage_1__2409_, data_stage_1__2408_, data_stage_1__2407_, data_stage_1__2406_, data_stage_1__2405_, data_stage_1__2404_, data_stage_1__2403_, data_stage_1__2402_, data_stage_1__2401_, data_stage_1__2400_, data_stage_1__2399_, data_stage_1__2398_, data_stage_1__2397_, data_stage_1__2396_, data_stage_1__2395_, data_stage_1__2394_, data_stage_1__2393_, data_stage_1__2392_, data_stage_1__2391_, data_stage_1__2390_, data_stage_1__2389_, data_stage_1__2388_, data_stage_1__2387_, data_stage_1__2386_, data_stage_1__2385_, data_stage_1__2384_, data_stage_1__2383_, data_stage_1__2382_, data_stage_1__2381_, data_stage_1__2380_, data_stage_1__2379_, data_stage_1__2378_, data_stage_1__2377_, data_stage_1__2376_, data_stage_1__2375_, data_stage_1__2374_, data_stage_1__2373_, data_stage_1__2372_, data_stage_1__2371_, data_stage_1__2370_, data_stage_1__2369_, data_stage_1__2368_, data_stage_1__2367_, data_stage_1__2366_, data_stage_1__2365_, data_stage_1__2364_, data_stage_1__2363_, data_stage_1__2362_, data_stage_1__2361_, data_stage_1__2360_, data_stage_1__2359_, data_stage_1__2358_, data_stage_1__2357_, data_stage_1__2356_, data_stage_1__2355_, data_stage_1__2354_, data_stage_1__2353_, data_stage_1__2352_, data_stage_1__2351_, data_stage_1__2350_, data_stage_1__2349_, data_stage_1__2348_, data_stage_1__2347_, data_stage_1__2346_, data_stage_1__2345_, data_stage_1__2344_, data_stage_1__2343_, data_stage_1__2342_, data_stage_1__2341_, data_stage_1__2340_, data_stage_1__2339_, data_stage_1__2338_, data_stage_1__2337_, data_stage_1__2336_, data_stage_1__2335_, data_stage_1__2334_, data_stage_1__2333_, data_stage_1__2332_, data_stage_1__2331_, data_stage_1__2330_, data_stage_1__2329_, data_stage_1__2328_, data_stage_1__2327_, data_stage_1__2326_, data_stage_1__2325_, data_stage_1__2324_, data_stage_1__2323_, data_stage_1__2322_, data_stage_1__2321_, data_stage_1__2320_, data_stage_1__2319_, data_stage_1__2318_, data_stage_1__2317_, data_stage_1__2316_, data_stage_1__2315_, data_stage_1__2314_, data_stage_1__2313_, data_stage_1__2312_, data_stage_1__2311_, data_stage_1__2310_, data_stage_1__2309_, data_stage_1__2308_, data_stage_1__2307_, data_stage_1__2306_, data_stage_1__2305_, data_stage_1__2304_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__2559_, data_stage_2__2558_, data_stage_2__2557_, data_stage_2__2556_, data_stage_2__2555_, data_stage_2__2554_, data_stage_2__2553_, data_stage_2__2552_, data_stage_2__2551_, data_stage_2__2550_, data_stage_2__2549_, data_stage_2__2548_, data_stage_2__2547_, data_stage_2__2546_, data_stage_2__2545_, data_stage_2__2544_, data_stage_2__2543_, data_stage_2__2542_, data_stage_2__2541_, data_stage_2__2540_, data_stage_2__2539_, data_stage_2__2538_, data_stage_2__2537_, data_stage_2__2536_, data_stage_2__2535_, data_stage_2__2534_, data_stage_2__2533_, data_stage_2__2532_, data_stage_2__2531_, data_stage_2__2530_, data_stage_2__2529_, data_stage_2__2528_, data_stage_2__2527_, data_stage_2__2526_, data_stage_2__2525_, data_stage_2__2524_, data_stage_2__2523_, data_stage_2__2522_, data_stage_2__2521_, data_stage_2__2520_, data_stage_2__2519_, data_stage_2__2518_, data_stage_2__2517_, data_stage_2__2516_, data_stage_2__2515_, data_stage_2__2514_, data_stage_2__2513_, data_stage_2__2512_, data_stage_2__2511_, data_stage_2__2510_, data_stage_2__2509_, data_stage_2__2508_, data_stage_2__2507_, data_stage_2__2506_, data_stage_2__2505_, data_stage_2__2504_, data_stage_2__2503_, data_stage_2__2502_, data_stage_2__2501_, data_stage_2__2500_, data_stage_2__2499_, data_stage_2__2498_, data_stage_2__2497_, data_stage_2__2496_, data_stage_2__2495_, data_stage_2__2494_, data_stage_2__2493_, data_stage_2__2492_, data_stage_2__2491_, data_stage_2__2490_, data_stage_2__2489_, data_stage_2__2488_, data_stage_2__2487_, data_stage_2__2486_, data_stage_2__2485_, data_stage_2__2484_, data_stage_2__2483_, data_stage_2__2482_, data_stage_2__2481_, data_stage_2__2480_, data_stage_2__2479_, data_stage_2__2478_, data_stage_2__2477_, data_stage_2__2476_, data_stage_2__2475_, data_stage_2__2474_, data_stage_2__2473_, data_stage_2__2472_, data_stage_2__2471_, data_stage_2__2470_, data_stage_2__2469_, data_stage_2__2468_, data_stage_2__2467_, data_stage_2__2466_, data_stage_2__2465_, data_stage_2__2464_, data_stage_2__2463_, data_stage_2__2462_, data_stage_2__2461_, data_stage_2__2460_, data_stage_2__2459_, data_stage_2__2458_, data_stage_2__2457_, data_stage_2__2456_, data_stage_2__2455_, data_stage_2__2454_, data_stage_2__2453_, data_stage_2__2452_, data_stage_2__2451_, data_stage_2__2450_, data_stage_2__2449_, data_stage_2__2448_, data_stage_2__2447_, data_stage_2__2446_, data_stage_2__2445_, data_stage_2__2444_, data_stage_2__2443_, data_stage_2__2442_, data_stage_2__2441_, data_stage_2__2440_, data_stage_2__2439_, data_stage_2__2438_, data_stage_2__2437_, data_stage_2__2436_, data_stage_2__2435_, data_stage_2__2434_, data_stage_2__2433_, data_stage_2__2432_, data_stage_2__2431_, data_stage_2__2430_, data_stage_2__2429_, data_stage_2__2428_, data_stage_2__2427_, data_stage_2__2426_, data_stage_2__2425_, data_stage_2__2424_, data_stage_2__2423_, data_stage_2__2422_, data_stage_2__2421_, data_stage_2__2420_, data_stage_2__2419_, data_stage_2__2418_, data_stage_2__2417_, data_stage_2__2416_, data_stage_2__2415_, data_stage_2__2414_, data_stage_2__2413_, data_stage_2__2412_, data_stage_2__2411_, data_stage_2__2410_, data_stage_2__2409_, data_stage_2__2408_, data_stage_2__2407_, data_stage_2__2406_, data_stage_2__2405_, data_stage_2__2404_, data_stage_2__2403_, data_stage_2__2402_, data_stage_2__2401_, data_stage_2__2400_, data_stage_2__2399_, data_stage_2__2398_, data_stage_2__2397_, data_stage_2__2396_, data_stage_2__2395_, data_stage_2__2394_, data_stage_2__2393_, data_stage_2__2392_, data_stage_2__2391_, data_stage_2__2390_, data_stage_2__2389_, data_stage_2__2388_, data_stage_2__2387_, data_stage_2__2386_, data_stage_2__2385_, data_stage_2__2384_, data_stage_2__2383_, data_stage_2__2382_, data_stage_2__2381_, data_stage_2__2380_, data_stage_2__2379_, data_stage_2__2378_, data_stage_2__2377_, data_stage_2__2376_, data_stage_2__2375_, data_stage_2__2374_, data_stage_2__2373_, data_stage_2__2372_, data_stage_2__2371_, data_stage_2__2370_, data_stage_2__2369_, data_stage_2__2368_, data_stage_2__2367_, data_stage_2__2366_, data_stage_2__2365_, data_stage_2__2364_, data_stage_2__2363_, data_stage_2__2362_, data_stage_2__2361_, data_stage_2__2360_, data_stage_2__2359_, data_stage_2__2358_, data_stage_2__2357_, data_stage_2__2356_, data_stage_2__2355_, data_stage_2__2354_, data_stage_2__2353_, data_stage_2__2352_, data_stage_2__2351_, data_stage_2__2350_, data_stage_2__2349_, data_stage_2__2348_, data_stage_2__2347_, data_stage_2__2346_, data_stage_2__2345_, data_stage_2__2344_, data_stage_2__2343_, data_stage_2__2342_, data_stage_2__2341_, data_stage_2__2340_, data_stage_2__2339_, data_stage_2__2338_, data_stage_2__2337_, data_stage_2__2336_, data_stage_2__2335_, data_stage_2__2334_, data_stage_2__2333_, data_stage_2__2332_, data_stage_2__2331_, data_stage_2__2330_, data_stage_2__2329_, data_stage_2__2328_, data_stage_2__2327_, data_stage_2__2326_, data_stage_2__2325_, data_stage_2__2324_, data_stage_2__2323_, data_stage_2__2322_, data_stage_2__2321_, data_stage_2__2320_, data_stage_2__2319_, data_stage_2__2318_, data_stage_2__2317_, data_stage_2__2316_, data_stage_2__2315_, data_stage_2__2314_, data_stage_2__2313_, data_stage_2__2312_, data_stage_2__2311_, data_stage_2__2310_, data_stage_2__2309_, data_stage_2__2308_, data_stage_2__2307_, data_stage_2__2306_, data_stage_2__2305_, data_stage_2__2304_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_10__swap_inst
  (
    .data_i({ data_stage_1__2815_, data_stage_1__2814_, data_stage_1__2813_, data_stage_1__2812_, data_stage_1__2811_, data_stage_1__2810_, data_stage_1__2809_, data_stage_1__2808_, data_stage_1__2807_, data_stage_1__2806_, data_stage_1__2805_, data_stage_1__2804_, data_stage_1__2803_, data_stage_1__2802_, data_stage_1__2801_, data_stage_1__2800_, data_stage_1__2799_, data_stage_1__2798_, data_stage_1__2797_, data_stage_1__2796_, data_stage_1__2795_, data_stage_1__2794_, data_stage_1__2793_, data_stage_1__2792_, data_stage_1__2791_, data_stage_1__2790_, data_stage_1__2789_, data_stage_1__2788_, data_stage_1__2787_, data_stage_1__2786_, data_stage_1__2785_, data_stage_1__2784_, data_stage_1__2783_, data_stage_1__2782_, data_stage_1__2781_, data_stage_1__2780_, data_stage_1__2779_, data_stage_1__2778_, data_stage_1__2777_, data_stage_1__2776_, data_stage_1__2775_, data_stage_1__2774_, data_stage_1__2773_, data_stage_1__2772_, data_stage_1__2771_, data_stage_1__2770_, data_stage_1__2769_, data_stage_1__2768_, data_stage_1__2767_, data_stage_1__2766_, data_stage_1__2765_, data_stage_1__2764_, data_stage_1__2763_, data_stage_1__2762_, data_stage_1__2761_, data_stage_1__2760_, data_stage_1__2759_, data_stage_1__2758_, data_stage_1__2757_, data_stage_1__2756_, data_stage_1__2755_, data_stage_1__2754_, data_stage_1__2753_, data_stage_1__2752_, data_stage_1__2751_, data_stage_1__2750_, data_stage_1__2749_, data_stage_1__2748_, data_stage_1__2747_, data_stage_1__2746_, data_stage_1__2745_, data_stage_1__2744_, data_stage_1__2743_, data_stage_1__2742_, data_stage_1__2741_, data_stage_1__2740_, data_stage_1__2739_, data_stage_1__2738_, data_stage_1__2737_, data_stage_1__2736_, data_stage_1__2735_, data_stage_1__2734_, data_stage_1__2733_, data_stage_1__2732_, data_stage_1__2731_, data_stage_1__2730_, data_stage_1__2729_, data_stage_1__2728_, data_stage_1__2727_, data_stage_1__2726_, data_stage_1__2725_, data_stage_1__2724_, data_stage_1__2723_, data_stage_1__2722_, data_stage_1__2721_, data_stage_1__2720_, data_stage_1__2719_, data_stage_1__2718_, data_stage_1__2717_, data_stage_1__2716_, data_stage_1__2715_, data_stage_1__2714_, data_stage_1__2713_, data_stage_1__2712_, data_stage_1__2711_, data_stage_1__2710_, data_stage_1__2709_, data_stage_1__2708_, data_stage_1__2707_, data_stage_1__2706_, data_stage_1__2705_, data_stage_1__2704_, data_stage_1__2703_, data_stage_1__2702_, data_stage_1__2701_, data_stage_1__2700_, data_stage_1__2699_, data_stage_1__2698_, data_stage_1__2697_, data_stage_1__2696_, data_stage_1__2695_, data_stage_1__2694_, data_stage_1__2693_, data_stage_1__2692_, data_stage_1__2691_, data_stage_1__2690_, data_stage_1__2689_, data_stage_1__2688_, data_stage_1__2687_, data_stage_1__2686_, data_stage_1__2685_, data_stage_1__2684_, data_stage_1__2683_, data_stage_1__2682_, data_stage_1__2681_, data_stage_1__2680_, data_stage_1__2679_, data_stage_1__2678_, data_stage_1__2677_, data_stage_1__2676_, data_stage_1__2675_, data_stage_1__2674_, data_stage_1__2673_, data_stage_1__2672_, data_stage_1__2671_, data_stage_1__2670_, data_stage_1__2669_, data_stage_1__2668_, data_stage_1__2667_, data_stage_1__2666_, data_stage_1__2665_, data_stage_1__2664_, data_stage_1__2663_, data_stage_1__2662_, data_stage_1__2661_, data_stage_1__2660_, data_stage_1__2659_, data_stage_1__2658_, data_stage_1__2657_, data_stage_1__2656_, data_stage_1__2655_, data_stage_1__2654_, data_stage_1__2653_, data_stage_1__2652_, data_stage_1__2651_, data_stage_1__2650_, data_stage_1__2649_, data_stage_1__2648_, data_stage_1__2647_, data_stage_1__2646_, data_stage_1__2645_, data_stage_1__2644_, data_stage_1__2643_, data_stage_1__2642_, data_stage_1__2641_, data_stage_1__2640_, data_stage_1__2639_, data_stage_1__2638_, data_stage_1__2637_, data_stage_1__2636_, data_stage_1__2635_, data_stage_1__2634_, data_stage_1__2633_, data_stage_1__2632_, data_stage_1__2631_, data_stage_1__2630_, data_stage_1__2629_, data_stage_1__2628_, data_stage_1__2627_, data_stage_1__2626_, data_stage_1__2625_, data_stage_1__2624_, data_stage_1__2623_, data_stage_1__2622_, data_stage_1__2621_, data_stage_1__2620_, data_stage_1__2619_, data_stage_1__2618_, data_stage_1__2617_, data_stage_1__2616_, data_stage_1__2615_, data_stage_1__2614_, data_stage_1__2613_, data_stage_1__2612_, data_stage_1__2611_, data_stage_1__2610_, data_stage_1__2609_, data_stage_1__2608_, data_stage_1__2607_, data_stage_1__2606_, data_stage_1__2605_, data_stage_1__2604_, data_stage_1__2603_, data_stage_1__2602_, data_stage_1__2601_, data_stage_1__2600_, data_stage_1__2599_, data_stage_1__2598_, data_stage_1__2597_, data_stage_1__2596_, data_stage_1__2595_, data_stage_1__2594_, data_stage_1__2593_, data_stage_1__2592_, data_stage_1__2591_, data_stage_1__2590_, data_stage_1__2589_, data_stage_1__2588_, data_stage_1__2587_, data_stage_1__2586_, data_stage_1__2585_, data_stage_1__2584_, data_stage_1__2583_, data_stage_1__2582_, data_stage_1__2581_, data_stage_1__2580_, data_stage_1__2579_, data_stage_1__2578_, data_stage_1__2577_, data_stage_1__2576_, data_stage_1__2575_, data_stage_1__2574_, data_stage_1__2573_, data_stage_1__2572_, data_stage_1__2571_, data_stage_1__2570_, data_stage_1__2569_, data_stage_1__2568_, data_stage_1__2567_, data_stage_1__2566_, data_stage_1__2565_, data_stage_1__2564_, data_stage_1__2563_, data_stage_1__2562_, data_stage_1__2561_, data_stage_1__2560_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__2815_, data_stage_2__2814_, data_stage_2__2813_, data_stage_2__2812_, data_stage_2__2811_, data_stage_2__2810_, data_stage_2__2809_, data_stage_2__2808_, data_stage_2__2807_, data_stage_2__2806_, data_stage_2__2805_, data_stage_2__2804_, data_stage_2__2803_, data_stage_2__2802_, data_stage_2__2801_, data_stage_2__2800_, data_stage_2__2799_, data_stage_2__2798_, data_stage_2__2797_, data_stage_2__2796_, data_stage_2__2795_, data_stage_2__2794_, data_stage_2__2793_, data_stage_2__2792_, data_stage_2__2791_, data_stage_2__2790_, data_stage_2__2789_, data_stage_2__2788_, data_stage_2__2787_, data_stage_2__2786_, data_stage_2__2785_, data_stage_2__2784_, data_stage_2__2783_, data_stage_2__2782_, data_stage_2__2781_, data_stage_2__2780_, data_stage_2__2779_, data_stage_2__2778_, data_stage_2__2777_, data_stage_2__2776_, data_stage_2__2775_, data_stage_2__2774_, data_stage_2__2773_, data_stage_2__2772_, data_stage_2__2771_, data_stage_2__2770_, data_stage_2__2769_, data_stage_2__2768_, data_stage_2__2767_, data_stage_2__2766_, data_stage_2__2765_, data_stage_2__2764_, data_stage_2__2763_, data_stage_2__2762_, data_stage_2__2761_, data_stage_2__2760_, data_stage_2__2759_, data_stage_2__2758_, data_stage_2__2757_, data_stage_2__2756_, data_stage_2__2755_, data_stage_2__2754_, data_stage_2__2753_, data_stage_2__2752_, data_stage_2__2751_, data_stage_2__2750_, data_stage_2__2749_, data_stage_2__2748_, data_stage_2__2747_, data_stage_2__2746_, data_stage_2__2745_, data_stage_2__2744_, data_stage_2__2743_, data_stage_2__2742_, data_stage_2__2741_, data_stage_2__2740_, data_stage_2__2739_, data_stage_2__2738_, data_stage_2__2737_, data_stage_2__2736_, data_stage_2__2735_, data_stage_2__2734_, data_stage_2__2733_, data_stage_2__2732_, data_stage_2__2731_, data_stage_2__2730_, data_stage_2__2729_, data_stage_2__2728_, data_stage_2__2727_, data_stage_2__2726_, data_stage_2__2725_, data_stage_2__2724_, data_stage_2__2723_, data_stage_2__2722_, data_stage_2__2721_, data_stage_2__2720_, data_stage_2__2719_, data_stage_2__2718_, data_stage_2__2717_, data_stage_2__2716_, data_stage_2__2715_, data_stage_2__2714_, data_stage_2__2713_, data_stage_2__2712_, data_stage_2__2711_, data_stage_2__2710_, data_stage_2__2709_, data_stage_2__2708_, data_stage_2__2707_, data_stage_2__2706_, data_stage_2__2705_, data_stage_2__2704_, data_stage_2__2703_, data_stage_2__2702_, data_stage_2__2701_, data_stage_2__2700_, data_stage_2__2699_, data_stage_2__2698_, data_stage_2__2697_, data_stage_2__2696_, data_stage_2__2695_, data_stage_2__2694_, data_stage_2__2693_, data_stage_2__2692_, data_stage_2__2691_, data_stage_2__2690_, data_stage_2__2689_, data_stage_2__2688_, data_stage_2__2687_, data_stage_2__2686_, data_stage_2__2685_, data_stage_2__2684_, data_stage_2__2683_, data_stage_2__2682_, data_stage_2__2681_, data_stage_2__2680_, data_stage_2__2679_, data_stage_2__2678_, data_stage_2__2677_, data_stage_2__2676_, data_stage_2__2675_, data_stage_2__2674_, data_stage_2__2673_, data_stage_2__2672_, data_stage_2__2671_, data_stage_2__2670_, data_stage_2__2669_, data_stage_2__2668_, data_stage_2__2667_, data_stage_2__2666_, data_stage_2__2665_, data_stage_2__2664_, data_stage_2__2663_, data_stage_2__2662_, data_stage_2__2661_, data_stage_2__2660_, data_stage_2__2659_, data_stage_2__2658_, data_stage_2__2657_, data_stage_2__2656_, data_stage_2__2655_, data_stage_2__2654_, data_stage_2__2653_, data_stage_2__2652_, data_stage_2__2651_, data_stage_2__2650_, data_stage_2__2649_, data_stage_2__2648_, data_stage_2__2647_, data_stage_2__2646_, data_stage_2__2645_, data_stage_2__2644_, data_stage_2__2643_, data_stage_2__2642_, data_stage_2__2641_, data_stage_2__2640_, data_stage_2__2639_, data_stage_2__2638_, data_stage_2__2637_, data_stage_2__2636_, data_stage_2__2635_, data_stage_2__2634_, data_stage_2__2633_, data_stage_2__2632_, data_stage_2__2631_, data_stage_2__2630_, data_stage_2__2629_, data_stage_2__2628_, data_stage_2__2627_, data_stage_2__2626_, data_stage_2__2625_, data_stage_2__2624_, data_stage_2__2623_, data_stage_2__2622_, data_stage_2__2621_, data_stage_2__2620_, data_stage_2__2619_, data_stage_2__2618_, data_stage_2__2617_, data_stage_2__2616_, data_stage_2__2615_, data_stage_2__2614_, data_stage_2__2613_, data_stage_2__2612_, data_stage_2__2611_, data_stage_2__2610_, data_stage_2__2609_, data_stage_2__2608_, data_stage_2__2607_, data_stage_2__2606_, data_stage_2__2605_, data_stage_2__2604_, data_stage_2__2603_, data_stage_2__2602_, data_stage_2__2601_, data_stage_2__2600_, data_stage_2__2599_, data_stage_2__2598_, data_stage_2__2597_, data_stage_2__2596_, data_stage_2__2595_, data_stage_2__2594_, data_stage_2__2593_, data_stage_2__2592_, data_stage_2__2591_, data_stage_2__2590_, data_stage_2__2589_, data_stage_2__2588_, data_stage_2__2587_, data_stage_2__2586_, data_stage_2__2585_, data_stage_2__2584_, data_stage_2__2583_, data_stage_2__2582_, data_stage_2__2581_, data_stage_2__2580_, data_stage_2__2579_, data_stage_2__2578_, data_stage_2__2577_, data_stage_2__2576_, data_stage_2__2575_, data_stage_2__2574_, data_stage_2__2573_, data_stage_2__2572_, data_stage_2__2571_, data_stage_2__2570_, data_stage_2__2569_, data_stage_2__2568_, data_stage_2__2567_, data_stage_2__2566_, data_stage_2__2565_, data_stage_2__2564_, data_stage_2__2563_, data_stage_2__2562_, data_stage_2__2561_, data_stage_2__2560_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_11__swap_inst
  (
    .data_i({ data_stage_1__3071_, data_stage_1__3070_, data_stage_1__3069_, data_stage_1__3068_, data_stage_1__3067_, data_stage_1__3066_, data_stage_1__3065_, data_stage_1__3064_, data_stage_1__3063_, data_stage_1__3062_, data_stage_1__3061_, data_stage_1__3060_, data_stage_1__3059_, data_stage_1__3058_, data_stage_1__3057_, data_stage_1__3056_, data_stage_1__3055_, data_stage_1__3054_, data_stage_1__3053_, data_stage_1__3052_, data_stage_1__3051_, data_stage_1__3050_, data_stage_1__3049_, data_stage_1__3048_, data_stage_1__3047_, data_stage_1__3046_, data_stage_1__3045_, data_stage_1__3044_, data_stage_1__3043_, data_stage_1__3042_, data_stage_1__3041_, data_stage_1__3040_, data_stage_1__3039_, data_stage_1__3038_, data_stage_1__3037_, data_stage_1__3036_, data_stage_1__3035_, data_stage_1__3034_, data_stage_1__3033_, data_stage_1__3032_, data_stage_1__3031_, data_stage_1__3030_, data_stage_1__3029_, data_stage_1__3028_, data_stage_1__3027_, data_stage_1__3026_, data_stage_1__3025_, data_stage_1__3024_, data_stage_1__3023_, data_stage_1__3022_, data_stage_1__3021_, data_stage_1__3020_, data_stage_1__3019_, data_stage_1__3018_, data_stage_1__3017_, data_stage_1__3016_, data_stage_1__3015_, data_stage_1__3014_, data_stage_1__3013_, data_stage_1__3012_, data_stage_1__3011_, data_stage_1__3010_, data_stage_1__3009_, data_stage_1__3008_, data_stage_1__3007_, data_stage_1__3006_, data_stage_1__3005_, data_stage_1__3004_, data_stage_1__3003_, data_stage_1__3002_, data_stage_1__3001_, data_stage_1__3000_, data_stage_1__2999_, data_stage_1__2998_, data_stage_1__2997_, data_stage_1__2996_, data_stage_1__2995_, data_stage_1__2994_, data_stage_1__2993_, data_stage_1__2992_, data_stage_1__2991_, data_stage_1__2990_, data_stage_1__2989_, data_stage_1__2988_, data_stage_1__2987_, data_stage_1__2986_, data_stage_1__2985_, data_stage_1__2984_, data_stage_1__2983_, data_stage_1__2982_, data_stage_1__2981_, data_stage_1__2980_, data_stage_1__2979_, data_stage_1__2978_, data_stage_1__2977_, data_stage_1__2976_, data_stage_1__2975_, data_stage_1__2974_, data_stage_1__2973_, data_stage_1__2972_, data_stage_1__2971_, data_stage_1__2970_, data_stage_1__2969_, data_stage_1__2968_, data_stage_1__2967_, data_stage_1__2966_, data_stage_1__2965_, data_stage_1__2964_, data_stage_1__2963_, data_stage_1__2962_, data_stage_1__2961_, data_stage_1__2960_, data_stage_1__2959_, data_stage_1__2958_, data_stage_1__2957_, data_stage_1__2956_, data_stage_1__2955_, data_stage_1__2954_, data_stage_1__2953_, data_stage_1__2952_, data_stage_1__2951_, data_stage_1__2950_, data_stage_1__2949_, data_stage_1__2948_, data_stage_1__2947_, data_stage_1__2946_, data_stage_1__2945_, data_stage_1__2944_, data_stage_1__2943_, data_stage_1__2942_, data_stage_1__2941_, data_stage_1__2940_, data_stage_1__2939_, data_stage_1__2938_, data_stage_1__2937_, data_stage_1__2936_, data_stage_1__2935_, data_stage_1__2934_, data_stage_1__2933_, data_stage_1__2932_, data_stage_1__2931_, data_stage_1__2930_, data_stage_1__2929_, data_stage_1__2928_, data_stage_1__2927_, data_stage_1__2926_, data_stage_1__2925_, data_stage_1__2924_, data_stage_1__2923_, data_stage_1__2922_, data_stage_1__2921_, data_stage_1__2920_, data_stage_1__2919_, data_stage_1__2918_, data_stage_1__2917_, data_stage_1__2916_, data_stage_1__2915_, data_stage_1__2914_, data_stage_1__2913_, data_stage_1__2912_, data_stage_1__2911_, data_stage_1__2910_, data_stage_1__2909_, data_stage_1__2908_, data_stage_1__2907_, data_stage_1__2906_, data_stage_1__2905_, data_stage_1__2904_, data_stage_1__2903_, data_stage_1__2902_, data_stage_1__2901_, data_stage_1__2900_, data_stage_1__2899_, data_stage_1__2898_, data_stage_1__2897_, data_stage_1__2896_, data_stage_1__2895_, data_stage_1__2894_, data_stage_1__2893_, data_stage_1__2892_, data_stage_1__2891_, data_stage_1__2890_, data_stage_1__2889_, data_stage_1__2888_, data_stage_1__2887_, data_stage_1__2886_, data_stage_1__2885_, data_stage_1__2884_, data_stage_1__2883_, data_stage_1__2882_, data_stage_1__2881_, data_stage_1__2880_, data_stage_1__2879_, data_stage_1__2878_, data_stage_1__2877_, data_stage_1__2876_, data_stage_1__2875_, data_stage_1__2874_, data_stage_1__2873_, data_stage_1__2872_, data_stage_1__2871_, data_stage_1__2870_, data_stage_1__2869_, data_stage_1__2868_, data_stage_1__2867_, data_stage_1__2866_, data_stage_1__2865_, data_stage_1__2864_, data_stage_1__2863_, data_stage_1__2862_, data_stage_1__2861_, data_stage_1__2860_, data_stage_1__2859_, data_stage_1__2858_, data_stage_1__2857_, data_stage_1__2856_, data_stage_1__2855_, data_stage_1__2854_, data_stage_1__2853_, data_stage_1__2852_, data_stage_1__2851_, data_stage_1__2850_, data_stage_1__2849_, data_stage_1__2848_, data_stage_1__2847_, data_stage_1__2846_, data_stage_1__2845_, data_stage_1__2844_, data_stage_1__2843_, data_stage_1__2842_, data_stage_1__2841_, data_stage_1__2840_, data_stage_1__2839_, data_stage_1__2838_, data_stage_1__2837_, data_stage_1__2836_, data_stage_1__2835_, data_stage_1__2834_, data_stage_1__2833_, data_stage_1__2832_, data_stage_1__2831_, data_stage_1__2830_, data_stage_1__2829_, data_stage_1__2828_, data_stage_1__2827_, data_stage_1__2826_, data_stage_1__2825_, data_stage_1__2824_, data_stage_1__2823_, data_stage_1__2822_, data_stage_1__2821_, data_stage_1__2820_, data_stage_1__2819_, data_stage_1__2818_, data_stage_1__2817_, data_stage_1__2816_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__3071_, data_stage_2__3070_, data_stage_2__3069_, data_stage_2__3068_, data_stage_2__3067_, data_stage_2__3066_, data_stage_2__3065_, data_stage_2__3064_, data_stage_2__3063_, data_stage_2__3062_, data_stage_2__3061_, data_stage_2__3060_, data_stage_2__3059_, data_stage_2__3058_, data_stage_2__3057_, data_stage_2__3056_, data_stage_2__3055_, data_stage_2__3054_, data_stage_2__3053_, data_stage_2__3052_, data_stage_2__3051_, data_stage_2__3050_, data_stage_2__3049_, data_stage_2__3048_, data_stage_2__3047_, data_stage_2__3046_, data_stage_2__3045_, data_stage_2__3044_, data_stage_2__3043_, data_stage_2__3042_, data_stage_2__3041_, data_stage_2__3040_, data_stage_2__3039_, data_stage_2__3038_, data_stage_2__3037_, data_stage_2__3036_, data_stage_2__3035_, data_stage_2__3034_, data_stage_2__3033_, data_stage_2__3032_, data_stage_2__3031_, data_stage_2__3030_, data_stage_2__3029_, data_stage_2__3028_, data_stage_2__3027_, data_stage_2__3026_, data_stage_2__3025_, data_stage_2__3024_, data_stage_2__3023_, data_stage_2__3022_, data_stage_2__3021_, data_stage_2__3020_, data_stage_2__3019_, data_stage_2__3018_, data_stage_2__3017_, data_stage_2__3016_, data_stage_2__3015_, data_stage_2__3014_, data_stage_2__3013_, data_stage_2__3012_, data_stage_2__3011_, data_stage_2__3010_, data_stage_2__3009_, data_stage_2__3008_, data_stage_2__3007_, data_stage_2__3006_, data_stage_2__3005_, data_stage_2__3004_, data_stage_2__3003_, data_stage_2__3002_, data_stage_2__3001_, data_stage_2__3000_, data_stage_2__2999_, data_stage_2__2998_, data_stage_2__2997_, data_stage_2__2996_, data_stage_2__2995_, data_stage_2__2994_, data_stage_2__2993_, data_stage_2__2992_, data_stage_2__2991_, data_stage_2__2990_, data_stage_2__2989_, data_stage_2__2988_, data_stage_2__2987_, data_stage_2__2986_, data_stage_2__2985_, data_stage_2__2984_, data_stage_2__2983_, data_stage_2__2982_, data_stage_2__2981_, data_stage_2__2980_, data_stage_2__2979_, data_stage_2__2978_, data_stage_2__2977_, data_stage_2__2976_, data_stage_2__2975_, data_stage_2__2974_, data_stage_2__2973_, data_stage_2__2972_, data_stage_2__2971_, data_stage_2__2970_, data_stage_2__2969_, data_stage_2__2968_, data_stage_2__2967_, data_stage_2__2966_, data_stage_2__2965_, data_stage_2__2964_, data_stage_2__2963_, data_stage_2__2962_, data_stage_2__2961_, data_stage_2__2960_, data_stage_2__2959_, data_stage_2__2958_, data_stage_2__2957_, data_stage_2__2956_, data_stage_2__2955_, data_stage_2__2954_, data_stage_2__2953_, data_stage_2__2952_, data_stage_2__2951_, data_stage_2__2950_, data_stage_2__2949_, data_stage_2__2948_, data_stage_2__2947_, data_stage_2__2946_, data_stage_2__2945_, data_stage_2__2944_, data_stage_2__2943_, data_stage_2__2942_, data_stage_2__2941_, data_stage_2__2940_, data_stage_2__2939_, data_stage_2__2938_, data_stage_2__2937_, data_stage_2__2936_, data_stage_2__2935_, data_stage_2__2934_, data_stage_2__2933_, data_stage_2__2932_, data_stage_2__2931_, data_stage_2__2930_, data_stage_2__2929_, data_stage_2__2928_, data_stage_2__2927_, data_stage_2__2926_, data_stage_2__2925_, data_stage_2__2924_, data_stage_2__2923_, data_stage_2__2922_, data_stage_2__2921_, data_stage_2__2920_, data_stage_2__2919_, data_stage_2__2918_, data_stage_2__2917_, data_stage_2__2916_, data_stage_2__2915_, data_stage_2__2914_, data_stage_2__2913_, data_stage_2__2912_, data_stage_2__2911_, data_stage_2__2910_, data_stage_2__2909_, data_stage_2__2908_, data_stage_2__2907_, data_stage_2__2906_, data_stage_2__2905_, data_stage_2__2904_, data_stage_2__2903_, data_stage_2__2902_, data_stage_2__2901_, data_stage_2__2900_, data_stage_2__2899_, data_stage_2__2898_, data_stage_2__2897_, data_stage_2__2896_, data_stage_2__2895_, data_stage_2__2894_, data_stage_2__2893_, data_stage_2__2892_, data_stage_2__2891_, data_stage_2__2890_, data_stage_2__2889_, data_stage_2__2888_, data_stage_2__2887_, data_stage_2__2886_, data_stage_2__2885_, data_stage_2__2884_, data_stage_2__2883_, data_stage_2__2882_, data_stage_2__2881_, data_stage_2__2880_, data_stage_2__2879_, data_stage_2__2878_, data_stage_2__2877_, data_stage_2__2876_, data_stage_2__2875_, data_stage_2__2874_, data_stage_2__2873_, data_stage_2__2872_, data_stage_2__2871_, data_stage_2__2870_, data_stage_2__2869_, data_stage_2__2868_, data_stage_2__2867_, data_stage_2__2866_, data_stage_2__2865_, data_stage_2__2864_, data_stage_2__2863_, data_stage_2__2862_, data_stage_2__2861_, data_stage_2__2860_, data_stage_2__2859_, data_stage_2__2858_, data_stage_2__2857_, data_stage_2__2856_, data_stage_2__2855_, data_stage_2__2854_, data_stage_2__2853_, data_stage_2__2852_, data_stage_2__2851_, data_stage_2__2850_, data_stage_2__2849_, data_stage_2__2848_, data_stage_2__2847_, data_stage_2__2846_, data_stage_2__2845_, data_stage_2__2844_, data_stage_2__2843_, data_stage_2__2842_, data_stage_2__2841_, data_stage_2__2840_, data_stage_2__2839_, data_stage_2__2838_, data_stage_2__2837_, data_stage_2__2836_, data_stage_2__2835_, data_stage_2__2834_, data_stage_2__2833_, data_stage_2__2832_, data_stage_2__2831_, data_stage_2__2830_, data_stage_2__2829_, data_stage_2__2828_, data_stage_2__2827_, data_stage_2__2826_, data_stage_2__2825_, data_stage_2__2824_, data_stage_2__2823_, data_stage_2__2822_, data_stage_2__2821_, data_stage_2__2820_, data_stage_2__2819_, data_stage_2__2818_, data_stage_2__2817_, data_stage_2__2816_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_12__swap_inst
  (
    .data_i({ data_stage_1__3327_, data_stage_1__3326_, data_stage_1__3325_, data_stage_1__3324_, data_stage_1__3323_, data_stage_1__3322_, data_stage_1__3321_, data_stage_1__3320_, data_stage_1__3319_, data_stage_1__3318_, data_stage_1__3317_, data_stage_1__3316_, data_stage_1__3315_, data_stage_1__3314_, data_stage_1__3313_, data_stage_1__3312_, data_stage_1__3311_, data_stage_1__3310_, data_stage_1__3309_, data_stage_1__3308_, data_stage_1__3307_, data_stage_1__3306_, data_stage_1__3305_, data_stage_1__3304_, data_stage_1__3303_, data_stage_1__3302_, data_stage_1__3301_, data_stage_1__3300_, data_stage_1__3299_, data_stage_1__3298_, data_stage_1__3297_, data_stage_1__3296_, data_stage_1__3295_, data_stage_1__3294_, data_stage_1__3293_, data_stage_1__3292_, data_stage_1__3291_, data_stage_1__3290_, data_stage_1__3289_, data_stage_1__3288_, data_stage_1__3287_, data_stage_1__3286_, data_stage_1__3285_, data_stage_1__3284_, data_stage_1__3283_, data_stage_1__3282_, data_stage_1__3281_, data_stage_1__3280_, data_stage_1__3279_, data_stage_1__3278_, data_stage_1__3277_, data_stage_1__3276_, data_stage_1__3275_, data_stage_1__3274_, data_stage_1__3273_, data_stage_1__3272_, data_stage_1__3271_, data_stage_1__3270_, data_stage_1__3269_, data_stage_1__3268_, data_stage_1__3267_, data_stage_1__3266_, data_stage_1__3265_, data_stage_1__3264_, data_stage_1__3263_, data_stage_1__3262_, data_stage_1__3261_, data_stage_1__3260_, data_stage_1__3259_, data_stage_1__3258_, data_stage_1__3257_, data_stage_1__3256_, data_stage_1__3255_, data_stage_1__3254_, data_stage_1__3253_, data_stage_1__3252_, data_stage_1__3251_, data_stage_1__3250_, data_stage_1__3249_, data_stage_1__3248_, data_stage_1__3247_, data_stage_1__3246_, data_stage_1__3245_, data_stage_1__3244_, data_stage_1__3243_, data_stage_1__3242_, data_stage_1__3241_, data_stage_1__3240_, data_stage_1__3239_, data_stage_1__3238_, data_stage_1__3237_, data_stage_1__3236_, data_stage_1__3235_, data_stage_1__3234_, data_stage_1__3233_, data_stage_1__3232_, data_stage_1__3231_, data_stage_1__3230_, data_stage_1__3229_, data_stage_1__3228_, data_stage_1__3227_, data_stage_1__3226_, data_stage_1__3225_, data_stage_1__3224_, data_stage_1__3223_, data_stage_1__3222_, data_stage_1__3221_, data_stage_1__3220_, data_stage_1__3219_, data_stage_1__3218_, data_stage_1__3217_, data_stage_1__3216_, data_stage_1__3215_, data_stage_1__3214_, data_stage_1__3213_, data_stage_1__3212_, data_stage_1__3211_, data_stage_1__3210_, data_stage_1__3209_, data_stage_1__3208_, data_stage_1__3207_, data_stage_1__3206_, data_stage_1__3205_, data_stage_1__3204_, data_stage_1__3203_, data_stage_1__3202_, data_stage_1__3201_, data_stage_1__3200_, data_stage_1__3199_, data_stage_1__3198_, data_stage_1__3197_, data_stage_1__3196_, data_stage_1__3195_, data_stage_1__3194_, data_stage_1__3193_, data_stage_1__3192_, data_stage_1__3191_, data_stage_1__3190_, data_stage_1__3189_, data_stage_1__3188_, data_stage_1__3187_, data_stage_1__3186_, data_stage_1__3185_, data_stage_1__3184_, data_stage_1__3183_, data_stage_1__3182_, data_stage_1__3181_, data_stage_1__3180_, data_stage_1__3179_, data_stage_1__3178_, data_stage_1__3177_, data_stage_1__3176_, data_stage_1__3175_, data_stage_1__3174_, data_stage_1__3173_, data_stage_1__3172_, data_stage_1__3171_, data_stage_1__3170_, data_stage_1__3169_, data_stage_1__3168_, data_stage_1__3167_, data_stage_1__3166_, data_stage_1__3165_, data_stage_1__3164_, data_stage_1__3163_, data_stage_1__3162_, data_stage_1__3161_, data_stage_1__3160_, data_stage_1__3159_, data_stage_1__3158_, data_stage_1__3157_, data_stage_1__3156_, data_stage_1__3155_, data_stage_1__3154_, data_stage_1__3153_, data_stage_1__3152_, data_stage_1__3151_, data_stage_1__3150_, data_stage_1__3149_, data_stage_1__3148_, data_stage_1__3147_, data_stage_1__3146_, data_stage_1__3145_, data_stage_1__3144_, data_stage_1__3143_, data_stage_1__3142_, data_stage_1__3141_, data_stage_1__3140_, data_stage_1__3139_, data_stage_1__3138_, data_stage_1__3137_, data_stage_1__3136_, data_stage_1__3135_, data_stage_1__3134_, data_stage_1__3133_, data_stage_1__3132_, data_stage_1__3131_, data_stage_1__3130_, data_stage_1__3129_, data_stage_1__3128_, data_stage_1__3127_, data_stage_1__3126_, data_stage_1__3125_, data_stage_1__3124_, data_stage_1__3123_, data_stage_1__3122_, data_stage_1__3121_, data_stage_1__3120_, data_stage_1__3119_, data_stage_1__3118_, data_stage_1__3117_, data_stage_1__3116_, data_stage_1__3115_, data_stage_1__3114_, data_stage_1__3113_, data_stage_1__3112_, data_stage_1__3111_, data_stage_1__3110_, data_stage_1__3109_, data_stage_1__3108_, data_stage_1__3107_, data_stage_1__3106_, data_stage_1__3105_, data_stage_1__3104_, data_stage_1__3103_, data_stage_1__3102_, data_stage_1__3101_, data_stage_1__3100_, data_stage_1__3099_, data_stage_1__3098_, data_stage_1__3097_, data_stage_1__3096_, data_stage_1__3095_, data_stage_1__3094_, data_stage_1__3093_, data_stage_1__3092_, data_stage_1__3091_, data_stage_1__3090_, data_stage_1__3089_, data_stage_1__3088_, data_stage_1__3087_, data_stage_1__3086_, data_stage_1__3085_, data_stage_1__3084_, data_stage_1__3083_, data_stage_1__3082_, data_stage_1__3081_, data_stage_1__3080_, data_stage_1__3079_, data_stage_1__3078_, data_stage_1__3077_, data_stage_1__3076_, data_stage_1__3075_, data_stage_1__3074_, data_stage_1__3073_, data_stage_1__3072_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__3327_, data_stage_2__3326_, data_stage_2__3325_, data_stage_2__3324_, data_stage_2__3323_, data_stage_2__3322_, data_stage_2__3321_, data_stage_2__3320_, data_stage_2__3319_, data_stage_2__3318_, data_stage_2__3317_, data_stage_2__3316_, data_stage_2__3315_, data_stage_2__3314_, data_stage_2__3313_, data_stage_2__3312_, data_stage_2__3311_, data_stage_2__3310_, data_stage_2__3309_, data_stage_2__3308_, data_stage_2__3307_, data_stage_2__3306_, data_stage_2__3305_, data_stage_2__3304_, data_stage_2__3303_, data_stage_2__3302_, data_stage_2__3301_, data_stage_2__3300_, data_stage_2__3299_, data_stage_2__3298_, data_stage_2__3297_, data_stage_2__3296_, data_stage_2__3295_, data_stage_2__3294_, data_stage_2__3293_, data_stage_2__3292_, data_stage_2__3291_, data_stage_2__3290_, data_stage_2__3289_, data_stage_2__3288_, data_stage_2__3287_, data_stage_2__3286_, data_stage_2__3285_, data_stage_2__3284_, data_stage_2__3283_, data_stage_2__3282_, data_stage_2__3281_, data_stage_2__3280_, data_stage_2__3279_, data_stage_2__3278_, data_stage_2__3277_, data_stage_2__3276_, data_stage_2__3275_, data_stage_2__3274_, data_stage_2__3273_, data_stage_2__3272_, data_stage_2__3271_, data_stage_2__3270_, data_stage_2__3269_, data_stage_2__3268_, data_stage_2__3267_, data_stage_2__3266_, data_stage_2__3265_, data_stage_2__3264_, data_stage_2__3263_, data_stage_2__3262_, data_stage_2__3261_, data_stage_2__3260_, data_stage_2__3259_, data_stage_2__3258_, data_stage_2__3257_, data_stage_2__3256_, data_stage_2__3255_, data_stage_2__3254_, data_stage_2__3253_, data_stage_2__3252_, data_stage_2__3251_, data_stage_2__3250_, data_stage_2__3249_, data_stage_2__3248_, data_stage_2__3247_, data_stage_2__3246_, data_stage_2__3245_, data_stage_2__3244_, data_stage_2__3243_, data_stage_2__3242_, data_stage_2__3241_, data_stage_2__3240_, data_stage_2__3239_, data_stage_2__3238_, data_stage_2__3237_, data_stage_2__3236_, data_stage_2__3235_, data_stage_2__3234_, data_stage_2__3233_, data_stage_2__3232_, data_stage_2__3231_, data_stage_2__3230_, data_stage_2__3229_, data_stage_2__3228_, data_stage_2__3227_, data_stage_2__3226_, data_stage_2__3225_, data_stage_2__3224_, data_stage_2__3223_, data_stage_2__3222_, data_stage_2__3221_, data_stage_2__3220_, data_stage_2__3219_, data_stage_2__3218_, data_stage_2__3217_, data_stage_2__3216_, data_stage_2__3215_, data_stage_2__3214_, data_stage_2__3213_, data_stage_2__3212_, data_stage_2__3211_, data_stage_2__3210_, data_stage_2__3209_, data_stage_2__3208_, data_stage_2__3207_, data_stage_2__3206_, data_stage_2__3205_, data_stage_2__3204_, data_stage_2__3203_, data_stage_2__3202_, data_stage_2__3201_, data_stage_2__3200_, data_stage_2__3199_, data_stage_2__3198_, data_stage_2__3197_, data_stage_2__3196_, data_stage_2__3195_, data_stage_2__3194_, data_stage_2__3193_, data_stage_2__3192_, data_stage_2__3191_, data_stage_2__3190_, data_stage_2__3189_, data_stage_2__3188_, data_stage_2__3187_, data_stage_2__3186_, data_stage_2__3185_, data_stage_2__3184_, data_stage_2__3183_, data_stage_2__3182_, data_stage_2__3181_, data_stage_2__3180_, data_stage_2__3179_, data_stage_2__3178_, data_stage_2__3177_, data_stage_2__3176_, data_stage_2__3175_, data_stage_2__3174_, data_stage_2__3173_, data_stage_2__3172_, data_stage_2__3171_, data_stage_2__3170_, data_stage_2__3169_, data_stage_2__3168_, data_stage_2__3167_, data_stage_2__3166_, data_stage_2__3165_, data_stage_2__3164_, data_stage_2__3163_, data_stage_2__3162_, data_stage_2__3161_, data_stage_2__3160_, data_stage_2__3159_, data_stage_2__3158_, data_stage_2__3157_, data_stage_2__3156_, data_stage_2__3155_, data_stage_2__3154_, data_stage_2__3153_, data_stage_2__3152_, data_stage_2__3151_, data_stage_2__3150_, data_stage_2__3149_, data_stage_2__3148_, data_stage_2__3147_, data_stage_2__3146_, data_stage_2__3145_, data_stage_2__3144_, data_stage_2__3143_, data_stage_2__3142_, data_stage_2__3141_, data_stage_2__3140_, data_stage_2__3139_, data_stage_2__3138_, data_stage_2__3137_, data_stage_2__3136_, data_stage_2__3135_, data_stage_2__3134_, data_stage_2__3133_, data_stage_2__3132_, data_stage_2__3131_, data_stage_2__3130_, data_stage_2__3129_, data_stage_2__3128_, data_stage_2__3127_, data_stage_2__3126_, data_stage_2__3125_, data_stage_2__3124_, data_stage_2__3123_, data_stage_2__3122_, data_stage_2__3121_, data_stage_2__3120_, data_stage_2__3119_, data_stage_2__3118_, data_stage_2__3117_, data_stage_2__3116_, data_stage_2__3115_, data_stage_2__3114_, data_stage_2__3113_, data_stage_2__3112_, data_stage_2__3111_, data_stage_2__3110_, data_stage_2__3109_, data_stage_2__3108_, data_stage_2__3107_, data_stage_2__3106_, data_stage_2__3105_, data_stage_2__3104_, data_stage_2__3103_, data_stage_2__3102_, data_stage_2__3101_, data_stage_2__3100_, data_stage_2__3099_, data_stage_2__3098_, data_stage_2__3097_, data_stage_2__3096_, data_stage_2__3095_, data_stage_2__3094_, data_stage_2__3093_, data_stage_2__3092_, data_stage_2__3091_, data_stage_2__3090_, data_stage_2__3089_, data_stage_2__3088_, data_stage_2__3087_, data_stage_2__3086_, data_stage_2__3085_, data_stage_2__3084_, data_stage_2__3083_, data_stage_2__3082_, data_stage_2__3081_, data_stage_2__3080_, data_stage_2__3079_, data_stage_2__3078_, data_stage_2__3077_, data_stage_2__3076_, data_stage_2__3075_, data_stage_2__3074_, data_stage_2__3073_, data_stage_2__3072_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_13__swap_inst
  (
    .data_i({ data_stage_1__3583_, data_stage_1__3582_, data_stage_1__3581_, data_stage_1__3580_, data_stage_1__3579_, data_stage_1__3578_, data_stage_1__3577_, data_stage_1__3576_, data_stage_1__3575_, data_stage_1__3574_, data_stage_1__3573_, data_stage_1__3572_, data_stage_1__3571_, data_stage_1__3570_, data_stage_1__3569_, data_stage_1__3568_, data_stage_1__3567_, data_stage_1__3566_, data_stage_1__3565_, data_stage_1__3564_, data_stage_1__3563_, data_stage_1__3562_, data_stage_1__3561_, data_stage_1__3560_, data_stage_1__3559_, data_stage_1__3558_, data_stage_1__3557_, data_stage_1__3556_, data_stage_1__3555_, data_stage_1__3554_, data_stage_1__3553_, data_stage_1__3552_, data_stage_1__3551_, data_stage_1__3550_, data_stage_1__3549_, data_stage_1__3548_, data_stage_1__3547_, data_stage_1__3546_, data_stage_1__3545_, data_stage_1__3544_, data_stage_1__3543_, data_stage_1__3542_, data_stage_1__3541_, data_stage_1__3540_, data_stage_1__3539_, data_stage_1__3538_, data_stage_1__3537_, data_stage_1__3536_, data_stage_1__3535_, data_stage_1__3534_, data_stage_1__3533_, data_stage_1__3532_, data_stage_1__3531_, data_stage_1__3530_, data_stage_1__3529_, data_stage_1__3528_, data_stage_1__3527_, data_stage_1__3526_, data_stage_1__3525_, data_stage_1__3524_, data_stage_1__3523_, data_stage_1__3522_, data_stage_1__3521_, data_stage_1__3520_, data_stage_1__3519_, data_stage_1__3518_, data_stage_1__3517_, data_stage_1__3516_, data_stage_1__3515_, data_stage_1__3514_, data_stage_1__3513_, data_stage_1__3512_, data_stage_1__3511_, data_stage_1__3510_, data_stage_1__3509_, data_stage_1__3508_, data_stage_1__3507_, data_stage_1__3506_, data_stage_1__3505_, data_stage_1__3504_, data_stage_1__3503_, data_stage_1__3502_, data_stage_1__3501_, data_stage_1__3500_, data_stage_1__3499_, data_stage_1__3498_, data_stage_1__3497_, data_stage_1__3496_, data_stage_1__3495_, data_stage_1__3494_, data_stage_1__3493_, data_stage_1__3492_, data_stage_1__3491_, data_stage_1__3490_, data_stage_1__3489_, data_stage_1__3488_, data_stage_1__3487_, data_stage_1__3486_, data_stage_1__3485_, data_stage_1__3484_, data_stage_1__3483_, data_stage_1__3482_, data_stage_1__3481_, data_stage_1__3480_, data_stage_1__3479_, data_stage_1__3478_, data_stage_1__3477_, data_stage_1__3476_, data_stage_1__3475_, data_stage_1__3474_, data_stage_1__3473_, data_stage_1__3472_, data_stage_1__3471_, data_stage_1__3470_, data_stage_1__3469_, data_stage_1__3468_, data_stage_1__3467_, data_stage_1__3466_, data_stage_1__3465_, data_stage_1__3464_, data_stage_1__3463_, data_stage_1__3462_, data_stage_1__3461_, data_stage_1__3460_, data_stage_1__3459_, data_stage_1__3458_, data_stage_1__3457_, data_stage_1__3456_, data_stage_1__3455_, data_stage_1__3454_, data_stage_1__3453_, data_stage_1__3452_, data_stage_1__3451_, data_stage_1__3450_, data_stage_1__3449_, data_stage_1__3448_, data_stage_1__3447_, data_stage_1__3446_, data_stage_1__3445_, data_stage_1__3444_, data_stage_1__3443_, data_stage_1__3442_, data_stage_1__3441_, data_stage_1__3440_, data_stage_1__3439_, data_stage_1__3438_, data_stage_1__3437_, data_stage_1__3436_, data_stage_1__3435_, data_stage_1__3434_, data_stage_1__3433_, data_stage_1__3432_, data_stage_1__3431_, data_stage_1__3430_, data_stage_1__3429_, data_stage_1__3428_, data_stage_1__3427_, data_stage_1__3426_, data_stage_1__3425_, data_stage_1__3424_, data_stage_1__3423_, data_stage_1__3422_, data_stage_1__3421_, data_stage_1__3420_, data_stage_1__3419_, data_stage_1__3418_, data_stage_1__3417_, data_stage_1__3416_, data_stage_1__3415_, data_stage_1__3414_, data_stage_1__3413_, data_stage_1__3412_, data_stage_1__3411_, data_stage_1__3410_, data_stage_1__3409_, data_stage_1__3408_, data_stage_1__3407_, data_stage_1__3406_, data_stage_1__3405_, data_stage_1__3404_, data_stage_1__3403_, data_stage_1__3402_, data_stage_1__3401_, data_stage_1__3400_, data_stage_1__3399_, data_stage_1__3398_, data_stage_1__3397_, data_stage_1__3396_, data_stage_1__3395_, data_stage_1__3394_, data_stage_1__3393_, data_stage_1__3392_, data_stage_1__3391_, data_stage_1__3390_, data_stage_1__3389_, data_stage_1__3388_, data_stage_1__3387_, data_stage_1__3386_, data_stage_1__3385_, data_stage_1__3384_, data_stage_1__3383_, data_stage_1__3382_, data_stage_1__3381_, data_stage_1__3380_, data_stage_1__3379_, data_stage_1__3378_, data_stage_1__3377_, data_stage_1__3376_, data_stage_1__3375_, data_stage_1__3374_, data_stage_1__3373_, data_stage_1__3372_, data_stage_1__3371_, data_stage_1__3370_, data_stage_1__3369_, data_stage_1__3368_, data_stage_1__3367_, data_stage_1__3366_, data_stage_1__3365_, data_stage_1__3364_, data_stage_1__3363_, data_stage_1__3362_, data_stage_1__3361_, data_stage_1__3360_, data_stage_1__3359_, data_stage_1__3358_, data_stage_1__3357_, data_stage_1__3356_, data_stage_1__3355_, data_stage_1__3354_, data_stage_1__3353_, data_stage_1__3352_, data_stage_1__3351_, data_stage_1__3350_, data_stage_1__3349_, data_stage_1__3348_, data_stage_1__3347_, data_stage_1__3346_, data_stage_1__3345_, data_stage_1__3344_, data_stage_1__3343_, data_stage_1__3342_, data_stage_1__3341_, data_stage_1__3340_, data_stage_1__3339_, data_stage_1__3338_, data_stage_1__3337_, data_stage_1__3336_, data_stage_1__3335_, data_stage_1__3334_, data_stage_1__3333_, data_stage_1__3332_, data_stage_1__3331_, data_stage_1__3330_, data_stage_1__3329_, data_stage_1__3328_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__3583_, data_stage_2__3582_, data_stage_2__3581_, data_stage_2__3580_, data_stage_2__3579_, data_stage_2__3578_, data_stage_2__3577_, data_stage_2__3576_, data_stage_2__3575_, data_stage_2__3574_, data_stage_2__3573_, data_stage_2__3572_, data_stage_2__3571_, data_stage_2__3570_, data_stage_2__3569_, data_stage_2__3568_, data_stage_2__3567_, data_stage_2__3566_, data_stage_2__3565_, data_stage_2__3564_, data_stage_2__3563_, data_stage_2__3562_, data_stage_2__3561_, data_stage_2__3560_, data_stage_2__3559_, data_stage_2__3558_, data_stage_2__3557_, data_stage_2__3556_, data_stage_2__3555_, data_stage_2__3554_, data_stage_2__3553_, data_stage_2__3552_, data_stage_2__3551_, data_stage_2__3550_, data_stage_2__3549_, data_stage_2__3548_, data_stage_2__3547_, data_stage_2__3546_, data_stage_2__3545_, data_stage_2__3544_, data_stage_2__3543_, data_stage_2__3542_, data_stage_2__3541_, data_stage_2__3540_, data_stage_2__3539_, data_stage_2__3538_, data_stage_2__3537_, data_stage_2__3536_, data_stage_2__3535_, data_stage_2__3534_, data_stage_2__3533_, data_stage_2__3532_, data_stage_2__3531_, data_stage_2__3530_, data_stage_2__3529_, data_stage_2__3528_, data_stage_2__3527_, data_stage_2__3526_, data_stage_2__3525_, data_stage_2__3524_, data_stage_2__3523_, data_stage_2__3522_, data_stage_2__3521_, data_stage_2__3520_, data_stage_2__3519_, data_stage_2__3518_, data_stage_2__3517_, data_stage_2__3516_, data_stage_2__3515_, data_stage_2__3514_, data_stage_2__3513_, data_stage_2__3512_, data_stage_2__3511_, data_stage_2__3510_, data_stage_2__3509_, data_stage_2__3508_, data_stage_2__3507_, data_stage_2__3506_, data_stage_2__3505_, data_stage_2__3504_, data_stage_2__3503_, data_stage_2__3502_, data_stage_2__3501_, data_stage_2__3500_, data_stage_2__3499_, data_stage_2__3498_, data_stage_2__3497_, data_stage_2__3496_, data_stage_2__3495_, data_stage_2__3494_, data_stage_2__3493_, data_stage_2__3492_, data_stage_2__3491_, data_stage_2__3490_, data_stage_2__3489_, data_stage_2__3488_, data_stage_2__3487_, data_stage_2__3486_, data_stage_2__3485_, data_stage_2__3484_, data_stage_2__3483_, data_stage_2__3482_, data_stage_2__3481_, data_stage_2__3480_, data_stage_2__3479_, data_stage_2__3478_, data_stage_2__3477_, data_stage_2__3476_, data_stage_2__3475_, data_stage_2__3474_, data_stage_2__3473_, data_stage_2__3472_, data_stage_2__3471_, data_stage_2__3470_, data_stage_2__3469_, data_stage_2__3468_, data_stage_2__3467_, data_stage_2__3466_, data_stage_2__3465_, data_stage_2__3464_, data_stage_2__3463_, data_stage_2__3462_, data_stage_2__3461_, data_stage_2__3460_, data_stage_2__3459_, data_stage_2__3458_, data_stage_2__3457_, data_stage_2__3456_, data_stage_2__3455_, data_stage_2__3454_, data_stage_2__3453_, data_stage_2__3452_, data_stage_2__3451_, data_stage_2__3450_, data_stage_2__3449_, data_stage_2__3448_, data_stage_2__3447_, data_stage_2__3446_, data_stage_2__3445_, data_stage_2__3444_, data_stage_2__3443_, data_stage_2__3442_, data_stage_2__3441_, data_stage_2__3440_, data_stage_2__3439_, data_stage_2__3438_, data_stage_2__3437_, data_stage_2__3436_, data_stage_2__3435_, data_stage_2__3434_, data_stage_2__3433_, data_stage_2__3432_, data_stage_2__3431_, data_stage_2__3430_, data_stage_2__3429_, data_stage_2__3428_, data_stage_2__3427_, data_stage_2__3426_, data_stage_2__3425_, data_stage_2__3424_, data_stage_2__3423_, data_stage_2__3422_, data_stage_2__3421_, data_stage_2__3420_, data_stage_2__3419_, data_stage_2__3418_, data_stage_2__3417_, data_stage_2__3416_, data_stage_2__3415_, data_stage_2__3414_, data_stage_2__3413_, data_stage_2__3412_, data_stage_2__3411_, data_stage_2__3410_, data_stage_2__3409_, data_stage_2__3408_, data_stage_2__3407_, data_stage_2__3406_, data_stage_2__3405_, data_stage_2__3404_, data_stage_2__3403_, data_stage_2__3402_, data_stage_2__3401_, data_stage_2__3400_, data_stage_2__3399_, data_stage_2__3398_, data_stage_2__3397_, data_stage_2__3396_, data_stage_2__3395_, data_stage_2__3394_, data_stage_2__3393_, data_stage_2__3392_, data_stage_2__3391_, data_stage_2__3390_, data_stage_2__3389_, data_stage_2__3388_, data_stage_2__3387_, data_stage_2__3386_, data_stage_2__3385_, data_stage_2__3384_, data_stage_2__3383_, data_stage_2__3382_, data_stage_2__3381_, data_stage_2__3380_, data_stage_2__3379_, data_stage_2__3378_, data_stage_2__3377_, data_stage_2__3376_, data_stage_2__3375_, data_stage_2__3374_, data_stage_2__3373_, data_stage_2__3372_, data_stage_2__3371_, data_stage_2__3370_, data_stage_2__3369_, data_stage_2__3368_, data_stage_2__3367_, data_stage_2__3366_, data_stage_2__3365_, data_stage_2__3364_, data_stage_2__3363_, data_stage_2__3362_, data_stage_2__3361_, data_stage_2__3360_, data_stage_2__3359_, data_stage_2__3358_, data_stage_2__3357_, data_stage_2__3356_, data_stage_2__3355_, data_stage_2__3354_, data_stage_2__3353_, data_stage_2__3352_, data_stage_2__3351_, data_stage_2__3350_, data_stage_2__3349_, data_stage_2__3348_, data_stage_2__3347_, data_stage_2__3346_, data_stage_2__3345_, data_stage_2__3344_, data_stage_2__3343_, data_stage_2__3342_, data_stage_2__3341_, data_stage_2__3340_, data_stage_2__3339_, data_stage_2__3338_, data_stage_2__3337_, data_stage_2__3336_, data_stage_2__3335_, data_stage_2__3334_, data_stage_2__3333_, data_stage_2__3332_, data_stage_2__3331_, data_stage_2__3330_, data_stage_2__3329_, data_stage_2__3328_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_14__swap_inst
  (
    .data_i({ data_stage_1__3839_, data_stage_1__3838_, data_stage_1__3837_, data_stage_1__3836_, data_stage_1__3835_, data_stage_1__3834_, data_stage_1__3833_, data_stage_1__3832_, data_stage_1__3831_, data_stage_1__3830_, data_stage_1__3829_, data_stage_1__3828_, data_stage_1__3827_, data_stage_1__3826_, data_stage_1__3825_, data_stage_1__3824_, data_stage_1__3823_, data_stage_1__3822_, data_stage_1__3821_, data_stage_1__3820_, data_stage_1__3819_, data_stage_1__3818_, data_stage_1__3817_, data_stage_1__3816_, data_stage_1__3815_, data_stage_1__3814_, data_stage_1__3813_, data_stage_1__3812_, data_stage_1__3811_, data_stage_1__3810_, data_stage_1__3809_, data_stage_1__3808_, data_stage_1__3807_, data_stage_1__3806_, data_stage_1__3805_, data_stage_1__3804_, data_stage_1__3803_, data_stage_1__3802_, data_stage_1__3801_, data_stage_1__3800_, data_stage_1__3799_, data_stage_1__3798_, data_stage_1__3797_, data_stage_1__3796_, data_stage_1__3795_, data_stage_1__3794_, data_stage_1__3793_, data_stage_1__3792_, data_stage_1__3791_, data_stage_1__3790_, data_stage_1__3789_, data_stage_1__3788_, data_stage_1__3787_, data_stage_1__3786_, data_stage_1__3785_, data_stage_1__3784_, data_stage_1__3783_, data_stage_1__3782_, data_stage_1__3781_, data_stage_1__3780_, data_stage_1__3779_, data_stage_1__3778_, data_stage_1__3777_, data_stage_1__3776_, data_stage_1__3775_, data_stage_1__3774_, data_stage_1__3773_, data_stage_1__3772_, data_stage_1__3771_, data_stage_1__3770_, data_stage_1__3769_, data_stage_1__3768_, data_stage_1__3767_, data_stage_1__3766_, data_stage_1__3765_, data_stage_1__3764_, data_stage_1__3763_, data_stage_1__3762_, data_stage_1__3761_, data_stage_1__3760_, data_stage_1__3759_, data_stage_1__3758_, data_stage_1__3757_, data_stage_1__3756_, data_stage_1__3755_, data_stage_1__3754_, data_stage_1__3753_, data_stage_1__3752_, data_stage_1__3751_, data_stage_1__3750_, data_stage_1__3749_, data_stage_1__3748_, data_stage_1__3747_, data_stage_1__3746_, data_stage_1__3745_, data_stage_1__3744_, data_stage_1__3743_, data_stage_1__3742_, data_stage_1__3741_, data_stage_1__3740_, data_stage_1__3739_, data_stage_1__3738_, data_stage_1__3737_, data_stage_1__3736_, data_stage_1__3735_, data_stage_1__3734_, data_stage_1__3733_, data_stage_1__3732_, data_stage_1__3731_, data_stage_1__3730_, data_stage_1__3729_, data_stage_1__3728_, data_stage_1__3727_, data_stage_1__3726_, data_stage_1__3725_, data_stage_1__3724_, data_stage_1__3723_, data_stage_1__3722_, data_stage_1__3721_, data_stage_1__3720_, data_stage_1__3719_, data_stage_1__3718_, data_stage_1__3717_, data_stage_1__3716_, data_stage_1__3715_, data_stage_1__3714_, data_stage_1__3713_, data_stage_1__3712_, data_stage_1__3711_, data_stage_1__3710_, data_stage_1__3709_, data_stage_1__3708_, data_stage_1__3707_, data_stage_1__3706_, data_stage_1__3705_, data_stage_1__3704_, data_stage_1__3703_, data_stage_1__3702_, data_stage_1__3701_, data_stage_1__3700_, data_stage_1__3699_, data_stage_1__3698_, data_stage_1__3697_, data_stage_1__3696_, data_stage_1__3695_, data_stage_1__3694_, data_stage_1__3693_, data_stage_1__3692_, data_stage_1__3691_, data_stage_1__3690_, data_stage_1__3689_, data_stage_1__3688_, data_stage_1__3687_, data_stage_1__3686_, data_stage_1__3685_, data_stage_1__3684_, data_stage_1__3683_, data_stage_1__3682_, data_stage_1__3681_, data_stage_1__3680_, data_stage_1__3679_, data_stage_1__3678_, data_stage_1__3677_, data_stage_1__3676_, data_stage_1__3675_, data_stage_1__3674_, data_stage_1__3673_, data_stage_1__3672_, data_stage_1__3671_, data_stage_1__3670_, data_stage_1__3669_, data_stage_1__3668_, data_stage_1__3667_, data_stage_1__3666_, data_stage_1__3665_, data_stage_1__3664_, data_stage_1__3663_, data_stage_1__3662_, data_stage_1__3661_, data_stage_1__3660_, data_stage_1__3659_, data_stage_1__3658_, data_stage_1__3657_, data_stage_1__3656_, data_stage_1__3655_, data_stage_1__3654_, data_stage_1__3653_, data_stage_1__3652_, data_stage_1__3651_, data_stage_1__3650_, data_stage_1__3649_, data_stage_1__3648_, data_stage_1__3647_, data_stage_1__3646_, data_stage_1__3645_, data_stage_1__3644_, data_stage_1__3643_, data_stage_1__3642_, data_stage_1__3641_, data_stage_1__3640_, data_stage_1__3639_, data_stage_1__3638_, data_stage_1__3637_, data_stage_1__3636_, data_stage_1__3635_, data_stage_1__3634_, data_stage_1__3633_, data_stage_1__3632_, data_stage_1__3631_, data_stage_1__3630_, data_stage_1__3629_, data_stage_1__3628_, data_stage_1__3627_, data_stage_1__3626_, data_stage_1__3625_, data_stage_1__3624_, data_stage_1__3623_, data_stage_1__3622_, data_stage_1__3621_, data_stage_1__3620_, data_stage_1__3619_, data_stage_1__3618_, data_stage_1__3617_, data_stage_1__3616_, data_stage_1__3615_, data_stage_1__3614_, data_stage_1__3613_, data_stage_1__3612_, data_stage_1__3611_, data_stage_1__3610_, data_stage_1__3609_, data_stage_1__3608_, data_stage_1__3607_, data_stage_1__3606_, data_stage_1__3605_, data_stage_1__3604_, data_stage_1__3603_, data_stage_1__3602_, data_stage_1__3601_, data_stage_1__3600_, data_stage_1__3599_, data_stage_1__3598_, data_stage_1__3597_, data_stage_1__3596_, data_stage_1__3595_, data_stage_1__3594_, data_stage_1__3593_, data_stage_1__3592_, data_stage_1__3591_, data_stage_1__3590_, data_stage_1__3589_, data_stage_1__3588_, data_stage_1__3587_, data_stage_1__3586_, data_stage_1__3585_, data_stage_1__3584_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__3839_, data_stage_2__3838_, data_stage_2__3837_, data_stage_2__3836_, data_stage_2__3835_, data_stage_2__3834_, data_stage_2__3833_, data_stage_2__3832_, data_stage_2__3831_, data_stage_2__3830_, data_stage_2__3829_, data_stage_2__3828_, data_stage_2__3827_, data_stage_2__3826_, data_stage_2__3825_, data_stage_2__3824_, data_stage_2__3823_, data_stage_2__3822_, data_stage_2__3821_, data_stage_2__3820_, data_stage_2__3819_, data_stage_2__3818_, data_stage_2__3817_, data_stage_2__3816_, data_stage_2__3815_, data_stage_2__3814_, data_stage_2__3813_, data_stage_2__3812_, data_stage_2__3811_, data_stage_2__3810_, data_stage_2__3809_, data_stage_2__3808_, data_stage_2__3807_, data_stage_2__3806_, data_stage_2__3805_, data_stage_2__3804_, data_stage_2__3803_, data_stage_2__3802_, data_stage_2__3801_, data_stage_2__3800_, data_stage_2__3799_, data_stage_2__3798_, data_stage_2__3797_, data_stage_2__3796_, data_stage_2__3795_, data_stage_2__3794_, data_stage_2__3793_, data_stage_2__3792_, data_stage_2__3791_, data_stage_2__3790_, data_stage_2__3789_, data_stage_2__3788_, data_stage_2__3787_, data_stage_2__3786_, data_stage_2__3785_, data_stage_2__3784_, data_stage_2__3783_, data_stage_2__3782_, data_stage_2__3781_, data_stage_2__3780_, data_stage_2__3779_, data_stage_2__3778_, data_stage_2__3777_, data_stage_2__3776_, data_stage_2__3775_, data_stage_2__3774_, data_stage_2__3773_, data_stage_2__3772_, data_stage_2__3771_, data_stage_2__3770_, data_stage_2__3769_, data_stage_2__3768_, data_stage_2__3767_, data_stage_2__3766_, data_stage_2__3765_, data_stage_2__3764_, data_stage_2__3763_, data_stage_2__3762_, data_stage_2__3761_, data_stage_2__3760_, data_stage_2__3759_, data_stage_2__3758_, data_stage_2__3757_, data_stage_2__3756_, data_stage_2__3755_, data_stage_2__3754_, data_stage_2__3753_, data_stage_2__3752_, data_stage_2__3751_, data_stage_2__3750_, data_stage_2__3749_, data_stage_2__3748_, data_stage_2__3747_, data_stage_2__3746_, data_stage_2__3745_, data_stage_2__3744_, data_stage_2__3743_, data_stage_2__3742_, data_stage_2__3741_, data_stage_2__3740_, data_stage_2__3739_, data_stage_2__3738_, data_stage_2__3737_, data_stage_2__3736_, data_stage_2__3735_, data_stage_2__3734_, data_stage_2__3733_, data_stage_2__3732_, data_stage_2__3731_, data_stage_2__3730_, data_stage_2__3729_, data_stage_2__3728_, data_stage_2__3727_, data_stage_2__3726_, data_stage_2__3725_, data_stage_2__3724_, data_stage_2__3723_, data_stage_2__3722_, data_stage_2__3721_, data_stage_2__3720_, data_stage_2__3719_, data_stage_2__3718_, data_stage_2__3717_, data_stage_2__3716_, data_stage_2__3715_, data_stage_2__3714_, data_stage_2__3713_, data_stage_2__3712_, data_stage_2__3711_, data_stage_2__3710_, data_stage_2__3709_, data_stage_2__3708_, data_stage_2__3707_, data_stage_2__3706_, data_stage_2__3705_, data_stage_2__3704_, data_stage_2__3703_, data_stage_2__3702_, data_stage_2__3701_, data_stage_2__3700_, data_stage_2__3699_, data_stage_2__3698_, data_stage_2__3697_, data_stage_2__3696_, data_stage_2__3695_, data_stage_2__3694_, data_stage_2__3693_, data_stage_2__3692_, data_stage_2__3691_, data_stage_2__3690_, data_stage_2__3689_, data_stage_2__3688_, data_stage_2__3687_, data_stage_2__3686_, data_stage_2__3685_, data_stage_2__3684_, data_stage_2__3683_, data_stage_2__3682_, data_stage_2__3681_, data_stage_2__3680_, data_stage_2__3679_, data_stage_2__3678_, data_stage_2__3677_, data_stage_2__3676_, data_stage_2__3675_, data_stage_2__3674_, data_stage_2__3673_, data_stage_2__3672_, data_stage_2__3671_, data_stage_2__3670_, data_stage_2__3669_, data_stage_2__3668_, data_stage_2__3667_, data_stage_2__3666_, data_stage_2__3665_, data_stage_2__3664_, data_stage_2__3663_, data_stage_2__3662_, data_stage_2__3661_, data_stage_2__3660_, data_stage_2__3659_, data_stage_2__3658_, data_stage_2__3657_, data_stage_2__3656_, data_stage_2__3655_, data_stage_2__3654_, data_stage_2__3653_, data_stage_2__3652_, data_stage_2__3651_, data_stage_2__3650_, data_stage_2__3649_, data_stage_2__3648_, data_stage_2__3647_, data_stage_2__3646_, data_stage_2__3645_, data_stage_2__3644_, data_stage_2__3643_, data_stage_2__3642_, data_stage_2__3641_, data_stage_2__3640_, data_stage_2__3639_, data_stage_2__3638_, data_stage_2__3637_, data_stage_2__3636_, data_stage_2__3635_, data_stage_2__3634_, data_stage_2__3633_, data_stage_2__3632_, data_stage_2__3631_, data_stage_2__3630_, data_stage_2__3629_, data_stage_2__3628_, data_stage_2__3627_, data_stage_2__3626_, data_stage_2__3625_, data_stage_2__3624_, data_stage_2__3623_, data_stage_2__3622_, data_stage_2__3621_, data_stage_2__3620_, data_stage_2__3619_, data_stage_2__3618_, data_stage_2__3617_, data_stage_2__3616_, data_stage_2__3615_, data_stage_2__3614_, data_stage_2__3613_, data_stage_2__3612_, data_stage_2__3611_, data_stage_2__3610_, data_stage_2__3609_, data_stage_2__3608_, data_stage_2__3607_, data_stage_2__3606_, data_stage_2__3605_, data_stage_2__3604_, data_stage_2__3603_, data_stage_2__3602_, data_stage_2__3601_, data_stage_2__3600_, data_stage_2__3599_, data_stage_2__3598_, data_stage_2__3597_, data_stage_2__3596_, data_stage_2__3595_, data_stage_2__3594_, data_stage_2__3593_, data_stage_2__3592_, data_stage_2__3591_, data_stage_2__3590_, data_stage_2__3589_, data_stage_2__3588_, data_stage_2__3587_, data_stage_2__3586_, data_stage_2__3585_, data_stage_2__3584_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_15__swap_inst
  (
    .data_i({ data_stage_1__4095_, data_stage_1__4094_, data_stage_1__4093_, data_stage_1__4092_, data_stage_1__4091_, data_stage_1__4090_, data_stage_1__4089_, data_stage_1__4088_, data_stage_1__4087_, data_stage_1__4086_, data_stage_1__4085_, data_stage_1__4084_, data_stage_1__4083_, data_stage_1__4082_, data_stage_1__4081_, data_stage_1__4080_, data_stage_1__4079_, data_stage_1__4078_, data_stage_1__4077_, data_stage_1__4076_, data_stage_1__4075_, data_stage_1__4074_, data_stage_1__4073_, data_stage_1__4072_, data_stage_1__4071_, data_stage_1__4070_, data_stage_1__4069_, data_stage_1__4068_, data_stage_1__4067_, data_stage_1__4066_, data_stage_1__4065_, data_stage_1__4064_, data_stage_1__4063_, data_stage_1__4062_, data_stage_1__4061_, data_stage_1__4060_, data_stage_1__4059_, data_stage_1__4058_, data_stage_1__4057_, data_stage_1__4056_, data_stage_1__4055_, data_stage_1__4054_, data_stage_1__4053_, data_stage_1__4052_, data_stage_1__4051_, data_stage_1__4050_, data_stage_1__4049_, data_stage_1__4048_, data_stage_1__4047_, data_stage_1__4046_, data_stage_1__4045_, data_stage_1__4044_, data_stage_1__4043_, data_stage_1__4042_, data_stage_1__4041_, data_stage_1__4040_, data_stage_1__4039_, data_stage_1__4038_, data_stage_1__4037_, data_stage_1__4036_, data_stage_1__4035_, data_stage_1__4034_, data_stage_1__4033_, data_stage_1__4032_, data_stage_1__4031_, data_stage_1__4030_, data_stage_1__4029_, data_stage_1__4028_, data_stage_1__4027_, data_stage_1__4026_, data_stage_1__4025_, data_stage_1__4024_, data_stage_1__4023_, data_stage_1__4022_, data_stage_1__4021_, data_stage_1__4020_, data_stage_1__4019_, data_stage_1__4018_, data_stage_1__4017_, data_stage_1__4016_, data_stage_1__4015_, data_stage_1__4014_, data_stage_1__4013_, data_stage_1__4012_, data_stage_1__4011_, data_stage_1__4010_, data_stage_1__4009_, data_stage_1__4008_, data_stage_1__4007_, data_stage_1__4006_, data_stage_1__4005_, data_stage_1__4004_, data_stage_1__4003_, data_stage_1__4002_, data_stage_1__4001_, data_stage_1__4000_, data_stage_1__3999_, data_stage_1__3998_, data_stage_1__3997_, data_stage_1__3996_, data_stage_1__3995_, data_stage_1__3994_, data_stage_1__3993_, data_stage_1__3992_, data_stage_1__3991_, data_stage_1__3990_, data_stage_1__3989_, data_stage_1__3988_, data_stage_1__3987_, data_stage_1__3986_, data_stage_1__3985_, data_stage_1__3984_, data_stage_1__3983_, data_stage_1__3982_, data_stage_1__3981_, data_stage_1__3980_, data_stage_1__3979_, data_stage_1__3978_, data_stage_1__3977_, data_stage_1__3976_, data_stage_1__3975_, data_stage_1__3974_, data_stage_1__3973_, data_stage_1__3972_, data_stage_1__3971_, data_stage_1__3970_, data_stage_1__3969_, data_stage_1__3968_, data_stage_1__3967_, data_stage_1__3966_, data_stage_1__3965_, data_stage_1__3964_, data_stage_1__3963_, data_stage_1__3962_, data_stage_1__3961_, data_stage_1__3960_, data_stage_1__3959_, data_stage_1__3958_, data_stage_1__3957_, data_stage_1__3956_, data_stage_1__3955_, data_stage_1__3954_, data_stage_1__3953_, data_stage_1__3952_, data_stage_1__3951_, data_stage_1__3950_, data_stage_1__3949_, data_stage_1__3948_, data_stage_1__3947_, data_stage_1__3946_, data_stage_1__3945_, data_stage_1__3944_, data_stage_1__3943_, data_stage_1__3942_, data_stage_1__3941_, data_stage_1__3940_, data_stage_1__3939_, data_stage_1__3938_, data_stage_1__3937_, data_stage_1__3936_, data_stage_1__3935_, data_stage_1__3934_, data_stage_1__3933_, data_stage_1__3932_, data_stage_1__3931_, data_stage_1__3930_, data_stage_1__3929_, data_stage_1__3928_, data_stage_1__3927_, data_stage_1__3926_, data_stage_1__3925_, data_stage_1__3924_, data_stage_1__3923_, data_stage_1__3922_, data_stage_1__3921_, data_stage_1__3920_, data_stage_1__3919_, data_stage_1__3918_, data_stage_1__3917_, data_stage_1__3916_, data_stage_1__3915_, data_stage_1__3914_, data_stage_1__3913_, data_stage_1__3912_, data_stage_1__3911_, data_stage_1__3910_, data_stage_1__3909_, data_stage_1__3908_, data_stage_1__3907_, data_stage_1__3906_, data_stage_1__3905_, data_stage_1__3904_, data_stage_1__3903_, data_stage_1__3902_, data_stage_1__3901_, data_stage_1__3900_, data_stage_1__3899_, data_stage_1__3898_, data_stage_1__3897_, data_stage_1__3896_, data_stage_1__3895_, data_stage_1__3894_, data_stage_1__3893_, data_stage_1__3892_, data_stage_1__3891_, data_stage_1__3890_, data_stage_1__3889_, data_stage_1__3888_, data_stage_1__3887_, data_stage_1__3886_, data_stage_1__3885_, data_stage_1__3884_, data_stage_1__3883_, data_stage_1__3882_, data_stage_1__3881_, data_stage_1__3880_, data_stage_1__3879_, data_stage_1__3878_, data_stage_1__3877_, data_stage_1__3876_, data_stage_1__3875_, data_stage_1__3874_, data_stage_1__3873_, data_stage_1__3872_, data_stage_1__3871_, data_stage_1__3870_, data_stage_1__3869_, data_stage_1__3868_, data_stage_1__3867_, data_stage_1__3866_, data_stage_1__3865_, data_stage_1__3864_, data_stage_1__3863_, data_stage_1__3862_, data_stage_1__3861_, data_stage_1__3860_, data_stage_1__3859_, data_stage_1__3858_, data_stage_1__3857_, data_stage_1__3856_, data_stage_1__3855_, data_stage_1__3854_, data_stage_1__3853_, data_stage_1__3852_, data_stage_1__3851_, data_stage_1__3850_, data_stage_1__3849_, data_stage_1__3848_, data_stage_1__3847_, data_stage_1__3846_, data_stage_1__3845_, data_stage_1__3844_, data_stage_1__3843_, data_stage_1__3842_, data_stage_1__3841_, data_stage_1__3840_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__4095_, data_stage_2__4094_, data_stage_2__4093_, data_stage_2__4092_, data_stage_2__4091_, data_stage_2__4090_, data_stage_2__4089_, data_stage_2__4088_, data_stage_2__4087_, data_stage_2__4086_, data_stage_2__4085_, data_stage_2__4084_, data_stage_2__4083_, data_stage_2__4082_, data_stage_2__4081_, data_stage_2__4080_, data_stage_2__4079_, data_stage_2__4078_, data_stage_2__4077_, data_stage_2__4076_, data_stage_2__4075_, data_stage_2__4074_, data_stage_2__4073_, data_stage_2__4072_, data_stage_2__4071_, data_stage_2__4070_, data_stage_2__4069_, data_stage_2__4068_, data_stage_2__4067_, data_stage_2__4066_, data_stage_2__4065_, data_stage_2__4064_, data_stage_2__4063_, data_stage_2__4062_, data_stage_2__4061_, data_stage_2__4060_, data_stage_2__4059_, data_stage_2__4058_, data_stage_2__4057_, data_stage_2__4056_, data_stage_2__4055_, data_stage_2__4054_, data_stage_2__4053_, data_stage_2__4052_, data_stage_2__4051_, data_stage_2__4050_, data_stage_2__4049_, data_stage_2__4048_, data_stage_2__4047_, data_stage_2__4046_, data_stage_2__4045_, data_stage_2__4044_, data_stage_2__4043_, data_stage_2__4042_, data_stage_2__4041_, data_stage_2__4040_, data_stage_2__4039_, data_stage_2__4038_, data_stage_2__4037_, data_stage_2__4036_, data_stage_2__4035_, data_stage_2__4034_, data_stage_2__4033_, data_stage_2__4032_, data_stage_2__4031_, data_stage_2__4030_, data_stage_2__4029_, data_stage_2__4028_, data_stage_2__4027_, data_stage_2__4026_, data_stage_2__4025_, data_stage_2__4024_, data_stage_2__4023_, data_stage_2__4022_, data_stage_2__4021_, data_stage_2__4020_, data_stage_2__4019_, data_stage_2__4018_, data_stage_2__4017_, data_stage_2__4016_, data_stage_2__4015_, data_stage_2__4014_, data_stage_2__4013_, data_stage_2__4012_, data_stage_2__4011_, data_stage_2__4010_, data_stage_2__4009_, data_stage_2__4008_, data_stage_2__4007_, data_stage_2__4006_, data_stage_2__4005_, data_stage_2__4004_, data_stage_2__4003_, data_stage_2__4002_, data_stage_2__4001_, data_stage_2__4000_, data_stage_2__3999_, data_stage_2__3998_, data_stage_2__3997_, data_stage_2__3996_, data_stage_2__3995_, data_stage_2__3994_, data_stage_2__3993_, data_stage_2__3992_, data_stage_2__3991_, data_stage_2__3990_, data_stage_2__3989_, data_stage_2__3988_, data_stage_2__3987_, data_stage_2__3986_, data_stage_2__3985_, data_stage_2__3984_, data_stage_2__3983_, data_stage_2__3982_, data_stage_2__3981_, data_stage_2__3980_, data_stage_2__3979_, data_stage_2__3978_, data_stage_2__3977_, data_stage_2__3976_, data_stage_2__3975_, data_stage_2__3974_, data_stage_2__3973_, data_stage_2__3972_, data_stage_2__3971_, data_stage_2__3970_, data_stage_2__3969_, data_stage_2__3968_, data_stage_2__3967_, data_stage_2__3966_, data_stage_2__3965_, data_stage_2__3964_, data_stage_2__3963_, data_stage_2__3962_, data_stage_2__3961_, data_stage_2__3960_, data_stage_2__3959_, data_stage_2__3958_, data_stage_2__3957_, data_stage_2__3956_, data_stage_2__3955_, data_stage_2__3954_, data_stage_2__3953_, data_stage_2__3952_, data_stage_2__3951_, data_stage_2__3950_, data_stage_2__3949_, data_stage_2__3948_, data_stage_2__3947_, data_stage_2__3946_, data_stage_2__3945_, data_stage_2__3944_, data_stage_2__3943_, data_stage_2__3942_, data_stage_2__3941_, data_stage_2__3940_, data_stage_2__3939_, data_stage_2__3938_, data_stage_2__3937_, data_stage_2__3936_, data_stage_2__3935_, data_stage_2__3934_, data_stage_2__3933_, data_stage_2__3932_, data_stage_2__3931_, data_stage_2__3930_, data_stage_2__3929_, data_stage_2__3928_, data_stage_2__3927_, data_stage_2__3926_, data_stage_2__3925_, data_stage_2__3924_, data_stage_2__3923_, data_stage_2__3922_, data_stage_2__3921_, data_stage_2__3920_, data_stage_2__3919_, data_stage_2__3918_, data_stage_2__3917_, data_stage_2__3916_, data_stage_2__3915_, data_stage_2__3914_, data_stage_2__3913_, data_stage_2__3912_, data_stage_2__3911_, data_stage_2__3910_, data_stage_2__3909_, data_stage_2__3908_, data_stage_2__3907_, data_stage_2__3906_, data_stage_2__3905_, data_stage_2__3904_, data_stage_2__3903_, data_stage_2__3902_, data_stage_2__3901_, data_stage_2__3900_, data_stage_2__3899_, data_stage_2__3898_, data_stage_2__3897_, data_stage_2__3896_, data_stage_2__3895_, data_stage_2__3894_, data_stage_2__3893_, data_stage_2__3892_, data_stage_2__3891_, data_stage_2__3890_, data_stage_2__3889_, data_stage_2__3888_, data_stage_2__3887_, data_stage_2__3886_, data_stage_2__3885_, data_stage_2__3884_, data_stage_2__3883_, data_stage_2__3882_, data_stage_2__3881_, data_stage_2__3880_, data_stage_2__3879_, data_stage_2__3878_, data_stage_2__3877_, data_stage_2__3876_, data_stage_2__3875_, data_stage_2__3874_, data_stage_2__3873_, data_stage_2__3872_, data_stage_2__3871_, data_stage_2__3870_, data_stage_2__3869_, data_stage_2__3868_, data_stage_2__3867_, data_stage_2__3866_, data_stage_2__3865_, data_stage_2__3864_, data_stage_2__3863_, data_stage_2__3862_, data_stage_2__3861_, data_stage_2__3860_, data_stage_2__3859_, data_stage_2__3858_, data_stage_2__3857_, data_stage_2__3856_, data_stage_2__3855_, data_stage_2__3854_, data_stage_2__3853_, data_stage_2__3852_, data_stage_2__3851_, data_stage_2__3850_, data_stage_2__3849_, data_stage_2__3848_, data_stage_2__3847_, data_stage_2__3846_, data_stage_2__3845_, data_stage_2__3844_, data_stage_2__3843_, data_stage_2__3842_, data_stage_2__3841_, data_stage_2__3840_ })
  );


  bsg_swap_width_p256
  mux_stage_2__mux_swap_0__swap_inst
  (
    .data_i({ data_stage_2__511_, data_stage_2__510_, data_stage_2__509_, data_stage_2__508_, data_stage_2__507_, data_stage_2__506_, data_stage_2__505_, data_stage_2__504_, data_stage_2__503_, data_stage_2__502_, data_stage_2__501_, data_stage_2__500_, data_stage_2__499_, data_stage_2__498_, data_stage_2__497_, data_stage_2__496_, data_stage_2__495_, data_stage_2__494_, data_stage_2__493_, data_stage_2__492_, data_stage_2__491_, data_stage_2__490_, data_stage_2__489_, data_stage_2__488_, data_stage_2__487_, data_stage_2__486_, data_stage_2__485_, data_stage_2__484_, data_stage_2__483_, data_stage_2__482_, data_stage_2__481_, data_stage_2__480_, data_stage_2__479_, data_stage_2__478_, data_stage_2__477_, data_stage_2__476_, data_stage_2__475_, data_stage_2__474_, data_stage_2__473_, data_stage_2__472_, data_stage_2__471_, data_stage_2__470_, data_stage_2__469_, data_stage_2__468_, data_stage_2__467_, data_stage_2__466_, data_stage_2__465_, data_stage_2__464_, data_stage_2__463_, data_stage_2__462_, data_stage_2__461_, data_stage_2__460_, data_stage_2__459_, data_stage_2__458_, data_stage_2__457_, data_stage_2__456_, data_stage_2__455_, data_stage_2__454_, data_stage_2__453_, data_stage_2__452_, data_stage_2__451_, data_stage_2__450_, data_stage_2__449_, data_stage_2__448_, data_stage_2__447_, data_stage_2__446_, data_stage_2__445_, data_stage_2__444_, data_stage_2__443_, data_stage_2__442_, data_stage_2__441_, data_stage_2__440_, data_stage_2__439_, data_stage_2__438_, data_stage_2__437_, data_stage_2__436_, data_stage_2__435_, data_stage_2__434_, data_stage_2__433_, data_stage_2__432_, data_stage_2__431_, data_stage_2__430_, data_stage_2__429_, data_stage_2__428_, data_stage_2__427_, data_stage_2__426_, data_stage_2__425_, data_stage_2__424_, data_stage_2__423_, data_stage_2__422_, data_stage_2__421_, data_stage_2__420_, data_stage_2__419_, data_stage_2__418_, data_stage_2__417_, data_stage_2__416_, data_stage_2__415_, data_stage_2__414_, data_stage_2__413_, data_stage_2__412_, data_stage_2__411_, data_stage_2__410_, data_stage_2__409_, data_stage_2__408_, data_stage_2__407_, data_stage_2__406_, data_stage_2__405_, data_stage_2__404_, data_stage_2__403_, data_stage_2__402_, data_stage_2__401_, data_stage_2__400_, data_stage_2__399_, data_stage_2__398_, data_stage_2__397_, data_stage_2__396_, data_stage_2__395_, data_stage_2__394_, data_stage_2__393_, data_stage_2__392_, data_stage_2__391_, data_stage_2__390_, data_stage_2__389_, data_stage_2__388_, data_stage_2__387_, data_stage_2__386_, data_stage_2__385_, data_stage_2__384_, data_stage_2__383_, data_stage_2__382_, data_stage_2__381_, data_stage_2__380_, data_stage_2__379_, data_stage_2__378_, data_stage_2__377_, data_stage_2__376_, data_stage_2__375_, data_stage_2__374_, data_stage_2__373_, data_stage_2__372_, data_stage_2__371_, data_stage_2__370_, data_stage_2__369_, data_stage_2__368_, data_stage_2__367_, data_stage_2__366_, data_stage_2__365_, data_stage_2__364_, data_stage_2__363_, data_stage_2__362_, data_stage_2__361_, data_stage_2__360_, data_stage_2__359_, data_stage_2__358_, data_stage_2__357_, data_stage_2__356_, data_stage_2__355_, data_stage_2__354_, data_stage_2__353_, data_stage_2__352_, data_stage_2__351_, data_stage_2__350_, data_stage_2__349_, data_stage_2__348_, data_stage_2__347_, data_stage_2__346_, data_stage_2__345_, data_stage_2__344_, data_stage_2__343_, data_stage_2__342_, data_stage_2__341_, data_stage_2__340_, data_stage_2__339_, data_stage_2__338_, data_stage_2__337_, data_stage_2__336_, data_stage_2__335_, data_stage_2__334_, data_stage_2__333_, data_stage_2__332_, data_stage_2__331_, data_stage_2__330_, data_stage_2__329_, data_stage_2__328_, data_stage_2__327_, data_stage_2__326_, data_stage_2__325_, data_stage_2__324_, data_stage_2__323_, data_stage_2__322_, data_stage_2__321_, data_stage_2__320_, data_stage_2__319_, data_stage_2__318_, data_stage_2__317_, data_stage_2__316_, data_stage_2__315_, data_stage_2__314_, data_stage_2__313_, data_stage_2__312_, data_stage_2__311_, data_stage_2__310_, data_stage_2__309_, data_stage_2__308_, data_stage_2__307_, data_stage_2__306_, data_stage_2__305_, data_stage_2__304_, data_stage_2__303_, data_stage_2__302_, data_stage_2__301_, data_stage_2__300_, data_stage_2__299_, data_stage_2__298_, data_stage_2__297_, data_stage_2__296_, data_stage_2__295_, data_stage_2__294_, data_stage_2__293_, data_stage_2__292_, data_stage_2__291_, data_stage_2__290_, data_stage_2__289_, data_stage_2__288_, data_stage_2__287_, data_stage_2__286_, data_stage_2__285_, data_stage_2__284_, data_stage_2__283_, data_stage_2__282_, data_stage_2__281_, data_stage_2__280_, data_stage_2__279_, data_stage_2__278_, data_stage_2__277_, data_stage_2__276_, data_stage_2__275_, data_stage_2__274_, data_stage_2__273_, data_stage_2__272_, data_stage_2__271_, data_stage_2__270_, data_stage_2__269_, data_stage_2__268_, data_stage_2__267_, data_stage_2__266_, data_stage_2__265_, data_stage_2__264_, data_stage_2__263_, data_stage_2__262_, data_stage_2__261_, data_stage_2__260_, data_stage_2__259_, data_stage_2__258_, data_stage_2__257_, data_stage_2__256_, data_stage_2__255_, data_stage_2__254_, data_stage_2__253_, data_stage_2__252_, data_stage_2__251_, data_stage_2__250_, data_stage_2__249_, data_stage_2__248_, data_stage_2__247_, data_stage_2__246_, data_stage_2__245_, data_stage_2__244_, data_stage_2__243_, data_stage_2__242_, data_stage_2__241_, data_stage_2__240_, data_stage_2__239_, data_stage_2__238_, data_stage_2__237_, data_stage_2__236_, data_stage_2__235_, data_stage_2__234_, data_stage_2__233_, data_stage_2__232_, data_stage_2__231_, data_stage_2__230_, data_stage_2__229_, data_stage_2__228_, data_stage_2__227_, data_stage_2__226_, data_stage_2__225_, data_stage_2__224_, data_stage_2__223_, data_stage_2__222_, data_stage_2__221_, data_stage_2__220_, data_stage_2__219_, data_stage_2__218_, data_stage_2__217_, data_stage_2__216_, data_stage_2__215_, data_stage_2__214_, data_stage_2__213_, data_stage_2__212_, data_stage_2__211_, data_stage_2__210_, data_stage_2__209_, data_stage_2__208_, data_stage_2__207_, data_stage_2__206_, data_stage_2__205_, data_stage_2__204_, data_stage_2__203_, data_stage_2__202_, data_stage_2__201_, data_stage_2__200_, data_stage_2__199_, data_stage_2__198_, data_stage_2__197_, data_stage_2__196_, data_stage_2__195_, data_stage_2__194_, data_stage_2__193_, data_stage_2__192_, data_stage_2__191_, data_stage_2__190_, data_stage_2__189_, data_stage_2__188_, data_stage_2__187_, data_stage_2__186_, data_stage_2__185_, data_stage_2__184_, data_stage_2__183_, data_stage_2__182_, data_stage_2__181_, data_stage_2__180_, data_stage_2__179_, data_stage_2__178_, data_stage_2__177_, data_stage_2__176_, data_stage_2__175_, data_stage_2__174_, data_stage_2__173_, data_stage_2__172_, data_stage_2__171_, data_stage_2__170_, data_stage_2__169_, data_stage_2__168_, data_stage_2__167_, data_stage_2__166_, data_stage_2__165_, data_stage_2__164_, data_stage_2__163_, data_stage_2__162_, data_stage_2__161_, data_stage_2__160_, data_stage_2__159_, data_stage_2__158_, data_stage_2__157_, data_stage_2__156_, data_stage_2__155_, data_stage_2__154_, data_stage_2__153_, data_stage_2__152_, data_stage_2__151_, data_stage_2__150_, data_stage_2__149_, data_stage_2__148_, data_stage_2__147_, data_stage_2__146_, data_stage_2__145_, data_stage_2__144_, data_stage_2__143_, data_stage_2__142_, data_stage_2__141_, data_stage_2__140_, data_stage_2__139_, data_stage_2__138_, data_stage_2__137_, data_stage_2__136_, data_stage_2__135_, data_stage_2__134_, data_stage_2__133_, data_stage_2__132_, data_stage_2__131_, data_stage_2__130_, data_stage_2__129_, data_stage_2__128_, data_stage_2__127_, data_stage_2__126_, data_stage_2__125_, data_stage_2__124_, data_stage_2__123_, data_stage_2__122_, data_stage_2__121_, data_stage_2__120_, data_stage_2__119_, data_stage_2__118_, data_stage_2__117_, data_stage_2__116_, data_stage_2__115_, data_stage_2__114_, data_stage_2__113_, data_stage_2__112_, data_stage_2__111_, data_stage_2__110_, data_stage_2__109_, data_stage_2__108_, data_stage_2__107_, data_stage_2__106_, data_stage_2__105_, data_stage_2__104_, data_stage_2__103_, data_stage_2__102_, data_stage_2__101_, data_stage_2__100_, data_stage_2__99_, data_stage_2__98_, data_stage_2__97_, data_stage_2__96_, data_stage_2__95_, data_stage_2__94_, data_stage_2__93_, data_stage_2__92_, data_stage_2__91_, data_stage_2__90_, data_stage_2__89_, data_stage_2__88_, data_stage_2__87_, data_stage_2__86_, data_stage_2__85_, data_stage_2__84_, data_stage_2__83_, data_stage_2__82_, data_stage_2__81_, data_stage_2__80_, data_stage_2__79_, data_stage_2__78_, data_stage_2__77_, data_stage_2__76_, data_stage_2__75_, data_stage_2__74_, data_stage_2__73_, data_stage_2__72_, data_stage_2__71_, data_stage_2__70_, data_stage_2__69_, data_stage_2__68_, data_stage_2__67_, data_stage_2__66_, data_stage_2__65_, data_stage_2__64_, data_stage_2__63_, data_stage_2__62_, data_stage_2__61_, data_stage_2__60_, data_stage_2__59_, data_stage_2__58_, data_stage_2__57_, data_stage_2__56_, data_stage_2__55_, data_stage_2__54_, data_stage_2__53_, data_stage_2__52_, data_stage_2__51_, data_stage_2__50_, data_stage_2__49_, data_stage_2__48_, data_stage_2__47_, data_stage_2__46_, data_stage_2__45_, data_stage_2__44_, data_stage_2__43_, data_stage_2__42_, data_stage_2__41_, data_stage_2__40_, data_stage_2__39_, data_stage_2__38_, data_stage_2__37_, data_stage_2__36_, data_stage_2__35_, data_stage_2__34_, data_stage_2__33_, data_stage_2__32_, data_stage_2__31_, data_stage_2__30_, data_stage_2__29_, data_stage_2__28_, data_stage_2__27_, data_stage_2__26_, data_stage_2__25_, data_stage_2__24_, data_stage_2__23_, data_stage_2__22_, data_stage_2__21_, data_stage_2__20_, data_stage_2__19_, data_stage_2__18_, data_stage_2__17_, data_stage_2__16_, data_stage_2__15_, data_stage_2__14_, data_stage_2__13_, data_stage_2__12_, data_stage_2__11_, data_stage_2__10_, data_stage_2__9_, data_stage_2__8_, data_stage_2__7_, data_stage_2__6_, data_stage_2__5_, data_stage_2__4_, data_stage_2__3_, data_stage_2__2_, data_stage_2__1_, data_stage_2__0_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__511_, data_stage_3__510_, data_stage_3__509_, data_stage_3__508_, data_stage_3__507_, data_stage_3__506_, data_stage_3__505_, data_stage_3__504_, data_stage_3__503_, data_stage_3__502_, data_stage_3__501_, data_stage_3__500_, data_stage_3__499_, data_stage_3__498_, data_stage_3__497_, data_stage_3__496_, data_stage_3__495_, data_stage_3__494_, data_stage_3__493_, data_stage_3__492_, data_stage_3__491_, data_stage_3__490_, data_stage_3__489_, data_stage_3__488_, data_stage_3__487_, data_stage_3__486_, data_stage_3__485_, data_stage_3__484_, data_stage_3__483_, data_stage_3__482_, data_stage_3__481_, data_stage_3__480_, data_stage_3__479_, data_stage_3__478_, data_stage_3__477_, data_stage_3__476_, data_stage_3__475_, data_stage_3__474_, data_stage_3__473_, data_stage_3__472_, data_stage_3__471_, data_stage_3__470_, data_stage_3__469_, data_stage_3__468_, data_stage_3__467_, data_stage_3__466_, data_stage_3__465_, data_stage_3__464_, data_stage_3__463_, data_stage_3__462_, data_stage_3__461_, data_stage_3__460_, data_stage_3__459_, data_stage_3__458_, data_stage_3__457_, data_stage_3__456_, data_stage_3__455_, data_stage_3__454_, data_stage_3__453_, data_stage_3__452_, data_stage_3__451_, data_stage_3__450_, data_stage_3__449_, data_stage_3__448_, data_stage_3__447_, data_stage_3__446_, data_stage_3__445_, data_stage_3__444_, data_stage_3__443_, data_stage_3__442_, data_stage_3__441_, data_stage_3__440_, data_stage_3__439_, data_stage_3__438_, data_stage_3__437_, data_stage_3__436_, data_stage_3__435_, data_stage_3__434_, data_stage_3__433_, data_stage_3__432_, data_stage_3__431_, data_stage_3__430_, data_stage_3__429_, data_stage_3__428_, data_stage_3__427_, data_stage_3__426_, data_stage_3__425_, data_stage_3__424_, data_stage_3__423_, data_stage_3__422_, data_stage_3__421_, data_stage_3__420_, data_stage_3__419_, data_stage_3__418_, data_stage_3__417_, data_stage_3__416_, data_stage_3__415_, data_stage_3__414_, data_stage_3__413_, data_stage_3__412_, data_stage_3__411_, data_stage_3__410_, data_stage_3__409_, data_stage_3__408_, data_stage_3__407_, data_stage_3__406_, data_stage_3__405_, data_stage_3__404_, data_stage_3__403_, data_stage_3__402_, data_stage_3__401_, data_stage_3__400_, data_stage_3__399_, data_stage_3__398_, data_stage_3__397_, data_stage_3__396_, data_stage_3__395_, data_stage_3__394_, data_stage_3__393_, data_stage_3__392_, data_stage_3__391_, data_stage_3__390_, data_stage_3__389_, data_stage_3__388_, data_stage_3__387_, data_stage_3__386_, data_stage_3__385_, data_stage_3__384_, data_stage_3__383_, data_stage_3__382_, data_stage_3__381_, data_stage_3__380_, data_stage_3__379_, data_stage_3__378_, data_stage_3__377_, data_stage_3__376_, data_stage_3__375_, data_stage_3__374_, data_stage_3__373_, data_stage_3__372_, data_stage_3__371_, data_stage_3__370_, data_stage_3__369_, data_stage_3__368_, data_stage_3__367_, data_stage_3__366_, data_stage_3__365_, data_stage_3__364_, data_stage_3__363_, data_stage_3__362_, data_stage_3__361_, data_stage_3__360_, data_stage_3__359_, data_stage_3__358_, data_stage_3__357_, data_stage_3__356_, data_stage_3__355_, data_stage_3__354_, data_stage_3__353_, data_stage_3__352_, data_stage_3__351_, data_stage_3__350_, data_stage_3__349_, data_stage_3__348_, data_stage_3__347_, data_stage_3__346_, data_stage_3__345_, data_stage_3__344_, data_stage_3__343_, data_stage_3__342_, data_stage_3__341_, data_stage_3__340_, data_stage_3__339_, data_stage_3__338_, data_stage_3__337_, data_stage_3__336_, data_stage_3__335_, data_stage_3__334_, data_stage_3__333_, data_stage_3__332_, data_stage_3__331_, data_stage_3__330_, data_stage_3__329_, data_stage_3__328_, data_stage_3__327_, data_stage_3__326_, data_stage_3__325_, data_stage_3__324_, data_stage_3__323_, data_stage_3__322_, data_stage_3__321_, data_stage_3__320_, data_stage_3__319_, data_stage_3__318_, data_stage_3__317_, data_stage_3__316_, data_stage_3__315_, data_stage_3__314_, data_stage_3__313_, data_stage_3__312_, data_stage_3__311_, data_stage_3__310_, data_stage_3__309_, data_stage_3__308_, data_stage_3__307_, data_stage_3__306_, data_stage_3__305_, data_stage_3__304_, data_stage_3__303_, data_stage_3__302_, data_stage_3__301_, data_stage_3__300_, data_stage_3__299_, data_stage_3__298_, data_stage_3__297_, data_stage_3__296_, data_stage_3__295_, data_stage_3__294_, data_stage_3__293_, data_stage_3__292_, data_stage_3__291_, data_stage_3__290_, data_stage_3__289_, data_stage_3__288_, data_stage_3__287_, data_stage_3__286_, data_stage_3__285_, data_stage_3__284_, data_stage_3__283_, data_stage_3__282_, data_stage_3__281_, data_stage_3__280_, data_stage_3__279_, data_stage_3__278_, data_stage_3__277_, data_stage_3__276_, data_stage_3__275_, data_stage_3__274_, data_stage_3__273_, data_stage_3__272_, data_stage_3__271_, data_stage_3__270_, data_stage_3__269_, data_stage_3__268_, data_stage_3__267_, data_stage_3__266_, data_stage_3__265_, data_stage_3__264_, data_stage_3__263_, data_stage_3__262_, data_stage_3__261_, data_stage_3__260_, data_stage_3__259_, data_stage_3__258_, data_stage_3__257_, data_stage_3__256_, data_stage_3__255_, data_stage_3__254_, data_stage_3__253_, data_stage_3__252_, data_stage_3__251_, data_stage_3__250_, data_stage_3__249_, data_stage_3__248_, data_stage_3__247_, data_stage_3__246_, data_stage_3__245_, data_stage_3__244_, data_stage_3__243_, data_stage_3__242_, data_stage_3__241_, data_stage_3__240_, data_stage_3__239_, data_stage_3__238_, data_stage_3__237_, data_stage_3__236_, data_stage_3__235_, data_stage_3__234_, data_stage_3__233_, data_stage_3__232_, data_stage_3__231_, data_stage_3__230_, data_stage_3__229_, data_stage_3__228_, data_stage_3__227_, data_stage_3__226_, data_stage_3__225_, data_stage_3__224_, data_stage_3__223_, data_stage_3__222_, data_stage_3__221_, data_stage_3__220_, data_stage_3__219_, data_stage_3__218_, data_stage_3__217_, data_stage_3__216_, data_stage_3__215_, data_stage_3__214_, data_stage_3__213_, data_stage_3__212_, data_stage_3__211_, data_stage_3__210_, data_stage_3__209_, data_stage_3__208_, data_stage_3__207_, data_stage_3__206_, data_stage_3__205_, data_stage_3__204_, data_stage_3__203_, data_stage_3__202_, data_stage_3__201_, data_stage_3__200_, data_stage_3__199_, data_stage_3__198_, data_stage_3__197_, data_stage_3__196_, data_stage_3__195_, data_stage_3__194_, data_stage_3__193_, data_stage_3__192_, data_stage_3__191_, data_stage_3__190_, data_stage_3__189_, data_stage_3__188_, data_stage_3__187_, data_stage_3__186_, data_stage_3__185_, data_stage_3__184_, data_stage_3__183_, data_stage_3__182_, data_stage_3__181_, data_stage_3__180_, data_stage_3__179_, data_stage_3__178_, data_stage_3__177_, data_stage_3__176_, data_stage_3__175_, data_stage_3__174_, data_stage_3__173_, data_stage_3__172_, data_stage_3__171_, data_stage_3__170_, data_stage_3__169_, data_stage_3__168_, data_stage_3__167_, data_stage_3__166_, data_stage_3__165_, data_stage_3__164_, data_stage_3__163_, data_stage_3__162_, data_stage_3__161_, data_stage_3__160_, data_stage_3__159_, data_stage_3__158_, data_stage_3__157_, data_stage_3__156_, data_stage_3__155_, data_stage_3__154_, data_stage_3__153_, data_stage_3__152_, data_stage_3__151_, data_stage_3__150_, data_stage_3__149_, data_stage_3__148_, data_stage_3__147_, data_stage_3__146_, data_stage_3__145_, data_stage_3__144_, data_stage_3__143_, data_stage_3__142_, data_stage_3__141_, data_stage_3__140_, data_stage_3__139_, data_stage_3__138_, data_stage_3__137_, data_stage_3__136_, data_stage_3__135_, data_stage_3__134_, data_stage_3__133_, data_stage_3__132_, data_stage_3__131_, data_stage_3__130_, data_stage_3__129_, data_stage_3__128_, data_stage_3__127_, data_stage_3__126_, data_stage_3__125_, data_stage_3__124_, data_stage_3__123_, data_stage_3__122_, data_stage_3__121_, data_stage_3__120_, data_stage_3__119_, data_stage_3__118_, data_stage_3__117_, data_stage_3__116_, data_stage_3__115_, data_stage_3__114_, data_stage_3__113_, data_stage_3__112_, data_stage_3__111_, data_stage_3__110_, data_stage_3__109_, data_stage_3__108_, data_stage_3__107_, data_stage_3__106_, data_stage_3__105_, data_stage_3__104_, data_stage_3__103_, data_stage_3__102_, data_stage_3__101_, data_stage_3__100_, data_stage_3__99_, data_stage_3__98_, data_stage_3__97_, data_stage_3__96_, data_stage_3__95_, data_stage_3__94_, data_stage_3__93_, data_stage_3__92_, data_stage_3__91_, data_stage_3__90_, data_stage_3__89_, data_stage_3__88_, data_stage_3__87_, data_stage_3__86_, data_stage_3__85_, data_stage_3__84_, data_stage_3__83_, data_stage_3__82_, data_stage_3__81_, data_stage_3__80_, data_stage_3__79_, data_stage_3__78_, data_stage_3__77_, data_stage_3__76_, data_stage_3__75_, data_stage_3__74_, data_stage_3__73_, data_stage_3__72_, data_stage_3__71_, data_stage_3__70_, data_stage_3__69_, data_stage_3__68_, data_stage_3__67_, data_stage_3__66_, data_stage_3__65_, data_stage_3__64_, data_stage_3__63_, data_stage_3__62_, data_stage_3__61_, data_stage_3__60_, data_stage_3__59_, data_stage_3__58_, data_stage_3__57_, data_stage_3__56_, data_stage_3__55_, data_stage_3__54_, data_stage_3__53_, data_stage_3__52_, data_stage_3__51_, data_stage_3__50_, data_stage_3__49_, data_stage_3__48_, data_stage_3__47_, data_stage_3__46_, data_stage_3__45_, data_stage_3__44_, data_stage_3__43_, data_stage_3__42_, data_stage_3__41_, data_stage_3__40_, data_stage_3__39_, data_stage_3__38_, data_stage_3__37_, data_stage_3__36_, data_stage_3__35_, data_stage_3__34_, data_stage_3__33_, data_stage_3__32_, data_stage_3__31_, data_stage_3__30_, data_stage_3__29_, data_stage_3__28_, data_stage_3__27_, data_stage_3__26_, data_stage_3__25_, data_stage_3__24_, data_stage_3__23_, data_stage_3__22_, data_stage_3__21_, data_stage_3__20_, data_stage_3__19_, data_stage_3__18_, data_stage_3__17_, data_stage_3__16_, data_stage_3__15_, data_stage_3__14_, data_stage_3__13_, data_stage_3__12_, data_stage_3__11_, data_stage_3__10_, data_stage_3__9_, data_stage_3__8_, data_stage_3__7_, data_stage_3__6_, data_stage_3__5_, data_stage_3__4_, data_stage_3__3_, data_stage_3__2_, data_stage_3__1_, data_stage_3__0_ })
  );


  bsg_swap_width_p256
  mux_stage_2__mux_swap_1__swap_inst
  (
    .data_i({ data_stage_2__1023_, data_stage_2__1022_, data_stage_2__1021_, data_stage_2__1020_, data_stage_2__1019_, data_stage_2__1018_, data_stage_2__1017_, data_stage_2__1016_, data_stage_2__1015_, data_stage_2__1014_, data_stage_2__1013_, data_stage_2__1012_, data_stage_2__1011_, data_stage_2__1010_, data_stage_2__1009_, data_stage_2__1008_, data_stage_2__1007_, data_stage_2__1006_, data_stage_2__1005_, data_stage_2__1004_, data_stage_2__1003_, data_stage_2__1002_, data_stage_2__1001_, data_stage_2__1000_, data_stage_2__999_, data_stage_2__998_, data_stage_2__997_, data_stage_2__996_, data_stage_2__995_, data_stage_2__994_, data_stage_2__993_, data_stage_2__992_, data_stage_2__991_, data_stage_2__990_, data_stage_2__989_, data_stage_2__988_, data_stage_2__987_, data_stage_2__986_, data_stage_2__985_, data_stage_2__984_, data_stage_2__983_, data_stage_2__982_, data_stage_2__981_, data_stage_2__980_, data_stage_2__979_, data_stage_2__978_, data_stage_2__977_, data_stage_2__976_, data_stage_2__975_, data_stage_2__974_, data_stage_2__973_, data_stage_2__972_, data_stage_2__971_, data_stage_2__970_, data_stage_2__969_, data_stage_2__968_, data_stage_2__967_, data_stage_2__966_, data_stage_2__965_, data_stage_2__964_, data_stage_2__963_, data_stage_2__962_, data_stage_2__961_, data_stage_2__960_, data_stage_2__959_, data_stage_2__958_, data_stage_2__957_, data_stage_2__956_, data_stage_2__955_, data_stage_2__954_, data_stage_2__953_, data_stage_2__952_, data_stage_2__951_, data_stage_2__950_, data_stage_2__949_, data_stage_2__948_, data_stage_2__947_, data_stage_2__946_, data_stage_2__945_, data_stage_2__944_, data_stage_2__943_, data_stage_2__942_, data_stage_2__941_, data_stage_2__940_, data_stage_2__939_, data_stage_2__938_, data_stage_2__937_, data_stage_2__936_, data_stage_2__935_, data_stage_2__934_, data_stage_2__933_, data_stage_2__932_, data_stage_2__931_, data_stage_2__930_, data_stage_2__929_, data_stage_2__928_, data_stage_2__927_, data_stage_2__926_, data_stage_2__925_, data_stage_2__924_, data_stage_2__923_, data_stage_2__922_, data_stage_2__921_, data_stage_2__920_, data_stage_2__919_, data_stage_2__918_, data_stage_2__917_, data_stage_2__916_, data_stage_2__915_, data_stage_2__914_, data_stage_2__913_, data_stage_2__912_, data_stage_2__911_, data_stage_2__910_, data_stage_2__909_, data_stage_2__908_, data_stage_2__907_, data_stage_2__906_, data_stage_2__905_, data_stage_2__904_, data_stage_2__903_, data_stage_2__902_, data_stage_2__901_, data_stage_2__900_, data_stage_2__899_, data_stage_2__898_, data_stage_2__897_, data_stage_2__896_, data_stage_2__895_, data_stage_2__894_, data_stage_2__893_, data_stage_2__892_, data_stage_2__891_, data_stage_2__890_, data_stage_2__889_, data_stage_2__888_, data_stage_2__887_, data_stage_2__886_, data_stage_2__885_, data_stage_2__884_, data_stage_2__883_, data_stage_2__882_, data_stage_2__881_, data_stage_2__880_, data_stage_2__879_, data_stage_2__878_, data_stage_2__877_, data_stage_2__876_, data_stage_2__875_, data_stage_2__874_, data_stage_2__873_, data_stage_2__872_, data_stage_2__871_, data_stage_2__870_, data_stage_2__869_, data_stage_2__868_, data_stage_2__867_, data_stage_2__866_, data_stage_2__865_, data_stage_2__864_, data_stage_2__863_, data_stage_2__862_, data_stage_2__861_, data_stage_2__860_, data_stage_2__859_, data_stage_2__858_, data_stage_2__857_, data_stage_2__856_, data_stage_2__855_, data_stage_2__854_, data_stage_2__853_, data_stage_2__852_, data_stage_2__851_, data_stage_2__850_, data_stage_2__849_, data_stage_2__848_, data_stage_2__847_, data_stage_2__846_, data_stage_2__845_, data_stage_2__844_, data_stage_2__843_, data_stage_2__842_, data_stage_2__841_, data_stage_2__840_, data_stage_2__839_, data_stage_2__838_, data_stage_2__837_, data_stage_2__836_, data_stage_2__835_, data_stage_2__834_, data_stage_2__833_, data_stage_2__832_, data_stage_2__831_, data_stage_2__830_, data_stage_2__829_, data_stage_2__828_, data_stage_2__827_, data_stage_2__826_, data_stage_2__825_, data_stage_2__824_, data_stage_2__823_, data_stage_2__822_, data_stage_2__821_, data_stage_2__820_, data_stage_2__819_, data_stage_2__818_, data_stage_2__817_, data_stage_2__816_, data_stage_2__815_, data_stage_2__814_, data_stage_2__813_, data_stage_2__812_, data_stage_2__811_, data_stage_2__810_, data_stage_2__809_, data_stage_2__808_, data_stage_2__807_, data_stage_2__806_, data_stage_2__805_, data_stage_2__804_, data_stage_2__803_, data_stage_2__802_, data_stage_2__801_, data_stage_2__800_, data_stage_2__799_, data_stage_2__798_, data_stage_2__797_, data_stage_2__796_, data_stage_2__795_, data_stage_2__794_, data_stage_2__793_, data_stage_2__792_, data_stage_2__791_, data_stage_2__790_, data_stage_2__789_, data_stage_2__788_, data_stage_2__787_, data_stage_2__786_, data_stage_2__785_, data_stage_2__784_, data_stage_2__783_, data_stage_2__782_, data_stage_2__781_, data_stage_2__780_, data_stage_2__779_, data_stage_2__778_, data_stage_2__777_, data_stage_2__776_, data_stage_2__775_, data_stage_2__774_, data_stage_2__773_, data_stage_2__772_, data_stage_2__771_, data_stage_2__770_, data_stage_2__769_, data_stage_2__768_, data_stage_2__767_, data_stage_2__766_, data_stage_2__765_, data_stage_2__764_, data_stage_2__763_, data_stage_2__762_, data_stage_2__761_, data_stage_2__760_, data_stage_2__759_, data_stage_2__758_, data_stage_2__757_, data_stage_2__756_, data_stage_2__755_, data_stage_2__754_, data_stage_2__753_, data_stage_2__752_, data_stage_2__751_, data_stage_2__750_, data_stage_2__749_, data_stage_2__748_, data_stage_2__747_, data_stage_2__746_, data_stage_2__745_, data_stage_2__744_, data_stage_2__743_, data_stage_2__742_, data_stage_2__741_, data_stage_2__740_, data_stage_2__739_, data_stage_2__738_, data_stage_2__737_, data_stage_2__736_, data_stage_2__735_, data_stage_2__734_, data_stage_2__733_, data_stage_2__732_, data_stage_2__731_, data_stage_2__730_, data_stage_2__729_, data_stage_2__728_, data_stage_2__727_, data_stage_2__726_, data_stage_2__725_, data_stage_2__724_, data_stage_2__723_, data_stage_2__722_, data_stage_2__721_, data_stage_2__720_, data_stage_2__719_, data_stage_2__718_, data_stage_2__717_, data_stage_2__716_, data_stage_2__715_, data_stage_2__714_, data_stage_2__713_, data_stage_2__712_, data_stage_2__711_, data_stage_2__710_, data_stage_2__709_, data_stage_2__708_, data_stage_2__707_, data_stage_2__706_, data_stage_2__705_, data_stage_2__704_, data_stage_2__703_, data_stage_2__702_, data_stage_2__701_, data_stage_2__700_, data_stage_2__699_, data_stage_2__698_, data_stage_2__697_, data_stage_2__696_, data_stage_2__695_, data_stage_2__694_, data_stage_2__693_, data_stage_2__692_, data_stage_2__691_, data_stage_2__690_, data_stage_2__689_, data_stage_2__688_, data_stage_2__687_, data_stage_2__686_, data_stage_2__685_, data_stage_2__684_, data_stage_2__683_, data_stage_2__682_, data_stage_2__681_, data_stage_2__680_, data_stage_2__679_, data_stage_2__678_, data_stage_2__677_, data_stage_2__676_, data_stage_2__675_, data_stage_2__674_, data_stage_2__673_, data_stage_2__672_, data_stage_2__671_, data_stage_2__670_, data_stage_2__669_, data_stage_2__668_, data_stage_2__667_, data_stage_2__666_, data_stage_2__665_, data_stage_2__664_, data_stage_2__663_, data_stage_2__662_, data_stage_2__661_, data_stage_2__660_, data_stage_2__659_, data_stage_2__658_, data_stage_2__657_, data_stage_2__656_, data_stage_2__655_, data_stage_2__654_, data_stage_2__653_, data_stage_2__652_, data_stage_2__651_, data_stage_2__650_, data_stage_2__649_, data_stage_2__648_, data_stage_2__647_, data_stage_2__646_, data_stage_2__645_, data_stage_2__644_, data_stage_2__643_, data_stage_2__642_, data_stage_2__641_, data_stage_2__640_, data_stage_2__639_, data_stage_2__638_, data_stage_2__637_, data_stage_2__636_, data_stage_2__635_, data_stage_2__634_, data_stage_2__633_, data_stage_2__632_, data_stage_2__631_, data_stage_2__630_, data_stage_2__629_, data_stage_2__628_, data_stage_2__627_, data_stage_2__626_, data_stage_2__625_, data_stage_2__624_, data_stage_2__623_, data_stage_2__622_, data_stage_2__621_, data_stage_2__620_, data_stage_2__619_, data_stage_2__618_, data_stage_2__617_, data_stage_2__616_, data_stage_2__615_, data_stage_2__614_, data_stage_2__613_, data_stage_2__612_, data_stage_2__611_, data_stage_2__610_, data_stage_2__609_, data_stage_2__608_, data_stage_2__607_, data_stage_2__606_, data_stage_2__605_, data_stage_2__604_, data_stage_2__603_, data_stage_2__602_, data_stage_2__601_, data_stage_2__600_, data_stage_2__599_, data_stage_2__598_, data_stage_2__597_, data_stage_2__596_, data_stage_2__595_, data_stage_2__594_, data_stage_2__593_, data_stage_2__592_, data_stage_2__591_, data_stage_2__590_, data_stage_2__589_, data_stage_2__588_, data_stage_2__587_, data_stage_2__586_, data_stage_2__585_, data_stage_2__584_, data_stage_2__583_, data_stage_2__582_, data_stage_2__581_, data_stage_2__580_, data_stage_2__579_, data_stage_2__578_, data_stage_2__577_, data_stage_2__576_, data_stage_2__575_, data_stage_2__574_, data_stage_2__573_, data_stage_2__572_, data_stage_2__571_, data_stage_2__570_, data_stage_2__569_, data_stage_2__568_, data_stage_2__567_, data_stage_2__566_, data_stage_2__565_, data_stage_2__564_, data_stage_2__563_, data_stage_2__562_, data_stage_2__561_, data_stage_2__560_, data_stage_2__559_, data_stage_2__558_, data_stage_2__557_, data_stage_2__556_, data_stage_2__555_, data_stage_2__554_, data_stage_2__553_, data_stage_2__552_, data_stage_2__551_, data_stage_2__550_, data_stage_2__549_, data_stage_2__548_, data_stage_2__547_, data_stage_2__546_, data_stage_2__545_, data_stage_2__544_, data_stage_2__543_, data_stage_2__542_, data_stage_2__541_, data_stage_2__540_, data_stage_2__539_, data_stage_2__538_, data_stage_2__537_, data_stage_2__536_, data_stage_2__535_, data_stage_2__534_, data_stage_2__533_, data_stage_2__532_, data_stage_2__531_, data_stage_2__530_, data_stage_2__529_, data_stage_2__528_, data_stage_2__527_, data_stage_2__526_, data_stage_2__525_, data_stage_2__524_, data_stage_2__523_, data_stage_2__522_, data_stage_2__521_, data_stage_2__520_, data_stage_2__519_, data_stage_2__518_, data_stage_2__517_, data_stage_2__516_, data_stage_2__515_, data_stage_2__514_, data_stage_2__513_, data_stage_2__512_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__1023_, data_stage_3__1022_, data_stage_3__1021_, data_stage_3__1020_, data_stage_3__1019_, data_stage_3__1018_, data_stage_3__1017_, data_stage_3__1016_, data_stage_3__1015_, data_stage_3__1014_, data_stage_3__1013_, data_stage_3__1012_, data_stage_3__1011_, data_stage_3__1010_, data_stage_3__1009_, data_stage_3__1008_, data_stage_3__1007_, data_stage_3__1006_, data_stage_3__1005_, data_stage_3__1004_, data_stage_3__1003_, data_stage_3__1002_, data_stage_3__1001_, data_stage_3__1000_, data_stage_3__999_, data_stage_3__998_, data_stage_3__997_, data_stage_3__996_, data_stage_3__995_, data_stage_3__994_, data_stage_3__993_, data_stage_3__992_, data_stage_3__991_, data_stage_3__990_, data_stage_3__989_, data_stage_3__988_, data_stage_3__987_, data_stage_3__986_, data_stage_3__985_, data_stage_3__984_, data_stage_3__983_, data_stage_3__982_, data_stage_3__981_, data_stage_3__980_, data_stage_3__979_, data_stage_3__978_, data_stage_3__977_, data_stage_3__976_, data_stage_3__975_, data_stage_3__974_, data_stage_3__973_, data_stage_3__972_, data_stage_3__971_, data_stage_3__970_, data_stage_3__969_, data_stage_3__968_, data_stage_3__967_, data_stage_3__966_, data_stage_3__965_, data_stage_3__964_, data_stage_3__963_, data_stage_3__962_, data_stage_3__961_, data_stage_3__960_, data_stage_3__959_, data_stage_3__958_, data_stage_3__957_, data_stage_3__956_, data_stage_3__955_, data_stage_3__954_, data_stage_3__953_, data_stage_3__952_, data_stage_3__951_, data_stage_3__950_, data_stage_3__949_, data_stage_3__948_, data_stage_3__947_, data_stage_3__946_, data_stage_3__945_, data_stage_3__944_, data_stage_3__943_, data_stage_3__942_, data_stage_3__941_, data_stage_3__940_, data_stage_3__939_, data_stage_3__938_, data_stage_3__937_, data_stage_3__936_, data_stage_3__935_, data_stage_3__934_, data_stage_3__933_, data_stage_3__932_, data_stage_3__931_, data_stage_3__930_, data_stage_3__929_, data_stage_3__928_, data_stage_3__927_, data_stage_3__926_, data_stage_3__925_, data_stage_3__924_, data_stage_3__923_, data_stage_3__922_, data_stage_3__921_, data_stage_3__920_, data_stage_3__919_, data_stage_3__918_, data_stage_3__917_, data_stage_3__916_, data_stage_3__915_, data_stage_3__914_, data_stage_3__913_, data_stage_3__912_, data_stage_3__911_, data_stage_3__910_, data_stage_3__909_, data_stage_3__908_, data_stage_3__907_, data_stage_3__906_, data_stage_3__905_, data_stage_3__904_, data_stage_3__903_, data_stage_3__902_, data_stage_3__901_, data_stage_3__900_, data_stage_3__899_, data_stage_3__898_, data_stage_3__897_, data_stage_3__896_, data_stage_3__895_, data_stage_3__894_, data_stage_3__893_, data_stage_3__892_, data_stage_3__891_, data_stage_3__890_, data_stage_3__889_, data_stage_3__888_, data_stage_3__887_, data_stage_3__886_, data_stage_3__885_, data_stage_3__884_, data_stage_3__883_, data_stage_3__882_, data_stage_3__881_, data_stage_3__880_, data_stage_3__879_, data_stage_3__878_, data_stage_3__877_, data_stage_3__876_, data_stage_3__875_, data_stage_3__874_, data_stage_3__873_, data_stage_3__872_, data_stage_3__871_, data_stage_3__870_, data_stage_3__869_, data_stage_3__868_, data_stage_3__867_, data_stage_3__866_, data_stage_3__865_, data_stage_3__864_, data_stage_3__863_, data_stage_3__862_, data_stage_3__861_, data_stage_3__860_, data_stage_3__859_, data_stage_3__858_, data_stage_3__857_, data_stage_3__856_, data_stage_3__855_, data_stage_3__854_, data_stage_3__853_, data_stage_3__852_, data_stage_3__851_, data_stage_3__850_, data_stage_3__849_, data_stage_3__848_, data_stage_3__847_, data_stage_3__846_, data_stage_3__845_, data_stage_3__844_, data_stage_3__843_, data_stage_3__842_, data_stage_3__841_, data_stage_3__840_, data_stage_3__839_, data_stage_3__838_, data_stage_3__837_, data_stage_3__836_, data_stage_3__835_, data_stage_3__834_, data_stage_3__833_, data_stage_3__832_, data_stage_3__831_, data_stage_3__830_, data_stage_3__829_, data_stage_3__828_, data_stage_3__827_, data_stage_3__826_, data_stage_3__825_, data_stage_3__824_, data_stage_3__823_, data_stage_3__822_, data_stage_3__821_, data_stage_3__820_, data_stage_3__819_, data_stage_3__818_, data_stage_3__817_, data_stage_3__816_, data_stage_3__815_, data_stage_3__814_, data_stage_3__813_, data_stage_3__812_, data_stage_3__811_, data_stage_3__810_, data_stage_3__809_, data_stage_3__808_, data_stage_3__807_, data_stage_3__806_, data_stage_3__805_, data_stage_3__804_, data_stage_3__803_, data_stage_3__802_, data_stage_3__801_, data_stage_3__800_, data_stage_3__799_, data_stage_3__798_, data_stage_3__797_, data_stage_3__796_, data_stage_3__795_, data_stage_3__794_, data_stage_3__793_, data_stage_3__792_, data_stage_3__791_, data_stage_3__790_, data_stage_3__789_, data_stage_3__788_, data_stage_3__787_, data_stage_3__786_, data_stage_3__785_, data_stage_3__784_, data_stage_3__783_, data_stage_3__782_, data_stage_3__781_, data_stage_3__780_, data_stage_3__779_, data_stage_3__778_, data_stage_3__777_, data_stage_3__776_, data_stage_3__775_, data_stage_3__774_, data_stage_3__773_, data_stage_3__772_, data_stage_3__771_, data_stage_3__770_, data_stage_3__769_, data_stage_3__768_, data_stage_3__767_, data_stage_3__766_, data_stage_3__765_, data_stage_3__764_, data_stage_3__763_, data_stage_3__762_, data_stage_3__761_, data_stage_3__760_, data_stage_3__759_, data_stage_3__758_, data_stage_3__757_, data_stage_3__756_, data_stage_3__755_, data_stage_3__754_, data_stage_3__753_, data_stage_3__752_, data_stage_3__751_, data_stage_3__750_, data_stage_3__749_, data_stage_3__748_, data_stage_3__747_, data_stage_3__746_, data_stage_3__745_, data_stage_3__744_, data_stage_3__743_, data_stage_3__742_, data_stage_3__741_, data_stage_3__740_, data_stage_3__739_, data_stage_3__738_, data_stage_3__737_, data_stage_3__736_, data_stage_3__735_, data_stage_3__734_, data_stage_3__733_, data_stage_3__732_, data_stage_3__731_, data_stage_3__730_, data_stage_3__729_, data_stage_3__728_, data_stage_3__727_, data_stage_3__726_, data_stage_3__725_, data_stage_3__724_, data_stage_3__723_, data_stage_3__722_, data_stage_3__721_, data_stage_3__720_, data_stage_3__719_, data_stage_3__718_, data_stage_3__717_, data_stage_3__716_, data_stage_3__715_, data_stage_3__714_, data_stage_3__713_, data_stage_3__712_, data_stage_3__711_, data_stage_3__710_, data_stage_3__709_, data_stage_3__708_, data_stage_3__707_, data_stage_3__706_, data_stage_3__705_, data_stage_3__704_, data_stage_3__703_, data_stage_3__702_, data_stage_3__701_, data_stage_3__700_, data_stage_3__699_, data_stage_3__698_, data_stage_3__697_, data_stage_3__696_, data_stage_3__695_, data_stage_3__694_, data_stage_3__693_, data_stage_3__692_, data_stage_3__691_, data_stage_3__690_, data_stage_3__689_, data_stage_3__688_, data_stage_3__687_, data_stage_3__686_, data_stage_3__685_, data_stage_3__684_, data_stage_3__683_, data_stage_3__682_, data_stage_3__681_, data_stage_3__680_, data_stage_3__679_, data_stage_3__678_, data_stage_3__677_, data_stage_3__676_, data_stage_3__675_, data_stage_3__674_, data_stage_3__673_, data_stage_3__672_, data_stage_3__671_, data_stage_3__670_, data_stage_3__669_, data_stage_3__668_, data_stage_3__667_, data_stage_3__666_, data_stage_3__665_, data_stage_3__664_, data_stage_3__663_, data_stage_3__662_, data_stage_3__661_, data_stage_3__660_, data_stage_3__659_, data_stage_3__658_, data_stage_3__657_, data_stage_3__656_, data_stage_3__655_, data_stage_3__654_, data_stage_3__653_, data_stage_3__652_, data_stage_3__651_, data_stage_3__650_, data_stage_3__649_, data_stage_3__648_, data_stage_3__647_, data_stage_3__646_, data_stage_3__645_, data_stage_3__644_, data_stage_3__643_, data_stage_3__642_, data_stage_3__641_, data_stage_3__640_, data_stage_3__639_, data_stage_3__638_, data_stage_3__637_, data_stage_3__636_, data_stage_3__635_, data_stage_3__634_, data_stage_3__633_, data_stage_3__632_, data_stage_3__631_, data_stage_3__630_, data_stage_3__629_, data_stage_3__628_, data_stage_3__627_, data_stage_3__626_, data_stage_3__625_, data_stage_3__624_, data_stage_3__623_, data_stage_3__622_, data_stage_3__621_, data_stage_3__620_, data_stage_3__619_, data_stage_3__618_, data_stage_3__617_, data_stage_3__616_, data_stage_3__615_, data_stage_3__614_, data_stage_3__613_, data_stage_3__612_, data_stage_3__611_, data_stage_3__610_, data_stage_3__609_, data_stage_3__608_, data_stage_3__607_, data_stage_3__606_, data_stage_3__605_, data_stage_3__604_, data_stage_3__603_, data_stage_3__602_, data_stage_3__601_, data_stage_3__600_, data_stage_3__599_, data_stage_3__598_, data_stage_3__597_, data_stage_3__596_, data_stage_3__595_, data_stage_3__594_, data_stage_3__593_, data_stage_3__592_, data_stage_3__591_, data_stage_3__590_, data_stage_3__589_, data_stage_3__588_, data_stage_3__587_, data_stage_3__586_, data_stage_3__585_, data_stage_3__584_, data_stage_3__583_, data_stage_3__582_, data_stage_3__581_, data_stage_3__580_, data_stage_3__579_, data_stage_3__578_, data_stage_3__577_, data_stage_3__576_, data_stage_3__575_, data_stage_3__574_, data_stage_3__573_, data_stage_3__572_, data_stage_3__571_, data_stage_3__570_, data_stage_3__569_, data_stage_3__568_, data_stage_3__567_, data_stage_3__566_, data_stage_3__565_, data_stage_3__564_, data_stage_3__563_, data_stage_3__562_, data_stage_3__561_, data_stage_3__560_, data_stage_3__559_, data_stage_3__558_, data_stage_3__557_, data_stage_3__556_, data_stage_3__555_, data_stage_3__554_, data_stage_3__553_, data_stage_3__552_, data_stage_3__551_, data_stage_3__550_, data_stage_3__549_, data_stage_3__548_, data_stage_3__547_, data_stage_3__546_, data_stage_3__545_, data_stage_3__544_, data_stage_3__543_, data_stage_3__542_, data_stage_3__541_, data_stage_3__540_, data_stage_3__539_, data_stage_3__538_, data_stage_3__537_, data_stage_3__536_, data_stage_3__535_, data_stage_3__534_, data_stage_3__533_, data_stage_3__532_, data_stage_3__531_, data_stage_3__530_, data_stage_3__529_, data_stage_3__528_, data_stage_3__527_, data_stage_3__526_, data_stage_3__525_, data_stage_3__524_, data_stage_3__523_, data_stage_3__522_, data_stage_3__521_, data_stage_3__520_, data_stage_3__519_, data_stage_3__518_, data_stage_3__517_, data_stage_3__516_, data_stage_3__515_, data_stage_3__514_, data_stage_3__513_, data_stage_3__512_ })
  );


  bsg_swap_width_p256
  mux_stage_2__mux_swap_2__swap_inst
  (
    .data_i({ data_stage_2__1535_, data_stage_2__1534_, data_stage_2__1533_, data_stage_2__1532_, data_stage_2__1531_, data_stage_2__1530_, data_stage_2__1529_, data_stage_2__1528_, data_stage_2__1527_, data_stage_2__1526_, data_stage_2__1525_, data_stage_2__1524_, data_stage_2__1523_, data_stage_2__1522_, data_stage_2__1521_, data_stage_2__1520_, data_stage_2__1519_, data_stage_2__1518_, data_stage_2__1517_, data_stage_2__1516_, data_stage_2__1515_, data_stage_2__1514_, data_stage_2__1513_, data_stage_2__1512_, data_stage_2__1511_, data_stage_2__1510_, data_stage_2__1509_, data_stage_2__1508_, data_stage_2__1507_, data_stage_2__1506_, data_stage_2__1505_, data_stage_2__1504_, data_stage_2__1503_, data_stage_2__1502_, data_stage_2__1501_, data_stage_2__1500_, data_stage_2__1499_, data_stage_2__1498_, data_stage_2__1497_, data_stage_2__1496_, data_stage_2__1495_, data_stage_2__1494_, data_stage_2__1493_, data_stage_2__1492_, data_stage_2__1491_, data_stage_2__1490_, data_stage_2__1489_, data_stage_2__1488_, data_stage_2__1487_, data_stage_2__1486_, data_stage_2__1485_, data_stage_2__1484_, data_stage_2__1483_, data_stage_2__1482_, data_stage_2__1481_, data_stage_2__1480_, data_stage_2__1479_, data_stage_2__1478_, data_stage_2__1477_, data_stage_2__1476_, data_stage_2__1475_, data_stage_2__1474_, data_stage_2__1473_, data_stage_2__1472_, data_stage_2__1471_, data_stage_2__1470_, data_stage_2__1469_, data_stage_2__1468_, data_stage_2__1467_, data_stage_2__1466_, data_stage_2__1465_, data_stage_2__1464_, data_stage_2__1463_, data_stage_2__1462_, data_stage_2__1461_, data_stage_2__1460_, data_stage_2__1459_, data_stage_2__1458_, data_stage_2__1457_, data_stage_2__1456_, data_stage_2__1455_, data_stage_2__1454_, data_stage_2__1453_, data_stage_2__1452_, data_stage_2__1451_, data_stage_2__1450_, data_stage_2__1449_, data_stage_2__1448_, data_stage_2__1447_, data_stage_2__1446_, data_stage_2__1445_, data_stage_2__1444_, data_stage_2__1443_, data_stage_2__1442_, data_stage_2__1441_, data_stage_2__1440_, data_stage_2__1439_, data_stage_2__1438_, data_stage_2__1437_, data_stage_2__1436_, data_stage_2__1435_, data_stage_2__1434_, data_stage_2__1433_, data_stage_2__1432_, data_stage_2__1431_, data_stage_2__1430_, data_stage_2__1429_, data_stage_2__1428_, data_stage_2__1427_, data_stage_2__1426_, data_stage_2__1425_, data_stage_2__1424_, data_stage_2__1423_, data_stage_2__1422_, data_stage_2__1421_, data_stage_2__1420_, data_stage_2__1419_, data_stage_2__1418_, data_stage_2__1417_, data_stage_2__1416_, data_stage_2__1415_, data_stage_2__1414_, data_stage_2__1413_, data_stage_2__1412_, data_stage_2__1411_, data_stage_2__1410_, data_stage_2__1409_, data_stage_2__1408_, data_stage_2__1407_, data_stage_2__1406_, data_stage_2__1405_, data_stage_2__1404_, data_stage_2__1403_, data_stage_2__1402_, data_stage_2__1401_, data_stage_2__1400_, data_stage_2__1399_, data_stage_2__1398_, data_stage_2__1397_, data_stage_2__1396_, data_stage_2__1395_, data_stage_2__1394_, data_stage_2__1393_, data_stage_2__1392_, data_stage_2__1391_, data_stage_2__1390_, data_stage_2__1389_, data_stage_2__1388_, data_stage_2__1387_, data_stage_2__1386_, data_stage_2__1385_, data_stage_2__1384_, data_stage_2__1383_, data_stage_2__1382_, data_stage_2__1381_, data_stage_2__1380_, data_stage_2__1379_, data_stage_2__1378_, data_stage_2__1377_, data_stage_2__1376_, data_stage_2__1375_, data_stage_2__1374_, data_stage_2__1373_, data_stage_2__1372_, data_stage_2__1371_, data_stage_2__1370_, data_stage_2__1369_, data_stage_2__1368_, data_stage_2__1367_, data_stage_2__1366_, data_stage_2__1365_, data_stage_2__1364_, data_stage_2__1363_, data_stage_2__1362_, data_stage_2__1361_, data_stage_2__1360_, data_stage_2__1359_, data_stage_2__1358_, data_stage_2__1357_, data_stage_2__1356_, data_stage_2__1355_, data_stage_2__1354_, data_stage_2__1353_, data_stage_2__1352_, data_stage_2__1351_, data_stage_2__1350_, data_stage_2__1349_, data_stage_2__1348_, data_stage_2__1347_, data_stage_2__1346_, data_stage_2__1345_, data_stage_2__1344_, data_stage_2__1343_, data_stage_2__1342_, data_stage_2__1341_, data_stage_2__1340_, data_stage_2__1339_, data_stage_2__1338_, data_stage_2__1337_, data_stage_2__1336_, data_stage_2__1335_, data_stage_2__1334_, data_stage_2__1333_, data_stage_2__1332_, data_stage_2__1331_, data_stage_2__1330_, data_stage_2__1329_, data_stage_2__1328_, data_stage_2__1327_, data_stage_2__1326_, data_stage_2__1325_, data_stage_2__1324_, data_stage_2__1323_, data_stage_2__1322_, data_stage_2__1321_, data_stage_2__1320_, data_stage_2__1319_, data_stage_2__1318_, data_stage_2__1317_, data_stage_2__1316_, data_stage_2__1315_, data_stage_2__1314_, data_stage_2__1313_, data_stage_2__1312_, data_stage_2__1311_, data_stage_2__1310_, data_stage_2__1309_, data_stage_2__1308_, data_stage_2__1307_, data_stage_2__1306_, data_stage_2__1305_, data_stage_2__1304_, data_stage_2__1303_, data_stage_2__1302_, data_stage_2__1301_, data_stage_2__1300_, data_stage_2__1299_, data_stage_2__1298_, data_stage_2__1297_, data_stage_2__1296_, data_stage_2__1295_, data_stage_2__1294_, data_stage_2__1293_, data_stage_2__1292_, data_stage_2__1291_, data_stage_2__1290_, data_stage_2__1289_, data_stage_2__1288_, data_stage_2__1287_, data_stage_2__1286_, data_stage_2__1285_, data_stage_2__1284_, data_stage_2__1283_, data_stage_2__1282_, data_stage_2__1281_, data_stage_2__1280_, data_stage_2__1279_, data_stage_2__1278_, data_stage_2__1277_, data_stage_2__1276_, data_stage_2__1275_, data_stage_2__1274_, data_stage_2__1273_, data_stage_2__1272_, data_stage_2__1271_, data_stage_2__1270_, data_stage_2__1269_, data_stage_2__1268_, data_stage_2__1267_, data_stage_2__1266_, data_stage_2__1265_, data_stage_2__1264_, data_stage_2__1263_, data_stage_2__1262_, data_stage_2__1261_, data_stage_2__1260_, data_stage_2__1259_, data_stage_2__1258_, data_stage_2__1257_, data_stage_2__1256_, data_stage_2__1255_, data_stage_2__1254_, data_stage_2__1253_, data_stage_2__1252_, data_stage_2__1251_, data_stage_2__1250_, data_stage_2__1249_, data_stage_2__1248_, data_stage_2__1247_, data_stage_2__1246_, data_stage_2__1245_, data_stage_2__1244_, data_stage_2__1243_, data_stage_2__1242_, data_stage_2__1241_, data_stage_2__1240_, data_stage_2__1239_, data_stage_2__1238_, data_stage_2__1237_, data_stage_2__1236_, data_stage_2__1235_, data_stage_2__1234_, data_stage_2__1233_, data_stage_2__1232_, data_stage_2__1231_, data_stage_2__1230_, data_stage_2__1229_, data_stage_2__1228_, data_stage_2__1227_, data_stage_2__1226_, data_stage_2__1225_, data_stage_2__1224_, data_stage_2__1223_, data_stage_2__1222_, data_stage_2__1221_, data_stage_2__1220_, data_stage_2__1219_, data_stage_2__1218_, data_stage_2__1217_, data_stage_2__1216_, data_stage_2__1215_, data_stage_2__1214_, data_stage_2__1213_, data_stage_2__1212_, data_stage_2__1211_, data_stage_2__1210_, data_stage_2__1209_, data_stage_2__1208_, data_stage_2__1207_, data_stage_2__1206_, data_stage_2__1205_, data_stage_2__1204_, data_stage_2__1203_, data_stage_2__1202_, data_stage_2__1201_, data_stage_2__1200_, data_stage_2__1199_, data_stage_2__1198_, data_stage_2__1197_, data_stage_2__1196_, data_stage_2__1195_, data_stage_2__1194_, data_stage_2__1193_, data_stage_2__1192_, data_stage_2__1191_, data_stage_2__1190_, data_stage_2__1189_, data_stage_2__1188_, data_stage_2__1187_, data_stage_2__1186_, data_stage_2__1185_, data_stage_2__1184_, data_stage_2__1183_, data_stage_2__1182_, data_stage_2__1181_, data_stage_2__1180_, data_stage_2__1179_, data_stage_2__1178_, data_stage_2__1177_, data_stage_2__1176_, data_stage_2__1175_, data_stage_2__1174_, data_stage_2__1173_, data_stage_2__1172_, data_stage_2__1171_, data_stage_2__1170_, data_stage_2__1169_, data_stage_2__1168_, data_stage_2__1167_, data_stage_2__1166_, data_stage_2__1165_, data_stage_2__1164_, data_stage_2__1163_, data_stage_2__1162_, data_stage_2__1161_, data_stage_2__1160_, data_stage_2__1159_, data_stage_2__1158_, data_stage_2__1157_, data_stage_2__1156_, data_stage_2__1155_, data_stage_2__1154_, data_stage_2__1153_, data_stage_2__1152_, data_stage_2__1151_, data_stage_2__1150_, data_stage_2__1149_, data_stage_2__1148_, data_stage_2__1147_, data_stage_2__1146_, data_stage_2__1145_, data_stage_2__1144_, data_stage_2__1143_, data_stage_2__1142_, data_stage_2__1141_, data_stage_2__1140_, data_stage_2__1139_, data_stage_2__1138_, data_stage_2__1137_, data_stage_2__1136_, data_stage_2__1135_, data_stage_2__1134_, data_stage_2__1133_, data_stage_2__1132_, data_stage_2__1131_, data_stage_2__1130_, data_stage_2__1129_, data_stage_2__1128_, data_stage_2__1127_, data_stage_2__1126_, data_stage_2__1125_, data_stage_2__1124_, data_stage_2__1123_, data_stage_2__1122_, data_stage_2__1121_, data_stage_2__1120_, data_stage_2__1119_, data_stage_2__1118_, data_stage_2__1117_, data_stage_2__1116_, data_stage_2__1115_, data_stage_2__1114_, data_stage_2__1113_, data_stage_2__1112_, data_stage_2__1111_, data_stage_2__1110_, data_stage_2__1109_, data_stage_2__1108_, data_stage_2__1107_, data_stage_2__1106_, data_stage_2__1105_, data_stage_2__1104_, data_stage_2__1103_, data_stage_2__1102_, data_stage_2__1101_, data_stage_2__1100_, data_stage_2__1099_, data_stage_2__1098_, data_stage_2__1097_, data_stage_2__1096_, data_stage_2__1095_, data_stage_2__1094_, data_stage_2__1093_, data_stage_2__1092_, data_stage_2__1091_, data_stage_2__1090_, data_stage_2__1089_, data_stage_2__1088_, data_stage_2__1087_, data_stage_2__1086_, data_stage_2__1085_, data_stage_2__1084_, data_stage_2__1083_, data_stage_2__1082_, data_stage_2__1081_, data_stage_2__1080_, data_stage_2__1079_, data_stage_2__1078_, data_stage_2__1077_, data_stage_2__1076_, data_stage_2__1075_, data_stage_2__1074_, data_stage_2__1073_, data_stage_2__1072_, data_stage_2__1071_, data_stage_2__1070_, data_stage_2__1069_, data_stage_2__1068_, data_stage_2__1067_, data_stage_2__1066_, data_stage_2__1065_, data_stage_2__1064_, data_stage_2__1063_, data_stage_2__1062_, data_stage_2__1061_, data_stage_2__1060_, data_stage_2__1059_, data_stage_2__1058_, data_stage_2__1057_, data_stage_2__1056_, data_stage_2__1055_, data_stage_2__1054_, data_stage_2__1053_, data_stage_2__1052_, data_stage_2__1051_, data_stage_2__1050_, data_stage_2__1049_, data_stage_2__1048_, data_stage_2__1047_, data_stage_2__1046_, data_stage_2__1045_, data_stage_2__1044_, data_stage_2__1043_, data_stage_2__1042_, data_stage_2__1041_, data_stage_2__1040_, data_stage_2__1039_, data_stage_2__1038_, data_stage_2__1037_, data_stage_2__1036_, data_stage_2__1035_, data_stage_2__1034_, data_stage_2__1033_, data_stage_2__1032_, data_stage_2__1031_, data_stage_2__1030_, data_stage_2__1029_, data_stage_2__1028_, data_stage_2__1027_, data_stage_2__1026_, data_stage_2__1025_, data_stage_2__1024_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__1535_, data_stage_3__1534_, data_stage_3__1533_, data_stage_3__1532_, data_stage_3__1531_, data_stage_3__1530_, data_stage_3__1529_, data_stage_3__1528_, data_stage_3__1527_, data_stage_3__1526_, data_stage_3__1525_, data_stage_3__1524_, data_stage_3__1523_, data_stage_3__1522_, data_stage_3__1521_, data_stage_3__1520_, data_stage_3__1519_, data_stage_3__1518_, data_stage_3__1517_, data_stage_3__1516_, data_stage_3__1515_, data_stage_3__1514_, data_stage_3__1513_, data_stage_3__1512_, data_stage_3__1511_, data_stage_3__1510_, data_stage_3__1509_, data_stage_3__1508_, data_stage_3__1507_, data_stage_3__1506_, data_stage_3__1505_, data_stage_3__1504_, data_stage_3__1503_, data_stage_3__1502_, data_stage_3__1501_, data_stage_3__1500_, data_stage_3__1499_, data_stage_3__1498_, data_stage_3__1497_, data_stage_3__1496_, data_stage_3__1495_, data_stage_3__1494_, data_stage_3__1493_, data_stage_3__1492_, data_stage_3__1491_, data_stage_3__1490_, data_stage_3__1489_, data_stage_3__1488_, data_stage_3__1487_, data_stage_3__1486_, data_stage_3__1485_, data_stage_3__1484_, data_stage_3__1483_, data_stage_3__1482_, data_stage_3__1481_, data_stage_3__1480_, data_stage_3__1479_, data_stage_3__1478_, data_stage_3__1477_, data_stage_3__1476_, data_stage_3__1475_, data_stage_3__1474_, data_stage_3__1473_, data_stage_3__1472_, data_stage_3__1471_, data_stage_3__1470_, data_stage_3__1469_, data_stage_3__1468_, data_stage_3__1467_, data_stage_3__1466_, data_stage_3__1465_, data_stage_3__1464_, data_stage_3__1463_, data_stage_3__1462_, data_stage_3__1461_, data_stage_3__1460_, data_stage_3__1459_, data_stage_3__1458_, data_stage_3__1457_, data_stage_3__1456_, data_stage_3__1455_, data_stage_3__1454_, data_stage_3__1453_, data_stage_3__1452_, data_stage_3__1451_, data_stage_3__1450_, data_stage_3__1449_, data_stage_3__1448_, data_stage_3__1447_, data_stage_3__1446_, data_stage_3__1445_, data_stage_3__1444_, data_stage_3__1443_, data_stage_3__1442_, data_stage_3__1441_, data_stage_3__1440_, data_stage_3__1439_, data_stage_3__1438_, data_stage_3__1437_, data_stage_3__1436_, data_stage_3__1435_, data_stage_3__1434_, data_stage_3__1433_, data_stage_3__1432_, data_stage_3__1431_, data_stage_3__1430_, data_stage_3__1429_, data_stage_3__1428_, data_stage_3__1427_, data_stage_3__1426_, data_stage_3__1425_, data_stage_3__1424_, data_stage_3__1423_, data_stage_3__1422_, data_stage_3__1421_, data_stage_3__1420_, data_stage_3__1419_, data_stage_3__1418_, data_stage_3__1417_, data_stage_3__1416_, data_stage_3__1415_, data_stage_3__1414_, data_stage_3__1413_, data_stage_3__1412_, data_stage_3__1411_, data_stage_3__1410_, data_stage_3__1409_, data_stage_3__1408_, data_stage_3__1407_, data_stage_3__1406_, data_stage_3__1405_, data_stage_3__1404_, data_stage_3__1403_, data_stage_3__1402_, data_stage_3__1401_, data_stage_3__1400_, data_stage_3__1399_, data_stage_3__1398_, data_stage_3__1397_, data_stage_3__1396_, data_stage_3__1395_, data_stage_3__1394_, data_stage_3__1393_, data_stage_3__1392_, data_stage_3__1391_, data_stage_3__1390_, data_stage_3__1389_, data_stage_3__1388_, data_stage_3__1387_, data_stage_3__1386_, data_stage_3__1385_, data_stage_3__1384_, data_stage_3__1383_, data_stage_3__1382_, data_stage_3__1381_, data_stage_3__1380_, data_stage_3__1379_, data_stage_3__1378_, data_stage_3__1377_, data_stage_3__1376_, data_stage_3__1375_, data_stage_3__1374_, data_stage_3__1373_, data_stage_3__1372_, data_stage_3__1371_, data_stage_3__1370_, data_stage_3__1369_, data_stage_3__1368_, data_stage_3__1367_, data_stage_3__1366_, data_stage_3__1365_, data_stage_3__1364_, data_stage_3__1363_, data_stage_3__1362_, data_stage_3__1361_, data_stage_3__1360_, data_stage_3__1359_, data_stage_3__1358_, data_stage_3__1357_, data_stage_3__1356_, data_stage_3__1355_, data_stage_3__1354_, data_stage_3__1353_, data_stage_3__1352_, data_stage_3__1351_, data_stage_3__1350_, data_stage_3__1349_, data_stage_3__1348_, data_stage_3__1347_, data_stage_3__1346_, data_stage_3__1345_, data_stage_3__1344_, data_stage_3__1343_, data_stage_3__1342_, data_stage_3__1341_, data_stage_3__1340_, data_stage_3__1339_, data_stage_3__1338_, data_stage_3__1337_, data_stage_3__1336_, data_stage_3__1335_, data_stage_3__1334_, data_stage_3__1333_, data_stage_3__1332_, data_stage_3__1331_, data_stage_3__1330_, data_stage_3__1329_, data_stage_3__1328_, data_stage_3__1327_, data_stage_3__1326_, data_stage_3__1325_, data_stage_3__1324_, data_stage_3__1323_, data_stage_3__1322_, data_stage_3__1321_, data_stage_3__1320_, data_stage_3__1319_, data_stage_3__1318_, data_stage_3__1317_, data_stage_3__1316_, data_stage_3__1315_, data_stage_3__1314_, data_stage_3__1313_, data_stage_3__1312_, data_stage_3__1311_, data_stage_3__1310_, data_stage_3__1309_, data_stage_3__1308_, data_stage_3__1307_, data_stage_3__1306_, data_stage_3__1305_, data_stage_3__1304_, data_stage_3__1303_, data_stage_3__1302_, data_stage_3__1301_, data_stage_3__1300_, data_stage_3__1299_, data_stage_3__1298_, data_stage_3__1297_, data_stage_3__1296_, data_stage_3__1295_, data_stage_3__1294_, data_stage_3__1293_, data_stage_3__1292_, data_stage_3__1291_, data_stage_3__1290_, data_stage_3__1289_, data_stage_3__1288_, data_stage_3__1287_, data_stage_3__1286_, data_stage_3__1285_, data_stage_3__1284_, data_stage_3__1283_, data_stage_3__1282_, data_stage_3__1281_, data_stage_3__1280_, data_stage_3__1279_, data_stage_3__1278_, data_stage_3__1277_, data_stage_3__1276_, data_stage_3__1275_, data_stage_3__1274_, data_stage_3__1273_, data_stage_3__1272_, data_stage_3__1271_, data_stage_3__1270_, data_stage_3__1269_, data_stage_3__1268_, data_stage_3__1267_, data_stage_3__1266_, data_stage_3__1265_, data_stage_3__1264_, data_stage_3__1263_, data_stage_3__1262_, data_stage_3__1261_, data_stage_3__1260_, data_stage_3__1259_, data_stage_3__1258_, data_stage_3__1257_, data_stage_3__1256_, data_stage_3__1255_, data_stage_3__1254_, data_stage_3__1253_, data_stage_3__1252_, data_stage_3__1251_, data_stage_3__1250_, data_stage_3__1249_, data_stage_3__1248_, data_stage_3__1247_, data_stage_3__1246_, data_stage_3__1245_, data_stage_3__1244_, data_stage_3__1243_, data_stage_3__1242_, data_stage_3__1241_, data_stage_3__1240_, data_stage_3__1239_, data_stage_3__1238_, data_stage_3__1237_, data_stage_3__1236_, data_stage_3__1235_, data_stage_3__1234_, data_stage_3__1233_, data_stage_3__1232_, data_stage_3__1231_, data_stage_3__1230_, data_stage_3__1229_, data_stage_3__1228_, data_stage_3__1227_, data_stage_3__1226_, data_stage_3__1225_, data_stage_3__1224_, data_stage_3__1223_, data_stage_3__1222_, data_stage_3__1221_, data_stage_3__1220_, data_stage_3__1219_, data_stage_3__1218_, data_stage_3__1217_, data_stage_3__1216_, data_stage_3__1215_, data_stage_3__1214_, data_stage_3__1213_, data_stage_3__1212_, data_stage_3__1211_, data_stage_3__1210_, data_stage_3__1209_, data_stage_3__1208_, data_stage_3__1207_, data_stage_3__1206_, data_stage_3__1205_, data_stage_3__1204_, data_stage_3__1203_, data_stage_3__1202_, data_stage_3__1201_, data_stage_3__1200_, data_stage_3__1199_, data_stage_3__1198_, data_stage_3__1197_, data_stage_3__1196_, data_stage_3__1195_, data_stage_3__1194_, data_stage_3__1193_, data_stage_3__1192_, data_stage_3__1191_, data_stage_3__1190_, data_stage_3__1189_, data_stage_3__1188_, data_stage_3__1187_, data_stage_3__1186_, data_stage_3__1185_, data_stage_3__1184_, data_stage_3__1183_, data_stage_3__1182_, data_stage_3__1181_, data_stage_3__1180_, data_stage_3__1179_, data_stage_3__1178_, data_stage_3__1177_, data_stage_3__1176_, data_stage_3__1175_, data_stage_3__1174_, data_stage_3__1173_, data_stage_3__1172_, data_stage_3__1171_, data_stage_3__1170_, data_stage_3__1169_, data_stage_3__1168_, data_stage_3__1167_, data_stage_3__1166_, data_stage_3__1165_, data_stage_3__1164_, data_stage_3__1163_, data_stage_3__1162_, data_stage_3__1161_, data_stage_3__1160_, data_stage_3__1159_, data_stage_3__1158_, data_stage_3__1157_, data_stage_3__1156_, data_stage_3__1155_, data_stage_3__1154_, data_stage_3__1153_, data_stage_3__1152_, data_stage_3__1151_, data_stage_3__1150_, data_stage_3__1149_, data_stage_3__1148_, data_stage_3__1147_, data_stage_3__1146_, data_stage_3__1145_, data_stage_3__1144_, data_stage_3__1143_, data_stage_3__1142_, data_stage_3__1141_, data_stage_3__1140_, data_stage_3__1139_, data_stage_3__1138_, data_stage_3__1137_, data_stage_3__1136_, data_stage_3__1135_, data_stage_3__1134_, data_stage_3__1133_, data_stage_3__1132_, data_stage_3__1131_, data_stage_3__1130_, data_stage_3__1129_, data_stage_3__1128_, data_stage_3__1127_, data_stage_3__1126_, data_stage_3__1125_, data_stage_3__1124_, data_stage_3__1123_, data_stage_3__1122_, data_stage_3__1121_, data_stage_3__1120_, data_stage_3__1119_, data_stage_3__1118_, data_stage_3__1117_, data_stage_3__1116_, data_stage_3__1115_, data_stage_3__1114_, data_stage_3__1113_, data_stage_3__1112_, data_stage_3__1111_, data_stage_3__1110_, data_stage_3__1109_, data_stage_3__1108_, data_stage_3__1107_, data_stage_3__1106_, data_stage_3__1105_, data_stage_3__1104_, data_stage_3__1103_, data_stage_3__1102_, data_stage_3__1101_, data_stage_3__1100_, data_stage_3__1099_, data_stage_3__1098_, data_stage_3__1097_, data_stage_3__1096_, data_stage_3__1095_, data_stage_3__1094_, data_stage_3__1093_, data_stage_3__1092_, data_stage_3__1091_, data_stage_3__1090_, data_stage_3__1089_, data_stage_3__1088_, data_stage_3__1087_, data_stage_3__1086_, data_stage_3__1085_, data_stage_3__1084_, data_stage_3__1083_, data_stage_3__1082_, data_stage_3__1081_, data_stage_3__1080_, data_stage_3__1079_, data_stage_3__1078_, data_stage_3__1077_, data_stage_3__1076_, data_stage_3__1075_, data_stage_3__1074_, data_stage_3__1073_, data_stage_3__1072_, data_stage_3__1071_, data_stage_3__1070_, data_stage_3__1069_, data_stage_3__1068_, data_stage_3__1067_, data_stage_3__1066_, data_stage_3__1065_, data_stage_3__1064_, data_stage_3__1063_, data_stage_3__1062_, data_stage_3__1061_, data_stage_3__1060_, data_stage_3__1059_, data_stage_3__1058_, data_stage_3__1057_, data_stage_3__1056_, data_stage_3__1055_, data_stage_3__1054_, data_stage_3__1053_, data_stage_3__1052_, data_stage_3__1051_, data_stage_3__1050_, data_stage_3__1049_, data_stage_3__1048_, data_stage_3__1047_, data_stage_3__1046_, data_stage_3__1045_, data_stage_3__1044_, data_stage_3__1043_, data_stage_3__1042_, data_stage_3__1041_, data_stage_3__1040_, data_stage_3__1039_, data_stage_3__1038_, data_stage_3__1037_, data_stage_3__1036_, data_stage_3__1035_, data_stage_3__1034_, data_stage_3__1033_, data_stage_3__1032_, data_stage_3__1031_, data_stage_3__1030_, data_stage_3__1029_, data_stage_3__1028_, data_stage_3__1027_, data_stage_3__1026_, data_stage_3__1025_, data_stage_3__1024_ })
  );


  bsg_swap_width_p256
  mux_stage_2__mux_swap_3__swap_inst
  (
    .data_i({ data_stage_2__2047_, data_stage_2__2046_, data_stage_2__2045_, data_stage_2__2044_, data_stage_2__2043_, data_stage_2__2042_, data_stage_2__2041_, data_stage_2__2040_, data_stage_2__2039_, data_stage_2__2038_, data_stage_2__2037_, data_stage_2__2036_, data_stage_2__2035_, data_stage_2__2034_, data_stage_2__2033_, data_stage_2__2032_, data_stage_2__2031_, data_stage_2__2030_, data_stage_2__2029_, data_stage_2__2028_, data_stage_2__2027_, data_stage_2__2026_, data_stage_2__2025_, data_stage_2__2024_, data_stage_2__2023_, data_stage_2__2022_, data_stage_2__2021_, data_stage_2__2020_, data_stage_2__2019_, data_stage_2__2018_, data_stage_2__2017_, data_stage_2__2016_, data_stage_2__2015_, data_stage_2__2014_, data_stage_2__2013_, data_stage_2__2012_, data_stage_2__2011_, data_stage_2__2010_, data_stage_2__2009_, data_stage_2__2008_, data_stage_2__2007_, data_stage_2__2006_, data_stage_2__2005_, data_stage_2__2004_, data_stage_2__2003_, data_stage_2__2002_, data_stage_2__2001_, data_stage_2__2000_, data_stage_2__1999_, data_stage_2__1998_, data_stage_2__1997_, data_stage_2__1996_, data_stage_2__1995_, data_stage_2__1994_, data_stage_2__1993_, data_stage_2__1992_, data_stage_2__1991_, data_stage_2__1990_, data_stage_2__1989_, data_stage_2__1988_, data_stage_2__1987_, data_stage_2__1986_, data_stage_2__1985_, data_stage_2__1984_, data_stage_2__1983_, data_stage_2__1982_, data_stage_2__1981_, data_stage_2__1980_, data_stage_2__1979_, data_stage_2__1978_, data_stage_2__1977_, data_stage_2__1976_, data_stage_2__1975_, data_stage_2__1974_, data_stage_2__1973_, data_stage_2__1972_, data_stage_2__1971_, data_stage_2__1970_, data_stage_2__1969_, data_stage_2__1968_, data_stage_2__1967_, data_stage_2__1966_, data_stage_2__1965_, data_stage_2__1964_, data_stage_2__1963_, data_stage_2__1962_, data_stage_2__1961_, data_stage_2__1960_, data_stage_2__1959_, data_stage_2__1958_, data_stage_2__1957_, data_stage_2__1956_, data_stage_2__1955_, data_stage_2__1954_, data_stage_2__1953_, data_stage_2__1952_, data_stage_2__1951_, data_stage_2__1950_, data_stage_2__1949_, data_stage_2__1948_, data_stage_2__1947_, data_stage_2__1946_, data_stage_2__1945_, data_stage_2__1944_, data_stage_2__1943_, data_stage_2__1942_, data_stage_2__1941_, data_stage_2__1940_, data_stage_2__1939_, data_stage_2__1938_, data_stage_2__1937_, data_stage_2__1936_, data_stage_2__1935_, data_stage_2__1934_, data_stage_2__1933_, data_stage_2__1932_, data_stage_2__1931_, data_stage_2__1930_, data_stage_2__1929_, data_stage_2__1928_, data_stage_2__1927_, data_stage_2__1926_, data_stage_2__1925_, data_stage_2__1924_, data_stage_2__1923_, data_stage_2__1922_, data_stage_2__1921_, data_stage_2__1920_, data_stage_2__1919_, data_stage_2__1918_, data_stage_2__1917_, data_stage_2__1916_, data_stage_2__1915_, data_stage_2__1914_, data_stage_2__1913_, data_stage_2__1912_, data_stage_2__1911_, data_stage_2__1910_, data_stage_2__1909_, data_stage_2__1908_, data_stage_2__1907_, data_stage_2__1906_, data_stage_2__1905_, data_stage_2__1904_, data_stage_2__1903_, data_stage_2__1902_, data_stage_2__1901_, data_stage_2__1900_, data_stage_2__1899_, data_stage_2__1898_, data_stage_2__1897_, data_stage_2__1896_, data_stage_2__1895_, data_stage_2__1894_, data_stage_2__1893_, data_stage_2__1892_, data_stage_2__1891_, data_stage_2__1890_, data_stage_2__1889_, data_stage_2__1888_, data_stage_2__1887_, data_stage_2__1886_, data_stage_2__1885_, data_stage_2__1884_, data_stage_2__1883_, data_stage_2__1882_, data_stage_2__1881_, data_stage_2__1880_, data_stage_2__1879_, data_stage_2__1878_, data_stage_2__1877_, data_stage_2__1876_, data_stage_2__1875_, data_stage_2__1874_, data_stage_2__1873_, data_stage_2__1872_, data_stage_2__1871_, data_stage_2__1870_, data_stage_2__1869_, data_stage_2__1868_, data_stage_2__1867_, data_stage_2__1866_, data_stage_2__1865_, data_stage_2__1864_, data_stage_2__1863_, data_stage_2__1862_, data_stage_2__1861_, data_stage_2__1860_, data_stage_2__1859_, data_stage_2__1858_, data_stage_2__1857_, data_stage_2__1856_, data_stage_2__1855_, data_stage_2__1854_, data_stage_2__1853_, data_stage_2__1852_, data_stage_2__1851_, data_stage_2__1850_, data_stage_2__1849_, data_stage_2__1848_, data_stage_2__1847_, data_stage_2__1846_, data_stage_2__1845_, data_stage_2__1844_, data_stage_2__1843_, data_stage_2__1842_, data_stage_2__1841_, data_stage_2__1840_, data_stage_2__1839_, data_stage_2__1838_, data_stage_2__1837_, data_stage_2__1836_, data_stage_2__1835_, data_stage_2__1834_, data_stage_2__1833_, data_stage_2__1832_, data_stage_2__1831_, data_stage_2__1830_, data_stage_2__1829_, data_stage_2__1828_, data_stage_2__1827_, data_stage_2__1826_, data_stage_2__1825_, data_stage_2__1824_, data_stage_2__1823_, data_stage_2__1822_, data_stage_2__1821_, data_stage_2__1820_, data_stage_2__1819_, data_stage_2__1818_, data_stage_2__1817_, data_stage_2__1816_, data_stage_2__1815_, data_stage_2__1814_, data_stage_2__1813_, data_stage_2__1812_, data_stage_2__1811_, data_stage_2__1810_, data_stage_2__1809_, data_stage_2__1808_, data_stage_2__1807_, data_stage_2__1806_, data_stage_2__1805_, data_stage_2__1804_, data_stage_2__1803_, data_stage_2__1802_, data_stage_2__1801_, data_stage_2__1800_, data_stage_2__1799_, data_stage_2__1798_, data_stage_2__1797_, data_stage_2__1796_, data_stage_2__1795_, data_stage_2__1794_, data_stage_2__1793_, data_stage_2__1792_, data_stage_2__1791_, data_stage_2__1790_, data_stage_2__1789_, data_stage_2__1788_, data_stage_2__1787_, data_stage_2__1786_, data_stage_2__1785_, data_stage_2__1784_, data_stage_2__1783_, data_stage_2__1782_, data_stage_2__1781_, data_stage_2__1780_, data_stage_2__1779_, data_stage_2__1778_, data_stage_2__1777_, data_stage_2__1776_, data_stage_2__1775_, data_stage_2__1774_, data_stage_2__1773_, data_stage_2__1772_, data_stage_2__1771_, data_stage_2__1770_, data_stage_2__1769_, data_stage_2__1768_, data_stage_2__1767_, data_stage_2__1766_, data_stage_2__1765_, data_stage_2__1764_, data_stage_2__1763_, data_stage_2__1762_, data_stage_2__1761_, data_stage_2__1760_, data_stage_2__1759_, data_stage_2__1758_, data_stage_2__1757_, data_stage_2__1756_, data_stage_2__1755_, data_stage_2__1754_, data_stage_2__1753_, data_stage_2__1752_, data_stage_2__1751_, data_stage_2__1750_, data_stage_2__1749_, data_stage_2__1748_, data_stage_2__1747_, data_stage_2__1746_, data_stage_2__1745_, data_stage_2__1744_, data_stage_2__1743_, data_stage_2__1742_, data_stage_2__1741_, data_stage_2__1740_, data_stage_2__1739_, data_stage_2__1738_, data_stage_2__1737_, data_stage_2__1736_, data_stage_2__1735_, data_stage_2__1734_, data_stage_2__1733_, data_stage_2__1732_, data_stage_2__1731_, data_stage_2__1730_, data_stage_2__1729_, data_stage_2__1728_, data_stage_2__1727_, data_stage_2__1726_, data_stage_2__1725_, data_stage_2__1724_, data_stage_2__1723_, data_stage_2__1722_, data_stage_2__1721_, data_stage_2__1720_, data_stage_2__1719_, data_stage_2__1718_, data_stage_2__1717_, data_stage_2__1716_, data_stage_2__1715_, data_stage_2__1714_, data_stage_2__1713_, data_stage_2__1712_, data_stage_2__1711_, data_stage_2__1710_, data_stage_2__1709_, data_stage_2__1708_, data_stage_2__1707_, data_stage_2__1706_, data_stage_2__1705_, data_stage_2__1704_, data_stage_2__1703_, data_stage_2__1702_, data_stage_2__1701_, data_stage_2__1700_, data_stage_2__1699_, data_stage_2__1698_, data_stage_2__1697_, data_stage_2__1696_, data_stage_2__1695_, data_stage_2__1694_, data_stage_2__1693_, data_stage_2__1692_, data_stage_2__1691_, data_stage_2__1690_, data_stage_2__1689_, data_stage_2__1688_, data_stage_2__1687_, data_stage_2__1686_, data_stage_2__1685_, data_stage_2__1684_, data_stage_2__1683_, data_stage_2__1682_, data_stage_2__1681_, data_stage_2__1680_, data_stage_2__1679_, data_stage_2__1678_, data_stage_2__1677_, data_stage_2__1676_, data_stage_2__1675_, data_stage_2__1674_, data_stage_2__1673_, data_stage_2__1672_, data_stage_2__1671_, data_stage_2__1670_, data_stage_2__1669_, data_stage_2__1668_, data_stage_2__1667_, data_stage_2__1666_, data_stage_2__1665_, data_stage_2__1664_, data_stage_2__1663_, data_stage_2__1662_, data_stage_2__1661_, data_stage_2__1660_, data_stage_2__1659_, data_stage_2__1658_, data_stage_2__1657_, data_stage_2__1656_, data_stage_2__1655_, data_stage_2__1654_, data_stage_2__1653_, data_stage_2__1652_, data_stage_2__1651_, data_stage_2__1650_, data_stage_2__1649_, data_stage_2__1648_, data_stage_2__1647_, data_stage_2__1646_, data_stage_2__1645_, data_stage_2__1644_, data_stage_2__1643_, data_stage_2__1642_, data_stage_2__1641_, data_stage_2__1640_, data_stage_2__1639_, data_stage_2__1638_, data_stage_2__1637_, data_stage_2__1636_, data_stage_2__1635_, data_stage_2__1634_, data_stage_2__1633_, data_stage_2__1632_, data_stage_2__1631_, data_stage_2__1630_, data_stage_2__1629_, data_stage_2__1628_, data_stage_2__1627_, data_stage_2__1626_, data_stage_2__1625_, data_stage_2__1624_, data_stage_2__1623_, data_stage_2__1622_, data_stage_2__1621_, data_stage_2__1620_, data_stage_2__1619_, data_stage_2__1618_, data_stage_2__1617_, data_stage_2__1616_, data_stage_2__1615_, data_stage_2__1614_, data_stage_2__1613_, data_stage_2__1612_, data_stage_2__1611_, data_stage_2__1610_, data_stage_2__1609_, data_stage_2__1608_, data_stage_2__1607_, data_stage_2__1606_, data_stage_2__1605_, data_stage_2__1604_, data_stage_2__1603_, data_stage_2__1602_, data_stage_2__1601_, data_stage_2__1600_, data_stage_2__1599_, data_stage_2__1598_, data_stage_2__1597_, data_stage_2__1596_, data_stage_2__1595_, data_stage_2__1594_, data_stage_2__1593_, data_stage_2__1592_, data_stage_2__1591_, data_stage_2__1590_, data_stage_2__1589_, data_stage_2__1588_, data_stage_2__1587_, data_stage_2__1586_, data_stage_2__1585_, data_stage_2__1584_, data_stage_2__1583_, data_stage_2__1582_, data_stage_2__1581_, data_stage_2__1580_, data_stage_2__1579_, data_stage_2__1578_, data_stage_2__1577_, data_stage_2__1576_, data_stage_2__1575_, data_stage_2__1574_, data_stage_2__1573_, data_stage_2__1572_, data_stage_2__1571_, data_stage_2__1570_, data_stage_2__1569_, data_stage_2__1568_, data_stage_2__1567_, data_stage_2__1566_, data_stage_2__1565_, data_stage_2__1564_, data_stage_2__1563_, data_stage_2__1562_, data_stage_2__1561_, data_stage_2__1560_, data_stage_2__1559_, data_stage_2__1558_, data_stage_2__1557_, data_stage_2__1556_, data_stage_2__1555_, data_stage_2__1554_, data_stage_2__1553_, data_stage_2__1552_, data_stage_2__1551_, data_stage_2__1550_, data_stage_2__1549_, data_stage_2__1548_, data_stage_2__1547_, data_stage_2__1546_, data_stage_2__1545_, data_stage_2__1544_, data_stage_2__1543_, data_stage_2__1542_, data_stage_2__1541_, data_stage_2__1540_, data_stage_2__1539_, data_stage_2__1538_, data_stage_2__1537_, data_stage_2__1536_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__2047_, data_stage_3__2046_, data_stage_3__2045_, data_stage_3__2044_, data_stage_3__2043_, data_stage_3__2042_, data_stage_3__2041_, data_stage_3__2040_, data_stage_3__2039_, data_stage_3__2038_, data_stage_3__2037_, data_stage_3__2036_, data_stage_3__2035_, data_stage_3__2034_, data_stage_3__2033_, data_stage_3__2032_, data_stage_3__2031_, data_stage_3__2030_, data_stage_3__2029_, data_stage_3__2028_, data_stage_3__2027_, data_stage_3__2026_, data_stage_3__2025_, data_stage_3__2024_, data_stage_3__2023_, data_stage_3__2022_, data_stage_3__2021_, data_stage_3__2020_, data_stage_3__2019_, data_stage_3__2018_, data_stage_3__2017_, data_stage_3__2016_, data_stage_3__2015_, data_stage_3__2014_, data_stage_3__2013_, data_stage_3__2012_, data_stage_3__2011_, data_stage_3__2010_, data_stage_3__2009_, data_stage_3__2008_, data_stage_3__2007_, data_stage_3__2006_, data_stage_3__2005_, data_stage_3__2004_, data_stage_3__2003_, data_stage_3__2002_, data_stage_3__2001_, data_stage_3__2000_, data_stage_3__1999_, data_stage_3__1998_, data_stage_3__1997_, data_stage_3__1996_, data_stage_3__1995_, data_stage_3__1994_, data_stage_3__1993_, data_stage_3__1992_, data_stage_3__1991_, data_stage_3__1990_, data_stage_3__1989_, data_stage_3__1988_, data_stage_3__1987_, data_stage_3__1986_, data_stage_3__1985_, data_stage_3__1984_, data_stage_3__1983_, data_stage_3__1982_, data_stage_3__1981_, data_stage_3__1980_, data_stage_3__1979_, data_stage_3__1978_, data_stage_3__1977_, data_stage_3__1976_, data_stage_3__1975_, data_stage_3__1974_, data_stage_3__1973_, data_stage_3__1972_, data_stage_3__1971_, data_stage_3__1970_, data_stage_3__1969_, data_stage_3__1968_, data_stage_3__1967_, data_stage_3__1966_, data_stage_3__1965_, data_stage_3__1964_, data_stage_3__1963_, data_stage_3__1962_, data_stage_3__1961_, data_stage_3__1960_, data_stage_3__1959_, data_stage_3__1958_, data_stage_3__1957_, data_stage_3__1956_, data_stage_3__1955_, data_stage_3__1954_, data_stage_3__1953_, data_stage_3__1952_, data_stage_3__1951_, data_stage_3__1950_, data_stage_3__1949_, data_stage_3__1948_, data_stage_3__1947_, data_stage_3__1946_, data_stage_3__1945_, data_stage_3__1944_, data_stage_3__1943_, data_stage_3__1942_, data_stage_3__1941_, data_stage_3__1940_, data_stage_3__1939_, data_stage_3__1938_, data_stage_3__1937_, data_stage_3__1936_, data_stage_3__1935_, data_stage_3__1934_, data_stage_3__1933_, data_stage_3__1932_, data_stage_3__1931_, data_stage_3__1930_, data_stage_3__1929_, data_stage_3__1928_, data_stage_3__1927_, data_stage_3__1926_, data_stage_3__1925_, data_stage_3__1924_, data_stage_3__1923_, data_stage_3__1922_, data_stage_3__1921_, data_stage_3__1920_, data_stage_3__1919_, data_stage_3__1918_, data_stage_3__1917_, data_stage_3__1916_, data_stage_3__1915_, data_stage_3__1914_, data_stage_3__1913_, data_stage_3__1912_, data_stage_3__1911_, data_stage_3__1910_, data_stage_3__1909_, data_stage_3__1908_, data_stage_3__1907_, data_stage_3__1906_, data_stage_3__1905_, data_stage_3__1904_, data_stage_3__1903_, data_stage_3__1902_, data_stage_3__1901_, data_stage_3__1900_, data_stage_3__1899_, data_stage_3__1898_, data_stage_3__1897_, data_stage_3__1896_, data_stage_3__1895_, data_stage_3__1894_, data_stage_3__1893_, data_stage_3__1892_, data_stage_3__1891_, data_stage_3__1890_, data_stage_3__1889_, data_stage_3__1888_, data_stage_3__1887_, data_stage_3__1886_, data_stage_3__1885_, data_stage_3__1884_, data_stage_3__1883_, data_stage_3__1882_, data_stage_3__1881_, data_stage_3__1880_, data_stage_3__1879_, data_stage_3__1878_, data_stage_3__1877_, data_stage_3__1876_, data_stage_3__1875_, data_stage_3__1874_, data_stage_3__1873_, data_stage_3__1872_, data_stage_3__1871_, data_stage_3__1870_, data_stage_3__1869_, data_stage_3__1868_, data_stage_3__1867_, data_stage_3__1866_, data_stage_3__1865_, data_stage_3__1864_, data_stage_3__1863_, data_stage_3__1862_, data_stage_3__1861_, data_stage_3__1860_, data_stage_3__1859_, data_stage_3__1858_, data_stage_3__1857_, data_stage_3__1856_, data_stage_3__1855_, data_stage_3__1854_, data_stage_3__1853_, data_stage_3__1852_, data_stage_3__1851_, data_stage_3__1850_, data_stage_3__1849_, data_stage_3__1848_, data_stage_3__1847_, data_stage_3__1846_, data_stage_3__1845_, data_stage_3__1844_, data_stage_3__1843_, data_stage_3__1842_, data_stage_3__1841_, data_stage_3__1840_, data_stage_3__1839_, data_stage_3__1838_, data_stage_3__1837_, data_stage_3__1836_, data_stage_3__1835_, data_stage_3__1834_, data_stage_3__1833_, data_stage_3__1832_, data_stage_3__1831_, data_stage_3__1830_, data_stage_3__1829_, data_stage_3__1828_, data_stage_3__1827_, data_stage_3__1826_, data_stage_3__1825_, data_stage_3__1824_, data_stage_3__1823_, data_stage_3__1822_, data_stage_3__1821_, data_stage_3__1820_, data_stage_3__1819_, data_stage_3__1818_, data_stage_3__1817_, data_stage_3__1816_, data_stage_3__1815_, data_stage_3__1814_, data_stage_3__1813_, data_stage_3__1812_, data_stage_3__1811_, data_stage_3__1810_, data_stage_3__1809_, data_stage_3__1808_, data_stage_3__1807_, data_stage_3__1806_, data_stage_3__1805_, data_stage_3__1804_, data_stage_3__1803_, data_stage_3__1802_, data_stage_3__1801_, data_stage_3__1800_, data_stage_3__1799_, data_stage_3__1798_, data_stage_3__1797_, data_stage_3__1796_, data_stage_3__1795_, data_stage_3__1794_, data_stage_3__1793_, data_stage_3__1792_, data_stage_3__1791_, data_stage_3__1790_, data_stage_3__1789_, data_stage_3__1788_, data_stage_3__1787_, data_stage_3__1786_, data_stage_3__1785_, data_stage_3__1784_, data_stage_3__1783_, data_stage_3__1782_, data_stage_3__1781_, data_stage_3__1780_, data_stage_3__1779_, data_stage_3__1778_, data_stage_3__1777_, data_stage_3__1776_, data_stage_3__1775_, data_stage_3__1774_, data_stage_3__1773_, data_stage_3__1772_, data_stage_3__1771_, data_stage_3__1770_, data_stage_3__1769_, data_stage_3__1768_, data_stage_3__1767_, data_stage_3__1766_, data_stage_3__1765_, data_stage_3__1764_, data_stage_3__1763_, data_stage_3__1762_, data_stage_3__1761_, data_stage_3__1760_, data_stage_3__1759_, data_stage_3__1758_, data_stage_3__1757_, data_stage_3__1756_, data_stage_3__1755_, data_stage_3__1754_, data_stage_3__1753_, data_stage_3__1752_, data_stage_3__1751_, data_stage_3__1750_, data_stage_3__1749_, data_stage_3__1748_, data_stage_3__1747_, data_stage_3__1746_, data_stage_3__1745_, data_stage_3__1744_, data_stage_3__1743_, data_stage_3__1742_, data_stage_3__1741_, data_stage_3__1740_, data_stage_3__1739_, data_stage_3__1738_, data_stage_3__1737_, data_stage_3__1736_, data_stage_3__1735_, data_stage_3__1734_, data_stage_3__1733_, data_stage_3__1732_, data_stage_3__1731_, data_stage_3__1730_, data_stage_3__1729_, data_stage_3__1728_, data_stage_3__1727_, data_stage_3__1726_, data_stage_3__1725_, data_stage_3__1724_, data_stage_3__1723_, data_stage_3__1722_, data_stage_3__1721_, data_stage_3__1720_, data_stage_3__1719_, data_stage_3__1718_, data_stage_3__1717_, data_stage_3__1716_, data_stage_3__1715_, data_stage_3__1714_, data_stage_3__1713_, data_stage_3__1712_, data_stage_3__1711_, data_stage_3__1710_, data_stage_3__1709_, data_stage_3__1708_, data_stage_3__1707_, data_stage_3__1706_, data_stage_3__1705_, data_stage_3__1704_, data_stage_3__1703_, data_stage_3__1702_, data_stage_3__1701_, data_stage_3__1700_, data_stage_3__1699_, data_stage_3__1698_, data_stage_3__1697_, data_stage_3__1696_, data_stage_3__1695_, data_stage_3__1694_, data_stage_3__1693_, data_stage_3__1692_, data_stage_3__1691_, data_stage_3__1690_, data_stage_3__1689_, data_stage_3__1688_, data_stage_3__1687_, data_stage_3__1686_, data_stage_3__1685_, data_stage_3__1684_, data_stage_3__1683_, data_stage_3__1682_, data_stage_3__1681_, data_stage_3__1680_, data_stage_3__1679_, data_stage_3__1678_, data_stage_3__1677_, data_stage_3__1676_, data_stage_3__1675_, data_stage_3__1674_, data_stage_3__1673_, data_stage_3__1672_, data_stage_3__1671_, data_stage_3__1670_, data_stage_3__1669_, data_stage_3__1668_, data_stage_3__1667_, data_stage_3__1666_, data_stage_3__1665_, data_stage_3__1664_, data_stage_3__1663_, data_stage_3__1662_, data_stage_3__1661_, data_stage_3__1660_, data_stage_3__1659_, data_stage_3__1658_, data_stage_3__1657_, data_stage_3__1656_, data_stage_3__1655_, data_stage_3__1654_, data_stage_3__1653_, data_stage_3__1652_, data_stage_3__1651_, data_stage_3__1650_, data_stage_3__1649_, data_stage_3__1648_, data_stage_3__1647_, data_stage_3__1646_, data_stage_3__1645_, data_stage_3__1644_, data_stage_3__1643_, data_stage_3__1642_, data_stage_3__1641_, data_stage_3__1640_, data_stage_3__1639_, data_stage_3__1638_, data_stage_3__1637_, data_stage_3__1636_, data_stage_3__1635_, data_stage_3__1634_, data_stage_3__1633_, data_stage_3__1632_, data_stage_3__1631_, data_stage_3__1630_, data_stage_3__1629_, data_stage_3__1628_, data_stage_3__1627_, data_stage_3__1626_, data_stage_3__1625_, data_stage_3__1624_, data_stage_3__1623_, data_stage_3__1622_, data_stage_3__1621_, data_stage_3__1620_, data_stage_3__1619_, data_stage_3__1618_, data_stage_3__1617_, data_stage_3__1616_, data_stage_3__1615_, data_stage_3__1614_, data_stage_3__1613_, data_stage_3__1612_, data_stage_3__1611_, data_stage_3__1610_, data_stage_3__1609_, data_stage_3__1608_, data_stage_3__1607_, data_stage_3__1606_, data_stage_3__1605_, data_stage_3__1604_, data_stage_3__1603_, data_stage_3__1602_, data_stage_3__1601_, data_stage_3__1600_, data_stage_3__1599_, data_stage_3__1598_, data_stage_3__1597_, data_stage_3__1596_, data_stage_3__1595_, data_stage_3__1594_, data_stage_3__1593_, data_stage_3__1592_, data_stage_3__1591_, data_stage_3__1590_, data_stage_3__1589_, data_stage_3__1588_, data_stage_3__1587_, data_stage_3__1586_, data_stage_3__1585_, data_stage_3__1584_, data_stage_3__1583_, data_stage_3__1582_, data_stage_3__1581_, data_stage_3__1580_, data_stage_3__1579_, data_stage_3__1578_, data_stage_3__1577_, data_stage_3__1576_, data_stage_3__1575_, data_stage_3__1574_, data_stage_3__1573_, data_stage_3__1572_, data_stage_3__1571_, data_stage_3__1570_, data_stage_3__1569_, data_stage_3__1568_, data_stage_3__1567_, data_stage_3__1566_, data_stage_3__1565_, data_stage_3__1564_, data_stage_3__1563_, data_stage_3__1562_, data_stage_3__1561_, data_stage_3__1560_, data_stage_3__1559_, data_stage_3__1558_, data_stage_3__1557_, data_stage_3__1556_, data_stage_3__1555_, data_stage_3__1554_, data_stage_3__1553_, data_stage_3__1552_, data_stage_3__1551_, data_stage_3__1550_, data_stage_3__1549_, data_stage_3__1548_, data_stage_3__1547_, data_stage_3__1546_, data_stage_3__1545_, data_stage_3__1544_, data_stage_3__1543_, data_stage_3__1542_, data_stage_3__1541_, data_stage_3__1540_, data_stage_3__1539_, data_stage_3__1538_, data_stage_3__1537_, data_stage_3__1536_ })
  );


  bsg_swap_width_p256
  mux_stage_2__mux_swap_4__swap_inst
  (
    .data_i({ data_stage_2__2559_, data_stage_2__2558_, data_stage_2__2557_, data_stage_2__2556_, data_stage_2__2555_, data_stage_2__2554_, data_stage_2__2553_, data_stage_2__2552_, data_stage_2__2551_, data_stage_2__2550_, data_stage_2__2549_, data_stage_2__2548_, data_stage_2__2547_, data_stage_2__2546_, data_stage_2__2545_, data_stage_2__2544_, data_stage_2__2543_, data_stage_2__2542_, data_stage_2__2541_, data_stage_2__2540_, data_stage_2__2539_, data_stage_2__2538_, data_stage_2__2537_, data_stage_2__2536_, data_stage_2__2535_, data_stage_2__2534_, data_stage_2__2533_, data_stage_2__2532_, data_stage_2__2531_, data_stage_2__2530_, data_stage_2__2529_, data_stage_2__2528_, data_stage_2__2527_, data_stage_2__2526_, data_stage_2__2525_, data_stage_2__2524_, data_stage_2__2523_, data_stage_2__2522_, data_stage_2__2521_, data_stage_2__2520_, data_stage_2__2519_, data_stage_2__2518_, data_stage_2__2517_, data_stage_2__2516_, data_stage_2__2515_, data_stage_2__2514_, data_stage_2__2513_, data_stage_2__2512_, data_stage_2__2511_, data_stage_2__2510_, data_stage_2__2509_, data_stage_2__2508_, data_stage_2__2507_, data_stage_2__2506_, data_stage_2__2505_, data_stage_2__2504_, data_stage_2__2503_, data_stage_2__2502_, data_stage_2__2501_, data_stage_2__2500_, data_stage_2__2499_, data_stage_2__2498_, data_stage_2__2497_, data_stage_2__2496_, data_stage_2__2495_, data_stage_2__2494_, data_stage_2__2493_, data_stage_2__2492_, data_stage_2__2491_, data_stage_2__2490_, data_stage_2__2489_, data_stage_2__2488_, data_stage_2__2487_, data_stage_2__2486_, data_stage_2__2485_, data_stage_2__2484_, data_stage_2__2483_, data_stage_2__2482_, data_stage_2__2481_, data_stage_2__2480_, data_stage_2__2479_, data_stage_2__2478_, data_stage_2__2477_, data_stage_2__2476_, data_stage_2__2475_, data_stage_2__2474_, data_stage_2__2473_, data_stage_2__2472_, data_stage_2__2471_, data_stage_2__2470_, data_stage_2__2469_, data_stage_2__2468_, data_stage_2__2467_, data_stage_2__2466_, data_stage_2__2465_, data_stage_2__2464_, data_stage_2__2463_, data_stage_2__2462_, data_stage_2__2461_, data_stage_2__2460_, data_stage_2__2459_, data_stage_2__2458_, data_stage_2__2457_, data_stage_2__2456_, data_stage_2__2455_, data_stage_2__2454_, data_stage_2__2453_, data_stage_2__2452_, data_stage_2__2451_, data_stage_2__2450_, data_stage_2__2449_, data_stage_2__2448_, data_stage_2__2447_, data_stage_2__2446_, data_stage_2__2445_, data_stage_2__2444_, data_stage_2__2443_, data_stage_2__2442_, data_stage_2__2441_, data_stage_2__2440_, data_stage_2__2439_, data_stage_2__2438_, data_stage_2__2437_, data_stage_2__2436_, data_stage_2__2435_, data_stage_2__2434_, data_stage_2__2433_, data_stage_2__2432_, data_stage_2__2431_, data_stage_2__2430_, data_stage_2__2429_, data_stage_2__2428_, data_stage_2__2427_, data_stage_2__2426_, data_stage_2__2425_, data_stage_2__2424_, data_stage_2__2423_, data_stage_2__2422_, data_stage_2__2421_, data_stage_2__2420_, data_stage_2__2419_, data_stage_2__2418_, data_stage_2__2417_, data_stage_2__2416_, data_stage_2__2415_, data_stage_2__2414_, data_stage_2__2413_, data_stage_2__2412_, data_stage_2__2411_, data_stage_2__2410_, data_stage_2__2409_, data_stage_2__2408_, data_stage_2__2407_, data_stage_2__2406_, data_stage_2__2405_, data_stage_2__2404_, data_stage_2__2403_, data_stage_2__2402_, data_stage_2__2401_, data_stage_2__2400_, data_stage_2__2399_, data_stage_2__2398_, data_stage_2__2397_, data_stage_2__2396_, data_stage_2__2395_, data_stage_2__2394_, data_stage_2__2393_, data_stage_2__2392_, data_stage_2__2391_, data_stage_2__2390_, data_stage_2__2389_, data_stage_2__2388_, data_stage_2__2387_, data_stage_2__2386_, data_stage_2__2385_, data_stage_2__2384_, data_stage_2__2383_, data_stage_2__2382_, data_stage_2__2381_, data_stage_2__2380_, data_stage_2__2379_, data_stage_2__2378_, data_stage_2__2377_, data_stage_2__2376_, data_stage_2__2375_, data_stage_2__2374_, data_stage_2__2373_, data_stage_2__2372_, data_stage_2__2371_, data_stage_2__2370_, data_stage_2__2369_, data_stage_2__2368_, data_stage_2__2367_, data_stage_2__2366_, data_stage_2__2365_, data_stage_2__2364_, data_stage_2__2363_, data_stage_2__2362_, data_stage_2__2361_, data_stage_2__2360_, data_stage_2__2359_, data_stage_2__2358_, data_stage_2__2357_, data_stage_2__2356_, data_stage_2__2355_, data_stage_2__2354_, data_stage_2__2353_, data_stage_2__2352_, data_stage_2__2351_, data_stage_2__2350_, data_stage_2__2349_, data_stage_2__2348_, data_stage_2__2347_, data_stage_2__2346_, data_stage_2__2345_, data_stage_2__2344_, data_stage_2__2343_, data_stage_2__2342_, data_stage_2__2341_, data_stage_2__2340_, data_stage_2__2339_, data_stage_2__2338_, data_stage_2__2337_, data_stage_2__2336_, data_stage_2__2335_, data_stage_2__2334_, data_stage_2__2333_, data_stage_2__2332_, data_stage_2__2331_, data_stage_2__2330_, data_stage_2__2329_, data_stage_2__2328_, data_stage_2__2327_, data_stage_2__2326_, data_stage_2__2325_, data_stage_2__2324_, data_stage_2__2323_, data_stage_2__2322_, data_stage_2__2321_, data_stage_2__2320_, data_stage_2__2319_, data_stage_2__2318_, data_stage_2__2317_, data_stage_2__2316_, data_stage_2__2315_, data_stage_2__2314_, data_stage_2__2313_, data_stage_2__2312_, data_stage_2__2311_, data_stage_2__2310_, data_stage_2__2309_, data_stage_2__2308_, data_stage_2__2307_, data_stage_2__2306_, data_stage_2__2305_, data_stage_2__2304_, data_stage_2__2303_, data_stage_2__2302_, data_stage_2__2301_, data_stage_2__2300_, data_stage_2__2299_, data_stage_2__2298_, data_stage_2__2297_, data_stage_2__2296_, data_stage_2__2295_, data_stage_2__2294_, data_stage_2__2293_, data_stage_2__2292_, data_stage_2__2291_, data_stage_2__2290_, data_stage_2__2289_, data_stage_2__2288_, data_stage_2__2287_, data_stage_2__2286_, data_stage_2__2285_, data_stage_2__2284_, data_stage_2__2283_, data_stage_2__2282_, data_stage_2__2281_, data_stage_2__2280_, data_stage_2__2279_, data_stage_2__2278_, data_stage_2__2277_, data_stage_2__2276_, data_stage_2__2275_, data_stage_2__2274_, data_stage_2__2273_, data_stage_2__2272_, data_stage_2__2271_, data_stage_2__2270_, data_stage_2__2269_, data_stage_2__2268_, data_stage_2__2267_, data_stage_2__2266_, data_stage_2__2265_, data_stage_2__2264_, data_stage_2__2263_, data_stage_2__2262_, data_stage_2__2261_, data_stage_2__2260_, data_stage_2__2259_, data_stage_2__2258_, data_stage_2__2257_, data_stage_2__2256_, data_stage_2__2255_, data_stage_2__2254_, data_stage_2__2253_, data_stage_2__2252_, data_stage_2__2251_, data_stage_2__2250_, data_stage_2__2249_, data_stage_2__2248_, data_stage_2__2247_, data_stage_2__2246_, data_stage_2__2245_, data_stage_2__2244_, data_stage_2__2243_, data_stage_2__2242_, data_stage_2__2241_, data_stage_2__2240_, data_stage_2__2239_, data_stage_2__2238_, data_stage_2__2237_, data_stage_2__2236_, data_stage_2__2235_, data_stage_2__2234_, data_stage_2__2233_, data_stage_2__2232_, data_stage_2__2231_, data_stage_2__2230_, data_stage_2__2229_, data_stage_2__2228_, data_stage_2__2227_, data_stage_2__2226_, data_stage_2__2225_, data_stage_2__2224_, data_stage_2__2223_, data_stage_2__2222_, data_stage_2__2221_, data_stage_2__2220_, data_stage_2__2219_, data_stage_2__2218_, data_stage_2__2217_, data_stage_2__2216_, data_stage_2__2215_, data_stage_2__2214_, data_stage_2__2213_, data_stage_2__2212_, data_stage_2__2211_, data_stage_2__2210_, data_stage_2__2209_, data_stage_2__2208_, data_stage_2__2207_, data_stage_2__2206_, data_stage_2__2205_, data_stage_2__2204_, data_stage_2__2203_, data_stage_2__2202_, data_stage_2__2201_, data_stage_2__2200_, data_stage_2__2199_, data_stage_2__2198_, data_stage_2__2197_, data_stage_2__2196_, data_stage_2__2195_, data_stage_2__2194_, data_stage_2__2193_, data_stage_2__2192_, data_stage_2__2191_, data_stage_2__2190_, data_stage_2__2189_, data_stage_2__2188_, data_stage_2__2187_, data_stage_2__2186_, data_stage_2__2185_, data_stage_2__2184_, data_stage_2__2183_, data_stage_2__2182_, data_stage_2__2181_, data_stage_2__2180_, data_stage_2__2179_, data_stage_2__2178_, data_stage_2__2177_, data_stage_2__2176_, data_stage_2__2175_, data_stage_2__2174_, data_stage_2__2173_, data_stage_2__2172_, data_stage_2__2171_, data_stage_2__2170_, data_stage_2__2169_, data_stage_2__2168_, data_stage_2__2167_, data_stage_2__2166_, data_stage_2__2165_, data_stage_2__2164_, data_stage_2__2163_, data_stage_2__2162_, data_stage_2__2161_, data_stage_2__2160_, data_stage_2__2159_, data_stage_2__2158_, data_stage_2__2157_, data_stage_2__2156_, data_stage_2__2155_, data_stage_2__2154_, data_stage_2__2153_, data_stage_2__2152_, data_stage_2__2151_, data_stage_2__2150_, data_stage_2__2149_, data_stage_2__2148_, data_stage_2__2147_, data_stage_2__2146_, data_stage_2__2145_, data_stage_2__2144_, data_stage_2__2143_, data_stage_2__2142_, data_stage_2__2141_, data_stage_2__2140_, data_stage_2__2139_, data_stage_2__2138_, data_stage_2__2137_, data_stage_2__2136_, data_stage_2__2135_, data_stage_2__2134_, data_stage_2__2133_, data_stage_2__2132_, data_stage_2__2131_, data_stage_2__2130_, data_stage_2__2129_, data_stage_2__2128_, data_stage_2__2127_, data_stage_2__2126_, data_stage_2__2125_, data_stage_2__2124_, data_stage_2__2123_, data_stage_2__2122_, data_stage_2__2121_, data_stage_2__2120_, data_stage_2__2119_, data_stage_2__2118_, data_stage_2__2117_, data_stage_2__2116_, data_stage_2__2115_, data_stage_2__2114_, data_stage_2__2113_, data_stage_2__2112_, data_stage_2__2111_, data_stage_2__2110_, data_stage_2__2109_, data_stage_2__2108_, data_stage_2__2107_, data_stage_2__2106_, data_stage_2__2105_, data_stage_2__2104_, data_stage_2__2103_, data_stage_2__2102_, data_stage_2__2101_, data_stage_2__2100_, data_stage_2__2099_, data_stage_2__2098_, data_stage_2__2097_, data_stage_2__2096_, data_stage_2__2095_, data_stage_2__2094_, data_stage_2__2093_, data_stage_2__2092_, data_stage_2__2091_, data_stage_2__2090_, data_stage_2__2089_, data_stage_2__2088_, data_stage_2__2087_, data_stage_2__2086_, data_stage_2__2085_, data_stage_2__2084_, data_stage_2__2083_, data_stage_2__2082_, data_stage_2__2081_, data_stage_2__2080_, data_stage_2__2079_, data_stage_2__2078_, data_stage_2__2077_, data_stage_2__2076_, data_stage_2__2075_, data_stage_2__2074_, data_stage_2__2073_, data_stage_2__2072_, data_stage_2__2071_, data_stage_2__2070_, data_stage_2__2069_, data_stage_2__2068_, data_stage_2__2067_, data_stage_2__2066_, data_stage_2__2065_, data_stage_2__2064_, data_stage_2__2063_, data_stage_2__2062_, data_stage_2__2061_, data_stage_2__2060_, data_stage_2__2059_, data_stage_2__2058_, data_stage_2__2057_, data_stage_2__2056_, data_stage_2__2055_, data_stage_2__2054_, data_stage_2__2053_, data_stage_2__2052_, data_stage_2__2051_, data_stage_2__2050_, data_stage_2__2049_, data_stage_2__2048_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__2559_, data_stage_3__2558_, data_stage_3__2557_, data_stage_3__2556_, data_stage_3__2555_, data_stage_3__2554_, data_stage_3__2553_, data_stage_3__2552_, data_stage_3__2551_, data_stage_3__2550_, data_stage_3__2549_, data_stage_3__2548_, data_stage_3__2547_, data_stage_3__2546_, data_stage_3__2545_, data_stage_3__2544_, data_stage_3__2543_, data_stage_3__2542_, data_stage_3__2541_, data_stage_3__2540_, data_stage_3__2539_, data_stage_3__2538_, data_stage_3__2537_, data_stage_3__2536_, data_stage_3__2535_, data_stage_3__2534_, data_stage_3__2533_, data_stage_3__2532_, data_stage_3__2531_, data_stage_3__2530_, data_stage_3__2529_, data_stage_3__2528_, data_stage_3__2527_, data_stage_3__2526_, data_stage_3__2525_, data_stage_3__2524_, data_stage_3__2523_, data_stage_3__2522_, data_stage_3__2521_, data_stage_3__2520_, data_stage_3__2519_, data_stage_3__2518_, data_stage_3__2517_, data_stage_3__2516_, data_stage_3__2515_, data_stage_3__2514_, data_stage_3__2513_, data_stage_3__2512_, data_stage_3__2511_, data_stage_3__2510_, data_stage_3__2509_, data_stage_3__2508_, data_stage_3__2507_, data_stage_3__2506_, data_stage_3__2505_, data_stage_3__2504_, data_stage_3__2503_, data_stage_3__2502_, data_stage_3__2501_, data_stage_3__2500_, data_stage_3__2499_, data_stage_3__2498_, data_stage_3__2497_, data_stage_3__2496_, data_stage_3__2495_, data_stage_3__2494_, data_stage_3__2493_, data_stage_3__2492_, data_stage_3__2491_, data_stage_3__2490_, data_stage_3__2489_, data_stage_3__2488_, data_stage_3__2487_, data_stage_3__2486_, data_stage_3__2485_, data_stage_3__2484_, data_stage_3__2483_, data_stage_3__2482_, data_stage_3__2481_, data_stage_3__2480_, data_stage_3__2479_, data_stage_3__2478_, data_stage_3__2477_, data_stage_3__2476_, data_stage_3__2475_, data_stage_3__2474_, data_stage_3__2473_, data_stage_3__2472_, data_stage_3__2471_, data_stage_3__2470_, data_stage_3__2469_, data_stage_3__2468_, data_stage_3__2467_, data_stage_3__2466_, data_stage_3__2465_, data_stage_3__2464_, data_stage_3__2463_, data_stage_3__2462_, data_stage_3__2461_, data_stage_3__2460_, data_stage_3__2459_, data_stage_3__2458_, data_stage_3__2457_, data_stage_3__2456_, data_stage_3__2455_, data_stage_3__2454_, data_stage_3__2453_, data_stage_3__2452_, data_stage_3__2451_, data_stage_3__2450_, data_stage_3__2449_, data_stage_3__2448_, data_stage_3__2447_, data_stage_3__2446_, data_stage_3__2445_, data_stage_3__2444_, data_stage_3__2443_, data_stage_3__2442_, data_stage_3__2441_, data_stage_3__2440_, data_stage_3__2439_, data_stage_3__2438_, data_stage_3__2437_, data_stage_3__2436_, data_stage_3__2435_, data_stage_3__2434_, data_stage_3__2433_, data_stage_3__2432_, data_stage_3__2431_, data_stage_3__2430_, data_stage_3__2429_, data_stage_3__2428_, data_stage_3__2427_, data_stage_3__2426_, data_stage_3__2425_, data_stage_3__2424_, data_stage_3__2423_, data_stage_3__2422_, data_stage_3__2421_, data_stage_3__2420_, data_stage_3__2419_, data_stage_3__2418_, data_stage_3__2417_, data_stage_3__2416_, data_stage_3__2415_, data_stage_3__2414_, data_stage_3__2413_, data_stage_3__2412_, data_stage_3__2411_, data_stage_3__2410_, data_stage_3__2409_, data_stage_3__2408_, data_stage_3__2407_, data_stage_3__2406_, data_stage_3__2405_, data_stage_3__2404_, data_stage_3__2403_, data_stage_3__2402_, data_stage_3__2401_, data_stage_3__2400_, data_stage_3__2399_, data_stage_3__2398_, data_stage_3__2397_, data_stage_3__2396_, data_stage_3__2395_, data_stage_3__2394_, data_stage_3__2393_, data_stage_3__2392_, data_stage_3__2391_, data_stage_3__2390_, data_stage_3__2389_, data_stage_3__2388_, data_stage_3__2387_, data_stage_3__2386_, data_stage_3__2385_, data_stage_3__2384_, data_stage_3__2383_, data_stage_3__2382_, data_stage_3__2381_, data_stage_3__2380_, data_stage_3__2379_, data_stage_3__2378_, data_stage_3__2377_, data_stage_3__2376_, data_stage_3__2375_, data_stage_3__2374_, data_stage_3__2373_, data_stage_3__2372_, data_stage_3__2371_, data_stage_3__2370_, data_stage_3__2369_, data_stage_3__2368_, data_stage_3__2367_, data_stage_3__2366_, data_stage_3__2365_, data_stage_3__2364_, data_stage_3__2363_, data_stage_3__2362_, data_stage_3__2361_, data_stage_3__2360_, data_stage_3__2359_, data_stage_3__2358_, data_stage_3__2357_, data_stage_3__2356_, data_stage_3__2355_, data_stage_3__2354_, data_stage_3__2353_, data_stage_3__2352_, data_stage_3__2351_, data_stage_3__2350_, data_stage_3__2349_, data_stage_3__2348_, data_stage_3__2347_, data_stage_3__2346_, data_stage_3__2345_, data_stage_3__2344_, data_stage_3__2343_, data_stage_3__2342_, data_stage_3__2341_, data_stage_3__2340_, data_stage_3__2339_, data_stage_3__2338_, data_stage_3__2337_, data_stage_3__2336_, data_stage_3__2335_, data_stage_3__2334_, data_stage_3__2333_, data_stage_3__2332_, data_stage_3__2331_, data_stage_3__2330_, data_stage_3__2329_, data_stage_3__2328_, data_stage_3__2327_, data_stage_3__2326_, data_stage_3__2325_, data_stage_3__2324_, data_stage_3__2323_, data_stage_3__2322_, data_stage_3__2321_, data_stage_3__2320_, data_stage_3__2319_, data_stage_3__2318_, data_stage_3__2317_, data_stage_3__2316_, data_stage_3__2315_, data_stage_3__2314_, data_stage_3__2313_, data_stage_3__2312_, data_stage_3__2311_, data_stage_3__2310_, data_stage_3__2309_, data_stage_3__2308_, data_stage_3__2307_, data_stage_3__2306_, data_stage_3__2305_, data_stage_3__2304_, data_stage_3__2303_, data_stage_3__2302_, data_stage_3__2301_, data_stage_3__2300_, data_stage_3__2299_, data_stage_3__2298_, data_stage_3__2297_, data_stage_3__2296_, data_stage_3__2295_, data_stage_3__2294_, data_stage_3__2293_, data_stage_3__2292_, data_stage_3__2291_, data_stage_3__2290_, data_stage_3__2289_, data_stage_3__2288_, data_stage_3__2287_, data_stage_3__2286_, data_stage_3__2285_, data_stage_3__2284_, data_stage_3__2283_, data_stage_3__2282_, data_stage_3__2281_, data_stage_3__2280_, data_stage_3__2279_, data_stage_3__2278_, data_stage_3__2277_, data_stage_3__2276_, data_stage_3__2275_, data_stage_3__2274_, data_stage_3__2273_, data_stage_3__2272_, data_stage_3__2271_, data_stage_3__2270_, data_stage_3__2269_, data_stage_3__2268_, data_stage_3__2267_, data_stage_3__2266_, data_stage_3__2265_, data_stage_3__2264_, data_stage_3__2263_, data_stage_3__2262_, data_stage_3__2261_, data_stage_3__2260_, data_stage_3__2259_, data_stage_3__2258_, data_stage_3__2257_, data_stage_3__2256_, data_stage_3__2255_, data_stage_3__2254_, data_stage_3__2253_, data_stage_3__2252_, data_stage_3__2251_, data_stage_3__2250_, data_stage_3__2249_, data_stage_3__2248_, data_stage_3__2247_, data_stage_3__2246_, data_stage_3__2245_, data_stage_3__2244_, data_stage_3__2243_, data_stage_3__2242_, data_stage_3__2241_, data_stage_3__2240_, data_stage_3__2239_, data_stage_3__2238_, data_stage_3__2237_, data_stage_3__2236_, data_stage_3__2235_, data_stage_3__2234_, data_stage_3__2233_, data_stage_3__2232_, data_stage_3__2231_, data_stage_3__2230_, data_stage_3__2229_, data_stage_3__2228_, data_stage_3__2227_, data_stage_3__2226_, data_stage_3__2225_, data_stage_3__2224_, data_stage_3__2223_, data_stage_3__2222_, data_stage_3__2221_, data_stage_3__2220_, data_stage_3__2219_, data_stage_3__2218_, data_stage_3__2217_, data_stage_3__2216_, data_stage_3__2215_, data_stage_3__2214_, data_stage_3__2213_, data_stage_3__2212_, data_stage_3__2211_, data_stage_3__2210_, data_stage_3__2209_, data_stage_3__2208_, data_stage_3__2207_, data_stage_3__2206_, data_stage_3__2205_, data_stage_3__2204_, data_stage_3__2203_, data_stage_3__2202_, data_stage_3__2201_, data_stage_3__2200_, data_stage_3__2199_, data_stage_3__2198_, data_stage_3__2197_, data_stage_3__2196_, data_stage_3__2195_, data_stage_3__2194_, data_stage_3__2193_, data_stage_3__2192_, data_stage_3__2191_, data_stage_3__2190_, data_stage_3__2189_, data_stage_3__2188_, data_stage_3__2187_, data_stage_3__2186_, data_stage_3__2185_, data_stage_3__2184_, data_stage_3__2183_, data_stage_3__2182_, data_stage_3__2181_, data_stage_3__2180_, data_stage_3__2179_, data_stage_3__2178_, data_stage_3__2177_, data_stage_3__2176_, data_stage_3__2175_, data_stage_3__2174_, data_stage_3__2173_, data_stage_3__2172_, data_stage_3__2171_, data_stage_3__2170_, data_stage_3__2169_, data_stage_3__2168_, data_stage_3__2167_, data_stage_3__2166_, data_stage_3__2165_, data_stage_3__2164_, data_stage_3__2163_, data_stage_3__2162_, data_stage_3__2161_, data_stage_3__2160_, data_stage_3__2159_, data_stage_3__2158_, data_stage_3__2157_, data_stage_3__2156_, data_stage_3__2155_, data_stage_3__2154_, data_stage_3__2153_, data_stage_3__2152_, data_stage_3__2151_, data_stage_3__2150_, data_stage_3__2149_, data_stage_3__2148_, data_stage_3__2147_, data_stage_3__2146_, data_stage_3__2145_, data_stage_3__2144_, data_stage_3__2143_, data_stage_3__2142_, data_stage_3__2141_, data_stage_3__2140_, data_stage_3__2139_, data_stage_3__2138_, data_stage_3__2137_, data_stage_3__2136_, data_stage_3__2135_, data_stage_3__2134_, data_stage_3__2133_, data_stage_3__2132_, data_stage_3__2131_, data_stage_3__2130_, data_stage_3__2129_, data_stage_3__2128_, data_stage_3__2127_, data_stage_3__2126_, data_stage_3__2125_, data_stage_3__2124_, data_stage_3__2123_, data_stage_3__2122_, data_stage_3__2121_, data_stage_3__2120_, data_stage_3__2119_, data_stage_3__2118_, data_stage_3__2117_, data_stage_3__2116_, data_stage_3__2115_, data_stage_3__2114_, data_stage_3__2113_, data_stage_3__2112_, data_stage_3__2111_, data_stage_3__2110_, data_stage_3__2109_, data_stage_3__2108_, data_stage_3__2107_, data_stage_3__2106_, data_stage_3__2105_, data_stage_3__2104_, data_stage_3__2103_, data_stage_3__2102_, data_stage_3__2101_, data_stage_3__2100_, data_stage_3__2099_, data_stage_3__2098_, data_stage_3__2097_, data_stage_3__2096_, data_stage_3__2095_, data_stage_3__2094_, data_stage_3__2093_, data_stage_3__2092_, data_stage_3__2091_, data_stage_3__2090_, data_stage_3__2089_, data_stage_3__2088_, data_stage_3__2087_, data_stage_3__2086_, data_stage_3__2085_, data_stage_3__2084_, data_stage_3__2083_, data_stage_3__2082_, data_stage_3__2081_, data_stage_3__2080_, data_stage_3__2079_, data_stage_3__2078_, data_stage_3__2077_, data_stage_3__2076_, data_stage_3__2075_, data_stage_3__2074_, data_stage_3__2073_, data_stage_3__2072_, data_stage_3__2071_, data_stage_3__2070_, data_stage_3__2069_, data_stage_3__2068_, data_stage_3__2067_, data_stage_3__2066_, data_stage_3__2065_, data_stage_3__2064_, data_stage_3__2063_, data_stage_3__2062_, data_stage_3__2061_, data_stage_3__2060_, data_stage_3__2059_, data_stage_3__2058_, data_stage_3__2057_, data_stage_3__2056_, data_stage_3__2055_, data_stage_3__2054_, data_stage_3__2053_, data_stage_3__2052_, data_stage_3__2051_, data_stage_3__2050_, data_stage_3__2049_, data_stage_3__2048_ })
  );


  bsg_swap_width_p256
  mux_stage_2__mux_swap_5__swap_inst
  (
    .data_i({ data_stage_2__3071_, data_stage_2__3070_, data_stage_2__3069_, data_stage_2__3068_, data_stage_2__3067_, data_stage_2__3066_, data_stage_2__3065_, data_stage_2__3064_, data_stage_2__3063_, data_stage_2__3062_, data_stage_2__3061_, data_stage_2__3060_, data_stage_2__3059_, data_stage_2__3058_, data_stage_2__3057_, data_stage_2__3056_, data_stage_2__3055_, data_stage_2__3054_, data_stage_2__3053_, data_stage_2__3052_, data_stage_2__3051_, data_stage_2__3050_, data_stage_2__3049_, data_stage_2__3048_, data_stage_2__3047_, data_stage_2__3046_, data_stage_2__3045_, data_stage_2__3044_, data_stage_2__3043_, data_stage_2__3042_, data_stage_2__3041_, data_stage_2__3040_, data_stage_2__3039_, data_stage_2__3038_, data_stage_2__3037_, data_stage_2__3036_, data_stage_2__3035_, data_stage_2__3034_, data_stage_2__3033_, data_stage_2__3032_, data_stage_2__3031_, data_stage_2__3030_, data_stage_2__3029_, data_stage_2__3028_, data_stage_2__3027_, data_stage_2__3026_, data_stage_2__3025_, data_stage_2__3024_, data_stage_2__3023_, data_stage_2__3022_, data_stage_2__3021_, data_stage_2__3020_, data_stage_2__3019_, data_stage_2__3018_, data_stage_2__3017_, data_stage_2__3016_, data_stage_2__3015_, data_stage_2__3014_, data_stage_2__3013_, data_stage_2__3012_, data_stage_2__3011_, data_stage_2__3010_, data_stage_2__3009_, data_stage_2__3008_, data_stage_2__3007_, data_stage_2__3006_, data_stage_2__3005_, data_stage_2__3004_, data_stage_2__3003_, data_stage_2__3002_, data_stage_2__3001_, data_stage_2__3000_, data_stage_2__2999_, data_stage_2__2998_, data_stage_2__2997_, data_stage_2__2996_, data_stage_2__2995_, data_stage_2__2994_, data_stage_2__2993_, data_stage_2__2992_, data_stage_2__2991_, data_stage_2__2990_, data_stage_2__2989_, data_stage_2__2988_, data_stage_2__2987_, data_stage_2__2986_, data_stage_2__2985_, data_stage_2__2984_, data_stage_2__2983_, data_stage_2__2982_, data_stage_2__2981_, data_stage_2__2980_, data_stage_2__2979_, data_stage_2__2978_, data_stage_2__2977_, data_stage_2__2976_, data_stage_2__2975_, data_stage_2__2974_, data_stage_2__2973_, data_stage_2__2972_, data_stage_2__2971_, data_stage_2__2970_, data_stage_2__2969_, data_stage_2__2968_, data_stage_2__2967_, data_stage_2__2966_, data_stage_2__2965_, data_stage_2__2964_, data_stage_2__2963_, data_stage_2__2962_, data_stage_2__2961_, data_stage_2__2960_, data_stage_2__2959_, data_stage_2__2958_, data_stage_2__2957_, data_stage_2__2956_, data_stage_2__2955_, data_stage_2__2954_, data_stage_2__2953_, data_stage_2__2952_, data_stage_2__2951_, data_stage_2__2950_, data_stage_2__2949_, data_stage_2__2948_, data_stage_2__2947_, data_stage_2__2946_, data_stage_2__2945_, data_stage_2__2944_, data_stage_2__2943_, data_stage_2__2942_, data_stage_2__2941_, data_stage_2__2940_, data_stage_2__2939_, data_stage_2__2938_, data_stage_2__2937_, data_stage_2__2936_, data_stage_2__2935_, data_stage_2__2934_, data_stage_2__2933_, data_stage_2__2932_, data_stage_2__2931_, data_stage_2__2930_, data_stage_2__2929_, data_stage_2__2928_, data_stage_2__2927_, data_stage_2__2926_, data_stage_2__2925_, data_stage_2__2924_, data_stage_2__2923_, data_stage_2__2922_, data_stage_2__2921_, data_stage_2__2920_, data_stage_2__2919_, data_stage_2__2918_, data_stage_2__2917_, data_stage_2__2916_, data_stage_2__2915_, data_stage_2__2914_, data_stage_2__2913_, data_stage_2__2912_, data_stage_2__2911_, data_stage_2__2910_, data_stage_2__2909_, data_stage_2__2908_, data_stage_2__2907_, data_stage_2__2906_, data_stage_2__2905_, data_stage_2__2904_, data_stage_2__2903_, data_stage_2__2902_, data_stage_2__2901_, data_stage_2__2900_, data_stage_2__2899_, data_stage_2__2898_, data_stage_2__2897_, data_stage_2__2896_, data_stage_2__2895_, data_stage_2__2894_, data_stage_2__2893_, data_stage_2__2892_, data_stage_2__2891_, data_stage_2__2890_, data_stage_2__2889_, data_stage_2__2888_, data_stage_2__2887_, data_stage_2__2886_, data_stage_2__2885_, data_stage_2__2884_, data_stage_2__2883_, data_stage_2__2882_, data_stage_2__2881_, data_stage_2__2880_, data_stage_2__2879_, data_stage_2__2878_, data_stage_2__2877_, data_stage_2__2876_, data_stage_2__2875_, data_stage_2__2874_, data_stage_2__2873_, data_stage_2__2872_, data_stage_2__2871_, data_stage_2__2870_, data_stage_2__2869_, data_stage_2__2868_, data_stage_2__2867_, data_stage_2__2866_, data_stage_2__2865_, data_stage_2__2864_, data_stage_2__2863_, data_stage_2__2862_, data_stage_2__2861_, data_stage_2__2860_, data_stage_2__2859_, data_stage_2__2858_, data_stage_2__2857_, data_stage_2__2856_, data_stage_2__2855_, data_stage_2__2854_, data_stage_2__2853_, data_stage_2__2852_, data_stage_2__2851_, data_stage_2__2850_, data_stage_2__2849_, data_stage_2__2848_, data_stage_2__2847_, data_stage_2__2846_, data_stage_2__2845_, data_stage_2__2844_, data_stage_2__2843_, data_stage_2__2842_, data_stage_2__2841_, data_stage_2__2840_, data_stage_2__2839_, data_stage_2__2838_, data_stage_2__2837_, data_stage_2__2836_, data_stage_2__2835_, data_stage_2__2834_, data_stage_2__2833_, data_stage_2__2832_, data_stage_2__2831_, data_stage_2__2830_, data_stage_2__2829_, data_stage_2__2828_, data_stage_2__2827_, data_stage_2__2826_, data_stage_2__2825_, data_stage_2__2824_, data_stage_2__2823_, data_stage_2__2822_, data_stage_2__2821_, data_stage_2__2820_, data_stage_2__2819_, data_stage_2__2818_, data_stage_2__2817_, data_stage_2__2816_, data_stage_2__2815_, data_stage_2__2814_, data_stage_2__2813_, data_stage_2__2812_, data_stage_2__2811_, data_stage_2__2810_, data_stage_2__2809_, data_stage_2__2808_, data_stage_2__2807_, data_stage_2__2806_, data_stage_2__2805_, data_stage_2__2804_, data_stage_2__2803_, data_stage_2__2802_, data_stage_2__2801_, data_stage_2__2800_, data_stage_2__2799_, data_stage_2__2798_, data_stage_2__2797_, data_stage_2__2796_, data_stage_2__2795_, data_stage_2__2794_, data_stage_2__2793_, data_stage_2__2792_, data_stage_2__2791_, data_stage_2__2790_, data_stage_2__2789_, data_stage_2__2788_, data_stage_2__2787_, data_stage_2__2786_, data_stage_2__2785_, data_stage_2__2784_, data_stage_2__2783_, data_stage_2__2782_, data_stage_2__2781_, data_stage_2__2780_, data_stage_2__2779_, data_stage_2__2778_, data_stage_2__2777_, data_stage_2__2776_, data_stage_2__2775_, data_stage_2__2774_, data_stage_2__2773_, data_stage_2__2772_, data_stage_2__2771_, data_stage_2__2770_, data_stage_2__2769_, data_stage_2__2768_, data_stage_2__2767_, data_stage_2__2766_, data_stage_2__2765_, data_stage_2__2764_, data_stage_2__2763_, data_stage_2__2762_, data_stage_2__2761_, data_stage_2__2760_, data_stage_2__2759_, data_stage_2__2758_, data_stage_2__2757_, data_stage_2__2756_, data_stage_2__2755_, data_stage_2__2754_, data_stage_2__2753_, data_stage_2__2752_, data_stage_2__2751_, data_stage_2__2750_, data_stage_2__2749_, data_stage_2__2748_, data_stage_2__2747_, data_stage_2__2746_, data_stage_2__2745_, data_stage_2__2744_, data_stage_2__2743_, data_stage_2__2742_, data_stage_2__2741_, data_stage_2__2740_, data_stage_2__2739_, data_stage_2__2738_, data_stage_2__2737_, data_stage_2__2736_, data_stage_2__2735_, data_stage_2__2734_, data_stage_2__2733_, data_stage_2__2732_, data_stage_2__2731_, data_stage_2__2730_, data_stage_2__2729_, data_stage_2__2728_, data_stage_2__2727_, data_stage_2__2726_, data_stage_2__2725_, data_stage_2__2724_, data_stage_2__2723_, data_stage_2__2722_, data_stage_2__2721_, data_stage_2__2720_, data_stage_2__2719_, data_stage_2__2718_, data_stage_2__2717_, data_stage_2__2716_, data_stage_2__2715_, data_stage_2__2714_, data_stage_2__2713_, data_stage_2__2712_, data_stage_2__2711_, data_stage_2__2710_, data_stage_2__2709_, data_stage_2__2708_, data_stage_2__2707_, data_stage_2__2706_, data_stage_2__2705_, data_stage_2__2704_, data_stage_2__2703_, data_stage_2__2702_, data_stage_2__2701_, data_stage_2__2700_, data_stage_2__2699_, data_stage_2__2698_, data_stage_2__2697_, data_stage_2__2696_, data_stage_2__2695_, data_stage_2__2694_, data_stage_2__2693_, data_stage_2__2692_, data_stage_2__2691_, data_stage_2__2690_, data_stage_2__2689_, data_stage_2__2688_, data_stage_2__2687_, data_stage_2__2686_, data_stage_2__2685_, data_stage_2__2684_, data_stage_2__2683_, data_stage_2__2682_, data_stage_2__2681_, data_stage_2__2680_, data_stage_2__2679_, data_stage_2__2678_, data_stage_2__2677_, data_stage_2__2676_, data_stage_2__2675_, data_stage_2__2674_, data_stage_2__2673_, data_stage_2__2672_, data_stage_2__2671_, data_stage_2__2670_, data_stage_2__2669_, data_stage_2__2668_, data_stage_2__2667_, data_stage_2__2666_, data_stage_2__2665_, data_stage_2__2664_, data_stage_2__2663_, data_stage_2__2662_, data_stage_2__2661_, data_stage_2__2660_, data_stage_2__2659_, data_stage_2__2658_, data_stage_2__2657_, data_stage_2__2656_, data_stage_2__2655_, data_stage_2__2654_, data_stage_2__2653_, data_stage_2__2652_, data_stage_2__2651_, data_stage_2__2650_, data_stage_2__2649_, data_stage_2__2648_, data_stage_2__2647_, data_stage_2__2646_, data_stage_2__2645_, data_stage_2__2644_, data_stage_2__2643_, data_stage_2__2642_, data_stage_2__2641_, data_stage_2__2640_, data_stage_2__2639_, data_stage_2__2638_, data_stage_2__2637_, data_stage_2__2636_, data_stage_2__2635_, data_stage_2__2634_, data_stage_2__2633_, data_stage_2__2632_, data_stage_2__2631_, data_stage_2__2630_, data_stage_2__2629_, data_stage_2__2628_, data_stage_2__2627_, data_stage_2__2626_, data_stage_2__2625_, data_stage_2__2624_, data_stage_2__2623_, data_stage_2__2622_, data_stage_2__2621_, data_stage_2__2620_, data_stage_2__2619_, data_stage_2__2618_, data_stage_2__2617_, data_stage_2__2616_, data_stage_2__2615_, data_stage_2__2614_, data_stage_2__2613_, data_stage_2__2612_, data_stage_2__2611_, data_stage_2__2610_, data_stage_2__2609_, data_stage_2__2608_, data_stage_2__2607_, data_stage_2__2606_, data_stage_2__2605_, data_stage_2__2604_, data_stage_2__2603_, data_stage_2__2602_, data_stage_2__2601_, data_stage_2__2600_, data_stage_2__2599_, data_stage_2__2598_, data_stage_2__2597_, data_stage_2__2596_, data_stage_2__2595_, data_stage_2__2594_, data_stage_2__2593_, data_stage_2__2592_, data_stage_2__2591_, data_stage_2__2590_, data_stage_2__2589_, data_stage_2__2588_, data_stage_2__2587_, data_stage_2__2586_, data_stage_2__2585_, data_stage_2__2584_, data_stage_2__2583_, data_stage_2__2582_, data_stage_2__2581_, data_stage_2__2580_, data_stage_2__2579_, data_stage_2__2578_, data_stage_2__2577_, data_stage_2__2576_, data_stage_2__2575_, data_stage_2__2574_, data_stage_2__2573_, data_stage_2__2572_, data_stage_2__2571_, data_stage_2__2570_, data_stage_2__2569_, data_stage_2__2568_, data_stage_2__2567_, data_stage_2__2566_, data_stage_2__2565_, data_stage_2__2564_, data_stage_2__2563_, data_stage_2__2562_, data_stage_2__2561_, data_stage_2__2560_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__3071_, data_stage_3__3070_, data_stage_3__3069_, data_stage_3__3068_, data_stage_3__3067_, data_stage_3__3066_, data_stage_3__3065_, data_stage_3__3064_, data_stage_3__3063_, data_stage_3__3062_, data_stage_3__3061_, data_stage_3__3060_, data_stage_3__3059_, data_stage_3__3058_, data_stage_3__3057_, data_stage_3__3056_, data_stage_3__3055_, data_stage_3__3054_, data_stage_3__3053_, data_stage_3__3052_, data_stage_3__3051_, data_stage_3__3050_, data_stage_3__3049_, data_stage_3__3048_, data_stage_3__3047_, data_stage_3__3046_, data_stage_3__3045_, data_stage_3__3044_, data_stage_3__3043_, data_stage_3__3042_, data_stage_3__3041_, data_stage_3__3040_, data_stage_3__3039_, data_stage_3__3038_, data_stage_3__3037_, data_stage_3__3036_, data_stage_3__3035_, data_stage_3__3034_, data_stage_3__3033_, data_stage_3__3032_, data_stage_3__3031_, data_stage_3__3030_, data_stage_3__3029_, data_stage_3__3028_, data_stage_3__3027_, data_stage_3__3026_, data_stage_3__3025_, data_stage_3__3024_, data_stage_3__3023_, data_stage_3__3022_, data_stage_3__3021_, data_stage_3__3020_, data_stage_3__3019_, data_stage_3__3018_, data_stage_3__3017_, data_stage_3__3016_, data_stage_3__3015_, data_stage_3__3014_, data_stage_3__3013_, data_stage_3__3012_, data_stage_3__3011_, data_stage_3__3010_, data_stage_3__3009_, data_stage_3__3008_, data_stage_3__3007_, data_stage_3__3006_, data_stage_3__3005_, data_stage_3__3004_, data_stage_3__3003_, data_stage_3__3002_, data_stage_3__3001_, data_stage_3__3000_, data_stage_3__2999_, data_stage_3__2998_, data_stage_3__2997_, data_stage_3__2996_, data_stage_3__2995_, data_stage_3__2994_, data_stage_3__2993_, data_stage_3__2992_, data_stage_3__2991_, data_stage_3__2990_, data_stage_3__2989_, data_stage_3__2988_, data_stage_3__2987_, data_stage_3__2986_, data_stage_3__2985_, data_stage_3__2984_, data_stage_3__2983_, data_stage_3__2982_, data_stage_3__2981_, data_stage_3__2980_, data_stage_3__2979_, data_stage_3__2978_, data_stage_3__2977_, data_stage_3__2976_, data_stage_3__2975_, data_stage_3__2974_, data_stage_3__2973_, data_stage_3__2972_, data_stage_3__2971_, data_stage_3__2970_, data_stage_3__2969_, data_stage_3__2968_, data_stage_3__2967_, data_stage_3__2966_, data_stage_3__2965_, data_stage_3__2964_, data_stage_3__2963_, data_stage_3__2962_, data_stage_3__2961_, data_stage_3__2960_, data_stage_3__2959_, data_stage_3__2958_, data_stage_3__2957_, data_stage_3__2956_, data_stage_3__2955_, data_stage_3__2954_, data_stage_3__2953_, data_stage_3__2952_, data_stage_3__2951_, data_stage_3__2950_, data_stage_3__2949_, data_stage_3__2948_, data_stage_3__2947_, data_stage_3__2946_, data_stage_3__2945_, data_stage_3__2944_, data_stage_3__2943_, data_stage_3__2942_, data_stage_3__2941_, data_stage_3__2940_, data_stage_3__2939_, data_stage_3__2938_, data_stage_3__2937_, data_stage_3__2936_, data_stage_3__2935_, data_stage_3__2934_, data_stage_3__2933_, data_stage_3__2932_, data_stage_3__2931_, data_stage_3__2930_, data_stage_3__2929_, data_stage_3__2928_, data_stage_3__2927_, data_stage_3__2926_, data_stage_3__2925_, data_stage_3__2924_, data_stage_3__2923_, data_stage_3__2922_, data_stage_3__2921_, data_stage_3__2920_, data_stage_3__2919_, data_stage_3__2918_, data_stage_3__2917_, data_stage_3__2916_, data_stage_3__2915_, data_stage_3__2914_, data_stage_3__2913_, data_stage_3__2912_, data_stage_3__2911_, data_stage_3__2910_, data_stage_3__2909_, data_stage_3__2908_, data_stage_3__2907_, data_stage_3__2906_, data_stage_3__2905_, data_stage_3__2904_, data_stage_3__2903_, data_stage_3__2902_, data_stage_3__2901_, data_stage_3__2900_, data_stage_3__2899_, data_stage_3__2898_, data_stage_3__2897_, data_stage_3__2896_, data_stage_3__2895_, data_stage_3__2894_, data_stage_3__2893_, data_stage_3__2892_, data_stage_3__2891_, data_stage_3__2890_, data_stage_3__2889_, data_stage_3__2888_, data_stage_3__2887_, data_stage_3__2886_, data_stage_3__2885_, data_stage_3__2884_, data_stage_3__2883_, data_stage_3__2882_, data_stage_3__2881_, data_stage_3__2880_, data_stage_3__2879_, data_stage_3__2878_, data_stage_3__2877_, data_stage_3__2876_, data_stage_3__2875_, data_stage_3__2874_, data_stage_3__2873_, data_stage_3__2872_, data_stage_3__2871_, data_stage_3__2870_, data_stage_3__2869_, data_stage_3__2868_, data_stage_3__2867_, data_stage_3__2866_, data_stage_3__2865_, data_stage_3__2864_, data_stage_3__2863_, data_stage_3__2862_, data_stage_3__2861_, data_stage_3__2860_, data_stage_3__2859_, data_stage_3__2858_, data_stage_3__2857_, data_stage_3__2856_, data_stage_3__2855_, data_stage_3__2854_, data_stage_3__2853_, data_stage_3__2852_, data_stage_3__2851_, data_stage_3__2850_, data_stage_3__2849_, data_stage_3__2848_, data_stage_3__2847_, data_stage_3__2846_, data_stage_3__2845_, data_stage_3__2844_, data_stage_3__2843_, data_stage_3__2842_, data_stage_3__2841_, data_stage_3__2840_, data_stage_3__2839_, data_stage_3__2838_, data_stage_3__2837_, data_stage_3__2836_, data_stage_3__2835_, data_stage_3__2834_, data_stage_3__2833_, data_stage_3__2832_, data_stage_3__2831_, data_stage_3__2830_, data_stage_3__2829_, data_stage_3__2828_, data_stage_3__2827_, data_stage_3__2826_, data_stage_3__2825_, data_stage_3__2824_, data_stage_3__2823_, data_stage_3__2822_, data_stage_3__2821_, data_stage_3__2820_, data_stage_3__2819_, data_stage_3__2818_, data_stage_3__2817_, data_stage_3__2816_, data_stage_3__2815_, data_stage_3__2814_, data_stage_3__2813_, data_stage_3__2812_, data_stage_3__2811_, data_stage_3__2810_, data_stage_3__2809_, data_stage_3__2808_, data_stage_3__2807_, data_stage_3__2806_, data_stage_3__2805_, data_stage_3__2804_, data_stage_3__2803_, data_stage_3__2802_, data_stage_3__2801_, data_stage_3__2800_, data_stage_3__2799_, data_stage_3__2798_, data_stage_3__2797_, data_stage_3__2796_, data_stage_3__2795_, data_stage_3__2794_, data_stage_3__2793_, data_stage_3__2792_, data_stage_3__2791_, data_stage_3__2790_, data_stage_3__2789_, data_stage_3__2788_, data_stage_3__2787_, data_stage_3__2786_, data_stage_3__2785_, data_stage_3__2784_, data_stage_3__2783_, data_stage_3__2782_, data_stage_3__2781_, data_stage_3__2780_, data_stage_3__2779_, data_stage_3__2778_, data_stage_3__2777_, data_stage_3__2776_, data_stage_3__2775_, data_stage_3__2774_, data_stage_3__2773_, data_stage_3__2772_, data_stage_3__2771_, data_stage_3__2770_, data_stage_3__2769_, data_stage_3__2768_, data_stage_3__2767_, data_stage_3__2766_, data_stage_3__2765_, data_stage_3__2764_, data_stage_3__2763_, data_stage_3__2762_, data_stage_3__2761_, data_stage_3__2760_, data_stage_3__2759_, data_stage_3__2758_, data_stage_3__2757_, data_stage_3__2756_, data_stage_3__2755_, data_stage_3__2754_, data_stage_3__2753_, data_stage_3__2752_, data_stage_3__2751_, data_stage_3__2750_, data_stage_3__2749_, data_stage_3__2748_, data_stage_3__2747_, data_stage_3__2746_, data_stage_3__2745_, data_stage_3__2744_, data_stage_3__2743_, data_stage_3__2742_, data_stage_3__2741_, data_stage_3__2740_, data_stage_3__2739_, data_stage_3__2738_, data_stage_3__2737_, data_stage_3__2736_, data_stage_3__2735_, data_stage_3__2734_, data_stage_3__2733_, data_stage_3__2732_, data_stage_3__2731_, data_stage_3__2730_, data_stage_3__2729_, data_stage_3__2728_, data_stage_3__2727_, data_stage_3__2726_, data_stage_3__2725_, data_stage_3__2724_, data_stage_3__2723_, data_stage_3__2722_, data_stage_3__2721_, data_stage_3__2720_, data_stage_3__2719_, data_stage_3__2718_, data_stage_3__2717_, data_stage_3__2716_, data_stage_3__2715_, data_stage_3__2714_, data_stage_3__2713_, data_stage_3__2712_, data_stage_3__2711_, data_stage_3__2710_, data_stage_3__2709_, data_stage_3__2708_, data_stage_3__2707_, data_stage_3__2706_, data_stage_3__2705_, data_stage_3__2704_, data_stage_3__2703_, data_stage_3__2702_, data_stage_3__2701_, data_stage_3__2700_, data_stage_3__2699_, data_stage_3__2698_, data_stage_3__2697_, data_stage_3__2696_, data_stage_3__2695_, data_stage_3__2694_, data_stage_3__2693_, data_stage_3__2692_, data_stage_3__2691_, data_stage_3__2690_, data_stage_3__2689_, data_stage_3__2688_, data_stage_3__2687_, data_stage_3__2686_, data_stage_3__2685_, data_stage_3__2684_, data_stage_3__2683_, data_stage_3__2682_, data_stage_3__2681_, data_stage_3__2680_, data_stage_3__2679_, data_stage_3__2678_, data_stage_3__2677_, data_stage_3__2676_, data_stage_3__2675_, data_stage_3__2674_, data_stage_3__2673_, data_stage_3__2672_, data_stage_3__2671_, data_stage_3__2670_, data_stage_3__2669_, data_stage_3__2668_, data_stage_3__2667_, data_stage_3__2666_, data_stage_3__2665_, data_stage_3__2664_, data_stage_3__2663_, data_stage_3__2662_, data_stage_3__2661_, data_stage_3__2660_, data_stage_3__2659_, data_stage_3__2658_, data_stage_3__2657_, data_stage_3__2656_, data_stage_3__2655_, data_stage_3__2654_, data_stage_3__2653_, data_stage_3__2652_, data_stage_3__2651_, data_stage_3__2650_, data_stage_3__2649_, data_stage_3__2648_, data_stage_3__2647_, data_stage_3__2646_, data_stage_3__2645_, data_stage_3__2644_, data_stage_3__2643_, data_stage_3__2642_, data_stage_3__2641_, data_stage_3__2640_, data_stage_3__2639_, data_stage_3__2638_, data_stage_3__2637_, data_stage_3__2636_, data_stage_3__2635_, data_stage_3__2634_, data_stage_3__2633_, data_stage_3__2632_, data_stage_3__2631_, data_stage_3__2630_, data_stage_3__2629_, data_stage_3__2628_, data_stage_3__2627_, data_stage_3__2626_, data_stage_3__2625_, data_stage_3__2624_, data_stage_3__2623_, data_stage_3__2622_, data_stage_3__2621_, data_stage_3__2620_, data_stage_3__2619_, data_stage_3__2618_, data_stage_3__2617_, data_stage_3__2616_, data_stage_3__2615_, data_stage_3__2614_, data_stage_3__2613_, data_stage_3__2612_, data_stage_3__2611_, data_stage_3__2610_, data_stage_3__2609_, data_stage_3__2608_, data_stage_3__2607_, data_stage_3__2606_, data_stage_3__2605_, data_stage_3__2604_, data_stage_3__2603_, data_stage_3__2602_, data_stage_3__2601_, data_stage_3__2600_, data_stage_3__2599_, data_stage_3__2598_, data_stage_3__2597_, data_stage_3__2596_, data_stage_3__2595_, data_stage_3__2594_, data_stage_3__2593_, data_stage_3__2592_, data_stage_3__2591_, data_stage_3__2590_, data_stage_3__2589_, data_stage_3__2588_, data_stage_3__2587_, data_stage_3__2586_, data_stage_3__2585_, data_stage_3__2584_, data_stage_3__2583_, data_stage_3__2582_, data_stage_3__2581_, data_stage_3__2580_, data_stage_3__2579_, data_stage_3__2578_, data_stage_3__2577_, data_stage_3__2576_, data_stage_3__2575_, data_stage_3__2574_, data_stage_3__2573_, data_stage_3__2572_, data_stage_3__2571_, data_stage_3__2570_, data_stage_3__2569_, data_stage_3__2568_, data_stage_3__2567_, data_stage_3__2566_, data_stage_3__2565_, data_stage_3__2564_, data_stage_3__2563_, data_stage_3__2562_, data_stage_3__2561_, data_stage_3__2560_ })
  );


  bsg_swap_width_p256
  mux_stage_2__mux_swap_6__swap_inst
  (
    .data_i({ data_stage_2__3583_, data_stage_2__3582_, data_stage_2__3581_, data_stage_2__3580_, data_stage_2__3579_, data_stage_2__3578_, data_stage_2__3577_, data_stage_2__3576_, data_stage_2__3575_, data_stage_2__3574_, data_stage_2__3573_, data_stage_2__3572_, data_stage_2__3571_, data_stage_2__3570_, data_stage_2__3569_, data_stage_2__3568_, data_stage_2__3567_, data_stage_2__3566_, data_stage_2__3565_, data_stage_2__3564_, data_stage_2__3563_, data_stage_2__3562_, data_stage_2__3561_, data_stage_2__3560_, data_stage_2__3559_, data_stage_2__3558_, data_stage_2__3557_, data_stage_2__3556_, data_stage_2__3555_, data_stage_2__3554_, data_stage_2__3553_, data_stage_2__3552_, data_stage_2__3551_, data_stage_2__3550_, data_stage_2__3549_, data_stage_2__3548_, data_stage_2__3547_, data_stage_2__3546_, data_stage_2__3545_, data_stage_2__3544_, data_stage_2__3543_, data_stage_2__3542_, data_stage_2__3541_, data_stage_2__3540_, data_stage_2__3539_, data_stage_2__3538_, data_stage_2__3537_, data_stage_2__3536_, data_stage_2__3535_, data_stage_2__3534_, data_stage_2__3533_, data_stage_2__3532_, data_stage_2__3531_, data_stage_2__3530_, data_stage_2__3529_, data_stage_2__3528_, data_stage_2__3527_, data_stage_2__3526_, data_stage_2__3525_, data_stage_2__3524_, data_stage_2__3523_, data_stage_2__3522_, data_stage_2__3521_, data_stage_2__3520_, data_stage_2__3519_, data_stage_2__3518_, data_stage_2__3517_, data_stage_2__3516_, data_stage_2__3515_, data_stage_2__3514_, data_stage_2__3513_, data_stage_2__3512_, data_stage_2__3511_, data_stage_2__3510_, data_stage_2__3509_, data_stage_2__3508_, data_stage_2__3507_, data_stage_2__3506_, data_stage_2__3505_, data_stage_2__3504_, data_stage_2__3503_, data_stage_2__3502_, data_stage_2__3501_, data_stage_2__3500_, data_stage_2__3499_, data_stage_2__3498_, data_stage_2__3497_, data_stage_2__3496_, data_stage_2__3495_, data_stage_2__3494_, data_stage_2__3493_, data_stage_2__3492_, data_stage_2__3491_, data_stage_2__3490_, data_stage_2__3489_, data_stage_2__3488_, data_stage_2__3487_, data_stage_2__3486_, data_stage_2__3485_, data_stage_2__3484_, data_stage_2__3483_, data_stage_2__3482_, data_stage_2__3481_, data_stage_2__3480_, data_stage_2__3479_, data_stage_2__3478_, data_stage_2__3477_, data_stage_2__3476_, data_stage_2__3475_, data_stage_2__3474_, data_stage_2__3473_, data_stage_2__3472_, data_stage_2__3471_, data_stage_2__3470_, data_stage_2__3469_, data_stage_2__3468_, data_stage_2__3467_, data_stage_2__3466_, data_stage_2__3465_, data_stage_2__3464_, data_stage_2__3463_, data_stage_2__3462_, data_stage_2__3461_, data_stage_2__3460_, data_stage_2__3459_, data_stage_2__3458_, data_stage_2__3457_, data_stage_2__3456_, data_stage_2__3455_, data_stage_2__3454_, data_stage_2__3453_, data_stage_2__3452_, data_stage_2__3451_, data_stage_2__3450_, data_stage_2__3449_, data_stage_2__3448_, data_stage_2__3447_, data_stage_2__3446_, data_stage_2__3445_, data_stage_2__3444_, data_stage_2__3443_, data_stage_2__3442_, data_stage_2__3441_, data_stage_2__3440_, data_stage_2__3439_, data_stage_2__3438_, data_stage_2__3437_, data_stage_2__3436_, data_stage_2__3435_, data_stage_2__3434_, data_stage_2__3433_, data_stage_2__3432_, data_stage_2__3431_, data_stage_2__3430_, data_stage_2__3429_, data_stage_2__3428_, data_stage_2__3427_, data_stage_2__3426_, data_stage_2__3425_, data_stage_2__3424_, data_stage_2__3423_, data_stage_2__3422_, data_stage_2__3421_, data_stage_2__3420_, data_stage_2__3419_, data_stage_2__3418_, data_stage_2__3417_, data_stage_2__3416_, data_stage_2__3415_, data_stage_2__3414_, data_stage_2__3413_, data_stage_2__3412_, data_stage_2__3411_, data_stage_2__3410_, data_stage_2__3409_, data_stage_2__3408_, data_stage_2__3407_, data_stage_2__3406_, data_stage_2__3405_, data_stage_2__3404_, data_stage_2__3403_, data_stage_2__3402_, data_stage_2__3401_, data_stage_2__3400_, data_stage_2__3399_, data_stage_2__3398_, data_stage_2__3397_, data_stage_2__3396_, data_stage_2__3395_, data_stage_2__3394_, data_stage_2__3393_, data_stage_2__3392_, data_stage_2__3391_, data_stage_2__3390_, data_stage_2__3389_, data_stage_2__3388_, data_stage_2__3387_, data_stage_2__3386_, data_stage_2__3385_, data_stage_2__3384_, data_stage_2__3383_, data_stage_2__3382_, data_stage_2__3381_, data_stage_2__3380_, data_stage_2__3379_, data_stage_2__3378_, data_stage_2__3377_, data_stage_2__3376_, data_stage_2__3375_, data_stage_2__3374_, data_stage_2__3373_, data_stage_2__3372_, data_stage_2__3371_, data_stage_2__3370_, data_stage_2__3369_, data_stage_2__3368_, data_stage_2__3367_, data_stage_2__3366_, data_stage_2__3365_, data_stage_2__3364_, data_stage_2__3363_, data_stage_2__3362_, data_stage_2__3361_, data_stage_2__3360_, data_stage_2__3359_, data_stage_2__3358_, data_stage_2__3357_, data_stage_2__3356_, data_stage_2__3355_, data_stage_2__3354_, data_stage_2__3353_, data_stage_2__3352_, data_stage_2__3351_, data_stage_2__3350_, data_stage_2__3349_, data_stage_2__3348_, data_stage_2__3347_, data_stage_2__3346_, data_stage_2__3345_, data_stage_2__3344_, data_stage_2__3343_, data_stage_2__3342_, data_stage_2__3341_, data_stage_2__3340_, data_stage_2__3339_, data_stage_2__3338_, data_stage_2__3337_, data_stage_2__3336_, data_stage_2__3335_, data_stage_2__3334_, data_stage_2__3333_, data_stage_2__3332_, data_stage_2__3331_, data_stage_2__3330_, data_stage_2__3329_, data_stage_2__3328_, data_stage_2__3327_, data_stage_2__3326_, data_stage_2__3325_, data_stage_2__3324_, data_stage_2__3323_, data_stage_2__3322_, data_stage_2__3321_, data_stage_2__3320_, data_stage_2__3319_, data_stage_2__3318_, data_stage_2__3317_, data_stage_2__3316_, data_stage_2__3315_, data_stage_2__3314_, data_stage_2__3313_, data_stage_2__3312_, data_stage_2__3311_, data_stage_2__3310_, data_stage_2__3309_, data_stage_2__3308_, data_stage_2__3307_, data_stage_2__3306_, data_stage_2__3305_, data_stage_2__3304_, data_stage_2__3303_, data_stage_2__3302_, data_stage_2__3301_, data_stage_2__3300_, data_stage_2__3299_, data_stage_2__3298_, data_stage_2__3297_, data_stage_2__3296_, data_stage_2__3295_, data_stage_2__3294_, data_stage_2__3293_, data_stage_2__3292_, data_stage_2__3291_, data_stage_2__3290_, data_stage_2__3289_, data_stage_2__3288_, data_stage_2__3287_, data_stage_2__3286_, data_stage_2__3285_, data_stage_2__3284_, data_stage_2__3283_, data_stage_2__3282_, data_stage_2__3281_, data_stage_2__3280_, data_stage_2__3279_, data_stage_2__3278_, data_stage_2__3277_, data_stage_2__3276_, data_stage_2__3275_, data_stage_2__3274_, data_stage_2__3273_, data_stage_2__3272_, data_stage_2__3271_, data_stage_2__3270_, data_stage_2__3269_, data_stage_2__3268_, data_stage_2__3267_, data_stage_2__3266_, data_stage_2__3265_, data_stage_2__3264_, data_stage_2__3263_, data_stage_2__3262_, data_stage_2__3261_, data_stage_2__3260_, data_stage_2__3259_, data_stage_2__3258_, data_stage_2__3257_, data_stage_2__3256_, data_stage_2__3255_, data_stage_2__3254_, data_stage_2__3253_, data_stage_2__3252_, data_stage_2__3251_, data_stage_2__3250_, data_stage_2__3249_, data_stage_2__3248_, data_stage_2__3247_, data_stage_2__3246_, data_stage_2__3245_, data_stage_2__3244_, data_stage_2__3243_, data_stage_2__3242_, data_stage_2__3241_, data_stage_2__3240_, data_stage_2__3239_, data_stage_2__3238_, data_stage_2__3237_, data_stage_2__3236_, data_stage_2__3235_, data_stage_2__3234_, data_stage_2__3233_, data_stage_2__3232_, data_stage_2__3231_, data_stage_2__3230_, data_stage_2__3229_, data_stage_2__3228_, data_stage_2__3227_, data_stage_2__3226_, data_stage_2__3225_, data_stage_2__3224_, data_stage_2__3223_, data_stage_2__3222_, data_stage_2__3221_, data_stage_2__3220_, data_stage_2__3219_, data_stage_2__3218_, data_stage_2__3217_, data_stage_2__3216_, data_stage_2__3215_, data_stage_2__3214_, data_stage_2__3213_, data_stage_2__3212_, data_stage_2__3211_, data_stage_2__3210_, data_stage_2__3209_, data_stage_2__3208_, data_stage_2__3207_, data_stage_2__3206_, data_stage_2__3205_, data_stage_2__3204_, data_stage_2__3203_, data_stage_2__3202_, data_stage_2__3201_, data_stage_2__3200_, data_stage_2__3199_, data_stage_2__3198_, data_stage_2__3197_, data_stage_2__3196_, data_stage_2__3195_, data_stage_2__3194_, data_stage_2__3193_, data_stage_2__3192_, data_stage_2__3191_, data_stage_2__3190_, data_stage_2__3189_, data_stage_2__3188_, data_stage_2__3187_, data_stage_2__3186_, data_stage_2__3185_, data_stage_2__3184_, data_stage_2__3183_, data_stage_2__3182_, data_stage_2__3181_, data_stage_2__3180_, data_stage_2__3179_, data_stage_2__3178_, data_stage_2__3177_, data_stage_2__3176_, data_stage_2__3175_, data_stage_2__3174_, data_stage_2__3173_, data_stage_2__3172_, data_stage_2__3171_, data_stage_2__3170_, data_stage_2__3169_, data_stage_2__3168_, data_stage_2__3167_, data_stage_2__3166_, data_stage_2__3165_, data_stage_2__3164_, data_stage_2__3163_, data_stage_2__3162_, data_stage_2__3161_, data_stage_2__3160_, data_stage_2__3159_, data_stage_2__3158_, data_stage_2__3157_, data_stage_2__3156_, data_stage_2__3155_, data_stage_2__3154_, data_stage_2__3153_, data_stage_2__3152_, data_stage_2__3151_, data_stage_2__3150_, data_stage_2__3149_, data_stage_2__3148_, data_stage_2__3147_, data_stage_2__3146_, data_stage_2__3145_, data_stage_2__3144_, data_stage_2__3143_, data_stage_2__3142_, data_stage_2__3141_, data_stage_2__3140_, data_stage_2__3139_, data_stage_2__3138_, data_stage_2__3137_, data_stage_2__3136_, data_stage_2__3135_, data_stage_2__3134_, data_stage_2__3133_, data_stage_2__3132_, data_stage_2__3131_, data_stage_2__3130_, data_stage_2__3129_, data_stage_2__3128_, data_stage_2__3127_, data_stage_2__3126_, data_stage_2__3125_, data_stage_2__3124_, data_stage_2__3123_, data_stage_2__3122_, data_stage_2__3121_, data_stage_2__3120_, data_stage_2__3119_, data_stage_2__3118_, data_stage_2__3117_, data_stage_2__3116_, data_stage_2__3115_, data_stage_2__3114_, data_stage_2__3113_, data_stage_2__3112_, data_stage_2__3111_, data_stage_2__3110_, data_stage_2__3109_, data_stage_2__3108_, data_stage_2__3107_, data_stage_2__3106_, data_stage_2__3105_, data_stage_2__3104_, data_stage_2__3103_, data_stage_2__3102_, data_stage_2__3101_, data_stage_2__3100_, data_stage_2__3099_, data_stage_2__3098_, data_stage_2__3097_, data_stage_2__3096_, data_stage_2__3095_, data_stage_2__3094_, data_stage_2__3093_, data_stage_2__3092_, data_stage_2__3091_, data_stage_2__3090_, data_stage_2__3089_, data_stage_2__3088_, data_stage_2__3087_, data_stage_2__3086_, data_stage_2__3085_, data_stage_2__3084_, data_stage_2__3083_, data_stage_2__3082_, data_stage_2__3081_, data_stage_2__3080_, data_stage_2__3079_, data_stage_2__3078_, data_stage_2__3077_, data_stage_2__3076_, data_stage_2__3075_, data_stage_2__3074_, data_stage_2__3073_, data_stage_2__3072_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__3583_, data_stage_3__3582_, data_stage_3__3581_, data_stage_3__3580_, data_stage_3__3579_, data_stage_3__3578_, data_stage_3__3577_, data_stage_3__3576_, data_stage_3__3575_, data_stage_3__3574_, data_stage_3__3573_, data_stage_3__3572_, data_stage_3__3571_, data_stage_3__3570_, data_stage_3__3569_, data_stage_3__3568_, data_stage_3__3567_, data_stage_3__3566_, data_stage_3__3565_, data_stage_3__3564_, data_stage_3__3563_, data_stage_3__3562_, data_stage_3__3561_, data_stage_3__3560_, data_stage_3__3559_, data_stage_3__3558_, data_stage_3__3557_, data_stage_3__3556_, data_stage_3__3555_, data_stage_3__3554_, data_stage_3__3553_, data_stage_3__3552_, data_stage_3__3551_, data_stage_3__3550_, data_stage_3__3549_, data_stage_3__3548_, data_stage_3__3547_, data_stage_3__3546_, data_stage_3__3545_, data_stage_3__3544_, data_stage_3__3543_, data_stage_3__3542_, data_stage_3__3541_, data_stage_3__3540_, data_stage_3__3539_, data_stage_3__3538_, data_stage_3__3537_, data_stage_3__3536_, data_stage_3__3535_, data_stage_3__3534_, data_stage_3__3533_, data_stage_3__3532_, data_stage_3__3531_, data_stage_3__3530_, data_stage_3__3529_, data_stage_3__3528_, data_stage_3__3527_, data_stage_3__3526_, data_stage_3__3525_, data_stage_3__3524_, data_stage_3__3523_, data_stage_3__3522_, data_stage_3__3521_, data_stage_3__3520_, data_stage_3__3519_, data_stage_3__3518_, data_stage_3__3517_, data_stage_3__3516_, data_stage_3__3515_, data_stage_3__3514_, data_stage_3__3513_, data_stage_3__3512_, data_stage_3__3511_, data_stage_3__3510_, data_stage_3__3509_, data_stage_3__3508_, data_stage_3__3507_, data_stage_3__3506_, data_stage_3__3505_, data_stage_3__3504_, data_stage_3__3503_, data_stage_3__3502_, data_stage_3__3501_, data_stage_3__3500_, data_stage_3__3499_, data_stage_3__3498_, data_stage_3__3497_, data_stage_3__3496_, data_stage_3__3495_, data_stage_3__3494_, data_stage_3__3493_, data_stage_3__3492_, data_stage_3__3491_, data_stage_3__3490_, data_stage_3__3489_, data_stage_3__3488_, data_stage_3__3487_, data_stage_3__3486_, data_stage_3__3485_, data_stage_3__3484_, data_stage_3__3483_, data_stage_3__3482_, data_stage_3__3481_, data_stage_3__3480_, data_stage_3__3479_, data_stage_3__3478_, data_stage_3__3477_, data_stage_3__3476_, data_stage_3__3475_, data_stage_3__3474_, data_stage_3__3473_, data_stage_3__3472_, data_stage_3__3471_, data_stage_3__3470_, data_stage_3__3469_, data_stage_3__3468_, data_stage_3__3467_, data_stage_3__3466_, data_stage_3__3465_, data_stage_3__3464_, data_stage_3__3463_, data_stage_3__3462_, data_stage_3__3461_, data_stage_3__3460_, data_stage_3__3459_, data_stage_3__3458_, data_stage_3__3457_, data_stage_3__3456_, data_stage_3__3455_, data_stage_3__3454_, data_stage_3__3453_, data_stage_3__3452_, data_stage_3__3451_, data_stage_3__3450_, data_stage_3__3449_, data_stage_3__3448_, data_stage_3__3447_, data_stage_3__3446_, data_stage_3__3445_, data_stage_3__3444_, data_stage_3__3443_, data_stage_3__3442_, data_stage_3__3441_, data_stage_3__3440_, data_stage_3__3439_, data_stage_3__3438_, data_stage_3__3437_, data_stage_3__3436_, data_stage_3__3435_, data_stage_3__3434_, data_stage_3__3433_, data_stage_3__3432_, data_stage_3__3431_, data_stage_3__3430_, data_stage_3__3429_, data_stage_3__3428_, data_stage_3__3427_, data_stage_3__3426_, data_stage_3__3425_, data_stage_3__3424_, data_stage_3__3423_, data_stage_3__3422_, data_stage_3__3421_, data_stage_3__3420_, data_stage_3__3419_, data_stage_3__3418_, data_stage_3__3417_, data_stage_3__3416_, data_stage_3__3415_, data_stage_3__3414_, data_stage_3__3413_, data_stage_3__3412_, data_stage_3__3411_, data_stage_3__3410_, data_stage_3__3409_, data_stage_3__3408_, data_stage_3__3407_, data_stage_3__3406_, data_stage_3__3405_, data_stage_3__3404_, data_stage_3__3403_, data_stage_3__3402_, data_stage_3__3401_, data_stage_3__3400_, data_stage_3__3399_, data_stage_3__3398_, data_stage_3__3397_, data_stage_3__3396_, data_stage_3__3395_, data_stage_3__3394_, data_stage_3__3393_, data_stage_3__3392_, data_stage_3__3391_, data_stage_3__3390_, data_stage_3__3389_, data_stage_3__3388_, data_stage_3__3387_, data_stage_3__3386_, data_stage_3__3385_, data_stage_3__3384_, data_stage_3__3383_, data_stage_3__3382_, data_stage_3__3381_, data_stage_3__3380_, data_stage_3__3379_, data_stage_3__3378_, data_stage_3__3377_, data_stage_3__3376_, data_stage_3__3375_, data_stage_3__3374_, data_stage_3__3373_, data_stage_3__3372_, data_stage_3__3371_, data_stage_3__3370_, data_stage_3__3369_, data_stage_3__3368_, data_stage_3__3367_, data_stage_3__3366_, data_stage_3__3365_, data_stage_3__3364_, data_stage_3__3363_, data_stage_3__3362_, data_stage_3__3361_, data_stage_3__3360_, data_stage_3__3359_, data_stage_3__3358_, data_stage_3__3357_, data_stage_3__3356_, data_stage_3__3355_, data_stage_3__3354_, data_stage_3__3353_, data_stage_3__3352_, data_stage_3__3351_, data_stage_3__3350_, data_stage_3__3349_, data_stage_3__3348_, data_stage_3__3347_, data_stage_3__3346_, data_stage_3__3345_, data_stage_3__3344_, data_stage_3__3343_, data_stage_3__3342_, data_stage_3__3341_, data_stage_3__3340_, data_stage_3__3339_, data_stage_3__3338_, data_stage_3__3337_, data_stage_3__3336_, data_stage_3__3335_, data_stage_3__3334_, data_stage_3__3333_, data_stage_3__3332_, data_stage_3__3331_, data_stage_3__3330_, data_stage_3__3329_, data_stage_3__3328_, data_stage_3__3327_, data_stage_3__3326_, data_stage_3__3325_, data_stage_3__3324_, data_stage_3__3323_, data_stage_3__3322_, data_stage_3__3321_, data_stage_3__3320_, data_stage_3__3319_, data_stage_3__3318_, data_stage_3__3317_, data_stage_3__3316_, data_stage_3__3315_, data_stage_3__3314_, data_stage_3__3313_, data_stage_3__3312_, data_stage_3__3311_, data_stage_3__3310_, data_stage_3__3309_, data_stage_3__3308_, data_stage_3__3307_, data_stage_3__3306_, data_stage_3__3305_, data_stage_3__3304_, data_stage_3__3303_, data_stage_3__3302_, data_stage_3__3301_, data_stage_3__3300_, data_stage_3__3299_, data_stage_3__3298_, data_stage_3__3297_, data_stage_3__3296_, data_stage_3__3295_, data_stage_3__3294_, data_stage_3__3293_, data_stage_3__3292_, data_stage_3__3291_, data_stage_3__3290_, data_stage_3__3289_, data_stage_3__3288_, data_stage_3__3287_, data_stage_3__3286_, data_stage_3__3285_, data_stage_3__3284_, data_stage_3__3283_, data_stage_3__3282_, data_stage_3__3281_, data_stage_3__3280_, data_stage_3__3279_, data_stage_3__3278_, data_stage_3__3277_, data_stage_3__3276_, data_stage_3__3275_, data_stage_3__3274_, data_stage_3__3273_, data_stage_3__3272_, data_stage_3__3271_, data_stage_3__3270_, data_stage_3__3269_, data_stage_3__3268_, data_stage_3__3267_, data_stage_3__3266_, data_stage_3__3265_, data_stage_3__3264_, data_stage_3__3263_, data_stage_3__3262_, data_stage_3__3261_, data_stage_3__3260_, data_stage_3__3259_, data_stage_3__3258_, data_stage_3__3257_, data_stage_3__3256_, data_stage_3__3255_, data_stage_3__3254_, data_stage_3__3253_, data_stage_3__3252_, data_stage_3__3251_, data_stage_3__3250_, data_stage_3__3249_, data_stage_3__3248_, data_stage_3__3247_, data_stage_3__3246_, data_stage_3__3245_, data_stage_3__3244_, data_stage_3__3243_, data_stage_3__3242_, data_stage_3__3241_, data_stage_3__3240_, data_stage_3__3239_, data_stage_3__3238_, data_stage_3__3237_, data_stage_3__3236_, data_stage_3__3235_, data_stage_3__3234_, data_stage_3__3233_, data_stage_3__3232_, data_stage_3__3231_, data_stage_3__3230_, data_stage_3__3229_, data_stage_3__3228_, data_stage_3__3227_, data_stage_3__3226_, data_stage_3__3225_, data_stage_3__3224_, data_stage_3__3223_, data_stage_3__3222_, data_stage_3__3221_, data_stage_3__3220_, data_stage_3__3219_, data_stage_3__3218_, data_stage_3__3217_, data_stage_3__3216_, data_stage_3__3215_, data_stage_3__3214_, data_stage_3__3213_, data_stage_3__3212_, data_stage_3__3211_, data_stage_3__3210_, data_stage_3__3209_, data_stage_3__3208_, data_stage_3__3207_, data_stage_3__3206_, data_stage_3__3205_, data_stage_3__3204_, data_stage_3__3203_, data_stage_3__3202_, data_stage_3__3201_, data_stage_3__3200_, data_stage_3__3199_, data_stage_3__3198_, data_stage_3__3197_, data_stage_3__3196_, data_stage_3__3195_, data_stage_3__3194_, data_stage_3__3193_, data_stage_3__3192_, data_stage_3__3191_, data_stage_3__3190_, data_stage_3__3189_, data_stage_3__3188_, data_stage_3__3187_, data_stage_3__3186_, data_stage_3__3185_, data_stage_3__3184_, data_stage_3__3183_, data_stage_3__3182_, data_stage_3__3181_, data_stage_3__3180_, data_stage_3__3179_, data_stage_3__3178_, data_stage_3__3177_, data_stage_3__3176_, data_stage_3__3175_, data_stage_3__3174_, data_stage_3__3173_, data_stage_3__3172_, data_stage_3__3171_, data_stage_3__3170_, data_stage_3__3169_, data_stage_3__3168_, data_stage_3__3167_, data_stage_3__3166_, data_stage_3__3165_, data_stage_3__3164_, data_stage_3__3163_, data_stage_3__3162_, data_stage_3__3161_, data_stage_3__3160_, data_stage_3__3159_, data_stage_3__3158_, data_stage_3__3157_, data_stage_3__3156_, data_stage_3__3155_, data_stage_3__3154_, data_stage_3__3153_, data_stage_3__3152_, data_stage_3__3151_, data_stage_3__3150_, data_stage_3__3149_, data_stage_3__3148_, data_stage_3__3147_, data_stage_3__3146_, data_stage_3__3145_, data_stage_3__3144_, data_stage_3__3143_, data_stage_3__3142_, data_stage_3__3141_, data_stage_3__3140_, data_stage_3__3139_, data_stage_3__3138_, data_stage_3__3137_, data_stage_3__3136_, data_stage_3__3135_, data_stage_3__3134_, data_stage_3__3133_, data_stage_3__3132_, data_stage_3__3131_, data_stage_3__3130_, data_stage_3__3129_, data_stage_3__3128_, data_stage_3__3127_, data_stage_3__3126_, data_stage_3__3125_, data_stage_3__3124_, data_stage_3__3123_, data_stage_3__3122_, data_stage_3__3121_, data_stage_3__3120_, data_stage_3__3119_, data_stage_3__3118_, data_stage_3__3117_, data_stage_3__3116_, data_stage_3__3115_, data_stage_3__3114_, data_stage_3__3113_, data_stage_3__3112_, data_stage_3__3111_, data_stage_3__3110_, data_stage_3__3109_, data_stage_3__3108_, data_stage_3__3107_, data_stage_3__3106_, data_stage_3__3105_, data_stage_3__3104_, data_stage_3__3103_, data_stage_3__3102_, data_stage_3__3101_, data_stage_3__3100_, data_stage_3__3099_, data_stage_3__3098_, data_stage_3__3097_, data_stage_3__3096_, data_stage_3__3095_, data_stage_3__3094_, data_stage_3__3093_, data_stage_3__3092_, data_stage_3__3091_, data_stage_3__3090_, data_stage_3__3089_, data_stage_3__3088_, data_stage_3__3087_, data_stage_3__3086_, data_stage_3__3085_, data_stage_3__3084_, data_stage_3__3083_, data_stage_3__3082_, data_stage_3__3081_, data_stage_3__3080_, data_stage_3__3079_, data_stage_3__3078_, data_stage_3__3077_, data_stage_3__3076_, data_stage_3__3075_, data_stage_3__3074_, data_stage_3__3073_, data_stage_3__3072_ })
  );


  bsg_swap_width_p256
  mux_stage_2__mux_swap_7__swap_inst
  (
    .data_i({ data_stage_2__4095_, data_stage_2__4094_, data_stage_2__4093_, data_stage_2__4092_, data_stage_2__4091_, data_stage_2__4090_, data_stage_2__4089_, data_stage_2__4088_, data_stage_2__4087_, data_stage_2__4086_, data_stage_2__4085_, data_stage_2__4084_, data_stage_2__4083_, data_stage_2__4082_, data_stage_2__4081_, data_stage_2__4080_, data_stage_2__4079_, data_stage_2__4078_, data_stage_2__4077_, data_stage_2__4076_, data_stage_2__4075_, data_stage_2__4074_, data_stage_2__4073_, data_stage_2__4072_, data_stage_2__4071_, data_stage_2__4070_, data_stage_2__4069_, data_stage_2__4068_, data_stage_2__4067_, data_stage_2__4066_, data_stage_2__4065_, data_stage_2__4064_, data_stage_2__4063_, data_stage_2__4062_, data_stage_2__4061_, data_stage_2__4060_, data_stage_2__4059_, data_stage_2__4058_, data_stage_2__4057_, data_stage_2__4056_, data_stage_2__4055_, data_stage_2__4054_, data_stage_2__4053_, data_stage_2__4052_, data_stage_2__4051_, data_stage_2__4050_, data_stage_2__4049_, data_stage_2__4048_, data_stage_2__4047_, data_stage_2__4046_, data_stage_2__4045_, data_stage_2__4044_, data_stage_2__4043_, data_stage_2__4042_, data_stage_2__4041_, data_stage_2__4040_, data_stage_2__4039_, data_stage_2__4038_, data_stage_2__4037_, data_stage_2__4036_, data_stage_2__4035_, data_stage_2__4034_, data_stage_2__4033_, data_stage_2__4032_, data_stage_2__4031_, data_stage_2__4030_, data_stage_2__4029_, data_stage_2__4028_, data_stage_2__4027_, data_stage_2__4026_, data_stage_2__4025_, data_stage_2__4024_, data_stage_2__4023_, data_stage_2__4022_, data_stage_2__4021_, data_stage_2__4020_, data_stage_2__4019_, data_stage_2__4018_, data_stage_2__4017_, data_stage_2__4016_, data_stage_2__4015_, data_stage_2__4014_, data_stage_2__4013_, data_stage_2__4012_, data_stage_2__4011_, data_stage_2__4010_, data_stage_2__4009_, data_stage_2__4008_, data_stage_2__4007_, data_stage_2__4006_, data_stage_2__4005_, data_stage_2__4004_, data_stage_2__4003_, data_stage_2__4002_, data_stage_2__4001_, data_stage_2__4000_, data_stage_2__3999_, data_stage_2__3998_, data_stage_2__3997_, data_stage_2__3996_, data_stage_2__3995_, data_stage_2__3994_, data_stage_2__3993_, data_stage_2__3992_, data_stage_2__3991_, data_stage_2__3990_, data_stage_2__3989_, data_stage_2__3988_, data_stage_2__3987_, data_stage_2__3986_, data_stage_2__3985_, data_stage_2__3984_, data_stage_2__3983_, data_stage_2__3982_, data_stage_2__3981_, data_stage_2__3980_, data_stage_2__3979_, data_stage_2__3978_, data_stage_2__3977_, data_stage_2__3976_, data_stage_2__3975_, data_stage_2__3974_, data_stage_2__3973_, data_stage_2__3972_, data_stage_2__3971_, data_stage_2__3970_, data_stage_2__3969_, data_stage_2__3968_, data_stage_2__3967_, data_stage_2__3966_, data_stage_2__3965_, data_stage_2__3964_, data_stage_2__3963_, data_stage_2__3962_, data_stage_2__3961_, data_stage_2__3960_, data_stage_2__3959_, data_stage_2__3958_, data_stage_2__3957_, data_stage_2__3956_, data_stage_2__3955_, data_stage_2__3954_, data_stage_2__3953_, data_stage_2__3952_, data_stage_2__3951_, data_stage_2__3950_, data_stage_2__3949_, data_stage_2__3948_, data_stage_2__3947_, data_stage_2__3946_, data_stage_2__3945_, data_stage_2__3944_, data_stage_2__3943_, data_stage_2__3942_, data_stage_2__3941_, data_stage_2__3940_, data_stage_2__3939_, data_stage_2__3938_, data_stage_2__3937_, data_stage_2__3936_, data_stage_2__3935_, data_stage_2__3934_, data_stage_2__3933_, data_stage_2__3932_, data_stage_2__3931_, data_stage_2__3930_, data_stage_2__3929_, data_stage_2__3928_, data_stage_2__3927_, data_stage_2__3926_, data_stage_2__3925_, data_stage_2__3924_, data_stage_2__3923_, data_stage_2__3922_, data_stage_2__3921_, data_stage_2__3920_, data_stage_2__3919_, data_stage_2__3918_, data_stage_2__3917_, data_stage_2__3916_, data_stage_2__3915_, data_stage_2__3914_, data_stage_2__3913_, data_stage_2__3912_, data_stage_2__3911_, data_stage_2__3910_, data_stage_2__3909_, data_stage_2__3908_, data_stage_2__3907_, data_stage_2__3906_, data_stage_2__3905_, data_stage_2__3904_, data_stage_2__3903_, data_stage_2__3902_, data_stage_2__3901_, data_stage_2__3900_, data_stage_2__3899_, data_stage_2__3898_, data_stage_2__3897_, data_stage_2__3896_, data_stage_2__3895_, data_stage_2__3894_, data_stage_2__3893_, data_stage_2__3892_, data_stage_2__3891_, data_stage_2__3890_, data_stage_2__3889_, data_stage_2__3888_, data_stage_2__3887_, data_stage_2__3886_, data_stage_2__3885_, data_stage_2__3884_, data_stage_2__3883_, data_stage_2__3882_, data_stage_2__3881_, data_stage_2__3880_, data_stage_2__3879_, data_stage_2__3878_, data_stage_2__3877_, data_stage_2__3876_, data_stage_2__3875_, data_stage_2__3874_, data_stage_2__3873_, data_stage_2__3872_, data_stage_2__3871_, data_stage_2__3870_, data_stage_2__3869_, data_stage_2__3868_, data_stage_2__3867_, data_stage_2__3866_, data_stage_2__3865_, data_stage_2__3864_, data_stage_2__3863_, data_stage_2__3862_, data_stage_2__3861_, data_stage_2__3860_, data_stage_2__3859_, data_stage_2__3858_, data_stage_2__3857_, data_stage_2__3856_, data_stage_2__3855_, data_stage_2__3854_, data_stage_2__3853_, data_stage_2__3852_, data_stage_2__3851_, data_stage_2__3850_, data_stage_2__3849_, data_stage_2__3848_, data_stage_2__3847_, data_stage_2__3846_, data_stage_2__3845_, data_stage_2__3844_, data_stage_2__3843_, data_stage_2__3842_, data_stage_2__3841_, data_stage_2__3840_, data_stage_2__3839_, data_stage_2__3838_, data_stage_2__3837_, data_stage_2__3836_, data_stage_2__3835_, data_stage_2__3834_, data_stage_2__3833_, data_stage_2__3832_, data_stage_2__3831_, data_stage_2__3830_, data_stage_2__3829_, data_stage_2__3828_, data_stage_2__3827_, data_stage_2__3826_, data_stage_2__3825_, data_stage_2__3824_, data_stage_2__3823_, data_stage_2__3822_, data_stage_2__3821_, data_stage_2__3820_, data_stage_2__3819_, data_stage_2__3818_, data_stage_2__3817_, data_stage_2__3816_, data_stage_2__3815_, data_stage_2__3814_, data_stage_2__3813_, data_stage_2__3812_, data_stage_2__3811_, data_stage_2__3810_, data_stage_2__3809_, data_stage_2__3808_, data_stage_2__3807_, data_stage_2__3806_, data_stage_2__3805_, data_stage_2__3804_, data_stage_2__3803_, data_stage_2__3802_, data_stage_2__3801_, data_stage_2__3800_, data_stage_2__3799_, data_stage_2__3798_, data_stage_2__3797_, data_stage_2__3796_, data_stage_2__3795_, data_stage_2__3794_, data_stage_2__3793_, data_stage_2__3792_, data_stage_2__3791_, data_stage_2__3790_, data_stage_2__3789_, data_stage_2__3788_, data_stage_2__3787_, data_stage_2__3786_, data_stage_2__3785_, data_stage_2__3784_, data_stage_2__3783_, data_stage_2__3782_, data_stage_2__3781_, data_stage_2__3780_, data_stage_2__3779_, data_stage_2__3778_, data_stage_2__3777_, data_stage_2__3776_, data_stage_2__3775_, data_stage_2__3774_, data_stage_2__3773_, data_stage_2__3772_, data_stage_2__3771_, data_stage_2__3770_, data_stage_2__3769_, data_stage_2__3768_, data_stage_2__3767_, data_stage_2__3766_, data_stage_2__3765_, data_stage_2__3764_, data_stage_2__3763_, data_stage_2__3762_, data_stage_2__3761_, data_stage_2__3760_, data_stage_2__3759_, data_stage_2__3758_, data_stage_2__3757_, data_stage_2__3756_, data_stage_2__3755_, data_stage_2__3754_, data_stage_2__3753_, data_stage_2__3752_, data_stage_2__3751_, data_stage_2__3750_, data_stage_2__3749_, data_stage_2__3748_, data_stage_2__3747_, data_stage_2__3746_, data_stage_2__3745_, data_stage_2__3744_, data_stage_2__3743_, data_stage_2__3742_, data_stage_2__3741_, data_stage_2__3740_, data_stage_2__3739_, data_stage_2__3738_, data_stage_2__3737_, data_stage_2__3736_, data_stage_2__3735_, data_stage_2__3734_, data_stage_2__3733_, data_stage_2__3732_, data_stage_2__3731_, data_stage_2__3730_, data_stage_2__3729_, data_stage_2__3728_, data_stage_2__3727_, data_stage_2__3726_, data_stage_2__3725_, data_stage_2__3724_, data_stage_2__3723_, data_stage_2__3722_, data_stage_2__3721_, data_stage_2__3720_, data_stage_2__3719_, data_stage_2__3718_, data_stage_2__3717_, data_stage_2__3716_, data_stage_2__3715_, data_stage_2__3714_, data_stage_2__3713_, data_stage_2__3712_, data_stage_2__3711_, data_stage_2__3710_, data_stage_2__3709_, data_stage_2__3708_, data_stage_2__3707_, data_stage_2__3706_, data_stage_2__3705_, data_stage_2__3704_, data_stage_2__3703_, data_stage_2__3702_, data_stage_2__3701_, data_stage_2__3700_, data_stage_2__3699_, data_stage_2__3698_, data_stage_2__3697_, data_stage_2__3696_, data_stage_2__3695_, data_stage_2__3694_, data_stage_2__3693_, data_stage_2__3692_, data_stage_2__3691_, data_stage_2__3690_, data_stage_2__3689_, data_stage_2__3688_, data_stage_2__3687_, data_stage_2__3686_, data_stage_2__3685_, data_stage_2__3684_, data_stage_2__3683_, data_stage_2__3682_, data_stage_2__3681_, data_stage_2__3680_, data_stage_2__3679_, data_stage_2__3678_, data_stage_2__3677_, data_stage_2__3676_, data_stage_2__3675_, data_stage_2__3674_, data_stage_2__3673_, data_stage_2__3672_, data_stage_2__3671_, data_stage_2__3670_, data_stage_2__3669_, data_stage_2__3668_, data_stage_2__3667_, data_stage_2__3666_, data_stage_2__3665_, data_stage_2__3664_, data_stage_2__3663_, data_stage_2__3662_, data_stage_2__3661_, data_stage_2__3660_, data_stage_2__3659_, data_stage_2__3658_, data_stage_2__3657_, data_stage_2__3656_, data_stage_2__3655_, data_stage_2__3654_, data_stage_2__3653_, data_stage_2__3652_, data_stage_2__3651_, data_stage_2__3650_, data_stage_2__3649_, data_stage_2__3648_, data_stage_2__3647_, data_stage_2__3646_, data_stage_2__3645_, data_stage_2__3644_, data_stage_2__3643_, data_stage_2__3642_, data_stage_2__3641_, data_stage_2__3640_, data_stage_2__3639_, data_stage_2__3638_, data_stage_2__3637_, data_stage_2__3636_, data_stage_2__3635_, data_stage_2__3634_, data_stage_2__3633_, data_stage_2__3632_, data_stage_2__3631_, data_stage_2__3630_, data_stage_2__3629_, data_stage_2__3628_, data_stage_2__3627_, data_stage_2__3626_, data_stage_2__3625_, data_stage_2__3624_, data_stage_2__3623_, data_stage_2__3622_, data_stage_2__3621_, data_stage_2__3620_, data_stage_2__3619_, data_stage_2__3618_, data_stage_2__3617_, data_stage_2__3616_, data_stage_2__3615_, data_stage_2__3614_, data_stage_2__3613_, data_stage_2__3612_, data_stage_2__3611_, data_stage_2__3610_, data_stage_2__3609_, data_stage_2__3608_, data_stage_2__3607_, data_stage_2__3606_, data_stage_2__3605_, data_stage_2__3604_, data_stage_2__3603_, data_stage_2__3602_, data_stage_2__3601_, data_stage_2__3600_, data_stage_2__3599_, data_stage_2__3598_, data_stage_2__3597_, data_stage_2__3596_, data_stage_2__3595_, data_stage_2__3594_, data_stage_2__3593_, data_stage_2__3592_, data_stage_2__3591_, data_stage_2__3590_, data_stage_2__3589_, data_stage_2__3588_, data_stage_2__3587_, data_stage_2__3586_, data_stage_2__3585_, data_stage_2__3584_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__4095_, data_stage_3__4094_, data_stage_3__4093_, data_stage_3__4092_, data_stage_3__4091_, data_stage_3__4090_, data_stage_3__4089_, data_stage_3__4088_, data_stage_3__4087_, data_stage_3__4086_, data_stage_3__4085_, data_stage_3__4084_, data_stage_3__4083_, data_stage_3__4082_, data_stage_3__4081_, data_stage_3__4080_, data_stage_3__4079_, data_stage_3__4078_, data_stage_3__4077_, data_stage_3__4076_, data_stage_3__4075_, data_stage_3__4074_, data_stage_3__4073_, data_stage_3__4072_, data_stage_3__4071_, data_stage_3__4070_, data_stage_3__4069_, data_stage_3__4068_, data_stage_3__4067_, data_stage_3__4066_, data_stage_3__4065_, data_stage_3__4064_, data_stage_3__4063_, data_stage_3__4062_, data_stage_3__4061_, data_stage_3__4060_, data_stage_3__4059_, data_stage_3__4058_, data_stage_3__4057_, data_stage_3__4056_, data_stage_3__4055_, data_stage_3__4054_, data_stage_3__4053_, data_stage_3__4052_, data_stage_3__4051_, data_stage_3__4050_, data_stage_3__4049_, data_stage_3__4048_, data_stage_3__4047_, data_stage_3__4046_, data_stage_3__4045_, data_stage_3__4044_, data_stage_3__4043_, data_stage_3__4042_, data_stage_3__4041_, data_stage_3__4040_, data_stage_3__4039_, data_stage_3__4038_, data_stage_3__4037_, data_stage_3__4036_, data_stage_3__4035_, data_stage_3__4034_, data_stage_3__4033_, data_stage_3__4032_, data_stage_3__4031_, data_stage_3__4030_, data_stage_3__4029_, data_stage_3__4028_, data_stage_3__4027_, data_stage_3__4026_, data_stage_3__4025_, data_stage_3__4024_, data_stage_3__4023_, data_stage_3__4022_, data_stage_3__4021_, data_stage_3__4020_, data_stage_3__4019_, data_stage_3__4018_, data_stage_3__4017_, data_stage_3__4016_, data_stage_3__4015_, data_stage_3__4014_, data_stage_3__4013_, data_stage_3__4012_, data_stage_3__4011_, data_stage_3__4010_, data_stage_3__4009_, data_stage_3__4008_, data_stage_3__4007_, data_stage_3__4006_, data_stage_3__4005_, data_stage_3__4004_, data_stage_3__4003_, data_stage_3__4002_, data_stage_3__4001_, data_stage_3__4000_, data_stage_3__3999_, data_stage_3__3998_, data_stage_3__3997_, data_stage_3__3996_, data_stage_3__3995_, data_stage_3__3994_, data_stage_3__3993_, data_stage_3__3992_, data_stage_3__3991_, data_stage_3__3990_, data_stage_3__3989_, data_stage_3__3988_, data_stage_3__3987_, data_stage_3__3986_, data_stage_3__3985_, data_stage_3__3984_, data_stage_3__3983_, data_stage_3__3982_, data_stage_3__3981_, data_stage_3__3980_, data_stage_3__3979_, data_stage_3__3978_, data_stage_3__3977_, data_stage_3__3976_, data_stage_3__3975_, data_stage_3__3974_, data_stage_3__3973_, data_stage_3__3972_, data_stage_3__3971_, data_stage_3__3970_, data_stage_3__3969_, data_stage_3__3968_, data_stage_3__3967_, data_stage_3__3966_, data_stage_3__3965_, data_stage_3__3964_, data_stage_3__3963_, data_stage_3__3962_, data_stage_3__3961_, data_stage_3__3960_, data_stage_3__3959_, data_stage_3__3958_, data_stage_3__3957_, data_stage_3__3956_, data_stage_3__3955_, data_stage_3__3954_, data_stage_3__3953_, data_stage_3__3952_, data_stage_3__3951_, data_stage_3__3950_, data_stage_3__3949_, data_stage_3__3948_, data_stage_3__3947_, data_stage_3__3946_, data_stage_3__3945_, data_stage_3__3944_, data_stage_3__3943_, data_stage_3__3942_, data_stage_3__3941_, data_stage_3__3940_, data_stage_3__3939_, data_stage_3__3938_, data_stage_3__3937_, data_stage_3__3936_, data_stage_3__3935_, data_stage_3__3934_, data_stage_3__3933_, data_stage_3__3932_, data_stage_3__3931_, data_stage_3__3930_, data_stage_3__3929_, data_stage_3__3928_, data_stage_3__3927_, data_stage_3__3926_, data_stage_3__3925_, data_stage_3__3924_, data_stage_3__3923_, data_stage_3__3922_, data_stage_3__3921_, data_stage_3__3920_, data_stage_3__3919_, data_stage_3__3918_, data_stage_3__3917_, data_stage_3__3916_, data_stage_3__3915_, data_stage_3__3914_, data_stage_3__3913_, data_stage_3__3912_, data_stage_3__3911_, data_stage_3__3910_, data_stage_3__3909_, data_stage_3__3908_, data_stage_3__3907_, data_stage_3__3906_, data_stage_3__3905_, data_stage_3__3904_, data_stage_3__3903_, data_stage_3__3902_, data_stage_3__3901_, data_stage_3__3900_, data_stage_3__3899_, data_stage_3__3898_, data_stage_3__3897_, data_stage_3__3896_, data_stage_3__3895_, data_stage_3__3894_, data_stage_3__3893_, data_stage_3__3892_, data_stage_3__3891_, data_stage_3__3890_, data_stage_3__3889_, data_stage_3__3888_, data_stage_3__3887_, data_stage_3__3886_, data_stage_3__3885_, data_stage_3__3884_, data_stage_3__3883_, data_stage_3__3882_, data_stage_3__3881_, data_stage_3__3880_, data_stage_3__3879_, data_stage_3__3878_, data_stage_3__3877_, data_stage_3__3876_, data_stage_3__3875_, data_stage_3__3874_, data_stage_3__3873_, data_stage_3__3872_, data_stage_3__3871_, data_stage_3__3870_, data_stage_3__3869_, data_stage_3__3868_, data_stage_3__3867_, data_stage_3__3866_, data_stage_3__3865_, data_stage_3__3864_, data_stage_3__3863_, data_stage_3__3862_, data_stage_3__3861_, data_stage_3__3860_, data_stage_3__3859_, data_stage_3__3858_, data_stage_3__3857_, data_stage_3__3856_, data_stage_3__3855_, data_stage_3__3854_, data_stage_3__3853_, data_stage_3__3852_, data_stage_3__3851_, data_stage_3__3850_, data_stage_3__3849_, data_stage_3__3848_, data_stage_3__3847_, data_stage_3__3846_, data_stage_3__3845_, data_stage_3__3844_, data_stage_3__3843_, data_stage_3__3842_, data_stage_3__3841_, data_stage_3__3840_, data_stage_3__3839_, data_stage_3__3838_, data_stage_3__3837_, data_stage_3__3836_, data_stage_3__3835_, data_stage_3__3834_, data_stage_3__3833_, data_stage_3__3832_, data_stage_3__3831_, data_stage_3__3830_, data_stage_3__3829_, data_stage_3__3828_, data_stage_3__3827_, data_stage_3__3826_, data_stage_3__3825_, data_stage_3__3824_, data_stage_3__3823_, data_stage_3__3822_, data_stage_3__3821_, data_stage_3__3820_, data_stage_3__3819_, data_stage_3__3818_, data_stage_3__3817_, data_stage_3__3816_, data_stage_3__3815_, data_stage_3__3814_, data_stage_3__3813_, data_stage_3__3812_, data_stage_3__3811_, data_stage_3__3810_, data_stage_3__3809_, data_stage_3__3808_, data_stage_3__3807_, data_stage_3__3806_, data_stage_3__3805_, data_stage_3__3804_, data_stage_3__3803_, data_stage_3__3802_, data_stage_3__3801_, data_stage_3__3800_, data_stage_3__3799_, data_stage_3__3798_, data_stage_3__3797_, data_stage_3__3796_, data_stage_3__3795_, data_stage_3__3794_, data_stage_3__3793_, data_stage_3__3792_, data_stage_3__3791_, data_stage_3__3790_, data_stage_3__3789_, data_stage_3__3788_, data_stage_3__3787_, data_stage_3__3786_, data_stage_3__3785_, data_stage_3__3784_, data_stage_3__3783_, data_stage_3__3782_, data_stage_3__3781_, data_stage_3__3780_, data_stage_3__3779_, data_stage_3__3778_, data_stage_3__3777_, data_stage_3__3776_, data_stage_3__3775_, data_stage_3__3774_, data_stage_3__3773_, data_stage_3__3772_, data_stage_3__3771_, data_stage_3__3770_, data_stage_3__3769_, data_stage_3__3768_, data_stage_3__3767_, data_stage_3__3766_, data_stage_3__3765_, data_stage_3__3764_, data_stage_3__3763_, data_stage_3__3762_, data_stage_3__3761_, data_stage_3__3760_, data_stage_3__3759_, data_stage_3__3758_, data_stage_3__3757_, data_stage_3__3756_, data_stage_3__3755_, data_stage_3__3754_, data_stage_3__3753_, data_stage_3__3752_, data_stage_3__3751_, data_stage_3__3750_, data_stage_3__3749_, data_stage_3__3748_, data_stage_3__3747_, data_stage_3__3746_, data_stage_3__3745_, data_stage_3__3744_, data_stage_3__3743_, data_stage_3__3742_, data_stage_3__3741_, data_stage_3__3740_, data_stage_3__3739_, data_stage_3__3738_, data_stage_3__3737_, data_stage_3__3736_, data_stage_3__3735_, data_stage_3__3734_, data_stage_3__3733_, data_stage_3__3732_, data_stage_3__3731_, data_stage_3__3730_, data_stage_3__3729_, data_stage_3__3728_, data_stage_3__3727_, data_stage_3__3726_, data_stage_3__3725_, data_stage_3__3724_, data_stage_3__3723_, data_stage_3__3722_, data_stage_3__3721_, data_stage_3__3720_, data_stage_3__3719_, data_stage_3__3718_, data_stage_3__3717_, data_stage_3__3716_, data_stage_3__3715_, data_stage_3__3714_, data_stage_3__3713_, data_stage_3__3712_, data_stage_3__3711_, data_stage_3__3710_, data_stage_3__3709_, data_stage_3__3708_, data_stage_3__3707_, data_stage_3__3706_, data_stage_3__3705_, data_stage_3__3704_, data_stage_3__3703_, data_stage_3__3702_, data_stage_3__3701_, data_stage_3__3700_, data_stage_3__3699_, data_stage_3__3698_, data_stage_3__3697_, data_stage_3__3696_, data_stage_3__3695_, data_stage_3__3694_, data_stage_3__3693_, data_stage_3__3692_, data_stage_3__3691_, data_stage_3__3690_, data_stage_3__3689_, data_stage_3__3688_, data_stage_3__3687_, data_stage_3__3686_, data_stage_3__3685_, data_stage_3__3684_, data_stage_3__3683_, data_stage_3__3682_, data_stage_3__3681_, data_stage_3__3680_, data_stage_3__3679_, data_stage_3__3678_, data_stage_3__3677_, data_stage_3__3676_, data_stage_3__3675_, data_stage_3__3674_, data_stage_3__3673_, data_stage_3__3672_, data_stage_3__3671_, data_stage_3__3670_, data_stage_3__3669_, data_stage_3__3668_, data_stage_3__3667_, data_stage_3__3666_, data_stage_3__3665_, data_stage_3__3664_, data_stage_3__3663_, data_stage_3__3662_, data_stage_3__3661_, data_stage_3__3660_, data_stage_3__3659_, data_stage_3__3658_, data_stage_3__3657_, data_stage_3__3656_, data_stage_3__3655_, data_stage_3__3654_, data_stage_3__3653_, data_stage_3__3652_, data_stage_3__3651_, data_stage_3__3650_, data_stage_3__3649_, data_stage_3__3648_, data_stage_3__3647_, data_stage_3__3646_, data_stage_3__3645_, data_stage_3__3644_, data_stage_3__3643_, data_stage_3__3642_, data_stage_3__3641_, data_stage_3__3640_, data_stage_3__3639_, data_stage_3__3638_, data_stage_3__3637_, data_stage_3__3636_, data_stage_3__3635_, data_stage_3__3634_, data_stage_3__3633_, data_stage_3__3632_, data_stage_3__3631_, data_stage_3__3630_, data_stage_3__3629_, data_stage_3__3628_, data_stage_3__3627_, data_stage_3__3626_, data_stage_3__3625_, data_stage_3__3624_, data_stage_3__3623_, data_stage_3__3622_, data_stage_3__3621_, data_stage_3__3620_, data_stage_3__3619_, data_stage_3__3618_, data_stage_3__3617_, data_stage_3__3616_, data_stage_3__3615_, data_stage_3__3614_, data_stage_3__3613_, data_stage_3__3612_, data_stage_3__3611_, data_stage_3__3610_, data_stage_3__3609_, data_stage_3__3608_, data_stage_3__3607_, data_stage_3__3606_, data_stage_3__3605_, data_stage_3__3604_, data_stage_3__3603_, data_stage_3__3602_, data_stage_3__3601_, data_stage_3__3600_, data_stage_3__3599_, data_stage_3__3598_, data_stage_3__3597_, data_stage_3__3596_, data_stage_3__3595_, data_stage_3__3594_, data_stage_3__3593_, data_stage_3__3592_, data_stage_3__3591_, data_stage_3__3590_, data_stage_3__3589_, data_stage_3__3588_, data_stage_3__3587_, data_stage_3__3586_, data_stage_3__3585_, data_stage_3__3584_ })
  );


  bsg_swap_width_p512
  mux_stage_3__mux_swap_0__swap_inst
  (
    .data_i({ data_stage_3__1023_, data_stage_3__1022_, data_stage_3__1021_, data_stage_3__1020_, data_stage_3__1019_, data_stage_3__1018_, data_stage_3__1017_, data_stage_3__1016_, data_stage_3__1015_, data_stage_3__1014_, data_stage_3__1013_, data_stage_3__1012_, data_stage_3__1011_, data_stage_3__1010_, data_stage_3__1009_, data_stage_3__1008_, data_stage_3__1007_, data_stage_3__1006_, data_stage_3__1005_, data_stage_3__1004_, data_stage_3__1003_, data_stage_3__1002_, data_stage_3__1001_, data_stage_3__1000_, data_stage_3__999_, data_stage_3__998_, data_stage_3__997_, data_stage_3__996_, data_stage_3__995_, data_stage_3__994_, data_stage_3__993_, data_stage_3__992_, data_stage_3__991_, data_stage_3__990_, data_stage_3__989_, data_stage_3__988_, data_stage_3__987_, data_stage_3__986_, data_stage_3__985_, data_stage_3__984_, data_stage_3__983_, data_stage_3__982_, data_stage_3__981_, data_stage_3__980_, data_stage_3__979_, data_stage_3__978_, data_stage_3__977_, data_stage_3__976_, data_stage_3__975_, data_stage_3__974_, data_stage_3__973_, data_stage_3__972_, data_stage_3__971_, data_stage_3__970_, data_stage_3__969_, data_stage_3__968_, data_stage_3__967_, data_stage_3__966_, data_stage_3__965_, data_stage_3__964_, data_stage_3__963_, data_stage_3__962_, data_stage_3__961_, data_stage_3__960_, data_stage_3__959_, data_stage_3__958_, data_stage_3__957_, data_stage_3__956_, data_stage_3__955_, data_stage_3__954_, data_stage_3__953_, data_stage_3__952_, data_stage_3__951_, data_stage_3__950_, data_stage_3__949_, data_stage_3__948_, data_stage_3__947_, data_stage_3__946_, data_stage_3__945_, data_stage_3__944_, data_stage_3__943_, data_stage_3__942_, data_stage_3__941_, data_stage_3__940_, data_stage_3__939_, data_stage_3__938_, data_stage_3__937_, data_stage_3__936_, data_stage_3__935_, data_stage_3__934_, data_stage_3__933_, data_stage_3__932_, data_stage_3__931_, data_stage_3__930_, data_stage_3__929_, data_stage_3__928_, data_stage_3__927_, data_stage_3__926_, data_stage_3__925_, data_stage_3__924_, data_stage_3__923_, data_stage_3__922_, data_stage_3__921_, data_stage_3__920_, data_stage_3__919_, data_stage_3__918_, data_stage_3__917_, data_stage_3__916_, data_stage_3__915_, data_stage_3__914_, data_stage_3__913_, data_stage_3__912_, data_stage_3__911_, data_stage_3__910_, data_stage_3__909_, data_stage_3__908_, data_stage_3__907_, data_stage_3__906_, data_stage_3__905_, data_stage_3__904_, data_stage_3__903_, data_stage_3__902_, data_stage_3__901_, data_stage_3__900_, data_stage_3__899_, data_stage_3__898_, data_stage_3__897_, data_stage_3__896_, data_stage_3__895_, data_stage_3__894_, data_stage_3__893_, data_stage_3__892_, data_stage_3__891_, data_stage_3__890_, data_stage_3__889_, data_stage_3__888_, data_stage_3__887_, data_stage_3__886_, data_stage_3__885_, data_stage_3__884_, data_stage_3__883_, data_stage_3__882_, data_stage_3__881_, data_stage_3__880_, data_stage_3__879_, data_stage_3__878_, data_stage_3__877_, data_stage_3__876_, data_stage_3__875_, data_stage_3__874_, data_stage_3__873_, data_stage_3__872_, data_stage_3__871_, data_stage_3__870_, data_stage_3__869_, data_stage_3__868_, data_stage_3__867_, data_stage_3__866_, data_stage_3__865_, data_stage_3__864_, data_stage_3__863_, data_stage_3__862_, data_stage_3__861_, data_stage_3__860_, data_stage_3__859_, data_stage_3__858_, data_stage_3__857_, data_stage_3__856_, data_stage_3__855_, data_stage_3__854_, data_stage_3__853_, data_stage_3__852_, data_stage_3__851_, data_stage_3__850_, data_stage_3__849_, data_stage_3__848_, data_stage_3__847_, data_stage_3__846_, data_stage_3__845_, data_stage_3__844_, data_stage_3__843_, data_stage_3__842_, data_stage_3__841_, data_stage_3__840_, data_stage_3__839_, data_stage_3__838_, data_stage_3__837_, data_stage_3__836_, data_stage_3__835_, data_stage_3__834_, data_stage_3__833_, data_stage_3__832_, data_stage_3__831_, data_stage_3__830_, data_stage_3__829_, data_stage_3__828_, data_stage_3__827_, data_stage_3__826_, data_stage_3__825_, data_stage_3__824_, data_stage_3__823_, data_stage_3__822_, data_stage_3__821_, data_stage_3__820_, data_stage_3__819_, data_stage_3__818_, data_stage_3__817_, data_stage_3__816_, data_stage_3__815_, data_stage_3__814_, data_stage_3__813_, data_stage_3__812_, data_stage_3__811_, data_stage_3__810_, data_stage_3__809_, data_stage_3__808_, data_stage_3__807_, data_stage_3__806_, data_stage_3__805_, data_stage_3__804_, data_stage_3__803_, data_stage_3__802_, data_stage_3__801_, data_stage_3__800_, data_stage_3__799_, data_stage_3__798_, data_stage_3__797_, data_stage_3__796_, data_stage_3__795_, data_stage_3__794_, data_stage_3__793_, data_stage_3__792_, data_stage_3__791_, data_stage_3__790_, data_stage_3__789_, data_stage_3__788_, data_stage_3__787_, data_stage_3__786_, data_stage_3__785_, data_stage_3__784_, data_stage_3__783_, data_stage_3__782_, data_stage_3__781_, data_stage_3__780_, data_stage_3__779_, data_stage_3__778_, data_stage_3__777_, data_stage_3__776_, data_stage_3__775_, data_stage_3__774_, data_stage_3__773_, data_stage_3__772_, data_stage_3__771_, data_stage_3__770_, data_stage_3__769_, data_stage_3__768_, data_stage_3__767_, data_stage_3__766_, data_stage_3__765_, data_stage_3__764_, data_stage_3__763_, data_stage_3__762_, data_stage_3__761_, data_stage_3__760_, data_stage_3__759_, data_stage_3__758_, data_stage_3__757_, data_stage_3__756_, data_stage_3__755_, data_stage_3__754_, data_stage_3__753_, data_stage_3__752_, data_stage_3__751_, data_stage_3__750_, data_stage_3__749_, data_stage_3__748_, data_stage_3__747_, data_stage_3__746_, data_stage_3__745_, data_stage_3__744_, data_stage_3__743_, data_stage_3__742_, data_stage_3__741_, data_stage_3__740_, data_stage_3__739_, data_stage_3__738_, data_stage_3__737_, data_stage_3__736_, data_stage_3__735_, data_stage_3__734_, data_stage_3__733_, data_stage_3__732_, data_stage_3__731_, data_stage_3__730_, data_stage_3__729_, data_stage_3__728_, data_stage_3__727_, data_stage_3__726_, data_stage_3__725_, data_stage_3__724_, data_stage_3__723_, data_stage_3__722_, data_stage_3__721_, data_stage_3__720_, data_stage_3__719_, data_stage_3__718_, data_stage_3__717_, data_stage_3__716_, data_stage_3__715_, data_stage_3__714_, data_stage_3__713_, data_stage_3__712_, data_stage_3__711_, data_stage_3__710_, data_stage_3__709_, data_stage_3__708_, data_stage_3__707_, data_stage_3__706_, data_stage_3__705_, data_stage_3__704_, data_stage_3__703_, data_stage_3__702_, data_stage_3__701_, data_stage_3__700_, data_stage_3__699_, data_stage_3__698_, data_stage_3__697_, data_stage_3__696_, data_stage_3__695_, data_stage_3__694_, data_stage_3__693_, data_stage_3__692_, data_stage_3__691_, data_stage_3__690_, data_stage_3__689_, data_stage_3__688_, data_stage_3__687_, data_stage_3__686_, data_stage_3__685_, data_stage_3__684_, data_stage_3__683_, data_stage_3__682_, data_stage_3__681_, data_stage_3__680_, data_stage_3__679_, data_stage_3__678_, data_stage_3__677_, data_stage_3__676_, data_stage_3__675_, data_stage_3__674_, data_stage_3__673_, data_stage_3__672_, data_stage_3__671_, data_stage_3__670_, data_stage_3__669_, data_stage_3__668_, data_stage_3__667_, data_stage_3__666_, data_stage_3__665_, data_stage_3__664_, data_stage_3__663_, data_stage_3__662_, data_stage_3__661_, data_stage_3__660_, data_stage_3__659_, data_stage_3__658_, data_stage_3__657_, data_stage_3__656_, data_stage_3__655_, data_stage_3__654_, data_stage_3__653_, data_stage_3__652_, data_stage_3__651_, data_stage_3__650_, data_stage_3__649_, data_stage_3__648_, data_stage_3__647_, data_stage_3__646_, data_stage_3__645_, data_stage_3__644_, data_stage_3__643_, data_stage_3__642_, data_stage_3__641_, data_stage_3__640_, data_stage_3__639_, data_stage_3__638_, data_stage_3__637_, data_stage_3__636_, data_stage_3__635_, data_stage_3__634_, data_stage_3__633_, data_stage_3__632_, data_stage_3__631_, data_stage_3__630_, data_stage_3__629_, data_stage_3__628_, data_stage_3__627_, data_stage_3__626_, data_stage_3__625_, data_stage_3__624_, data_stage_3__623_, data_stage_3__622_, data_stage_3__621_, data_stage_3__620_, data_stage_3__619_, data_stage_3__618_, data_stage_3__617_, data_stage_3__616_, data_stage_3__615_, data_stage_3__614_, data_stage_3__613_, data_stage_3__612_, data_stage_3__611_, data_stage_3__610_, data_stage_3__609_, data_stage_3__608_, data_stage_3__607_, data_stage_3__606_, data_stage_3__605_, data_stage_3__604_, data_stage_3__603_, data_stage_3__602_, data_stage_3__601_, data_stage_3__600_, data_stage_3__599_, data_stage_3__598_, data_stage_3__597_, data_stage_3__596_, data_stage_3__595_, data_stage_3__594_, data_stage_3__593_, data_stage_3__592_, data_stage_3__591_, data_stage_3__590_, data_stage_3__589_, data_stage_3__588_, data_stage_3__587_, data_stage_3__586_, data_stage_3__585_, data_stage_3__584_, data_stage_3__583_, data_stage_3__582_, data_stage_3__581_, data_stage_3__580_, data_stage_3__579_, data_stage_3__578_, data_stage_3__577_, data_stage_3__576_, data_stage_3__575_, data_stage_3__574_, data_stage_3__573_, data_stage_3__572_, data_stage_3__571_, data_stage_3__570_, data_stage_3__569_, data_stage_3__568_, data_stage_3__567_, data_stage_3__566_, data_stage_3__565_, data_stage_3__564_, data_stage_3__563_, data_stage_3__562_, data_stage_3__561_, data_stage_3__560_, data_stage_3__559_, data_stage_3__558_, data_stage_3__557_, data_stage_3__556_, data_stage_3__555_, data_stage_3__554_, data_stage_3__553_, data_stage_3__552_, data_stage_3__551_, data_stage_3__550_, data_stage_3__549_, data_stage_3__548_, data_stage_3__547_, data_stage_3__546_, data_stage_3__545_, data_stage_3__544_, data_stage_3__543_, data_stage_3__542_, data_stage_3__541_, data_stage_3__540_, data_stage_3__539_, data_stage_3__538_, data_stage_3__537_, data_stage_3__536_, data_stage_3__535_, data_stage_3__534_, data_stage_3__533_, data_stage_3__532_, data_stage_3__531_, data_stage_3__530_, data_stage_3__529_, data_stage_3__528_, data_stage_3__527_, data_stage_3__526_, data_stage_3__525_, data_stage_3__524_, data_stage_3__523_, data_stage_3__522_, data_stage_3__521_, data_stage_3__520_, data_stage_3__519_, data_stage_3__518_, data_stage_3__517_, data_stage_3__516_, data_stage_3__515_, data_stage_3__514_, data_stage_3__513_, data_stage_3__512_, data_stage_3__511_, data_stage_3__510_, data_stage_3__509_, data_stage_3__508_, data_stage_3__507_, data_stage_3__506_, data_stage_3__505_, data_stage_3__504_, data_stage_3__503_, data_stage_3__502_, data_stage_3__501_, data_stage_3__500_, data_stage_3__499_, data_stage_3__498_, data_stage_3__497_, data_stage_3__496_, data_stage_3__495_, data_stage_3__494_, data_stage_3__493_, data_stage_3__492_, data_stage_3__491_, data_stage_3__490_, data_stage_3__489_, data_stage_3__488_, data_stage_3__487_, data_stage_3__486_, data_stage_3__485_, data_stage_3__484_, data_stage_3__483_, data_stage_3__482_, data_stage_3__481_, data_stage_3__480_, data_stage_3__479_, data_stage_3__478_, data_stage_3__477_, data_stage_3__476_, data_stage_3__475_, data_stage_3__474_, data_stage_3__473_, data_stage_3__472_, data_stage_3__471_, data_stage_3__470_, data_stage_3__469_, data_stage_3__468_, data_stage_3__467_, data_stage_3__466_, data_stage_3__465_, data_stage_3__464_, data_stage_3__463_, data_stage_3__462_, data_stage_3__461_, data_stage_3__460_, data_stage_3__459_, data_stage_3__458_, data_stage_3__457_, data_stage_3__456_, data_stage_3__455_, data_stage_3__454_, data_stage_3__453_, data_stage_3__452_, data_stage_3__451_, data_stage_3__450_, data_stage_3__449_, data_stage_3__448_, data_stage_3__447_, data_stage_3__446_, data_stage_3__445_, data_stage_3__444_, data_stage_3__443_, data_stage_3__442_, data_stage_3__441_, data_stage_3__440_, data_stage_3__439_, data_stage_3__438_, data_stage_3__437_, data_stage_3__436_, data_stage_3__435_, data_stage_3__434_, data_stage_3__433_, data_stage_3__432_, data_stage_3__431_, data_stage_3__430_, data_stage_3__429_, data_stage_3__428_, data_stage_3__427_, data_stage_3__426_, data_stage_3__425_, data_stage_3__424_, data_stage_3__423_, data_stage_3__422_, data_stage_3__421_, data_stage_3__420_, data_stage_3__419_, data_stage_3__418_, data_stage_3__417_, data_stage_3__416_, data_stage_3__415_, data_stage_3__414_, data_stage_3__413_, data_stage_3__412_, data_stage_3__411_, data_stage_3__410_, data_stage_3__409_, data_stage_3__408_, data_stage_3__407_, data_stage_3__406_, data_stage_3__405_, data_stage_3__404_, data_stage_3__403_, data_stage_3__402_, data_stage_3__401_, data_stage_3__400_, data_stage_3__399_, data_stage_3__398_, data_stage_3__397_, data_stage_3__396_, data_stage_3__395_, data_stage_3__394_, data_stage_3__393_, data_stage_3__392_, data_stage_3__391_, data_stage_3__390_, data_stage_3__389_, data_stage_3__388_, data_stage_3__387_, data_stage_3__386_, data_stage_3__385_, data_stage_3__384_, data_stage_3__383_, data_stage_3__382_, data_stage_3__381_, data_stage_3__380_, data_stage_3__379_, data_stage_3__378_, data_stage_3__377_, data_stage_3__376_, data_stage_3__375_, data_stage_3__374_, data_stage_3__373_, data_stage_3__372_, data_stage_3__371_, data_stage_3__370_, data_stage_3__369_, data_stage_3__368_, data_stage_3__367_, data_stage_3__366_, data_stage_3__365_, data_stage_3__364_, data_stage_3__363_, data_stage_3__362_, data_stage_3__361_, data_stage_3__360_, data_stage_3__359_, data_stage_3__358_, data_stage_3__357_, data_stage_3__356_, data_stage_3__355_, data_stage_3__354_, data_stage_3__353_, data_stage_3__352_, data_stage_3__351_, data_stage_3__350_, data_stage_3__349_, data_stage_3__348_, data_stage_3__347_, data_stage_3__346_, data_stage_3__345_, data_stage_3__344_, data_stage_3__343_, data_stage_3__342_, data_stage_3__341_, data_stage_3__340_, data_stage_3__339_, data_stage_3__338_, data_stage_3__337_, data_stage_3__336_, data_stage_3__335_, data_stage_3__334_, data_stage_3__333_, data_stage_3__332_, data_stage_3__331_, data_stage_3__330_, data_stage_3__329_, data_stage_3__328_, data_stage_3__327_, data_stage_3__326_, data_stage_3__325_, data_stage_3__324_, data_stage_3__323_, data_stage_3__322_, data_stage_3__321_, data_stage_3__320_, data_stage_3__319_, data_stage_3__318_, data_stage_3__317_, data_stage_3__316_, data_stage_3__315_, data_stage_3__314_, data_stage_3__313_, data_stage_3__312_, data_stage_3__311_, data_stage_3__310_, data_stage_3__309_, data_stage_3__308_, data_stage_3__307_, data_stage_3__306_, data_stage_3__305_, data_stage_3__304_, data_stage_3__303_, data_stage_3__302_, data_stage_3__301_, data_stage_3__300_, data_stage_3__299_, data_stage_3__298_, data_stage_3__297_, data_stage_3__296_, data_stage_3__295_, data_stage_3__294_, data_stage_3__293_, data_stage_3__292_, data_stage_3__291_, data_stage_3__290_, data_stage_3__289_, data_stage_3__288_, data_stage_3__287_, data_stage_3__286_, data_stage_3__285_, data_stage_3__284_, data_stage_3__283_, data_stage_3__282_, data_stage_3__281_, data_stage_3__280_, data_stage_3__279_, data_stage_3__278_, data_stage_3__277_, data_stage_3__276_, data_stage_3__275_, data_stage_3__274_, data_stage_3__273_, data_stage_3__272_, data_stage_3__271_, data_stage_3__270_, data_stage_3__269_, data_stage_3__268_, data_stage_3__267_, data_stage_3__266_, data_stage_3__265_, data_stage_3__264_, data_stage_3__263_, data_stage_3__262_, data_stage_3__261_, data_stage_3__260_, data_stage_3__259_, data_stage_3__258_, data_stage_3__257_, data_stage_3__256_, data_stage_3__255_, data_stage_3__254_, data_stage_3__253_, data_stage_3__252_, data_stage_3__251_, data_stage_3__250_, data_stage_3__249_, data_stage_3__248_, data_stage_3__247_, data_stage_3__246_, data_stage_3__245_, data_stage_3__244_, data_stage_3__243_, data_stage_3__242_, data_stage_3__241_, data_stage_3__240_, data_stage_3__239_, data_stage_3__238_, data_stage_3__237_, data_stage_3__236_, data_stage_3__235_, data_stage_3__234_, data_stage_3__233_, data_stage_3__232_, data_stage_3__231_, data_stage_3__230_, data_stage_3__229_, data_stage_3__228_, data_stage_3__227_, data_stage_3__226_, data_stage_3__225_, data_stage_3__224_, data_stage_3__223_, data_stage_3__222_, data_stage_3__221_, data_stage_3__220_, data_stage_3__219_, data_stage_3__218_, data_stage_3__217_, data_stage_3__216_, data_stage_3__215_, data_stage_3__214_, data_stage_3__213_, data_stage_3__212_, data_stage_3__211_, data_stage_3__210_, data_stage_3__209_, data_stage_3__208_, data_stage_3__207_, data_stage_3__206_, data_stage_3__205_, data_stage_3__204_, data_stage_3__203_, data_stage_3__202_, data_stage_3__201_, data_stage_3__200_, data_stage_3__199_, data_stage_3__198_, data_stage_3__197_, data_stage_3__196_, data_stage_3__195_, data_stage_3__194_, data_stage_3__193_, data_stage_3__192_, data_stage_3__191_, data_stage_3__190_, data_stage_3__189_, data_stage_3__188_, data_stage_3__187_, data_stage_3__186_, data_stage_3__185_, data_stage_3__184_, data_stage_3__183_, data_stage_3__182_, data_stage_3__181_, data_stage_3__180_, data_stage_3__179_, data_stage_3__178_, data_stage_3__177_, data_stage_3__176_, data_stage_3__175_, data_stage_3__174_, data_stage_3__173_, data_stage_3__172_, data_stage_3__171_, data_stage_3__170_, data_stage_3__169_, data_stage_3__168_, data_stage_3__167_, data_stage_3__166_, data_stage_3__165_, data_stage_3__164_, data_stage_3__163_, data_stage_3__162_, data_stage_3__161_, data_stage_3__160_, data_stage_3__159_, data_stage_3__158_, data_stage_3__157_, data_stage_3__156_, data_stage_3__155_, data_stage_3__154_, data_stage_3__153_, data_stage_3__152_, data_stage_3__151_, data_stage_3__150_, data_stage_3__149_, data_stage_3__148_, data_stage_3__147_, data_stage_3__146_, data_stage_3__145_, data_stage_3__144_, data_stage_3__143_, data_stage_3__142_, data_stage_3__141_, data_stage_3__140_, data_stage_3__139_, data_stage_3__138_, data_stage_3__137_, data_stage_3__136_, data_stage_3__135_, data_stage_3__134_, data_stage_3__133_, data_stage_3__132_, data_stage_3__131_, data_stage_3__130_, data_stage_3__129_, data_stage_3__128_, data_stage_3__127_, data_stage_3__126_, data_stage_3__125_, data_stage_3__124_, data_stage_3__123_, data_stage_3__122_, data_stage_3__121_, data_stage_3__120_, data_stage_3__119_, data_stage_3__118_, data_stage_3__117_, data_stage_3__116_, data_stage_3__115_, data_stage_3__114_, data_stage_3__113_, data_stage_3__112_, data_stage_3__111_, data_stage_3__110_, data_stage_3__109_, data_stage_3__108_, data_stage_3__107_, data_stage_3__106_, data_stage_3__105_, data_stage_3__104_, data_stage_3__103_, data_stage_3__102_, data_stage_3__101_, data_stage_3__100_, data_stage_3__99_, data_stage_3__98_, data_stage_3__97_, data_stage_3__96_, data_stage_3__95_, data_stage_3__94_, data_stage_3__93_, data_stage_3__92_, data_stage_3__91_, data_stage_3__90_, data_stage_3__89_, data_stage_3__88_, data_stage_3__87_, data_stage_3__86_, data_stage_3__85_, data_stage_3__84_, data_stage_3__83_, data_stage_3__82_, data_stage_3__81_, data_stage_3__80_, data_stage_3__79_, data_stage_3__78_, data_stage_3__77_, data_stage_3__76_, data_stage_3__75_, data_stage_3__74_, data_stage_3__73_, data_stage_3__72_, data_stage_3__71_, data_stage_3__70_, data_stage_3__69_, data_stage_3__68_, data_stage_3__67_, data_stage_3__66_, data_stage_3__65_, data_stage_3__64_, data_stage_3__63_, data_stage_3__62_, data_stage_3__61_, data_stage_3__60_, data_stage_3__59_, data_stage_3__58_, data_stage_3__57_, data_stage_3__56_, data_stage_3__55_, data_stage_3__54_, data_stage_3__53_, data_stage_3__52_, data_stage_3__51_, data_stage_3__50_, data_stage_3__49_, data_stage_3__48_, data_stage_3__47_, data_stage_3__46_, data_stage_3__45_, data_stage_3__44_, data_stage_3__43_, data_stage_3__42_, data_stage_3__41_, data_stage_3__40_, data_stage_3__39_, data_stage_3__38_, data_stage_3__37_, data_stage_3__36_, data_stage_3__35_, data_stage_3__34_, data_stage_3__33_, data_stage_3__32_, data_stage_3__31_, data_stage_3__30_, data_stage_3__29_, data_stage_3__28_, data_stage_3__27_, data_stage_3__26_, data_stage_3__25_, data_stage_3__24_, data_stage_3__23_, data_stage_3__22_, data_stage_3__21_, data_stage_3__20_, data_stage_3__19_, data_stage_3__18_, data_stage_3__17_, data_stage_3__16_, data_stage_3__15_, data_stage_3__14_, data_stage_3__13_, data_stage_3__12_, data_stage_3__11_, data_stage_3__10_, data_stage_3__9_, data_stage_3__8_, data_stage_3__7_, data_stage_3__6_, data_stage_3__5_, data_stage_3__4_, data_stage_3__3_, data_stage_3__2_, data_stage_3__1_, data_stage_3__0_ }),
    .swap_i(sel_i[3]),
    .data_o({ data_stage_4__1023_, data_stage_4__1022_, data_stage_4__1021_, data_stage_4__1020_, data_stage_4__1019_, data_stage_4__1018_, data_stage_4__1017_, data_stage_4__1016_, data_stage_4__1015_, data_stage_4__1014_, data_stage_4__1013_, data_stage_4__1012_, data_stage_4__1011_, data_stage_4__1010_, data_stage_4__1009_, data_stage_4__1008_, data_stage_4__1007_, data_stage_4__1006_, data_stage_4__1005_, data_stage_4__1004_, data_stage_4__1003_, data_stage_4__1002_, data_stage_4__1001_, data_stage_4__1000_, data_stage_4__999_, data_stage_4__998_, data_stage_4__997_, data_stage_4__996_, data_stage_4__995_, data_stage_4__994_, data_stage_4__993_, data_stage_4__992_, data_stage_4__991_, data_stage_4__990_, data_stage_4__989_, data_stage_4__988_, data_stage_4__987_, data_stage_4__986_, data_stage_4__985_, data_stage_4__984_, data_stage_4__983_, data_stage_4__982_, data_stage_4__981_, data_stage_4__980_, data_stage_4__979_, data_stage_4__978_, data_stage_4__977_, data_stage_4__976_, data_stage_4__975_, data_stage_4__974_, data_stage_4__973_, data_stage_4__972_, data_stage_4__971_, data_stage_4__970_, data_stage_4__969_, data_stage_4__968_, data_stage_4__967_, data_stage_4__966_, data_stage_4__965_, data_stage_4__964_, data_stage_4__963_, data_stage_4__962_, data_stage_4__961_, data_stage_4__960_, data_stage_4__959_, data_stage_4__958_, data_stage_4__957_, data_stage_4__956_, data_stage_4__955_, data_stage_4__954_, data_stage_4__953_, data_stage_4__952_, data_stage_4__951_, data_stage_4__950_, data_stage_4__949_, data_stage_4__948_, data_stage_4__947_, data_stage_4__946_, data_stage_4__945_, data_stage_4__944_, data_stage_4__943_, data_stage_4__942_, data_stage_4__941_, data_stage_4__940_, data_stage_4__939_, data_stage_4__938_, data_stage_4__937_, data_stage_4__936_, data_stage_4__935_, data_stage_4__934_, data_stage_4__933_, data_stage_4__932_, data_stage_4__931_, data_stage_4__930_, data_stage_4__929_, data_stage_4__928_, data_stage_4__927_, data_stage_4__926_, data_stage_4__925_, data_stage_4__924_, data_stage_4__923_, data_stage_4__922_, data_stage_4__921_, data_stage_4__920_, data_stage_4__919_, data_stage_4__918_, data_stage_4__917_, data_stage_4__916_, data_stage_4__915_, data_stage_4__914_, data_stage_4__913_, data_stage_4__912_, data_stage_4__911_, data_stage_4__910_, data_stage_4__909_, data_stage_4__908_, data_stage_4__907_, data_stage_4__906_, data_stage_4__905_, data_stage_4__904_, data_stage_4__903_, data_stage_4__902_, data_stage_4__901_, data_stage_4__900_, data_stage_4__899_, data_stage_4__898_, data_stage_4__897_, data_stage_4__896_, data_stage_4__895_, data_stage_4__894_, data_stage_4__893_, data_stage_4__892_, data_stage_4__891_, data_stage_4__890_, data_stage_4__889_, data_stage_4__888_, data_stage_4__887_, data_stage_4__886_, data_stage_4__885_, data_stage_4__884_, data_stage_4__883_, data_stage_4__882_, data_stage_4__881_, data_stage_4__880_, data_stage_4__879_, data_stage_4__878_, data_stage_4__877_, data_stage_4__876_, data_stage_4__875_, data_stage_4__874_, data_stage_4__873_, data_stage_4__872_, data_stage_4__871_, data_stage_4__870_, data_stage_4__869_, data_stage_4__868_, data_stage_4__867_, data_stage_4__866_, data_stage_4__865_, data_stage_4__864_, data_stage_4__863_, data_stage_4__862_, data_stage_4__861_, data_stage_4__860_, data_stage_4__859_, data_stage_4__858_, data_stage_4__857_, data_stage_4__856_, data_stage_4__855_, data_stage_4__854_, data_stage_4__853_, data_stage_4__852_, data_stage_4__851_, data_stage_4__850_, data_stage_4__849_, data_stage_4__848_, data_stage_4__847_, data_stage_4__846_, data_stage_4__845_, data_stage_4__844_, data_stage_4__843_, data_stage_4__842_, data_stage_4__841_, data_stage_4__840_, data_stage_4__839_, data_stage_4__838_, data_stage_4__837_, data_stage_4__836_, data_stage_4__835_, data_stage_4__834_, data_stage_4__833_, data_stage_4__832_, data_stage_4__831_, data_stage_4__830_, data_stage_4__829_, data_stage_4__828_, data_stage_4__827_, data_stage_4__826_, data_stage_4__825_, data_stage_4__824_, data_stage_4__823_, data_stage_4__822_, data_stage_4__821_, data_stage_4__820_, data_stage_4__819_, data_stage_4__818_, data_stage_4__817_, data_stage_4__816_, data_stage_4__815_, data_stage_4__814_, data_stage_4__813_, data_stage_4__812_, data_stage_4__811_, data_stage_4__810_, data_stage_4__809_, data_stage_4__808_, data_stage_4__807_, data_stage_4__806_, data_stage_4__805_, data_stage_4__804_, data_stage_4__803_, data_stage_4__802_, data_stage_4__801_, data_stage_4__800_, data_stage_4__799_, data_stage_4__798_, data_stage_4__797_, data_stage_4__796_, data_stage_4__795_, data_stage_4__794_, data_stage_4__793_, data_stage_4__792_, data_stage_4__791_, data_stage_4__790_, data_stage_4__789_, data_stage_4__788_, data_stage_4__787_, data_stage_4__786_, data_stage_4__785_, data_stage_4__784_, data_stage_4__783_, data_stage_4__782_, data_stage_4__781_, data_stage_4__780_, data_stage_4__779_, data_stage_4__778_, data_stage_4__777_, data_stage_4__776_, data_stage_4__775_, data_stage_4__774_, data_stage_4__773_, data_stage_4__772_, data_stage_4__771_, data_stage_4__770_, data_stage_4__769_, data_stage_4__768_, data_stage_4__767_, data_stage_4__766_, data_stage_4__765_, data_stage_4__764_, data_stage_4__763_, data_stage_4__762_, data_stage_4__761_, data_stage_4__760_, data_stage_4__759_, data_stage_4__758_, data_stage_4__757_, data_stage_4__756_, data_stage_4__755_, data_stage_4__754_, data_stage_4__753_, data_stage_4__752_, data_stage_4__751_, data_stage_4__750_, data_stage_4__749_, data_stage_4__748_, data_stage_4__747_, data_stage_4__746_, data_stage_4__745_, data_stage_4__744_, data_stage_4__743_, data_stage_4__742_, data_stage_4__741_, data_stage_4__740_, data_stage_4__739_, data_stage_4__738_, data_stage_4__737_, data_stage_4__736_, data_stage_4__735_, data_stage_4__734_, data_stage_4__733_, data_stage_4__732_, data_stage_4__731_, data_stage_4__730_, data_stage_4__729_, data_stage_4__728_, data_stage_4__727_, data_stage_4__726_, data_stage_4__725_, data_stage_4__724_, data_stage_4__723_, data_stage_4__722_, data_stage_4__721_, data_stage_4__720_, data_stage_4__719_, data_stage_4__718_, data_stage_4__717_, data_stage_4__716_, data_stage_4__715_, data_stage_4__714_, data_stage_4__713_, data_stage_4__712_, data_stage_4__711_, data_stage_4__710_, data_stage_4__709_, data_stage_4__708_, data_stage_4__707_, data_stage_4__706_, data_stage_4__705_, data_stage_4__704_, data_stage_4__703_, data_stage_4__702_, data_stage_4__701_, data_stage_4__700_, data_stage_4__699_, data_stage_4__698_, data_stage_4__697_, data_stage_4__696_, data_stage_4__695_, data_stage_4__694_, data_stage_4__693_, data_stage_4__692_, data_stage_4__691_, data_stage_4__690_, data_stage_4__689_, data_stage_4__688_, data_stage_4__687_, data_stage_4__686_, data_stage_4__685_, data_stage_4__684_, data_stage_4__683_, data_stage_4__682_, data_stage_4__681_, data_stage_4__680_, data_stage_4__679_, data_stage_4__678_, data_stage_4__677_, data_stage_4__676_, data_stage_4__675_, data_stage_4__674_, data_stage_4__673_, data_stage_4__672_, data_stage_4__671_, data_stage_4__670_, data_stage_4__669_, data_stage_4__668_, data_stage_4__667_, data_stage_4__666_, data_stage_4__665_, data_stage_4__664_, data_stage_4__663_, data_stage_4__662_, data_stage_4__661_, data_stage_4__660_, data_stage_4__659_, data_stage_4__658_, data_stage_4__657_, data_stage_4__656_, data_stage_4__655_, data_stage_4__654_, data_stage_4__653_, data_stage_4__652_, data_stage_4__651_, data_stage_4__650_, data_stage_4__649_, data_stage_4__648_, data_stage_4__647_, data_stage_4__646_, data_stage_4__645_, data_stage_4__644_, data_stage_4__643_, data_stage_4__642_, data_stage_4__641_, data_stage_4__640_, data_stage_4__639_, data_stage_4__638_, data_stage_4__637_, data_stage_4__636_, data_stage_4__635_, data_stage_4__634_, data_stage_4__633_, data_stage_4__632_, data_stage_4__631_, data_stage_4__630_, data_stage_4__629_, data_stage_4__628_, data_stage_4__627_, data_stage_4__626_, data_stage_4__625_, data_stage_4__624_, data_stage_4__623_, data_stage_4__622_, data_stage_4__621_, data_stage_4__620_, data_stage_4__619_, data_stage_4__618_, data_stage_4__617_, data_stage_4__616_, data_stage_4__615_, data_stage_4__614_, data_stage_4__613_, data_stage_4__612_, data_stage_4__611_, data_stage_4__610_, data_stage_4__609_, data_stage_4__608_, data_stage_4__607_, data_stage_4__606_, data_stage_4__605_, data_stage_4__604_, data_stage_4__603_, data_stage_4__602_, data_stage_4__601_, data_stage_4__600_, data_stage_4__599_, data_stage_4__598_, data_stage_4__597_, data_stage_4__596_, data_stage_4__595_, data_stage_4__594_, data_stage_4__593_, data_stage_4__592_, data_stage_4__591_, data_stage_4__590_, data_stage_4__589_, data_stage_4__588_, data_stage_4__587_, data_stage_4__586_, data_stage_4__585_, data_stage_4__584_, data_stage_4__583_, data_stage_4__582_, data_stage_4__581_, data_stage_4__580_, data_stage_4__579_, data_stage_4__578_, data_stage_4__577_, data_stage_4__576_, data_stage_4__575_, data_stage_4__574_, data_stage_4__573_, data_stage_4__572_, data_stage_4__571_, data_stage_4__570_, data_stage_4__569_, data_stage_4__568_, data_stage_4__567_, data_stage_4__566_, data_stage_4__565_, data_stage_4__564_, data_stage_4__563_, data_stage_4__562_, data_stage_4__561_, data_stage_4__560_, data_stage_4__559_, data_stage_4__558_, data_stage_4__557_, data_stage_4__556_, data_stage_4__555_, data_stage_4__554_, data_stage_4__553_, data_stage_4__552_, data_stage_4__551_, data_stage_4__550_, data_stage_4__549_, data_stage_4__548_, data_stage_4__547_, data_stage_4__546_, data_stage_4__545_, data_stage_4__544_, data_stage_4__543_, data_stage_4__542_, data_stage_4__541_, data_stage_4__540_, data_stage_4__539_, data_stage_4__538_, data_stage_4__537_, data_stage_4__536_, data_stage_4__535_, data_stage_4__534_, data_stage_4__533_, data_stage_4__532_, data_stage_4__531_, data_stage_4__530_, data_stage_4__529_, data_stage_4__528_, data_stage_4__527_, data_stage_4__526_, data_stage_4__525_, data_stage_4__524_, data_stage_4__523_, data_stage_4__522_, data_stage_4__521_, data_stage_4__520_, data_stage_4__519_, data_stage_4__518_, data_stage_4__517_, data_stage_4__516_, data_stage_4__515_, data_stage_4__514_, data_stage_4__513_, data_stage_4__512_, data_stage_4__511_, data_stage_4__510_, data_stage_4__509_, data_stage_4__508_, data_stage_4__507_, data_stage_4__506_, data_stage_4__505_, data_stage_4__504_, data_stage_4__503_, data_stage_4__502_, data_stage_4__501_, data_stage_4__500_, data_stage_4__499_, data_stage_4__498_, data_stage_4__497_, data_stage_4__496_, data_stage_4__495_, data_stage_4__494_, data_stage_4__493_, data_stage_4__492_, data_stage_4__491_, data_stage_4__490_, data_stage_4__489_, data_stage_4__488_, data_stage_4__487_, data_stage_4__486_, data_stage_4__485_, data_stage_4__484_, data_stage_4__483_, data_stage_4__482_, data_stage_4__481_, data_stage_4__480_, data_stage_4__479_, data_stage_4__478_, data_stage_4__477_, data_stage_4__476_, data_stage_4__475_, data_stage_4__474_, data_stage_4__473_, data_stage_4__472_, data_stage_4__471_, data_stage_4__470_, data_stage_4__469_, data_stage_4__468_, data_stage_4__467_, data_stage_4__466_, data_stage_4__465_, data_stage_4__464_, data_stage_4__463_, data_stage_4__462_, data_stage_4__461_, data_stage_4__460_, data_stage_4__459_, data_stage_4__458_, data_stage_4__457_, data_stage_4__456_, data_stage_4__455_, data_stage_4__454_, data_stage_4__453_, data_stage_4__452_, data_stage_4__451_, data_stage_4__450_, data_stage_4__449_, data_stage_4__448_, data_stage_4__447_, data_stage_4__446_, data_stage_4__445_, data_stage_4__444_, data_stage_4__443_, data_stage_4__442_, data_stage_4__441_, data_stage_4__440_, data_stage_4__439_, data_stage_4__438_, data_stage_4__437_, data_stage_4__436_, data_stage_4__435_, data_stage_4__434_, data_stage_4__433_, data_stage_4__432_, data_stage_4__431_, data_stage_4__430_, data_stage_4__429_, data_stage_4__428_, data_stage_4__427_, data_stage_4__426_, data_stage_4__425_, data_stage_4__424_, data_stage_4__423_, data_stage_4__422_, data_stage_4__421_, data_stage_4__420_, data_stage_4__419_, data_stage_4__418_, data_stage_4__417_, data_stage_4__416_, data_stage_4__415_, data_stage_4__414_, data_stage_4__413_, data_stage_4__412_, data_stage_4__411_, data_stage_4__410_, data_stage_4__409_, data_stage_4__408_, data_stage_4__407_, data_stage_4__406_, data_stage_4__405_, data_stage_4__404_, data_stage_4__403_, data_stage_4__402_, data_stage_4__401_, data_stage_4__400_, data_stage_4__399_, data_stage_4__398_, data_stage_4__397_, data_stage_4__396_, data_stage_4__395_, data_stage_4__394_, data_stage_4__393_, data_stage_4__392_, data_stage_4__391_, data_stage_4__390_, data_stage_4__389_, data_stage_4__388_, data_stage_4__387_, data_stage_4__386_, data_stage_4__385_, data_stage_4__384_, data_stage_4__383_, data_stage_4__382_, data_stage_4__381_, data_stage_4__380_, data_stage_4__379_, data_stage_4__378_, data_stage_4__377_, data_stage_4__376_, data_stage_4__375_, data_stage_4__374_, data_stage_4__373_, data_stage_4__372_, data_stage_4__371_, data_stage_4__370_, data_stage_4__369_, data_stage_4__368_, data_stage_4__367_, data_stage_4__366_, data_stage_4__365_, data_stage_4__364_, data_stage_4__363_, data_stage_4__362_, data_stage_4__361_, data_stage_4__360_, data_stage_4__359_, data_stage_4__358_, data_stage_4__357_, data_stage_4__356_, data_stage_4__355_, data_stage_4__354_, data_stage_4__353_, data_stage_4__352_, data_stage_4__351_, data_stage_4__350_, data_stage_4__349_, data_stage_4__348_, data_stage_4__347_, data_stage_4__346_, data_stage_4__345_, data_stage_4__344_, data_stage_4__343_, data_stage_4__342_, data_stage_4__341_, data_stage_4__340_, data_stage_4__339_, data_stage_4__338_, data_stage_4__337_, data_stage_4__336_, data_stage_4__335_, data_stage_4__334_, data_stage_4__333_, data_stage_4__332_, data_stage_4__331_, data_stage_4__330_, data_stage_4__329_, data_stage_4__328_, data_stage_4__327_, data_stage_4__326_, data_stage_4__325_, data_stage_4__324_, data_stage_4__323_, data_stage_4__322_, data_stage_4__321_, data_stage_4__320_, data_stage_4__319_, data_stage_4__318_, data_stage_4__317_, data_stage_4__316_, data_stage_4__315_, data_stage_4__314_, data_stage_4__313_, data_stage_4__312_, data_stage_4__311_, data_stage_4__310_, data_stage_4__309_, data_stage_4__308_, data_stage_4__307_, data_stage_4__306_, data_stage_4__305_, data_stage_4__304_, data_stage_4__303_, data_stage_4__302_, data_stage_4__301_, data_stage_4__300_, data_stage_4__299_, data_stage_4__298_, data_stage_4__297_, data_stage_4__296_, data_stage_4__295_, data_stage_4__294_, data_stage_4__293_, data_stage_4__292_, data_stage_4__291_, data_stage_4__290_, data_stage_4__289_, data_stage_4__288_, data_stage_4__287_, data_stage_4__286_, data_stage_4__285_, data_stage_4__284_, data_stage_4__283_, data_stage_4__282_, data_stage_4__281_, data_stage_4__280_, data_stage_4__279_, data_stage_4__278_, data_stage_4__277_, data_stage_4__276_, data_stage_4__275_, data_stage_4__274_, data_stage_4__273_, data_stage_4__272_, data_stage_4__271_, data_stage_4__270_, data_stage_4__269_, data_stage_4__268_, data_stage_4__267_, data_stage_4__266_, data_stage_4__265_, data_stage_4__264_, data_stage_4__263_, data_stage_4__262_, data_stage_4__261_, data_stage_4__260_, data_stage_4__259_, data_stage_4__258_, data_stage_4__257_, data_stage_4__256_, data_stage_4__255_, data_stage_4__254_, data_stage_4__253_, data_stage_4__252_, data_stage_4__251_, data_stage_4__250_, data_stage_4__249_, data_stage_4__248_, data_stage_4__247_, data_stage_4__246_, data_stage_4__245_, data_stage_4__244_, data_stage_4__243_, data_stage_4__242_, data_stage_4__241_, data_stage_4__240_, data_stage_4__239_, data_stage_4__238_, data_stage_4__237_, data_stage_4__236_, data_stage_4__235_, data_stage_4__234_, data_stage_4__233_, data_stage_4__232_, data_stage_4__231_, data_stage_4__230_, data_stage_4__229_, data_stage_4__228_, data_stage_4__227_, data_stage_4__226_, data_stage_4__225_, data_stage_4__224_, data_stage_4__223_, data_stage_4__222_, data_stage_4__221_, data_stage_4__220_, data_stage_4__219_, data_stage_4__218_, data_stage_4__217_, data_stage_4__216_, data_stage_4__215_, data_stage_4__214_, data_stage_4__213_, data_stage_4__212_, data_stage_4__211_, data_stage_4__210_, data_stage_4__209_, data_stage_4__208_, data_stage_4__207_, data_stage_4__206_, data_stage_4__205_, data_stage_4__204_, data_stage_4__203_, data_stage_4__202_, data_stage_4__201_, data_stage_4__200_, data_stage_4__199_, data_stage_4__198_, data_stage_4__197_, data_stage_4__196_, data_stage_4__195_, data_stage_4__194_, data_stage_4__193_, data_stage_4__192_, data_stage_4__191_, data_stage_4__190_, data_stage_4__189_, data_stage_4__188_, data_stage_4__187_, data_stage_4__186_, data_stage_4__185_, data_stage_4__184_, data_stage_4__183_, data_stage_4__182_, data_stage_4__181_, data_stage_4__180_, data_stage_4__179_, data_stage_4__178_, data_stage_4__177_, data_stage_4__176_, data_stage_4__175_, data_stage_4__174_, data_stage_4__173_, data_stage_4__172_, data_stage_4__171_, data_stage_4__170_, data_stage_4__169_, data_stage_4__168_, data_stage_4__167_, data_stage_4__166_, data_stage_4__165_, data_stage_4__164_, data_stage_4__163_, data_stage_4__162_, data_stage_4__161_, data_stage_4__160_, data_stage_4__159_, data_stage_4__158_, data_stage_4__157_, data_stage_4__156_, data_stage_4__155_, data_stage_4__154_, data_stage_4__153_, data_stage_4__152_, data_stage_4__151_, data_stage_4__150_, data_stage_4__149_, data_stage_4__148_, data_stage_4__147_, data_stage_4__146_, data_stage_4__145_, data_stage_4__144_, data_stage_4__143_, data_stage_4__142_, data_stage_4__141_, data_stage_4__140_, data_stage_4__139_, data_stage_4__138_, data_stage_4__137_, data_stage_4__136_, data_stage_4__135_, data_stage_4__134_, data_stage_4__133_, data_stage_4__132_, data_stage_4__131_, data_stage_4__130_, data_stage_4__129_, data_stage_4__128_, data_stage_4__127_, data_stage_4__126_, data_stage_4__125_, data_stage_4__124_, data_stage_4__123_, data_stage_4__122_, data_stage_4__121_, data_stage_4__120_, data_stage_4__119_, data_stage_4__118_, data_stage_4__117_, data_stage_4__116_, data_stage_4__115_, data_stage_4__114_, data_stage_4__113_, data_stage_4__112_, data_stage_4__111_, data_stage_4__110_, data_stage_4__109_, data_stage_4__108_, data_stage_4__107_, data_stage_4__106_, data_stage_4__105_, data_stage_4__104_, data_stage_4__103_, data_stage_4__102_, data_stage_4__101_, data_stage_4__100_, data_stage_4__99_, data_stage_4__98_, data_stage_4__97_, data_stage_4__96_, data_stage_4__95_, data_stage_4__94_, data_stage_4__93_, data_stage_4__92_, data_stage_4__91_, data_stage_4__90_, data_stage_4__89_, data_stage_4__88_, data_stage_4__87_, data_stage_4__86_, data_stage_4__85_, data_stage_4__84_, data_stage_4__83_, data_stage_4__82_, data_stage_4__81_, data_stage_4__80_, data_stage_4__79_, data_stage_4__78_, data_stage_4__77_, data_stage_4__76_, data_stage_4__75_, data_stage_4__74_, data_stage_4__73_, data_stage_4__72_, data_stage_4__71_, data_stage_4__70_, data_stage_4__69_, data_stage_4__68_, data_stage_4__67_, data_stage_4__66_, data_stage_4__65_, data_stage_4__64_, data_stage_4__63_, data_stage_4__62_, data_stage_4__61_, data_stage_4__60_, data_stage_4__59_, data_stage_4__58_, data_stage_4__57_, data_stage_4__56_, data_stage_4__55_, data_stage_4__54_, data_stage_4__53_, data_stage_4__52_, data_stage_4__51_, data_stage_4__50_, data_stage_4__49_, data_stage_4__48_, data_stage_4__47_, data_stage_4__46_, data_stage_4__45_, data_stage_4__44_, data_stage_4__43_, data_stage_4__42_, data_stage_4__41_, data_stage_4__40_, data_stage_4__39_, data_stage_4__38_, data_stage_4__37_, data_stage_4__36_, data_stage_4__35_, data_stage_4__34_, data_stage_4__33_, data_stage_4__32_, data_stage_4__31_, data_stage_4__30_, data_stage_4__29_, data_stage_4__28_, data_stage_4__27_, data_stage_4__26_, data_stage_4__25_, data_stage_4__24_, data_stage_4__23_, data_stage_4__22_, data_stage_4__21_, data_stage_4__20_, data_stage_4__19_, data_stage_4__18_, data_stage_4__17_, data_stage_4__16_, data_stage_4__15_, data_stage_4__14_, data_stage_4__13_, data_stage_4__12_, data_stage_4__11_, data_stage_4__10_, data_stage_4__9_, data_stage_4__8_, data_stage_4__7_, data_stage_4__6_, data_stage_4__5_, data_stage_4__4_, data_stage_4__3_, data_stage_4__2_, data_stage_4__1_, data_stage_4__0_ })
  );


  bsg_swap_width_p512
  mux_stage_3__mux_swap_1__swap_inst
  (
    .data_i({ data_stage_3__2047_, data_stage_3__2046_, data_stage_3__2045_, data_stage_3__2044_, data_stage_3__2043_, data_stage_3__2042_, data_stage_3__2041_, data_stage_3__2040_, data_stage_3__2039_, data_stage_3__2038_, data_stage_3__2037_, data_stage_3__2036_, data_stage_3__2035_, data_stage_3__2034_, data_stage_3__2033_, data_stage_3__2032_, data_stage_3__2031_, data_stage_3__2030_, data_stage_3__2029_, data_stage_3__2028_, data_stage_3__2027_, data_stage_3__2026_, data_stage_3__2025_, data_stage_3__2024_, data_stage_3__2023_, data_stage_3__2022_, data_stage_3__2021_, data_stage_3__2020_, data_stage_3__2019_, data_stage_3__2018_, data_stage_3__2017_, data_stage_3__2016_, data_stage_3__2015_, data_stage_3__2014_, data_stage_3__2013_, data_stage_3__2012_, data_stage_3__2011_, data_stage_3__2010_, data_stage_3__2009_, data_stage_3__2008_, data_stage_3__2007_, data_stage_3__2006_, data_stage_3__2005_, data_stage_3__2004_, data_stage_3__2003_, data_stage_3__2002_, data_stage_3__2001_, data_stage_3__2000_, data_stage_3__1999_, data_stage_3__1998_, data_stage_3__1997_, data_stage_3__1996_, data_stage_3__1995_, data_stage_3__1994_, data_stage_3__1993_, data_stage_3__1992_, data_stage_3__1991_, data_stage_3__1990_, data_stage_3__1989_, data_stage_3__1988_, data_stage_3__1987_, data_stage_3__1986_, data_stage_3__1985_, data_stage_3__1984_, data_stage_3__1983_, data_stage_3__1982_, data_stage_3__1981_, data_stage_3__1980_, data_stage_3__1979_, data_stage_3__1978_, data_stage_3__1977_, data_stage_3__1976_, data_stage_3__1975_, data_stage_3__1974_, data_stage_3__1973_, data_stage_3__1972_, data_stage_3__1971_, data_stage_3__1970_, data_stage_3__1969_, data_stage_3__1968_, data_stage_3__1967_, data_stage_3__1966_, data_stage_3__1965_, data_stage_3__1964_, data_stage_3__1963_, data_stage_3__1962_, data_stage_3__1961_, data_stage_3__1960_, data_stage_3__1959_, data_stage_3__1958_, data_stage_3__1957_, data_stage_3__1956_, data_stage_3__1955_, data_stage_3__1954_, data_stage_3__1953_, data_stage_3__1952_, data_stage_3__1951_, data_stage_3__1950_, data_stage_3__1949_, data_stage_3__1948_, data_stage_3__1947_, data_stage_3__1946_, data_stage_3__1945_, data_stage_3__1944_, data_stage_3__1943_, data_stage_3__1942_, data_stage_3__1941_, data_stage_3__1940_, data_stage_3__1939_, data_stage_3__1938_, data_stage_3__1937_, data_stage_3__1936_, data_stage_3__1935_, data_stage_3__1934_, data_stage_3__1933_, data_stage_3__1932_, data_stage_3__1931_, data_stage_3__1930_, data_stage_3__1929_, data_stage_3__1928_, data_stage_3__1927_, data_stage_3__1926_, data_stage_3__1925_, data_stage_3__1924_, data_stage_3__1923_, data_stage_3__1922_, data_stage_3__1921_, data_stage_3__1920_, data_stage_3__1919_, data_stage_3__1918_, data_stage_3__1917_, data_stage_3__1916_, data_stage_3__1915_, data_stage_3__1914_, data_stage_3__1913_, data_stage_3__1912_, data_stage_3__1911_, data_stage_3__1910_, data_stage_3__1909_, data_stage_3__1908_, data_stage_3__1907_, data_stage_3__1906_, data_stage_3__1905_, data_stage_3__1904_, data_stage_3__1903_, data_stage_3__1902_, data_stage_3__1901_, data_stage_3__1900_, data_stage_3__1899_, data_stage_3__1898_, data_stage_3__1897_, data_stage_3__1896_, data_stage_3__1895_, data_stage_3__1894_, data_stage_3__1893_, data_stage_3__1892_, data_stage_3__1891_, data_stage_3__1890_, data_stage_3__1889_, data_stage_3__1888_, data_stage_3__1887_, data_stage_3__1886_, data_stage_3__1885_, data_stage_3__1884_, data_stage_3__1883_, data_stage_3__1882_, data_stage_3__1881_, data_stage_3__1880_, data_stage_3__1879_, data_stage_3__1878_, data_stage_3__1877_, data_stage_3__1876_, data_stage_3__1875_, data_stage_3__1874_, data_stage_3__1873_, data_stage_3__1872_, data_stage_3__1871_, data_stage_3__1870_, data_stage_3__1869_, data_stage_3__1868_, data_stage_3__1867_, data_stage_3__1866_, data_stage_3__1865_, data_stage_3__1864_, data_stage_3__1863_, data_stage_3__1862_, data_stage_3__1861_, data_stage_3__1860_, data_stage_3__1859_, data_stage_3__1858_, data_stage_3__1857_, data_stage_3__1856_, data_stage_3__1855_, data_stage_3__1854_, data_stage_3__1853_, data_stage_3__1852_, data_stage_3__1851_, data_stage_3__1850_, data_stage_3__1849_, data_stage_3__1848_, data_stage_3__1847_, data_stage_3__1846_, data_stage_3__1845_, data_stage_3__1844_, data_stage_3__1843_, data_stage_3__1842_, data_stage_3__1841_, data_stage_3__1840_, data_stage_3__1839_, data_stage_3__1838_, data_stage_3__1837_, data_stage_3__1836_, data_stage_3__1835_, data_stage_3__1834_, data_stage_3__1833_, data_stage_3__1832_, data_stage_3__1831_, data_stage_3__1830_, data_stage_3__1829_, data_stage_3__1828_, data_stage_3__1827_, data_stage_3__1826_, data_stage_3__1825_, data_stage_3__1824_, data_stage_3__1823_, data_stage_3__1822_, data_stage_3__1821_, data_stage_3__1820_, data_stage_3__1819_, data_stage_3__1818_, data_stage_3__1817_, data_stage_3__1816_, data_stage_3__1815_, data_stage_3__1814_, data_stage_3__1813_, data_stage_3__1812_, data_stage_3__1811_, data_stage_3__1810_, data_stage_3__1809_, data_stage_3__1808_, data_stage_3__1807_, data_stage_3__1806_, data_stage_3__1805_, data_stage_3__1804_, data_stage_3__1803_, data_stage_3__1802_, data_stage_3__1801_, data_stage_3__1800_, data_stage_3__1799_, data_stage_3__1798_, data_stage_3__1797_, data_stage_3__1796_, data_stage_3__1795_, data_stage_3__1794_, data_stage_3__1793_, data_stage_3__1792_, data_stage_3__1791_, data_stage_3__1790_, data_stage_3__1789_, data_stage_3__1788_, data_stage_3__1787_, data_stage_3__1786_, data_stage_3__1785_, data_stage_3__1784_, data_stage_3__1783_, data_stage_3__1782_, data_stage_3__1781_, data_stage_3__1780_, data_stage_3__1779_, data_stage_3__1778_, data_stage_3__1777_, data_stage_3__1776_, data_stage_3__1775_, data_stage_3__1774_, data_stage_3__1773_, data_stage_3__1772_, data_stage_3__1771_, data_stage_3__1770_, data_stage_3__1769_, data_stage_3__1768_, data_stage_3__1767_, data_stage_3__1766_, data_stage_3__1765_, data_stage_3__1764_, data_stage_3__1763_, data_stage_3__1762_, data_stage_3__1761_, data_stage_3__1760_, data_stage_3__1759_, data_stage_3__1758_, data_stage_3__1757_, data_stage_3__1756_, data_stage_3__1755_, data_stage_3__1754_, data_stage_3__1753_, data_stage_3__1752_, data_stage_3__1751_, data_stage_3__1750_, data_stage_3__1749_, data_stage_3__1748_, data_stage_3__1747_, data_stage_3__1746_, data_stage_3__1745_, data_stage_3__1744_, data_stage_3__1743_, data_stage_3__1742_, data_stage_3__1741_, data_stage_3__1740_, data_stage_3__1739_, data_stage_3__1738_, data_stage_3__1737_, data_stage_3__1736_, data_stage_3__1735_, data_stage_3__1734_, data_stage_3__1733_, data_stage_3__1732_, data_stage_3__1731_, data_stage_3__1730_, data_stage_3__1729_, data_stage_3__1728_, data_stage_3__1727_, data_stage_3__1726_, data_stage_3__1725_, data_stage_3__1724_, data_stage_3__1723_, data_stage_3__1722_, data_stage_3__1721_, data_stage_3__1720_, data_stage_3__1719_, data_stage_3__1718_, data_stage_3__1717_, data_stage_3__1716_, data_stage_3__1715_, data_stage_3__1714_, data_stage_3__1713_, data_stage_3__1712_, data_stage_3__1711_, data_stage_3__1710_, data_stage_3__1709_, data_stage_3__1708_, data_stage_3__1707_, data_stage_3__1706_, data_stage_3__1705_, data_stage_3__1704_, data_stage_3__1703_, data_stage_3__1702_, data_stage_3__1701_, data_stage_3__1700_, data_stage_3__1699_, data_stage_3__1698_, data_stage_3__1697_, data_stage_3__1696_, data_stage_3__1695_, data_stage_3__1694_, data_stage_3__1693_, data_stage_3__1692_, data_stage_3__1691_, data_stage_3__1690_, data_stage_3__1689_, data_stage_3__1688_, data_stage_3__1687_, data_stage_3__1686_, data_stage_3__1685_, data_stage_3__1684_, data_stage_3__1683_, data_stage_3__1682_, data_stage_3__1681_, data_stage_3__1680_, data_stage_3__1679_, data_stage_3__1678_, data_stage_3__1677_, data_stage_3__1676_, data_stage_3__1675_, data_stage_3__1674_, data_stage_3__1673_, data_stage_3__1672_, data_stage_3__1671_, data_stage_3__1670_, data_stage_3__1669_, data_stage_3__1668_, data_stage_3__1667_, data_stage_3__1666_, data_stage_3__1665_, data_stage_3__1664_, data_stage_3__1663_, data_stage_3__1662_, data_stage_3__1661_, data_stage_3__1660_, data_stage_3__1659_, data_stage_3__1658_, data_stage_3__1657_, data_stage_3__1656_, data_stage_3__1655_, data_stage_3__1654_, data_stage_3__1653_, data_stage_3__1652_, data_stage_3__1651_, data_stage_3__1650_, data_stage_3__1649_, data_stage_3__1648_, data_stage_3__1647_, data_stage_3__1646_, data_stage_3__1645_, data_stage_3__1644_, data_stage_3__1643_, data_stage_3__1642_, data_stage_3__1641_, data_stage_3__1640_, data_stage_3__1639_, data_stage_3__1638_, data_stage_3__1637_, data_stage_3__1636_, data_stage_3__1635_, data_stage_3__1634_, data_stage_3__1633_, data_stage_3__1632_, data_stage_3__1631_, data_stage_3__1630_, data_stage_3__1629_, data_stage_3__1628_, data_stage_3__1627_, data_stage_3__1626_, data_stage_3__1625_, data_stage_3__1624_, data_stage_3__1623_, data_stage_3__1622_, data_stage_3__1621_, data_stage_3__1620_, data_stage_3__1619_, data_stage_3__1618_, data_stage_3__1617_, data_stage_3__1616_, data_stage_3__1615_, data_stage_3__1614_, data_stage_3__1613_, data_stage_3__1612_, data_stage_3__1611_, data_stage_3__1610_, data_stage_3__1609_, data_stage_3__1608_, data_stage_3__1607_, data_stage_3__1606_, data_stage_3__1605_, data_stage_3__1604_, data_stage_3__1603_, data_stage_3__1602_, data_stage_3__1601_, data_stage_3__1600_, data_stage_3__1599_, data_stage_3__1598_, data_stage_3__1597_, data_stage_3__1596_, data_stage_3__1595_, data_stage_3__1594_, data_stage_3__1593_, data_stage_3__1592_, data_stage_3__1591_, data_stage_3__1590_, data_stage_3__1589_, data_stage_3__1588_, data_stage_3__1587_, data_stage_3__1586_, data_stage_3__1585_, data_stage_3__1584_, data_stage_3__1583_, data_stage_3__1582_, data_stage_3__1581_, data_stage_3__1580_, data_stage_3__1579_, data_stage_3__1578_, data_stage_3__1577_, data_stage_3__1576_, data_stage_3__1575_, data_stage_3__1574_, data_stage_3__1573_, data_stage_3__1572_, data_stage_3__1571_, data_stage_3__1570_, data_stage_3__1569_, data_stage_3__1568_, data_stage_3__1567_, data_stage_3__1566_, data_stage_3__1565_, data_stage_3__1564_, data_stage_3__1563_, data_stage_3__1562_, data_stage_3__1561_, data_stage_3__1560_, data_stage_3__1559_, data_stage_3__1558_, data_stage_3__1557_, data_stage_3__1556_, data_stage_3__1555_, data_stage_3__1554_, data_stage_3__1553_, data_stage_3__1552_, data_stage_3__1551_, data_stage_3__1550_, data_stage_3__1549_, data_stage_3__1548_, data_stage_3__1547_, data_stage_3__1546_, data_stage_3__1545_, data_stage_3__1544_, data_stage_3__1543_, data_stage_3__1542_, data_stage_3__1541_, data_stage_3__1540_, data_stage_3__1539_, data_stage_3__1538_, data_stage_3__1537_, data_stage_3__1536_, data_stage_3__1535_, data_stage_3__1534_, data_stage_3__1533_, data_stage_3__1532_, data_stage_3__1531_, data_stage_3__1530_, data_stage_3__1529_, data_stage_3__1528_, data_stage_3__1527_, data_stage_3__1526_, data_stage_3__1525_, data_stage_3__1524_, data_stage_3__1523_, data_stage_3__1522_, data_stage_3__1521_, data_stage_3__1520_, data_stage_3__1519_, data_stage_3__1518_, data_stage_3__1517_, data_stage_3__1516_, data_stage_3__1515_, data_stage_3__1514_, data_stage_3__1513_, data_stage_3__1512_, data_stage_3__1511_, data_stage_3__1510_, data_stage_3__1509_, data_stage_3__1508_, data_stage_3__1507_, data_stage_3__1506_, data_stage_3__1505_, data_stage_3__1504_, data_stage_3__1503_, data_stage_3__1502_, data_stage_3__1501_, data_stage_3__1500_, data_stage_3__1499_, data_stage_3__1498_, data_stage_3__1497_, data_stage_3__1496_, data_stage_3__1495_, data_stage_3__1494_, data_stage_3__1493_, data_stage_3__1492_, data_stage_3__1491_, data_stage_3__1490_, data_stage_3__1489_, data_stage_3__1488_, data_stage_3__1487_, data_stage_3__1486_, data_stage_3__1485_, data_stage_3__1484_, data_stage_3__1483_, data_stage_3__1482_, data_stage_3__1481_, data_stage_3__1480_, data_stage_3__1479_, data_stage_3__1478_, data_stage_3__1477_, data_stage_3__1476_, data_stage_3__1475_, data_stage_3__1474_, data_stage_3__1473_, data_stage_3__1472_, data_stage_3__1471_, data_stage_3__1470_, data_stage_3__1469_, data_stage_3__1468_, data_stage_3__1467_, data_stage_3__1466_, data_stage_3__1465_, data_stage_3__1464_, data_stage_3__1463_, data_stage_3__1462_, data_stage_3__1461_, data_stage_3__1460_, data_stage_3__1459_, data_stage_3__1458_, data_stage_3__1457_, data_stage_3__1456_, data_stage_3__1455_, data_stage_3__1454_, data_stage_3__1453_, data_stage_3__1452_, data_stage_3__1451_, data_stage_3__1450_, data_stage_3__1449_, data_stage_3__1448_, data_stage_3__1447_, data_stage_3__1446_, data_stage_3__1445_, data_stage_3__1444_, data_stage_3__1443_, data_stage_3__1442_, data_stage_3__1441_, data_stage_3__1440_, data_stage_3__1439_, data_stage_3__1438_, data_stage_3__1437_, data_stage_3__1436_, data_stage_3__1435_, data_stage_3__1434_, data_stage_3__1433_, data_stage_3__1432_, data_stage_3__1431_, data_stage_3__1430_, data_stage_3__1429_, data_stage_3__1428_, data_stage_3__1427_, data_stage_3__1426_, data_stage_3__1425_, data_stage_3__1424_, data_stage_3__1423_, data_stage_3__1422_, data_stage_3__1421_, data_stage_3__1420_, data_stage_3__1419_, data_stage_3__1418_, data_stage_3__1417_, data_stage_3__1416_, data_stage_3__1415_, data_stage_3__1414_, data_stage_3__1413_, data_stage_3__1412_, data_stage_3__1411_, data_stage_3__1410_, data_stage_3__1409_, data_stage_3__1408_, data_stage_3__1407_, data_stage_3__1406_, data_stage_3__1405_, data_stage_3__1404_, data_stage_3__1403_, data_stage_3__1402_, data_stage_3__1401_, data_stage_3__1400_, data_stage_3__1399_, data_stage_3__1398_, data_stage_3__1397_, data_stage_3__1396_, data_stage_3__1395_, data_stage_3__1394_, data_stage_3__1393_, data_stage_3__1392_, data_stage_3__1391_, data_stage_3__1390_, data_stage_3__1389_, data_stage_3__1388_, data_stage_3__1387_, data_stage_3__1386_, data_stage_3__1385_, data_stage_3__1384_, data_stage_3__1383_, data_stage_3__1382_, data_stage_3__1381_, data_stage_3__1380_, data_stage_3__1379_, data_stage_3__1378_, data_stage_3__1377_, data_stage_3__1376_, data_stage_3__1375_, data_stage_3__1374_, data_stage_3__1373_, data_stage_3__1372_, data_stage_3__1371_, data_stage_3__1370_, data_stage_3__1369_, data_stage_3__1368_, data_stage_3__1367_, data_stage_3__1366_, data_stage_3__1365_, data_stage_3__1364_, data_stage_3__1363_, data_stage_3__1362_, data_stage_3__1361_, data_stage_3__1360_, data_stage_3__1359_, data_stage_3__1358_, data_stage_3__1357_, data_stage_3__1356_, data_stage_3__1355_, data_stage_3__1354_, data_stage_3__1353_, data_stage_3__1352_, data_stage_3__1351_, data_stage_3__1350_, data_stage_3__1349_, data_stage_3__1348_, data_stage_3__1347_, data_stage_3__1346_, data_stage_3__1345_, data_stage_3__1344_, data_stage_3__1343_, data_stage_3__1342_, data_stage_3__1341_, data_stage_3__1340_, data_stage_3__1339_, data_stage_3__1338_, data_stage_3__1337_, data_stage_3__1336_, data_stage_3__1335_, data_stage_3__1334_, data_stage_3__1333_, data_stage_3__1332_, data_stage_3__1331_, data_stage_3__1330_, data_stage_3__1329_, data_stage_3__1328_, data_stage_3__1327_, data_stage_3__1326_, data_stage_3__1325_, data_stage_3__1324_, data_stage_3__1323_, data_stage_3__1322_, data_stage_3__1321_, data_stage_3__1320_, data_stage_3__1319_, data_stage_3__1318_, data_stage_3__1317_, data_stage_3__1316_, data_stage_3__1315_, data_stage_3__1314_, data_stage_3__1313_, data_stage_3__1312_, data_stage_3__1311_, data_stage_3__1310_, data_stage_3__1309_, data_stage_3__1308_, data_stage_3__1307_, data_stage_3__1306_, data_stage_3__1305_, data_stage_3__1304_, data_stage_3__1303_, data_stage_3__1302_, data_stage_3__1301_, data_stage_3__1300_, data_stage_3__1299_, data_stage_3__1298_, data_stage_3__1297_, data_stage_3__1296_, data_stage_3__1295_, data_stage_3__1294_, data_stage_3__1293_, data_stage_3__1292_, data_stage_3__1291_, data_stage_3__1290_, data_stage_3__1289_, data_stage_3__1288_, data_stage_3__1287_, data_stage_3__1286_, data_stage_3__1285_, data_stage_3__1284_, data_stage_3__1283_, data_stage_3__1282_, data_stage_3__1281_, data_stage_3__1280_, data_stage_3__1279_, data_stage_3__1278_, data_stage_3__1277_, data_stage_3__1276_, data_stage_3__1275_, data_stage_3__1274_, data_stage_3__1273_, data_stage_3__1272_, data_stage_3__1271_, data_stage_3__1270_, data_stage_3__1269_, data_stage_3__1268_, data_stage_3__1267_, data_stage_3__1266_, data_stage_3__1265_, data_stage_3__1264_, data_stage_3__1263_, data_stage_3__1262_, data_stage_3__1261_, data_stage_3__1260_, data_stage_3__1259_, data_stage_3__1258_, data_stage_3__1257_, data_stage_3__1256_, data_stage_3__1255_, data_stage_3__1254_, data_stage_3__1253_, data_stage_3__1252_, data_stage_3__1251_, data_stage_3__1250_, data_stage_3__1249_, data_stage_3__1248_, data_stage_3__1247_, data_stage_3__1246_, data_stage_3__1245_, data_stage_3__1244_, data_stage_3__1243_, data_stage_3__1242_, data_stage_3__1241_, data_stage_3__1240_, data_stage_3__1239_, data_stage_3__1238_, data_stage_3__1237_, data_stage_3__1236_, data_stage_3__1235_, data_stage_3__1234_, data_stage_3__1233_, data_stage_3__1232_, data_stage_3__1231_, data_stage_3__1230_, data_stage_3__1229_, data_stage_3__1228_, data_stage_3__1227_, data_stage_3__1226_, data_stage_3__1225_, data_stage_3__1224_, data_stage_3__1223_, data_stage_3__1222_, data_stage_3__1221_, data_stage_3__1220_, data_stage_3__1219_, data_stage_3__1218_, data_stage_3__1217_, data_stage_3__1216_, data_stage_3__1215_, data_stage_3__1214_, data_stage_3__1213_, data_stage_3__1212_, data_stage_3__1211_, data_stage_3__1210_, data_stage_3__1209_, data_stage_3__1208_, data_stage_3__1207_, data_stage_3__1206_, data_stage_3__1205_, data_stage_3__1204_, data_stage_3__1203_, data_stage_3__1202_, data_stage_3__1201_, data_stage_3__1200_, data_stage_3__1199_, data_stage_3__1198_, data_stage_3__1197_, data_stage_3__1196_, data_stage_3__1195_, data_stage_3__1194_, data_stage_3__1193_, data_stage_3__1192_, data_stage_3__1191_, data_stage_3__1190_, data_stage_3__1189_, data_stage_3__1188_, data_stage_3__1187_, data_stage_3__1186_, data_stage_3__1185_, data_stage_3__1184_, data_stage_3__1183_, data_stage_3__1182_, data_stage_3__1181_, data_stage_3__1180_, data_stage_3__1179_, data_stage_3__1178_, data_stage_3__1177_, data_stage_3__1176_, data_stage_3__1175_, data_stage_3__1174_, data_stage_3__1173_, data_stage_3__1172_, data_stage_3__1171_, data_stage_3__1170_, data_stage_3__1169_, data_stage_3__1168_, data_stage_3__1167_, data_stage_3__1166_, data_stage_3__1165_, data_stage_3__1164_, data_stage_3__1163_, data_stage_3__1162_, data_stage_3__1161_, data_stage_3__1160_, data_stage_3__1159_, data_stage_3__1158_, data_stage_3__1157_, data_stage_3__1156_, data_stage_3__1155_, data_stage_3__1154_, data_stage_3__1153_, data_stage_3__1152_, data_stage_3__1151_, data_stage_3__1150_, data_stage_3__1149_, data_stage_3__1148_, data_stage_3__1147_, data_stage_3__1146_, data_stage_3__1145_, data_stage_3__1144_, data_stage_3__1143_, data_stage_3__1142_, data_stage_3__1141_, data_stage_3__1140_, data_stage_3__1139_, data_stage_3__1138_, data_stage_3__1137_, data_stage_3__1136_, data_stage_3__1135_, data_stage_3__1134_, data_stage_3__1133_, data_stage_3__1132_, data_stage_3__1131_, data_stage_3__1130_, data_stage_3__1129_, data_stage_3__1128_, data_stage_3__1127_, data_stage_3__1126_, data_stage_3__1125_, data_stage_3__1124_, data_stage_3__1123_, data_stage_3__1122_, data_stage_3__1121_, data_stage_3__1120_, data_stage_3__1119_, data_stage_3__1118_, data_stage_3__1117_, data_stage_3__1116_, data_stage_3__1115_, data_stage_3__1114_, data_stage_3__1113_, data_stage_3__1112_, data_stage_3__1111_, data_stage_3__1110_, data_stage_3__1109_, data_stage_3__1108_, data_stage_3__1107_, data_stage_3__1106_, data_stage_3__1105_, data_stage_3__1104_, data_stage_3__1103_, data_stage_3__1102_, data_stage_3__1101_, data_stage_3__1100_, data_stage_3__1099_, data_stage_3__1098_, data_stage_3__1097_, data_stage_3__1096_, data_stage_3__1095_, data_stage_3__1094_, data_stage_3__1093_, data_stage_3__1092_, data_stage_3__1091_, data_stage_3__1090_, data_stage_3__1089_, data_stage_3__1088_, data_stage_3__1087_, data_stage_3__1086_, data_stage_3__1085_, data_stage_3__1084_, data_stage_3__1083_, data_stage_3__1082_, data_stage_3__1081_, data_stage_3__1080_, data_stage_3__1079_, data_stage_3__1078_, data_stage_3__1077_, data_stage_3__1076_, data_stage_3__1075_, data_stage_3__1074_, data_stage_3__1073_, data_stage_3__1072_, data_stage_3__1071_, data_stage_3__1070_, data_stage_3__1069_, data_stage_3__1068_, data_stage_3__1067_, data_stage_3__1066_, data_stage_3__1065_, data_stage_3__1064_, data_stage_3__1063_, data_stage_3__1062_, data_stage_3__1061_, data_stage_3__1060_, data_stage_3__1059_, data_stage_3__1058_, data_stage_3__1057_, data_stage_3__1056_, data_stage_3__1055_, data_stage_3__1054_, data_stage_3__1053_, data_stage_3__1052_, data_stage_3__1051_, data_stage_3__1050_, data_stage_3__1049_, data_stage_3__1048_, data_stage_3__1047_, data_stage_3__1046_, data_stage_3__1045_, data_stage_3__1044_, data_stage_3__1043_, data_stage_3__1042_, data_stage_3__1041_, data_stage_3__1040_, data_stage_3__1039_, data_stage_3__1038_, data_stage_3__1037_, data_stage_3__1036_, data_stage_3__1035_, data_stage_3__1034_, data_stage_3__1033_, data_stage_3__1032_, data_stage_3__1031_, data_stage_3__1030_, data_stage_3__1029_, data_stage_3__1028_, data_stage_3__1027_, data_stage_3__1026_, data_stage_3__1025_, data_stage_3__1024_ }),
    .swap_i(sel_i[3]),
    .data_o({ data_stage_4__2047_, data_stage_4__2046_, data_stage_4__2045_, data_stage_4__2044_, data_stage_4__2043_, data_stage_4__2042_, data_stage_4__2041_, data_stage_4__2040_, data_stage_4__2039_, data_stage_4__2038_, data_stage_4__2037_, data_stage_4__2036_, data_stage_4__2035_, data_stage_4__2034_, data_stage_4__2033_, data_stage_4__2032_, data_stage_4__2031_, data_stage_4__2030_, data_stage_4__2029_, data_stage_4__2028_, data_stage_4__2027_, data_stage_4__2026_, data_stage_4__2025_, data_stage_4__2024_, data_stage_4__2023_, data_stage_4__2022_, data_stage_4__2021_, data_stage_4__2020_, data_stage_4__2019_, data_stage_4__2018_, data_stage_4__2017_, data_stage_4__2016_, data_stage_4__2015_, data_stage_4__2014_, data_stage_4__2013_, data_stage_4__2012_, data_stage_4__2011_, data_stage_4__2010_, data_stage_4__2009_, data_stage_4__2008_, data_stage_4__2007_, data_stage_4__2006_, data_stage_4__2005_, data_stage_4__2004_, data_stage_4__2003_, data_stage_4__2002_, data_stage_4__2001_, data_stage_4__2000_, data_stage_4__1999_, data_stage_4__1998_, data_stage_4__1997_, data_stage_4__1996_, data_stage_4__1995_, data_stage_4__1994_, data_stage_4__1993_, data_stage_4__1992_, data_stage_4__1991_, data_stage_4__1990_, data_stage_4__1989_, data_stage_4__1988_, data_stage_4__1987_, data_stage_4__1986_, data_stage_4__1985_, data_stage_4__1984_, data_stage_4__1983_, data_stage_4__1982_, data_stage_4__1981_, data_stage_4__1980_, data_stage_4__1979_, data_stage_4__1978_, data_stage_4__1977_, data_stage_4__1976_, data_stage_4__1975_, data_stage_4__1974_, data_stage_4__1973_, data_stage_4__1972_, data_stage_4__1971_, data_stage_4__1970_, data_stage_4__1969_, data_stage_4__1968_, data_stage_4__1967_, data_stage_4__1966_, data_stage_4__1965_, data_stage_4__1964_, data_stage_4__1963_, data_stage_4__1962_, data_stage_4__1961_, data_stage_4__1960_, data_stage_4__1959_, data_stage_4__1958_, data_stage_4__1957_, data_stage_4__1956_, data_stage_4__1955_, data_stage_4__1954_, data_stage_4__1953_, data_stage_4__1952_, data_stage_4__1951_, data_stage_4__1950_, data_stage_4__1949_, data_stage_4__1948_, data_stage_4__1947_, data_stage_4__1946_, data_stage_4__1945_, data_stage_4__1944_, data_stage_4__1943_, data_stage_4__1942_, data_stage_4__1941_, data_stage_4__1940_, data_stage_4__1939_, data_stage_4__1938_, data_stage_4__1937_, data_stage_4__1936_, data_stage_4__1935_, data_stage_4__1934_, data_stage_4__1933_, data_stage_4__1932_, data_stage_4__1931_, data_stage_4__1930_, data_stage_4__1929_, data_stage_4__1928_, data_stage_4__1927_, data_stage_4__1926_, data_stage_4__1925_, data_stage_4__1924_, data_stage_4__1923_, data_stage_4__1922_, data_stage_4__1921_, data_stage_4__1920_, data_stage_4__1919_, data_stage_4__1918_, data_stage_4__1917_, data_stage_4__1916_, data_stage_4__1915_, data_stage_4__1914_, data_stage_4__1913_, data_stage_4__1912_, data_stage_4__1911_, data_stage_4__1910_, data_stage_4__1909_, data_stage_4__1908_, data_stage_4__1907_, data_stage_4__1906_, data_stage_4__1905_, data_stage_4__1904_, data_stage_4__1903_, data_stage_4__1902_, data_stage_4__1901_, data_stage_4__1900_, data_stage_4__1899_, data_stage_4__1898_, data_stage_4__1897_, data_stage_4__1896_, data_stage_4__1895_, data_stage_4__1894_, data_stage_4__1893_, data_stage_4__1892_, data_stage_4__1891_, data_stage_4__1890_, data_stage_4__1889_, data_stage_4__1888_, data_stage_4__1887_, data_stage_4__1886_, data_stage_4__1885_, data_stage_4__1884_, data_stage_4__1883_, data_stage_4__1882_, data_stage_4__1881_, data_stage_4__1880_, data_stage_4__1879_, data_stage_4__1878_, data_stage_4__1877_, data_stage_4__1876_, data_stage_4__1875_, data_stage_4__1874_, data_stage_4__1873_, data_stage_4__1872_, data_stage_4__1871_, data_stage_4__1870_, data_stage_4__1869_, data_stage_4__1868_, data_stage_4__1867_, data_stage_4__1866_, data_stage_4__1865_, data_stage_4__1864_, data_stage_4__1863_, data_stage_4__1862_, data_stage_4__1861_, data_stage_4__1860_, data_stage_4__1859_, data_stage_4__1858_, data_stage_4__1857_, data_stage_4__1856_, data_stage_4__1855_, data_stage_4__1854_, data_stage_4__1853_, data_stage_4__1852_, data_stage_4__1851_, data_stage_4__1850_, data_stage_4__1849_, data_stage_4__1848_, data_stage_4__1847_, data_stage_4__1846_, data_stage_4__1845_, data_stage_4__1844_, data_stage_4__1843_, data_stage_4__1842_, data_stage_4__1841_, data_stage_4__1840_, data_stage_4__1839_, data_stage_4__1838_, data_stage_4__1837_, data_stage_4__1836_, data_stage_4__1835_, data_stage_4__1834_, data_stage_4__1833_, data_stage_4__1832_, data_stage_4__1831_, data_stage_4__1830_, data_stage_4__1829_, data_stage_4__1828_, data_stage_4__1827_, data_stage_4__1826_, data_stage_4__1825_, data_stage_4__1824_, data_stage_4__1823_, data_stage_4__1822_, data_stage_4__1821_, data_stage_4__1820_, data_stage_4__1819_, data_stage_4__1818_, data_stage_4__1817_, data_stage_4__1816_, data_stage_4__1815_, data_stage_4__1814_, data_stage_4__1813_, data_stage_4__1812_, data_stage_4__1811_, data_stage_4__1810_, data_stage_4__1809_, data_stage_4__1808_, data_stage_4__1807_, data_stage_4__1806_, data_stage_4__1805_, data_stage_4__1804_, data_stage_4__1803_, data_stage_4__1802_, data_stage_4__1801_, data_stage_4__1800_, data_stage_4__1799_, data_stage_4__1798_, data_stage_4__1797_, data_stage_4__1796_, data_stage_4__1795_, data_stage_4__1794_, data_stage_4__1793_, data_stage_4__1792_, data_stage_4__1791_, data_stage_4__1790_, data_stage_4__1789_, data_stage_4__1788_, data_stage_4__1787_, data_stage_4__1786_, data_stage_4__1785_, data_stage_4__1784_, data_stage_4__1783_, data_stage_4__1782_, data_stage_4__1781_, data_stage_4__1780_, data_stage_4__1779_, data_stage_4__1778_, data_stage_4__1777_, data_stage_4__1776_, data_stage_4__1775_, data_stage_4__1774_, data_stage_4__1773_, data_stage_4__1772_, data_stage_4__1771_, data_stage_4__1770_, data_stage_4__1769_, data_stage_4__1768_, data_stage_4__1767_, data_stage_4__1766_, data_stage_4__1765_, data_stage_4__1764_, data_stage_4__1763_, data_stage_4__1762_, data_stage_4__1761_, data_stage_4__1760_, data_stage_4__1759_, data_stage_4__1758_, data_stage_4__1757_, data_stage_4__1756_, data_stage_4__1755_, data_stage_4__1754_, data_stage_4__1753_, data_stage_4__1752_, data_stage_4__1751_, data_stage_4__1750_, data_stage_4__1749_, data_stage_4__1748_, data_stage_4__1747_, data_stage_4__1746_, data_stage_4__1745_, data_stage_4__1744_, data_stage_4__1743_, data_stage_4__1742_, data_stage_4__1741_, data_stage_4__1740_, data_stage_4__1739_, data_stage_4__1738_, data_stage_4__1737_, data_stage_4__1736_, data_stage_4__1735_, data_stage_4__1734_, data_stage_4__1733_, data_stage_4__1732_, data_stage_4__1731_, data_stage_4__1730_, data_stage_4__1729_, data_stage_4__1728_, data_stage_4__1727_, data_stage_4__1726_, data_stage_4__1725_, data_stage_4__1724_, data_stage_4__1723_, data_stage_4__1722_, data_stage_4__1721_, data_stage_4__1720_, data_stage_4__1719_, data_stage_4__1718_, data_stage_4__1717_, data_stage_4__1716_, data_stage_4__1715_, data_stage_4__1714_, data_stage_4__1713_, data_stage_4__1712_, data_stage_4__1711_, data_stage_4__1710_, data_stage_4__1709_, data_stage_4__1708_, data_stage_4__1707_, data_stage_4__1706_, data_stage_4__1705_, data_stage_4__1704_, data_stage_4__1703_, data_stage_4__1702_, data_stage_4__1701_, data_stage_4__1700_, data_stage_4__1699_, data_stage_4__1698_, data_stage_4__1697_, data_stage_4__1696_, data_stage_4__1695_, data_stage_4__1694_, data_stage_4__1693_, data_stage_4__1692_, data_stage_4__1691_, data_stage_4__1690_, data_stage_4__1689_, data_stage_4__1688_, data_stage_4__1687_, data_stage_4__1686_, data_stage_4__1685_, data_stage_4__1684_, data_stage_4__1683_, data_stage_4__1682_, data_stage_4__1681_, data_stage_4__1680_, data_stage_4__1679_, data_stage_4__1678_, data_stage_4__1677_, data_stage_4__1676_, data_stage_4__1675_, data_stage_4__1674_, data_stage_4__1673_, data_stage_4__1672_, data_stage_4__1671_, data_stage_4__1670_, data_stage_4__1669_, data_stage_4__1668_, data_stage_4__1667_, data_stage_4__1666_, data_stage_4__1665_, data_stage_4__1664_, data_stage_4__1663_, data_stage_4__1662_, data_stage_4__1661_, data_stage_4__1660_, data_stage_4__1659_, data_stage_4__1658_, data_stage_4__1657_, data_stage_4__1656_, data_stage_4__1655_, data_stage_4__1654_, data_stage_4__1653_, data_stage_4__1652_, data_stage_4__1651_, data_stage_4__1650_, data_stage_4__1649_, data_stage_4__1648_, data_stage_4__1647_, data_stage_4__1646_, data_stage_4__1645_, data_stage_4__1644_, data_stage_4__1643_, data_stage_4__1642_, data_stage_4__1641_, data_stage_4__1640_, data_stage_4__1639_, data_stage_4__1638_, data_stage_4__1637_, data_stage_4__1636_, data_stage_4__1635_, data_stage_4__1634_, data_stage_4__1633_, data_stage_4__1632_, data_stage_4__1631_, data_stage_4__1630_, data_stage_4__1629_, data_stage_4__1628_, data_stage_4__1627_, data_stage_4__1626_, data_stage_4__1625_, data_stage_4__1624_, data_stage_4__1623_, data_stage_4__1622_, data_stage_4__1621_, data_stage_4__1620_, data_stage_4__1619_, data_stage_4__1618_, data_stage_4__1617_, data_stage_4__1616_, data_stage_4__1615_, data_stage_4__1614_, data_stage_4__1613_, data_stage_4__1612_, data_stage_4__1611_, data_stage_4__1610_, data_stage_4__1609_, data_stage_4__1608_, data_stage_4__1607_, data_stage_4__1606_, data_stage_4__1605_, data_stage_4__1604_, data_stage_4__1603_, data_stage_4__1602_, data_stage_4__1601_, data_stage_4__1600_, data_stage_4__1599_, data_stage_4__1598_, data_stage_4__1597_, data_stage_4__1596_, data_stage_4__1595_, data_stage_4__1594_, data_stage_4__1593_, data_stage_4__1592_, data_stage_4__1591_, data_stage_4__1590_, data_stage_4__1589_, data_stage_4__1588_, data_stage_4__1587_, data_stage_4__1586_, data_stage_4__1585_, data_stage_4__1584_, data_stage_4__1583_, data_stage_4__1582_, data_stage_4__1581_, data_stage_4__1580_, data_stage_4__1579_, data_stage_4__1578_, data_stage_4__1577_, data_stage_4__1576_, data_stage_4__1575_, data_stage_4__1574_, data_stage_4__1573_, data_stage_4__1572_, data_stage_4__1571_, data_stage_4__1570_, data_stage_4__1569_, data_stage_4__1568_, data_stage_4__1567_, data_stage_4__1566_, data_stage_4__1565_, data_stage_4__1564_, data_stage_4__1563_, data_stage_4__1562_, data_stage_4__1561_, data_stage_4__1560_, data_stage_4__1559_, data_stage_4__1558_, data_stage_4__1557_, data_stage_4__1556_, data_stage_4__1555_, data_stage_4__1554_, data_stage_4__1553_, data_stage_4__1552_, data_stage_4__1551_, data_stage_4__1550_, data_stage_4__1549_, data_stage_4__1548_, data_stage_4__1547_, data_stage_4__1546_, data_stage_4__1545_, data_stage_4__1544_, data_stage_4__1543_, data_stage_4__1542_, data_stage_4__1541_, data_stage_4__1540_, data_stage_4__1539_, data_stage_4__1538_, data_stage_4__1537_, data_stage_4__1536_, data_stage_4__1535_, data_stage_4__1534_, data_stage_4__1533_, data_stage_4__1532_, data_stage_4__1531_, data_stage_4__1530_, data_stage_4__1529_, data_stage_4__1528_, data_stage_4__1527_, data_stage_4__1526_, data_stage_4__1525_, data_stage_4__1524_, data_stage_4__1523_, data_stage_4__1522_, data_stage_4__1521_, data_stage_4__1520_, data_stage_4__1519_, data_stage_4__1518_, data_stage_4__1517_, data_stage_4__1516_, data_stage_4__1515_, data_stage_4__1514_, data_stage_4__1513_, data_stage_4__1512_, data_stage_4__1511_, data_stage_4__1510_, data_stage_4__1509_, data_stage_4__1508_, data_stage_4__1507_, data_stage_4__1506_, data_stage_4__1505_, data_stage_4__1504_, data_stage_4__1503_, data_stage_4__1502_, data_stage_4__1501_, data_stage_4__1500_, data_stage_4__1499_, data_stage_4__1498_, data_stage_4__1497_, data_stage_4__1496_, data_stage_4__1495_, data_stage_4__1494_, data_stage_4__1493_, data_stage_4__1492_, data_stage_4__1491_, data_stage_4__1490_, data_stage_4__1489_, data_stage_4__1488_, data_stage_4__1487_, data_stage_4__1486_, data_stage_4__1485_, data_stage_4__1484_, data_stage_4__1483_, data_stage_4__1482_, data_stage_4__1481_, data_stage_4__1480_, data_stage_4__1479_, data_stage_4__1478_, data_stage_4__1477_, data_stage_4__1476_, data_stage_4__1475_, data_stage_4__1474_, data_stage_4__1473_, data_stage_4__1472_, data_stage_4__1471_, data_stage_4__1470_, data_stage_4__1469_, data_stage_4__1468_, data_stage_4__1467_, data_stage_4__1466_, data_stage_4__1465_, data_stage_4__1464_, data_stage_4__1463_, data_stage_4__1462_, data_stage_4__1461_, data_stage_4__1460_, data_stage_4__1459_, data_stage_4__1458_, data_stage_4__1457_, data_stage_4__1456_, data_stage_4__1455_, data_stage_4__1454_, data_stage_4__1453_, data_stage_4__1452_, data_stage_4__1451_, data_stage_4__1450_, data_stage_4__1449_, data_stage_4__1448_, data_stage_4__1447_, data_stage_4__1446_, data_stage_4__1445_, data_stage_4__1444_, data_stage_4__1443_, data_stage_4__1442_, data_stage_4__1441_, data_stage_4__1440_, data_stage_4__1439_, data_stage_4__1438_, data_stage_4__1437_, data_stage_4__1436_, data_stage_4__1435_, data_stage_4__1434_, data_stage_4__1433_, data_stage_4__1432_, data_stage_4__1431_, data_stage_4__1430_, data_stage_4__1429_, data_stage_4__1428_, data_stage_4__1427_, data_stage_4__1426_, data_stage_4__1425_, data_stage_4__1424_, data_stage_4__1423_, data_stage_4__1422_, data_stage_4__1421_, data_stage_4__1420_, data_stage_4__1419_, data_stage_4__1418_, data_stage_4__1417_, data_stage_4__1416_, data_stage_4__1415_, data_stage_4__1414_, data_stage_4__1413_, data_stage_4__1412_, data_stage_4__1411_, data_stage_4__1410_, data_stage_4__1409_, data_stage_4__1408_, data_stage_4__1407_, data_stage_4__1406_, data_stage_4__1405_, data_stage_4__1404_, data_stage_4__1403_, data_stage_4__1402_, data_stage_4__1401_, data_stage_4__1400_, data_stage_4__1399_, data_stage_4__1398_, data_stage_4__1397_, data_stage_4__1396_, data_stage_4__1395_, data_stage_4__1394_, data_stage_4__1393_, data_stage_4__1392_, data_stage_4__1391_, data_stage_4__1390_, data_stage_4__1389_, data_stage_4__1388_, data_stage_4__1387_, data_stage_4__1386_, data_stage_4__1385_, data_stage_4__1384_, data_stage_4__1383_, data_stage_4__1382_, data_stage_4__1381_, data_stage_4__1380_, data_stage_4__1379_, data_stage_4__1378_, data_stage_4__1377_, data_stage_4__1376_, data_stage_4__1375_, data_stage_4__1374_, data_stage_4__1373_, data_stage_4__1372_, data_stage_4__1371_, data_stage_4__1370_, data_stage_4__1369_, data_stage_4__1368_, data_stage_4__1367_, data_stage_4__1366_, data_stage_4__1365_, data_stage_4__1364_, data_stage_4__1363_, data_stage_4__1362_, data_stage_4__1361_, data_stage_4__1360_, data_stage_4__1359_, data_stage_4__1358_, data_stage_4__1357_, data_stage_4__1356_, data_stage_4__1355_, data_stage_4__1354_, data_stage_4__1353_, data_stage_4__1352_, data_stage_4__1351_, data_stage_4__1350_, data_stage_4__1349_, data_stage_4__1348_, data_stage_4__1347_, data_stage_4__1346_, data_stage_4__1345_, data_stage_4__1344_, data_stage_4__1343_, data_stage_4__1342_, data_stage_4__1341_, data_stage_4__1340_, data_stage_4__1339_, data_stage_4__1338_, data_stage_4__1337_, data_stage_4__1336_, data_stage_4__1335_, data_stage_4__1334_, data_stage_4__1333_, data_stage_4__1332_, data_stage_4__1331_, data_stage_4__1330_, data_stage_4__1329_, data_stage_4__1328_, data_stage_4__1327_, data_stage_4__1326_, data_stage_4__1325_, data_stage_4__1324_, data_stage_4__1323_, data_stage_4__1322_, data_stage_4__1321_, data_stage_4__1320_, data_stage_4__1319_, data_stage_4__1318_, data_stage_4__1317_, data_stage_4__1316_, data_stage_4__1315_, data_stage_4__1314_, data_stage_4__1313_, data_stage_4__1312_, data_stage_4__1311_, data_stage_4__1310_, data_stage_4__1309_, data_stage_4__1308_, data_stage_4__1307_, data_stage_4__1306_, data_stage_4__1305_, data_stage_4__1304_, data_stage_4__1303_, data_stage_4__1302_, data_stage_4__1301_, data_stage_4__1300_, data_stage_4__1299_, data_stage_4__1298_, data_stage_4__1297_, data_stage_4__1296_, data_stage_4__1295_, data_stage_4__1294_, data_stage_4__1293_, data_stage_4__1292_, data_stage_4__1291_, data_stage_4__1290_, data_stage_4__1289_, data_stage_4__1288_, data_stage_4__1287_, data_stage_4__1286_, data_stage_4__1285_, data_stage_4__1284_, data_stage_4__1283_, data_stage_4__1282_, data_stage_4__1281_, data_stage_4__1280_, data_stage_4__1279_, data_stage_4__1278_, data_stage_4__1277_, data_stage_4__1276_, data_stage_4__1275_, data_stage_4__1274_, data_stage_4__1273_, data_stage_4__1272_, data_stage_4__1271_, data_stage_4__1270_, data_stage_4__1269_, data_stage_4__1268_, data_stage_4__1267_, data_stage_4__1266_, data_stage_4__1265_, data_stage_4__1264_, data_stage_4__1263_, data_stage_4__1262_, data_stage_4__1261_, data_stage_4__1260_, data_stage_4__1259_, data_stage_4__1258_, data_stage_4__1257_, data_stage_4__1256_, data_stage_4__1255_, data_stage_4__1254_, data_stage_4__1253_, data_stage_4__1252_, data_stage_4__1251_, data_stage_4__1250_, data_stage_4__1249_, data_stage_4__1248_, data_stage_4__1247_, data_stage_4__1246_, data_stage_4__1245_, data_stage_4__1244_, data_stage_4__1243_, data_stage_4__1242_, data_stage_4__1241_, data_stage_4__1240_, data_stage_4__1239_, data_stage_4__1238_, data_stage_4__1237_, data_stage_4__1236_, data_stage_4__1235_, data_stage_4__1234_, data_stage_4__1233_, data_stage_4__1232_, data_stage_4__1231_, data_stage_4__1230_, data_stage_4__1229_, data_stage_4__1228_, data_stage_4__1227_, data_stage_4__1226_, data_stage_4__1225_, data_stage_4__1224_, data_stage_4__1223_, data_stage_4__1222_, data_stage_4__1221_, data_stage_4__1220_, data_stage_4__1219_, data_stage_4__1218_, data_stage_4__1217_, data_stage_4__1216_, data_stage_4__1215_, data_stage_4__1214_, data_stage_4__1213_, data_stage_4__1212_, data_stage_4__1211_, data_stage_4__1210_, data_stage_4__1209_, data_stage_4__1208_, data_stage_4__1207_, data_stage_4__1206_, data_stage_4__1205_, data_stage_4__1204_, data_stage_4__1203_, data_stage_4__1202_, data_stage_4__1201_, data_stage_4__1200_, data_stage_4__1199_, data_stage_4__1198_, data_stage_4__1197_, data_stage_4__1196_, data_stage_4__1195_, data_stage_4__1194_, data_stage_4__1193_, data_stage_4__1192_, data_stage_4__1191_, data_stage_4__1190_, data_stage_4__1189_, data_stage_4__1188_, data_stage_4__1187_, data_stage_4__1186_, data_stage_4__1185_, data_stage_4__1184_, data_stage_4__1183_, data_stage_4__1182_, data_stage_4__1181_, data_stage_4__1180_, data_stage_4__1179_, data_stage_4__1178_, data_stage_4__1177_, data_stage_4__1176_, data_stage_4__1175_, data_stage_4__1174_, data_stage_4__1173_, data_stage_4__1172_, data_stage_4__1171_, data_stage_4__1170_, data_stage_4__1169_, data_stage_4__1168_, data_stage_4__1167_, data_stage_4__1166_, data_stage_4__1165_, data_stage_4__1164_, data_stage_4__1163_, data_stage_4__1162_, data_stage_4__1161_, data_stage_4__1160_, data_stage_4__1159_, data_stage_4__1158_, data_stage_4__1157_, data_stage_4__1156_, data_stage_4__1155_, data_stage_4__1154_, data_stage_4__1153_, data_stage_4__1152_, data_stage_4__1151_, data_stage_4__1150_, data_stage_4__1149_, data_stage_4__1148_, data_stage_4__1147_, data_stage_4__1146_, data_stage_4__1145_, data_stage_4__1144_, data_stage_4__1143_, data_stage_4__1142_, data_stage_4__1141_, data_stage_4__1140_, data_stage_4__1139_, data_stage_4__1138_, data_stage_4__1137_, data_stage_4__1136_, data_stage_4__1135_, data_stage_4__1134_, data_stage_4__1133_, data_stage_4__1132_, data_stage_4__1131_, data_stage_4__1130_, data_stage_4__1129_, data_stage_4__1128_, data_stage_4__1127_, data_stage_4__1126_, data_stage_4__1125_, data_stage_4__1124_, data_stage_4__1123_, data_stage_4__1122_, data_stage_4__1121_, data_stage_4__1120_, data_stage_4__1119_, data_stage_4__1118_, data_stage_4__1117_, data_stage_4__1116_, data_stage_4__1115_, data_stage_4__1114_, data_stage_4__1113_, data_stage_4__1112_, data_stage_4__1111_, data_stage_4__1110_, data_stage_4__1109_, data_stage_4__1108_, data_stage_4__1107_, data_stage_4__1106_, data_stage_4__1105_, data_stage_4__1104_, data_stage_4__1103_, data_stage_4__1102_, data_stage_4__1101_, data_stage_4__1100_, data_stage_4__1099_, data_stage_4__1098_, data_stage_4__1097_, data_stage_4__1096_, data_stage_4__1095_, data_stage_4__1094_, data_stage_4__1093_, data_stage_4__1092_, data_stage_4__1091_, data_stage_4__1090_, data_stage_4__1089_, data_stage_4__1088_, data_stage_4__1087_, data_stage_4__1086_, data_stage_4__1085_, data_stage_4__1084_, data_stage_4__1083_, data_stage_4__1082_, data_stage_4__1081_, data_stage_4__1080_, data_stage_4__1079_, data_stage_4__1078_, data_stage_4__1077_, data_stage_4__1076_, data_stage_4__1075_, data_stage_4__1074_, data_stage_4__1073_, data_stage_4__1072_, data_stage_4__1071_, data_stage_4__1070_, data_stage_4__1069_, data_stage_4__1068_, data_stage_4__1067_, data_stage_4__1066_, data_stage_4__1065_, data_stage_4__1064_, data_stage_4__1063_, data_stage_4__1062_, data_stage_4__1061_, data_stage_4__1060_, data_stage_4__1059_, data_stage_4__1058_, data_stage_4__1057_, data_stage_4__1056_, data_stage_4__1055_, data_stage_4__1054_, data_stage_4__1053_, data_stage_4__1052_, data_stage_4__1051_, data_stage_4__1050_, data_stage_4__1049_, data_stage_4__1048_, data_stage_4__1047_, data_stage_4__1046_, data_stage_4__1045_, data_stage_4__1044_, data_stage_4__1043_, data_stage_4__1042_, data_stage_4__1041_, data_stage_4__1040_, data_stage_4__1039_, data_stage_4__1038_, data_stage_4__1037_, data_stage_4__1036_, data_stage_4__1035_, data_stage_4__1034_, data_stage_4__1033_, data_stage_4__1032_, data_stage_4__1031_, data_stage_4__1030_, data_stage_4__1029_, data_stage_4__1028_, data_stage_4__1027_, data_stage_4__1026_, data_stage_4__1025_, data_stage_4__1024_ })
  );


  bsg_swap_width_p512
  mux_stage_3__mux_swap_2__swap_inst
  (
    .data_i({ data_stage_3__3071_, data_stage_3__3070_, data_stage_3__3069_, data_stage_3__3068_, data_stage_3__3067_, data_stage_3__3066_, data_stage_3__3065_, data_stage_3__3064_, data_stage_3__3063_, data_stage_3__3062_, data_stage_3__3061_, data_stage_3__3060_, data_stage_3__3059_, data_stage_3__3058_, data_stage_3__3057_, data_stage_3__3056_, data_stage_3__3055_, data_stage_3__3054_, data_stage_3__3053_, data_stage_3__3052_, data_stage_3__3051_, data_stage_3__3050_, data_stage_3__3049_, data_stage_3__3048_, data_stage_3__3047_, data_stage_3__3046_, data_stage_3__3045_, data_stage_3__3044_, data_stage_3__3043_, data_stage_3__3042_, data_stage_3__3041_, data_stage_3__3040_, data_stage_3__3039_, data_stage_3__3038_, data_stage_3__3037_, data_stage_3__3036_, data_stage_3__3035_, data_stage_3__3034_, data_stage_3__3033_, data_stage_3__3032_, data_stage_3__3031_, data_stage_3__3030_, data_stage_3__3029_, data_stage_3__3028_, data_stage_3__3027_, data_stage_3__3026_, data_stage_3__3025_, data_stage_3__3024_, data_stage_3__3023_, data_stage_3__3022_, data_stage_3__3021_, data_stage_3__3020_, data_stage_3__3019_, data_stage_3__3018_, data_stage_3__3017_, data_stage_3__3016_, data_stage_3__3015_, data_stage_3__3014_, data_stage_3__3013_, data_stage_3__3012_, data_stage_3__3011_, data_stage_3__3010_, data_stage_3__3009_, data_stage_3__3008_, data_stage_3__3007_, data_stage_3__3006_, data_stage_3__3005_, data_stage_3__3004_, data_stage_3__3003_, data_stage_3__3002_, data_stage_3__3001_, data_stage_3__3000_, data_stage_3__2999_, data_stage_3__2998_, data_stage_3__2997_, data_stage_3__2996_, data_stage_3__2995_, data_stage_3__2994_, data_stage_3__2993_, data_stage_3__2992_, data_stage_3__2991_, data_stage_3__2990_, data_stage_3__2989_, data_stage_3__2988_, data_stage_3__2987_, data_stage_3__2986_, data_stage_3__2985_, data_stage_3__2984_, data_stage_3__2983_, data_stage_3__2982_, data_stage_3__2981_, data_stage_3__2980_, data_stage_3__2979_, data_stage_3__2978_, data_stage_3__2977_, data_stage_3__2976_, data_stage_3__2975_, data_stage_3__2974_, data_stage_3__2973_, data_stage_3__2972_, data_stage_3__2971_, data_stage_3__2970_, data_stage_3__2969_, data_stage_3__2968_, data_stage_3__2967_, data_stage_3__2966_, data_stage_3__2965_, data_stage_3__2964_, data_stage_3__2963_, data_stage_3__2962_, data_stage_3__2961_, data_stage_3__2960_, data_stage_3__2959_, data_stage_3__2958_, data_stage_3__2957_, data_stage_3__2956_, data_stage_3__2955_, data_stage_3__2954_, data_stage_3__2953_, data_stage_3__2952_, data_stage_3__2951_, data_stage_3__2950_, data_stage_3__2949_, data_stage_3__2948_, data_stage_3__2947_, data_stage_3__2946_, data_stage_3__2945_, data_stage_3__2944_, data_stage_3__2943_, data_stage_3__2942_, data_stage_3__2941_, data_stage_3__2940_, data_stage_3__2939_, data_stage_3__2938_, data_stage_3__2937_, data_stage_3__2936_, data_stage_3__2935_, data_stage_3__2934_, data_stage_3__2933_, data_stage_3__2932_, data_stage_3__2931_, data_stage_3__2930_, data_stage_3__2929_, data_stage_3__2928_, data_stage_3__2927_, data_stage_3__2926_, data_stage_3__2925_, data_stage_3__2924_, data_stage_3__2923_, data_stage_3__2922_, data_stage_3__2921_, data_stage_3__2920_, data_stage_3__2919_, data_stage_3__2918_, data_stage_3__2917_, data_stage_3__2916_, data_stage_3__2915_, data_stage_3__2914_, data_stage_3__2913_, data_stage_3__2912_, data_stage_3__2911_, data_stage_3__2910_, data_stage_3__2909_, data_stage_3__2908_, data_stage_3__2907_, data_stage_3__2906_, data_stage_3__2905_, data_stage_3__2904_, data_stage_3__2903_, data_stage_3__2902_, data_stage_3__2901_, data_stage_3__2900_, data_stage_3__2899_, data_stage_3__2898_, data_stage_3__2897_, data_stage_3__2896_, data_stage_3__2895_, data_stage_3__2894_, data_stage_3__2893_, data_stage_3__2892_, data_stage_3__2891_, data_stage_3__2890_, data_stage_3__2889_, data_stage_3__2888_, data_stage_3__2887_, data_stage_3__2886_, data_stage_3__2885_, data_stage_3__2884_, data_stage_3__2883_, data_stage_3__2882_, data_stage_3__2881_, data_stage_3__2880_, data_stage_3__2879_, data_stage_3__2878_, data_stage_3__2877_, data_stage_3__2876_, data_stage_3__2875_, data_stage_3__2874_, data_stage_3__2873_, data_stage_3__2872_, data_stage_3__2871_, data_stage_3__2870_, data_stage_3__2869_, data_stage_3__2868_, data_stage_3__2867_, data_stage_3__2866_, data_stage_3__2865_, data_stage_3__2864_, data_stage_3__2863_, data_stage_3__2862_, data_stage_3__2861_, data_stage_3__2860_, data_stage_3__2859_, data_stage_3__2858_, data_stage_3__2857_, data_stage_3__2856_, data_stage_3__2855_, data_stage_3__2854_, data_stage_3__2853_, data_stage_3__2852_, data_stage_3__2851_, data_stage_3__2850_, data_stage_3__2849_, data_stage_3__2848_, data_stage_3__2847_, data_stage_3__2846_, data_stage_3__2845_, data_stage_3__2844_, data_stage_3__2843_, data_stage_3__2842_, data_stage_3__2841_, data_stage_3__2840_, data_stage_3__2839_, data_stage_3__2838_, data_stage_3__2837_, data_stage_3__2836_, data_stage_3__2835_, data_stage_3__2834_, data_stage_3__2833_, data_stage_3__2832_, data_stage_3__2831_, data_stage_3__2830_, data_stage_3__2829_, data_stage_3__2828_, data_stage_3__2827_, data_stage_3__2826_, data_stage_3__2825_, data_stage_3__2824_, data_stage_3__2823_, data_stage_3__2822_, data_stage_3__2821_, data_stage_3__2820_, data_stage_3__2819_, data_stage_3__2818_, data_stage_3__2817_, data_stage_3__2816_, data_stage_3__2815_, data_stage_3__2814_, data_stage_3__2813_, data_stage_3__2812_, data_stage_3__2811_, data_stage_3__2810_, data_stage_3__2809_, data_stage_3__2808_, data_stage_3__2807_, data_stage_3__2806_, data_stage_3__2805_, data_stage_3__2804_, data_stage_3__2803_, data_stage_3__2802_, data_stage_3__2801_, data_stage_3__2800_, data_stage_3__2799_, data_stage_3__2798_, data_stage_3__2797_, data_stage_3__2796_, data_stage_3__2795_, data_stage_3__2794_, data_stage_3__2793_, data_stage_3__2792_, data_stage_3__2791_, data_stage_3__2790_, data_stage_3__2789_, data_stage_3__2788_, data_stage_3__2787_, data_stage_3__2786_, data_stage_3__2785_, data_stage_3__2784_, data_stage_3__2783_, data_stage_3__2782_, data_stage_3__2781_, data_stage_3__2780_, data_stage_3__2779_, data_stage_3__2778_, data_stage_3__2777_, data_stage_3__2776_, data_stage_3__2775_, data_stage_3__2774_, data_stage_3__2773_, data_stage_3__2772_, data_stage_3__2771_, data_stage_3__2770_, data_stage_3__2769_, data_stage_3__2768_, data_stage_3__2767_, data_stage_3__2766_, data_stage_3__2765_, data_stage_3__2764_, data_stage_3__2763_, data_stage_3__2762_, data_stage_3__2761_, data_stage_3__2760_, data_stage_3__2759_, data_stage_3__2758_, data_stage_3__2757_, data_stage_3__2756_, data_stage_3__2755_, data_stage_3__2754_, data_stage_3__2753_, data_stage_3__2752_, data_stage_3__2751_, data_stage_3__2750_, data_stage_3__2749_, data_stage_3__2748_, data_stage_3__2747_, data_stage_3__2746_, data_stage_3__2745_, data_stage_3__2744_, data_stage_3__2743_, data_stage_3__2742_, data_stage_3__2741_, data_stage_3__2740_, data_stage_3__2739_, data_stage_3__2738_, data_stage_3__2737_, data_stage_3__2736_, data_stage_3__2735_, data_stage_3__2734_, data_stage_3__2733_, data_stage_3__2732_, data_stage_3__2731_, data_stage_3__2730_, data_stage_3__2729_, data_stage_3__2728_, data_stage_3__2727_, data_stage_3__2726_, data_stage_3__2725_, data_stage_3__2724_, data_stage_3__2723_, data_stage_3__2722_, data_stage_3__2721_, data_stage_3__2720_, data_stage_3__2719_, data_stage_3__2718_, data_stage_3__2717_, data_stage_3__2716_, data_stage_3__2715_, data_stage_3__2714_, data_stage_3__2713_, data_stage_3__2712_, data_stage_3__2711_, data_stage_3__2710_, data_stage_3__2709_, data_stage_3__2708_, data_stage_3__2707_, data_stage_3__2706_, data_stage_3__2705_, data_stage_3__2704_, data_stage_3__2703_, data_stage_3__2702_, data_stage_3__2701_, data_stage_3__2700_, data_stage_3__2699_, data_stage_3__2698_, data_stage_3__2697_, data_stage_3__2696_, data_stage_3__2695_, data_stage_3__2694_, data_stage_3__2693_, data_stage_3__2692_, data_stage_3__2691_, data_stage_3__2690_, data_stage_3__2689_, data_stage_3__2688_, data_stage_3__2687_, data_stage_3__2686_, data_stage_3__2685_, data_stage_3__2684_, data_stage_3__2683_, data_stage_3__2682_, data_stage_3__2681_, data_stage_3__2680_, data_stage_3__2679_, data_stage_3__2678_, data_stage_3__2677_, data_stage_3__2676_, data_stage_3__2675_, data_stage_3__2674_, data_stage_3__2673_, data_stage_3__2672_, data_stage_3__2671_, data_stage_3__2670_, data_stage_3__2669_, data_stage_3__2668_, data_stage_3__2667_, data_stage_3__2666_, data_stage_3__2665_, data_stage_3__2664_, data_stage_3__2663_, data_stage_3__2662_, data_stage_3__2661_, data_stage_3__2660_, data_stage_3__2659_, data_stage_3__2658_, data_stage_3__2657_, data_stage_3__2656_, data_stage_3__2655_, data_stage_3__2654_, data_stage_3__2653_, data_stage_3__2652_, data_stage_3__2651_, data_stage_3__2650_, data_stage_3__2649_, data_stage_3__2648_, data_stage_3__2647_, data_stage_3__2646_, data_stage_3__2645_, data_stage_3__2644_, data_stage_3__2643_, data_stage_3__2642_, data_stage_3__2641_, data_stage_3__2640_, data_stage_3__2639_, data_stage_3__2638_, data_stage_3__2637_, data_stage_3__2636_, data_stage_3__2635_, data_stage_3__2634_, data_stage_3__2633_, data_stage_3__2632_, data_stage_3__2631_, data_stage_3__2630_, data_stage_3__2629_, data_stage_3__2628_, data_stage_3__2627_, data_stage_3__2626_, data_stage_3__2625_, data_stage_3__2624_, data_stage_3__2623_, data_stage_3__2622_, data_stage_3__2621_, data_stage_3__2620_, data_stage_3__2619_, data_stage_3__2618_, data_stage_3__2617_, data_stage_3__2616_, data_stage_3__2615_, data_stage_3__2614_, data_stage_3__2613_, data_stage_3__2612_, data_stage_3__2611_, data_stage_3__2610_, data_stage_3__2609_, data_stage_3__2608_, data_stage_3__2607_, data_stage_3__2606_, data_stage_3__2605_, data_stage_3__2604_, data_stage_3__2603_, data_stage_3__2602_, data_stage_3__2601_, data_stage_3__2600_, data_stage_3__2599_, data_stage_3__2598_, data_stage_3__2597_, data_stage_3__2596_, data_stage_3__2595_, data_stage_3__2594_, data_stage_3__2593_, data_stage_3__2592_, data_stage_3__2591_, data_stage_3__2590_, data_stage_3__2589_, data_stage_3__2588_, data_stage_3__2587_, data_stage_3__2586_, data_stage_3__2585_, data_stage_3__2584_, data_stage_3__2583_, data_stage_3__2582_, data_stage_3__2581_, data_stage_3__2580_, data_stage_3__2579_, data_stage_3__2578_, data_stage_3__2577_, data_stage_3__2576_, data_stage_3__2575_, data_stage_3__2574_, data_stage_3__2573_, data_stage_3__2572_, data_stage_3__2571_, data_stage_3__2570_, data_stage_3__2569_, data_stage_3__2568_, data_stage_3__2567_, data_stage_3__2566_, data_stage_3__2565_, data_stage_3__2564_, data_stage_3__2563_, data_stage_3__2562_, data_stage_3__2561_, data_stage_3__2560_, data_stage_3__2559_, data_stage_3__2558_, data_stage_3__2557_, data_stage_3__2556_, data_stage_3__2555_, data_stage_3__2554_, data_stage_3__2553_, data_stage_3__2552_, data_stage_3__2551_, data_stage_3__2550_, data_stage_3__2549_, data_stage_3__2548_, data_stage_3__2547_, data_stage_3__2546_, data_stage_3__2545_, data_stage_3__2544_, data_stage_3__2543_, data_stage_3__2542_, data_stage_3__2541_, data_stage_3__2540_, data_stage_3__2539_, data_stage_3__2538_, data_stage_3__2537_, data_stage_3__2536_, data_stage_3__2535_, data_stage_3__2534_, data_stage_3__2533_, data_stage_3__2532_, data_stage_3__2531_, data_stage_3__2530_, data_stage_3__2529_, data_stage_3__2528_, data_stage_3__2527_, data_stage_3__2526_, data_stage_3__2525_, data_stage_3__2524_, data_stage_3__2523_, data_stage_3__2522_, data_stage_3__2521_, data_stage_3__2520_, data_stage_3__2519_, data_stage_3__2518_, data_stage_3__2517_, data_stage_3__2516_, data_stage_3__2515_, data_stage_3__2514_, data_stage_3__2513_, data_stage_3__2512_, data_stage_3__2511_, data_stage_3__2510_, data_stage_3__2509_, data_stage_3__2508_, data_stage_3__2507_, data_stage_3__2506_, data_stage_3__2505_, data_stage_3__2504_, data_stage_3__2503_, data_stage_3__2502_, data_stage_3__2501_, data_stage_3__2500_, data_stage_3__2499_, data_stage_3__2498_, data_stage_3__2497_, data_stage_3__2496_, data_stage_3__2495_, data_stage_3__2494_, data_stage_3__2493_, data_stage_3__2492_, data_stage_3__2491_, data_stage_3__2490_, data_stage_3__2489_, data_stage_3__2488_, data_stage_3__2487_, data_stage_3__2486_, data_stage_3__2485_, data_stage_3__2484_, data_stage_3__2483_, data_stage_3__2482_, data_stage_3__2481_, data_stage_3__2480_, data_stage_3__2479_, data_stage_3__2478_, data_stage_3__2477_, data_stage_3__2476_, data_stage_3__2475_, data_stage_3__2474_, data_stage_3__2473_, data_stage_3__2472_, data_stage_3__2471_, data_stage_3__2470_, data_stage_3__2469_, data_stage_3__2468_, data_stage_3__2467_, data_stage_3__2466_, data_stage_3__2465_, data_stage_3__2464_, data_stage_3__2463_, data_stage_3__2462_, data_stage_3__2461_, data_stage_3__2460_, data_stage_3__2459_, data_stage_3__2458_, data_stage_3__2457_, data_stage_3__2456_, data_stage_3__2455_, data_stage_3__2454_, data_stage_3__2453_, data_stage_3__2452_, data_stage_3__2451_, data_stage_3__2450_, data_stage_3__2449_, data_stage_3__2448_, data_stage_3__2447_, data_stage_3__2446_, data_stage_3__2445_, data_stage_3__2444_, data_stage_3__2443_, data_stage_3__2442_, data_stage_3__2441_, data_stage_3__2440_, data_stage_3__2439_, data_stage_3__2438_, data_stage_3__2437_, data_stage_3__2436_, data_stage_3__2435_, data_stage_3__2434_, data_stage_3__2433_, data_stage_3__2432_, data_stage_3__2431_, data_stage_3__2430_, data_stage_3__2429_, data_stage_3__2428_, data_stage_3__2427_, data_stage_3__2426_, data_stage_3__2425_, data_stage_3__2424_, data_stage_3__2423_, data_stage_3__2422_, data_stage_3__2421_, data_stage_3__2420_, data_stage_3__2419_, data_stage_3__2418_, data_stage_3__2417_, data_stage_3__2416_, data_stage_3__2415_, data_stage_3__2414_, data_stage_3__2413_, data_stage_3__2412_, data_stage_3__2411_, data_stage_3__2410_, data_stage_3__2409_, data_stage_3__2408_, data_stage_3__2407_, data_stage_3__2406_, data_stage_3__2405_, data_stage_3__2404_, data_stage_3__2403_, data_stage_3__2402_, data_stage_3__2401_, data_stage_3__2400_, data_stage_3__2399_, data_stage_3__2398_, data_stage_3__2397_, data_stage_3__2396_, data_stage_3__2395_, data_stage_3__2394_, data_stage_3__2393_, data_stage_3__2392_, data_stage_3__2391_, data_stage_3__2390_, data_stage_3__2389_, data_stage_3__2388_, data_stage_3__2387_, data_stage_3__2386_, data_stage_3__2385_, data_stage_3__2384_, data_stage_3__2383_, data_stage_3__2382_, data_stage_3__2381_, data_stage_3__2380_, data_stage_3__2379_, data_stage_3__2378_, data_stage_3__2377_, data_stage_3__2376_, data_stage_3__2375_, data_stage_3__2374_, data_stage_3__2373_, data_stage_3__2372_, data_stage_3__2371_, data_stage_3__2370_, data_stage_3__2369_, data_stage_3__2368_, data_stage_3__2367_, data_stage_3__2366_, data_stage_3__2365_, data_stage_3__2364_, data_stage_3__2363_, data_stage_3__2362_, data_stage_3__2361_, data_stage_3__2360_, data_stage_3__2359_, data_stage_3__2358_, data_stage_3__2357_, data_stage_3__2356_, data_stage_3__2355_, data_stage_3__2354_, data_stage_3__2353_, data_stage_3__2352_, data_stage_3__2351_, data_stage_3__2350_, data_stage_3__2349_, data_stage_3__2348_, data_stage_3__2347_, data_stage_3__2346_, data_stage_3__2345_, data_stage_3__2344_, data_stage_3__2343_, data_stage_3__2342_, data_stage_3__2341_, data_stage_3__2340_, data_stage_3__2339_, data_stage_3__2338_, data_stage_3__2337_, data_stage_3__2336_, data_stage_3__2335_, data_stage_3__2334_, data_stage_3__2333_, data_stage_3__2332_, data_stage_3__2331_, data_stage_3__2330_, data_stage_3__2329_, data_stage_3__2328_, data_stage_3__2327_, data_stage_3__2326_, data_stage_3__2325_, data_stage_3__2324_, data_stage_3__2323_, data_stage_3__2322_, data_stage_3__2321_, data_stage_3__2320_, data_stage_3__2319_, data_stage_3__2318_, data_stage_3__2317_, data_stage_3__2316_, data_stage_3__2315_, data_stage_3__2314_, data_stage_3__2313_, data_stage_3__2312_, data_stage_3__2311_, data_stage_3__2310_, data_stage_3__2309_, data_stage_3__2308_, data_stage_3__2307_, data_stage_3__2306_, data_stage_3__2305_, data_stage_3__2304_, data_stage_3__2303_, data_stage_3__2302_, data_stage_3__2301_, data_stage_3__2300_, data_stage_3__2299_, data_stage_3__2298_, data_stage_3__2297_, data_stage_3__2296_, data_stage_3__2295_, data_stage_3__2294_, data_stage_3__2293_, data_stage_3__2292_, data_stage_3__2291_, data_stage_3__2290_, data_stage_3__2289_, data_stage_3__2288_, data_stage_3__2287_, data_stage_3__2286_, data_stage_3__2285_, data_stage_3__2284_, data_stage_3__2283_, data_stage_3__2282_, data_stage_3__2281_, data_stage_3__2280_, data_stage_3__2279_, data_stage_3__2278_, data_stage_3__2277_, data_stage_3__2276_, data_stage_3__2275_, data_stage_3__2274_, data_stage_3__2273_, data_stage_3__2272_, data_stage_3__2271_, data_stage_3__2270_, data_stage_3__2269_, data_stage_3__2268_, data_stage_3__2267_, data_stage_3__2266_, data_stage_3__2265_, data_stage_3__2264_, data_stage_3__2263_, data_stage_3__2262_, data_stage_3__2261_, data_stage_3__2260_, data_stage_3__2259_, data_stage_3__2258_, data_stage_3__2257_, data_stage_3__2256_, data_stage_3__2255_, data_stage_3__2254_, data_stage_3__2253_, data_stage_3__2252_, data_stage_3__2251_, data_stage_3__2250_, data_stage_3__2249_, data_stage_3__2248_, data_stage_3__2247_, data_stage_3__2246_, data_stage_3__2245_, data_stage_3__2244_, data_stage_3__2243_, data_stage_3__2242_, data_stage_3__2241_, data_stage_3__2240_, data_stage_3__2239_, data_stage_3__2238_, data_stage_3__2237_, data_stage_3__2236_, data_stage_3__2235_, data_stage_3__2234_, data_stage_3__2233_, data_stage_3__2232_, data_stage_3__2231_, data_stage_3__2230_, data_stage_3__2229_, data_stage_3__2228_, data_stage_3__2227_, data_stage_3__2226_, data_stage_3__2225_, data_stage_3__2224_, data_stage_3__2223_, data_stage_3__2222_, data_stage_3__2221_, data_stage_3__2220_, data_stage_3__2219_, data_stage_3__2218_, data_stage_3__2217_, data_stage_3__2216_, data_stage_3__2215_, data_stage_3__2214_, data_stage_3__2213_, data_stage_3__2212_, data_stage_3__2211_, data_stage_3__2210_, data_stage_3__2209_, data_stage_3__2208_, data_stage_3__2207_, data_stage_3__2206_, data_stage_3__2205_, data_stage_3__2204_, data_stage_3__2203_, data_stage_3__2202_, data_stage_3__2201_, data_stage_3__2200_, data_stage_3__2199_, data_stage_3__2198_, data_stage_3__2197_, data_stage_3__2196_, data_stage_3__2195_, data_stage_3__2194_, data_stage_3__2193_, data_stage_3__2192_, data_stage_3__2191_, data_stage_3__2190_, data_stage_3__2189_, data_stage_3__2188_, data_stage_3__2187_, data_stage_3__2186_, data_stage_3__2185_, data_stage_3__2184_, data_stage_3__2183_, data_stage_3__2182_, data_stage_3__2181_, data_stage_3__2180_, data_stage_3__2179_, data_stage_3__2178_, data_stage_3__2177_, data_stage_3__2176_, data_stage_3__2175_, data_stage_3__2174_, data_stage_3__2173_, data_stage_3__2172_, data_stage_3__2171_, data_stage_3__2170_, data_stage_3__2169_, data_stage_3__2168_, data_stage_3__2167_, data_stage_3__2166_, data_stage_3__2165_, data_stage_3__2164_, data_stage_3__2163_, data_stage_3__2162_, data_stage_3__2161_, data_stage_3__2160_, data_stage_3__2159_, data_stage_3__2158_, data_stage_3__2157_, data_stage_3__2156_, data_stage_3__2155_, data_stage_3__2154_, data_stage_3__2153_, data_stage_3__2152_, data_stage_3__2151_, data_stage_3__2150_, data_stage_3__2149_, data_stage_3__2148_, data_stage_3__2147_, data_stage_3__2146_, data_stage_3__2145_, data_stage_3__2144_, data_stage_3__2143_, data_stage_3__2142_, data_stage_3__2141_, data_stage_3__2140_, data_stage_3__2139_, data_stage_3__2138_, data_stage_3__2137_, data_stage_3__2136_, data_stage_3__2135_, data_stage_3__2134_, data_stage_3__2133_, data_stage_3__2132_, data_stage_3__2131_, data_stage_3__2130_, data_stage_3__2129_, data_stage_3__2128_, data_stage_3__2127_, data_stage_3__2126_, data_stage_3__2125_, data_stage_3__2124_, data_stage_3__2123_, data_stage_3__2122_, data_stage_3__2121_, data_stage_3__2120_, data_stage_3__2119_, data_stage_3__2118_, data_stage_3__2117_, data_stage_3__2116_, data_stage_3__2115_, data_stage_3__2114_, data_stage_3__2113_, data_stage_3__2112_, data_stage_3__2111_, data_stage_3__2110_, data_stage_3__2109_, data_stage_3__2108_, data_stage_3__2107_, data_stage_3__2106_, data_stage_3__2105_, data_stage_3__2104_, data_stage_3__2103_, data_stage_3__2102_, data_stage_3__2101_, data_stage_3__2100_, data_stage_3__2099_, data_stage_3__2098_, data_stage_3__2097_, data_stage_3__2096_, data_stage_3__2095_, data_stage_3__2094_, data_stage_3__2093_, data_stage_3__2092_, data_stage_3__2091_, data_stage_3__2090_, data_stage_3__2089_, data_stage_3__2088_, data_stage_3__2087_, data_stage_3__2086_, data_stage_3__2085_, data_stage_3__2084_, data_stage_3__2083_, data_stage_3__2082_, data_stage_3__2081_, data_stage_3__2080_, data_stage_3__2079_, data_stage_3__2078_, data_stage_3__2077_, data_stage_3__2076_, data_stage_3__2075_, data_stage_3__2074_, data_stage_3__2073_, data_stage_3__2072_, data_stage_3__2071_, data_stage_3__2070_, data_stage_3__2069_, data_stage_3__2068_, data_stage_3__2067_, data_stage_3__2066_, data_stage_3__2065_, data_stage_3__2064_, data_stage_3__2063_, data_stage_3__2062_, data_stage_3__2061_, data_stage_3__2060_, data_stage_3__2059_, data_stage_3__2058_, data_stage_3__2057_, data_stage_3__2056_, data_stage_3__2055_, data_stage_3__2054_, data_stage_3__2053_, data_stage_3__2052_, data_stage_3__2051_, data_stage_3__2050_, data_stage_3__2049_, data_stage_3__2048_ }),
    .swap_i(sel_i[3]),
    .data_o({ data_stage_4__3071_, data_stage_4__3070_, data_stage_4__3069_, data_stage_4__3068_, data_stage_4__3067_, data_stage_4__3066_, data_stage_4__3065_, data_stage_4__3064_, data_stage_4__3063_, data_stage_4__3062_, data_stage_4__3061_, data_stage_4__3060_, data_stage_4__3059_, data_stage_4__3058_, data_stage_4__3057_, data_stage_4__3056_, data_stage_4__3055_, data_stage_4__3054_, data_stage_4__3053_, data_stage_4__3052_, data_stage_4__3051_, data_stage_4__3050_, data_stage_4__3049_, data_stage_4__3048_, data_stage_4__3047_, data_stage_4__3046_, data_stage_4__3045_, data_stage_4__3044_, data_stage_4__3043_, data_stage_4__3042_, data_stage_4__3041_, data_stage_4__3040_, data_stage_4__3039_, data_stage_4__3038_, data_stage_4__3037_, data_stage_4__3036_, data_stage_4__3035_, data_stage_4__3034_, data_stage_4__3033_, data_stage_4__3032_, data_stage_4__3031_, data_stage_4__3030_, data_stage_4__3029_, data_stage_4__3028_, data_stage_4__3027_, data_stage_4__3026_, data_stage_4__3025_, data_stage_4__3024_, data_stage_4__3023_, data_stage_4__3022_, data_stage_4__3021_, data_stage_4__3020_, data_stage_4__3019_, data_stage_4__3018_, data_stage_4__3017_, data_stage_4__3016_, data_stage_4__3015_, data_stage_4__3014_, data_stage_4__3013_, data_stage_4__3012_, data_stage_4__3011_, data_stage_4__3010_, data_stage_4__3009_, data_stage_4__3008_, data_stage_4__3007_, data_stage_4__3006_, data_stage_4__3005_, data_stage_4__3004_, data_stage_4__3003_, data_stage_4__3002_, data_stage_4__3001_, data_stage_4__3000_, data_stage_4__2999_, data_stage_4__2998_, data_stage_4__2997_, data_stage_4__2996_, data_stage_4__2995_, data_stage_4__2994_, data_stage_4__2993_, data_stage_4__2992_, data_stage_4__2991_, data_stage_4__2990_, data_stage_4__2989_, data_stage_4__2988_, data_stage_4__2987_, data_stage_4__2986_, data_stage_4__2985_, data_stage_4__2984_, data_stage_4__2983_, data_stage_4__2982_, data_stage_4__2981_, data_stage_4__2980_, data_stage_4__2979_, data_stage_4__2978_, data_stage_4__2977_, data_stage_4__2976_, data_stage_4__2975_, data_stage_4__2974_, data_stage_4__2973_, data_stage_4__2972_, data_stage_4__2971_, data_stage_4__2970_, data_stage_4__2969_, data_stage_4__2968_, data_stage_4__2967_, data_stage_4__2966_, data_stage_4__2965_, data_stage_4__2964_, data_stage_4__2963_, data_stage_4__2962_, data_stage_4__2961_, data_stage_4__2960_, data_stage_4__2959_, data_stage_4__2958_, data_stage_4__2957_, data_stage_4__2956_, data_stage_4__2955_, data_stage_4__2954_, data_stage_4__2953_, data_stage_4__2952_, data_stage_4__2951_, data_stage_4__2950_, data_stage_4__2949_, data_stage_4__2948_, data_stage_4__2947_, data_stage_4__2946_, data_stage_4__2945_, data_stage_4__2944_, data_stage_4__2943_, data_stage_4__2942_, data_stage_4__2941_, data_stage_4__2940_, data_stage_4__2939_, data_stage_4__2938_, data_stage_4__2937_, data_stage_4__2936_, data_stage_4__2935_, data_stage_4__2934_, data_stage_4__2933_, data_stage_4__2932_, data_stage_4__2931_, data_stage_4__2930_, data_stage_4__2929_, data_stage_4__2928_, data_stage_4__2927_, data_stage_4__2926_, data_stage_4__2925_, data_stage_4__2924_, data_stage_4__2923_, data_stage_4__2922_, data_stage_4__2921_, data_stage_4__2920_, data_stage_4__2919_, data_stage_4__2918_, data_stage_4__2917_, data_stage_4__2916_, data_stage_4__2915_, data_stage_4__2914_, data_stage_4__2913_, data_stage_4__2912_, data_stage_4__2911_, data_stage_4__2910_, data_stage_4__2909_, data_stage_4__2908_, data_stage_4__2907_, data_stage_4__2906_, data_stage_4__2905_, data_stage_4__2904_, data_stage_4__2903_, data_stage_4__2902_, data_stage_4__2901_, data_stage_4__2900_, data_stage_4__2899_, data_stage_4__2898_, data_stage_4__2897_, data_stage_4__2896_, data_stage_4__2895_, data_stage_4__2894_, data_stage_4__2893_, data_stage_4__2892_, data_stage_4__2891_, data_stage_4__2890_, data_stage_4__2889_, data_stage_4__2888_, data_stage_4__2887_, data_stage_4__2886_, data_stage_4__2885_, data_stage_4__2884_, data_stage_4__2883_, data_stage_4__2882_, data_stage_4__2881_, data_stage_4__2880_, data_stage_4__2879_, data_stage_4__2878_, data_stage_4__2877_, data_stage_4__2876_, data_stage_4__2875_, data_stage_4__2874_, data_stage_4__2873_, data_stage_4__2872_, data_stage_4__2871_, data_stage_4__2870_, data_stage_4__2869_, data_stage_4__2868_, data_stage_4__2867_, data_stage_4__2866_, data_stage_4__2865_, data_stage_4__2864_, data_stage_4__2863_, data_stage_4__2862_, data_stage_4__2861_, data_stage_4__2860_, data_stage_4__2859_, data_stage_4__2858_, data_stage_4__2857_, data_stage_4__2856_, data_stage_4__2855_, data_stage_4__2854_, data_stage_4__2853_, data_stage_4__2852_, data_stage_4__2851_, data_stage_4__2850_, data_stage_4__2849_, data_stage_4__2848_, data_stage_4__2847_, data_stage_4__2846_, data_stage_4__2845_, data_stage_4__2844_, data_stage_4__2843_, data_stage_4__2842_, data_stage_4__2841_, data_stage_4__2840_, data_stage_4__2839_, data_stage_4__2838_, data_stage_4__2837_, data_stage_4__2836_, data_stage_4__2835_, data_stage_4__2834_, data_stage_4__2833_, data_stage_4__2832_, data_stage_4__2831_, data_stage_4__2830_, data_stage_4__2829_, data_stage_4__2828_, data_stage_4__2827_, data_stage_4__2826_, data_stage_4__2825_, data_stage_4__2824_, data_stage_4__2823_, data_stage_4__2822_, data_stage_4__2821_, data_stage_4__2820_, data_stage_4__2819_, data_stage_4__2818_, data_stage_4__2817_, data_stage_4__2816_, data_stage_4__2815_, data_stage_4__2814_, data_stage_4__2813_, data_stage_4__2812_, data_stage_4__2811_, data_stage_4__2810_, data_stage_4__2809_, data_stage_4__2808_, data_stage_4__2807_, data_stage_4__2806_, data_stage_4__2805_, data_stage_4__2804_, data_stage_4__2803_, data_stage_4__2802_, data_stage_4__2801_, data_stage_4__2800_, data_stage_4__2799_, data_stage_4__2798_, data_stage_4__2797_, data_stage_4__2796_, data_stage_4__2795_, data_stage_4__2794_, data_stage_4__2793_, data_stage_4__2792_, data_stage_4__2791_, data_stage_4__2790_, data_stage_4__2789_, data_stage_4__2788_, data_stage_4__2787_, data_stage_4__2786_, data_stage_4__2785_, data_stage_4__2784_, data_stage_4__2783_, data_stage_4__2782_, data_stage_4__2781_, data_stage_4__2780_, data_stage_4__2779_, data_stage_4__2778_, data_stage_4__2777_, data_stage_4__2776_, data_stage_4__2775_, data_stage_4__2774_, data_stage_4__2773_, data_stage_4__2772_, data_stage_4__2771_, data_stage_4__2770_, data_stage_4__2769_, data_stage_4__2768_, data_stage_4__2767_, data_stage_4__2766_, data_stage_4__2765_, data_stage_4__2764_, data_stage_4__2763_, data_stage_4__2762_, data_stage_4__2761_, data_stage_4__2760_, data_stage_4__2759_, data_stage_4__2758_, data_stage_4__2757_, data_stage_4__2756_, data_stage_4__2755_, data_stage_4__2754_, data_stage_4__2753_, data_stage_4__2752_, data_stage_4__2751_, data_stage_4__2750_, data_stage_4__2749_, data_stage_4__2748_, data_stage_4__2747_, data_stage_4__2746_, data_stage_4__2745_, data_stage_4__2744_, data_stage_4__2743_, data_stage_4__2742_, data_stage_4__2741_, data_stage_4__2740_, data_stage_4__2739_, data_stage_4__2738_, data_stage_4__2737_, data_stage_4__2736_, data_stage_4__2735_, data_stage_4__2734_, data_stage_4__2733_, data_stage_4__2732_, data_stage_4__2731_, data_stage_4__2730_, data_stage_4__2729_, data_stage_4__2728_, data_stage_4__2727_, data_stage_4__2726_, data_stage_4__2725_, data_stage_4__2724_, data_stage_4__2723_, data_stage_4__2722_, data_stage_4__2721_, data_stage_4__2720_, data_stage_4__2719_, data_stage_4__2718_, data_stage_4__2717_, data_stage_4__2716_, data_stage_4__2715_, data_stage_4__2714_, data_stage_4__2713_, data_stage_4__2712_, data_stage_4__2711_, data_stage_4__2710_, data_stage_4__2709_, data_stage_4__2708_, data_stage_4__2707_, data_stage_4__2706_, data_stage_4__2705_, data_stage_4__2704_, data_stage_4__2703_, data_stage_4__2702_, data_stage_4__2701_, data_stage_4__2700_, data_stage_4__2699_, data_stage_4__2698_, data_stage_4__2697_, data_stage_4__2696_, data_stage_4__2695_, data_stage_4__2694_, data_stage_4__2693_, data_stage_4__2692_, data_stage_4__2691_, data_stage_4__2690_, data_stage_4__2689_, data_stage_4__2688_, data_stage_4__2687_, data_stage_4__2686_, data_stage_4__2685_, data_stage_4__2684_, data_stage_4__2683_, data_stage_4__2682_, data_stage_4__2681_, data_stage_4__2680_, data_stage_4__2679_, data_stage_4__2678_, data_stage_4__2677_, data_stage_4__2676_, data_stage_4__2675_, data_stage_4__2674_, data_stage_4__2673_, data_stage_4__2672_, data_stage_4__2671_, data_stage_4__2670_, data_stage_4__2669_, data_stage_4__2668_, data_stage_4__2667_, data_stage_4__2666_, data_stage_4__2665_, data_stage_4__2664_, data_stage_4__2663_, data_stage_4__2662_, data_stage_4__2661_, data_stage_4__2660_, data_stage_4__2659_, data_stage_4__2658_, data_stage_4__2657_, data_stage_4__2656_, data_stage_4__2655_, data_stage_4__2654_, data_stage_4__2653_, data_stage_4__2652_, data_stage_4__2651_, data_stage_4__2650_, data_stage_4__2649_, data_stage_4__2648_, data_stage_4__2647_, data_stage_4__2646_, data_stage_4__2645_, data_stage_4__2644_, data_stage_4__2643_, data_stage_4__2642_, data_stage_4__2641_, data_stage_4__2640_, data_stage_4__2639_, data_stage_4__2638_, data_stage_4__2637_, data_stage_4__2636_, data_stage_4__2635_, data_stage_4__2634_, data_stage_4__2633_, data_stage_4__2632_, data_stage_4__2631_, data_stage_4__2630_, data_stage_4__2629_, data_stage_4__2628_, data_stage_4__2627_, data_stage_4__2626_, data_stage_4__2625_, data_stage_4__2624_, data_stage_4__2623_, data_stage_4__2622_, data_stage_4__2621_, data_stage_4__2620_, data_stage_4__2619_, data_stage_4__2618_, data_stage_4__2617_, data_stage_4__2616_, data_stage_4__2615_, data_stage_4__2614_, data_stage_4__2613_, data_stage_4__2612_, data_stage_4__2611_, data_stage_4__2610_, data_stage_4__2609_, data_stage_4__2608_, data_stage_4__2607_, data_stage_4__2606_, data_stage_4__2605_, data_stage_4__2604_, data_stage_4__2603_, data_stage_4__2602_, data_stage_4__2601_, data_stage_4__2600_, data_stage_4__2599_, data_stage_4__2598_, data_stage_4__2597_, data_stage_4__2596_, data_stage_4__2595_, data_stage_4__2594_, data_stage_4__2593_, data_stage_4__2592_, data_stage_4__2591_, data_stage_4__2590_, data_stage_4__2589_, data_stage_4__2588_, data_stage_4__2587_, data_stage_4__2586_, data_stage_4__2585_, data_stage_4__2584_, data_stage_4__2583_, data_stage_4__2582_, data_stage_4__2581_, data_stage_4__2580_, data_stage_4__2579_, data_stage_4__2578_, data_stage_4__2577_, data_stage_4__2576_, data_stage_4__2575_, data_stage_4__2574_, data_stage_4__2573_, data_stage_4__2572_, data_stage_4__2571_, data_stage_4__2570_, data_stage_4__2569_, data_stage_4__2568_, data_stage_4__2567_, data_stage_4__2566_, data_stage_4__2565_, data_stage_4__2564_, data_stage_4__2563_, data_stage_4__2562_, data_stage_4__2561_, data_stage_4__2560_, data_stage_4__2559_, data_stage_4__2558_, data_stage_4__2557_, data_stage_4__2556_, data_stage_4__2555_, data_stage_4__2554_, data_stage_4__2553_, data_stage_4__2552_, data_stage_4__2551_, data_stage_4__2550_, data_stage_4__2549_, data_stage_4__2548_, data_stage_4__2547_, data_stage_4__2546_, data_stage_4__2545_, data_stage_4__2544_, data_stage_4__2543_, data_stage_4__2542_, data_stage_4__2541_, data_stage_4__2540_, data_stage_4__2539_, data_stage_4__2538_, data_stage_4__2537_, data_stage_4__2536_, data_stage_4__2535_, data_stage_4__2534_, data_stage_4__2533_, data_stage_4__2532_, data_stage_4__2531_, data_stage_4__2530_, data_stage_4__2529_, data_stage_4__2528_, data_stage_4__2527_, data_stage_4__2526_, data_stage_4__2525_, data_stage_4__2524_, data_stage_4__2523_, data_stage_4__2522_, data_stage_4__2521_, data_stage_4__2520_, data_stage_4__2519_, data_stage_4__2518_, data_stage_4__2517_, data_stage_4__2516_, data_stage_4__2515_, data_stage_4__2514_, data_stage_4__2513_, data_stage_4__2512_, data_stage_4__2511_, data_stage_4__2510_, data_stage_4__2509_, data_stage_4__2508_, data_stage_4__2507_, data_stage_4__2506_, data_stage_4__2505_, data_stage_4__2504_, data_stage_4__2503_, data_stage_4__2502_, data_stage_4__2501_, data_stage_4__2500_, data_stage_4__2499_, data_stage_4__2498_, data_stage_4__2497_, data_stage_4__2496_, data_stage_4__2495_, data_stage_4__2494_, data_stage_4__2493_, data_stage_4__2492_, data_stage_4__2491_, data_stage_4__2490_, data_stage_4__2489_, data_stage_4__2488_, data_stage_4__2487_, data_stage_4__2486_, data_stage_4__2485_, data_stage_4__2484_, data_stage_4__2483_, data_stage_4__2482_, data_stage_4__2481_, data_stage_4__2480_, data_stage_4__2479_, data_stage_4__2478_, data_stage_4__2477_, data_stage_4__2476_, data_stage_4__2475_, data_stage_4__2474_, data_stage_4__2473_, data_stage_4__2472_, data_stage_4__2471_, data_stage_4__2470_, data_stage_4__2469_, data_stage_4__2468_, data_stage_4__2467_, data_stage_4__2466_, data_stage_4__2465_, data_stage_4__2464_, data_stage_4__2463_, data_stage_4__2462_, data_stage_4__2461_, data_stage_4__2460_, data_stage_4__2459_, data_stage_4__2458_, data_stage_4__2457_, data_stage_4__2456_, data_stage_4__2455_, data_stage_4__2454_, data_stage_4__2453_, data_stage_4__2452_, data_stage_4__2451_, data_stage_4__2450_, data_stage_4__2449_, data_stage_4__2448_, data_stage_4__2447_, data_stage_4__2446_, data_stage_4__2445_, data_stage_4__2444_, data_stage_4__2443_, data_stage_4__2442_, data_stage_4__2441_, data_stage_4__2440_, data_stage_4__2439_, data_stage_4__2438_, data_stage_4__2437_, data_stage_4__2436_, data_stage_4__2435_, data_stage_4__2434_, data_stage_4__2433_, data_stage_4__2432_, data_stage_4__2431_, data_stage_4__2430_, data_stage_4__2429_, data_stage_4__2428_, data_stage_4__2427_, data_stage_4__2426_, data_stage_4__2425_, data_stage_4__2424_, data_stage_4__2423_, data_stage_4__2422_, data_stage_4__2421_, data_stage_4__2420_, data_stage_4__2419_, data_stage_4__2418_, data_stage_4__2417_, data_stage_4__2416_, data_stage_4__2415_, data_stage_4__2414_, data_stage_4__2413_, data_stage_4__2412_, data_stage_4__2411_, data_stage_4__2410_, data_stage_4__2409_, data_stage_4__2408_, data_stage_4__2407_, data_stage_4__2406_, data_stage_4__2405_, data_stage_4__2404_, data_stage_4__2403_, data_stage_4__2402_, data_stage_4__2401_, data_stage_4__2400_, data_stage_4__2399_, data_stage_4__2398_, data_stage_4__2397_, data_stage_4__2396_, data_stage_4__2395_, data_stage_4__2394_, data_stage_4__2393_, data_stage_4__2392_, data_stage_4__2391_, data_stage_4__2390_, data_stage_4__2389_, data_stage_4__2388_, data_stage_4__2387_, data_stage_4__2386_, data_stage_4__2385_, data_stage_4__2384_, data_stage_4__2383_, data_stage_4__2382_, data_stage_4__2381_, data_stage_4__2380_, data_stage_4__2379_, data_stage_4__2378_, data_stage_4__2377_, data_stage_4__2376_, data_stage_4__2375_, data_stage_4__2374_, data_stage_4__2373_, data_stage_4__2372_, data_stage_4__2371_, data_stage_4__2370_, data_stage_4__2369_, data_stage_4__2368_, data_stage_4__2367_, data_stage_4__2366_, data_stage_4__2365_, data_stage_4__2364_, data_stage_4__2363_, data_stage_4__2362_, data_stage_4__2361_, data_stage_4__2360_, data_stage_4__2359_, data_stage_4__2358_, data_stage_4__2357_, data_stage_4__2356_, data_stage_4__2355_, data_stage_4__2354_, data_stage_4__2353_, data_stage_4__2352_, data_stage_4__2351_, data_stage_4__2350_, data_stage_4__2349_, data_stage_4__2348_, data_stage_4__2347_, data_stage_4__2346_, data_stage_4__2345_, data_stage_4__2344_, data_stage_4__2343_, data_stage_4__2342_, data_stage_4__2341_, data_stage_4__2340_, data_stage_4__2339_, data_stage_4__2338_, data_stage_4__2337_, data_stage_4__2336_, data_stage_4__2335_, data_stage_4__2334_, data_stage_4__2333_, data_stage_4__2332_, data_stage_4__2331_, data_stage_4__2330_, data_stage_4__2329_, data_stage_4__2328_, data_stage_4__2327_, data_stage_4__2326_, data_stage_4__2325_, data_stage_4__2324_, data_stage_4__2323_, data_stage_4__2322_, data_stage_4__2321_, data_stage_4__2320_, data_stage_4__2319_, data_stage_4__2318_, data_stage_4__2317_, data_stage_4__2316_, data_stage_4__2315_, data_stage_4__2314_, data_stage_4__2313_, data_stage_4__2312_, data_stage_4__2311_, data_stage_4__2310_, data_stage_4__2309_, data_stage_4__2308_, data_stage_4__2307_, data_stage_4__2306_, data_stage_4__2305_, data_stage_4__2304_, data_stage_4__2303_, data_stage_4__2302_, data_stage_4__2301_, data_stage_4__2300_, data_stage_4__2299_, data_stage_4__2298_, data_stage_4__2297_, data_stage_4__2296_, data_stage_4__2295_, data_stage_4__2294_, data_stage_4__2293_, data_stage_4__2292_, data_stage_4__2291_, data_stage_4__2290_, data_stage_4__2289_, data_stage_4__2288_, data_stage_4__2287_, data_stage_4__2286_, data_stage_4__2285_, data_stage_4__2284_, data_stage_4__2283_, data_stage_4__2282_, data_stage_4__2281_, data_stage_4__2280_, data_stage_4__2279_, data_stage_4__2278_, data_stage_4__2277_, data_stage_4__2276_, data_stage_4__2275_, data_stage_4__2274_, data_stage_4__2273_, data_stage_4__2272_, data_stage_4__2271_, data_stage_4__2270_, data_stage_4__2269_, data_stage_4__2268_, data_stage_4__2267_, data_stage_4__2266_, data_stage_4__2265_, data_stage_4__2264_, data_stage_4__2263_, data_stage_4__2262_, data_stage_4__2261_, data_stage_4__2260_, data_stage_4__2259_, data_stage_4__2258_, data_stage_4__2257_, data_stage_4__2256_, data_stage_4__2255_, data_stage_4__2254_, data_stage_4__2253_, data_stage_4__2252_, data_stage_4__2251_, data_stage_4__2250_, data_stage_4__2249_, data_stage_4__2248_, data_stage_4__2247_, data_stage_4__2246_, data_stage_4__2245_, data_stage_4__2244_, data_stage_4__2243_, data_stage_4__2242_, data_stage_4__2241_, data_stage_4__2240_, data_stage_4__2239_, data_stage_4__2238_, data_stage_4__2237_, data_stage_4__2236_, data_stage_4__2235_, data_stage_4__2234_, data_stage_4__2233_, data_stage_4__2232_, data_stage_4__2231_, data_stage_4__2230_, data_stage_4__2229_, data_stage_4__2228_, data_stage_4__2227_, data_stage_4__2226_, data_stage_4__2225_, data_stage_4__2224_, data_stage_4__2223_, data_stage_4__2222_, data_stage_4__2221_, data_stage_4__2220_, data_stage_4__2219_, data_stage_4__2218_, data_stage_4__2217_, data_stage_4__2216_, data_stage_4__2215_, data_stage_4__2214_, data_stage_4__2213_, data_stage_4__2212_, data_stage_4__2211_, data_stage_4__2210_, data_stage_4__2209_, data_stage_4__2208_, data_stage_4__2207_, data_stage_4__2206_, data_stage_4__2205_, data_stage_4__2204_, data_stage_4__2203_, data_stage_4__2202_, data_stage_4__2201_, data_stage_4__2200_, data_stage_4__2199_, data_stage_4__2198_, data_stage_4__2197_, data_stage_4__2196_, data_stage_4__2195_, data_stage_4__2194_, data_stage_4__2193_, data_stage_4__2192_, data_stage_4__2191_, data_stage_4__2190_, data_stage_4__2189_, data_stage_4__2188_, data_stage_4__2187_, data_stage_4__2186_, data_stage_4__2185_, data_stage_4__2184_, data_stage_4__2183_, data_stage_4__2182_, data_stage_4__2181_, data_stage_4__2180_, data_stage_4__2179_, data_stage_4__2178_, data_stage_4__2177_, data_stage_4__2176_, data_stage_4__2175_, data_stage_4__2174_, data_stage_4__2173_, data_stage_4__2172_, data_stage_4__2171_, data_stage_4__2170_, data_stage_4__2169_, data_stage_4__2168_, data_stage_4__2167_, data_stage_4__2166_, data_stage_4__2165_, data_stage_4__2164_, data_stage_4__2163_, data_stage_4__2162_, data_stage_4__2161_, data_stage_4__2160_, data_stage_4__2159_, data_stage_4__2158_, data_stage_4__2157_, data_stage_4__2156_, data_stage_4__2155_, data_stage_4__2154_, data_stage_4__2153_, data_stage_4__2152_, data_stage_4__2151_, data_stage_4__2150_, data_stage_4__2149_, data_stage_4__2148_, data_stage_4__2147_, data_stage_4__2146_, data_stage_4__2145_, data_stage_4__2144_, data_stage_4__2143_, data_stage_4__2142_, data_stage_4__2141_, data_stage_4__2140_, data_stage_4__2139_, data_stage_4__2138_, data_stage_4__2137_, data_stage_4__2136_, data_stage_4__2135_, data_stage_4__2134_, data_stage_4__2133_, data_stage_4__2132_, data_stage_4__2131_, data_stage_4__2130_, data_stage_4__2129_, data_stage_4__2128_, data_stage_4__2127_, data_stage_4__2126_, data_stage_4__2125_, data_stage_4__2124_, data_stage_4__2123_, data_stage_4__2122_, data_stage_4__2121_, data_stage_4__2120_, data_stage_4__2119_, data_stage_4__2118_, data_stage_4__2117_, data_stage_4__2116_, data_stage_4__2115_, data_stage_4__2114_, data_stage_4__2113_, data_stage_4__2112_, data_stage_4__2111_, data_stage_4__2110_, data_stage_4__2109_, data_stage_4__2108_, data_stage_4__2107_, data_stage_4__2106_, data_stage_4__2105_, data_stage_4__2104_, data_stage_4__2103_, data_stage_4__2102_, data_stage_4__2101_, data_stage_4__2100_, data_stage_4__2099_, data_stage_4__2098_, data_stage_4__2097_, data_stage_4__2096_, data_stage_4__2095_, data_stage_4__2094_, data_stage_4__2093_, data_stage_4__2092_, data_stage_4__2091_, data_stage_4__2090_, data_stage_4__2089_, data_stage_4__2088_, data_stage_4__2087_, data_stage_4__2086_, data_stage_4__2085_, data_stage_4__2084_, data_stage_4__2083_, data_stage_4__2082_, data_stage_4__2081_, data_stage_4__2080_, data_stage_4__2079_, data_stage_4__2078_, data_stage_4__2077_, data_stage_4__2076_, data_stage_4__2075_, data_stage_4__2074_, data_stage_4__2073_, data_stage_4__2072_, data_stage_4__2071_, data_stage_4__2070_, data_stage_4__2069_, data_stage_4__2068_, data_stage_4__2067_, data_stage_4__2066_, data_stage_4__2065_, data_stage_4__2064_, data_stage_4__2063_, data_stage_4__2062_, data_stage_4__2061_, data_stage_4__2060_, data_stage_4__2059_, data_stage_4__2058_, data_stage_4__2057_, data_stage_4__2056_, data_stage_4__2055_, data_stage_4__2054_, data_stage_4__2053_, data_stage_4__2052_, data_stage_4__2051_, data_stage_4__2050_, data_stage_4__2049_, data_stage_4__2048_ })
  );


  bsg_swap_width_p512
  mux_stage_3__mux_swap_3__swap_inst
  (
    .data_i({ data_stage_3__4095_, data_stage_3__4094_, data_stage_3__4093_, data_stage_3__4092_, data_stage_3__4091_, data_stage_3__4090_, data_stage_3__4089_, data_stage_3__4088_, data_stage_3__4087_, data_stage_3__4086_, data_stage_3__4085_, data_stage_3__4084_, data_stage_3__4083_, data_stage_3__4082_, data_stage_3__4081_, data_stage_3__4080_, data_stage_3__4079_, data_stage_3__4078_, data_stage_3__4077_, data_stage_3__4076_, data_stage_3__4075_, data_stage_3__4074_, data_stage_3__4073_, data_stage_3__4072_, data_stage_3__4071_, data_stage_3__4070_, data_stage_3__4069_, data_stage_3__4068_, data_stage_3__4067_, data_stage_3__4066_, data_stage_3__4065_, data_stage_3__4064_, data_stage_3__4063_, data_stage_3__4062_, data_stage_3__4061_, data_stage_3__4060_, data_stage_3__4059_, data_stage_3__4058_, data_stage_3__4057_, data_stage_3__4056_, data_stage_3__4055_, data_stage_3__4054_, data_stage_3__4053_, data_stage_3__4052_, data_stage_3__4051_, data_stage_3__4050_, data_stage_3__4049_, data_stage_3__4048_, data_stage_3__4047_, data_stage_3__4046_, data_stage_3__4045_, data_stage_3__4044_, data_stage_3__4043_, data_stage_3__4042_, data_stage_3__4041_, data_stage_3__4040_, data_stage_3__4039_, data_stage_3__4038_, data_stage_3__4037_, data_stage_3__4036_, data_stage_3__4035_, data_stage_3__4034_, data_stage_3__4033_, data_stage_3__4032_, data_stage_3__4031_, data_stage_3__4030_, data_stage_3__4029_, data_stage_3__4028_, data_stage_3__4027_, data_stage_3__4026_, data_stage_3__4025_, data_stage_3__4024_, data_stage_3__4023_, data_stage_3__4022_, data_stage_3__4021_, data_stage_3__4020_, data_stage_3__4019_, data_stage_3__4018_, data_stage_3__4017_, data_stage_3__4016_, data_stage_3__4015_, data_stage_3__4014_, data_stage_3__4013_, data_stage_3__4012_, data_stage_3__4011_, data_stage_3__4010_, data_stage_3__4009_, data_stage_3__4008_, data_stage_3__4007_, data_stage_3__4006_, data_stage_3__4005_, data_stage_3__4004_, data_stage_3__4003_, data_stage_3__4002_, data_stage_3__4001_, data_stage_3__4000_, data_stage_3__3999_, data_stage_3__3998_, data_stage_3__3997_, data_stage_3__3996_, data_stage_3__3995_, data_stage_3__3994_, data_stage_3__3993_, data_stage_3__3992_, data_stage_3__3991_, data_stage_3__3990_, data_stage_3__3989_, data_stage_3__3988_, data_stage_3__3987_, data_stage_3__3986_, data_stage_3__3985_, data_stage_3__3984_, data_stage_3__3983_, data_stage_3__3982_, data_stage_3__3981_, data_stage_3__3980_, data_stage_3__3979_, data_stage_3__3978_, data_stage_3__3977_, data_stage_3__3976_, data_stage_3__3975_, data_stage_3__3974_, data_stage_3__3973_, data_stage_3__3972_, data_stage_3__3971_, data_stage_3__3970_, data_stage_3__3969_, data_stage_3__3968_, data_stage_3__3967_, data_stage_3__3966_, data_stage_3__3965_, data_stage_3__3964_, data_stage_3__3963_, data_stage_3__3962_, data_stage_3__3961_, data_stage_3__3960_, data_stage_3__3959_, data_stage_3__3958_, data_stage_3__3957_, data_stage_3__3956_, data_stage_3__3955_, data_stage_3__3954_, data_stage_3__3953_, data_stage_3__3952_, data_stage_3__3951_, data_stage_3__3950_, data_stage_3__3949_, data_stage_3__3948_, data_stage_3__3947_, data_stage_3__3946_, data_stage_3__3945_, data_stage_3__3944_, data_stage_3__3943_, data_stage_3__3942_, data_stage_3__3941_, data_stage_3__3940_, data_stage_3__3939_, data_stage_3__3938_, data_stage_3__3937_, data_stage_3__3936_, data_stage_3__3935_, data_stage_3__3934_, data_stage_3__3933_, data_stage_3__3932_, data_stage_3__3931_, data_stage_3__3930_, data_stage_3__3929_, data_stage_3__3928_, data_stage_3__3927_, data_stage_3__3926_, data_stage_3__3925_, data_stage_3__3924_, data_stage_3__3923_, data_stage_3__3922_, data_stage_3__3921_, data_stage_3__3920_, data_stage_3__3919_, data_stage_3__3918_, data_stage_3__3917_, data_stage_3__3916_, data_stage_3__3915_, data_stage_3__3914_, data_stage_3__3913_, data_stage_3__3912_, data_stage_3__3911_, data_stage_3__3910_, data_stage_3__3909_, data_stage_3__3908_, data_stage_3__3907_, data_stage_3__3906_, data_stage_3__3905_, data_stage_3__3904_, data_stage_3__3903_, data_stage_3__3902_, data_stage_3__3901_, data_stage_3__3900_, data_stage_3__3899_, data_stage_3__3898_, data_stage_3__3897_, data_stage_3__3896_, data_stage_3__3895_, data_stage_3__3894_, data_stage_3__3893_, data_stage_3__3892_, data_stage_3__3891_, data_stage_3__3890_, data_stage_3__3889_, data_stage_3__3888_, data_stage_3__3887_, data_stage_3__3886_, data_stage_3__3885_, data_stage_3__3884_, data_stage_3__3883_, data_stage_3__3882_, data_stage_3__3881_, data_stage_3__3880_, data_stage_3__3879_, data_stage_3__3878_, data_stage_3__3877_, data_stage_3__3876_, data_stage_3__3875_, data_stage_3__3874_, data_stage_3__3873_, data_stage_3__3872_, data_stage_3__3871_, data_stage_3__3870_, data_stage_3__3869_, data_stage_3__3868_, data_stage_3__3867_, data_stage_3__3866_, data_stage_3__3865_, data_stage_3__3864_, data_stage_3__3863_, data_stage_3__3862_, data_stage_3__3861_, data_stage_3__3860_, data_stage_3__3859_, data_stage_3__3858_, data_stage_3__3857_, data_stage_3__3856_, data_stage_3__3855_, data_stage_3__3854_, data_stage_3__3853_, data_stage_3__3852_, data_stage_3__3851_, data_stage_3__3850_, data_stage_3__3849_, data_stage_3__3848_, data_stage_3__3847_, data_stage_3__3846_, data_stage_3__3845_, data_stage_3__3844_, data_stage_3__3843_, data_stage_3__3842_, data_stage_3__3841_, data_stage_3__3840_, data_stage_3__3839_, data_stage_3__3838_, data_stage_3__3837_, data_stage_3__3836_, data_stage_3__3835_, data_stage_3__3834_, data_stage_3__3833_, data_stage_3__3832_, data_stage_3__3831_, data_stage_3__3830_, data_stage_3__3829_, data_stage_3__3828_, data_stage_3__3827_, data_stage_3__3826_, data_stage_3__3825_, data_stage_3__3824_, data_stage_3__3823_, data_stage_3__3822_, data_stage_3__3821_, data_stage_3__3820_, data_stage_3__3819_, data_stage_3__3818_, data_stage_3__3817_, data_stage_3__3816_, data_stage_3__3815_, data_stage_3__3814_, data_stage_3__3813_, data_stage_3__3812_, data_stage_3__3811_, data_stage_3__3810_, data_stage_3__3809_, data_stage_3__3808_, data_stage_3__3807_, data_stage_3__3806_, data_stage_3__3805_, data_stage_3__3804_, data_stage_3__3803_, data_stage_3__3802_, data_stage_3__3801_, data_stage_3__3800_, data_stage_3__3799_, data_stage_3__3798_, data_stage_3__3797_, data_stage_3__3796_, data_stage_3__3795_, data_stage_3__3794_, data_stage_3__3793_, data_stage_3__3792_, data_stage_3__3791_, data_stage_3__3790_, data_stage_3__3789_, data_stage_3__3788_, data_stage_3__3787_, data_stage_3__3786_, data_stage_3__3785_, data_stage_3__3784_, data_stage_3__3783_, data_stage_3__3782_, data_stage_3__3781_, data_stage_3__3780_, data_stage_3__3779_, data_stage_3__3778_, data_stage_3__3777_, data_stage_3__3776_, data_stage_3__3775_, data_stage_3__3774_, data_stage_3__3773_, data_stage_3__3772_, data_stage_3__3771_, data_stage_3__3770_, data_stage_3__3769_, data_stage_3__3768_, data_stage_3__3767_, data_stage_3__3766_, data_stage_3__3765_, data_stage_3__3764_, data_stage_3__3763_, data_stage_3__3762_, data_stage_3__3761_, data_stage_3__3760_, data_stage_3__3759_, data_stage_3__3758_, data_stage_3__3757_, data_stage_3__3756_, data_stage_3__3755_, data_stage_3__3754_, data_stage_3__3753_, data_stage_3__3752_, data_stage_3__3751_, data_stage_3__3750_, data_stage_3__3749_, data_stage_3__3748_, data_stage_3__3747_, data_stage_3__3746_, data_stage_3__3745_, data_stage_3__3744_, data_stage_3__3743_, data_stage_3__3742_, data_stage_3__3741_, data_stage_3__3740_, data_stage_3__3739_, data_stage_3__3738_, data_stage_3__3737_, data_stage_3__3736_, data_stage_3__3735_, data_stage_3__3734_, data_stage_3__3733_, data_stage_3__3732_, data_stage_3__3731_, data_stage_3__3730_, data_stage_3__3729_, data_stage_3__3728_, data_stage_3__3727_, data_stage_3__3726_, data_stage_3__3725_, data_stage_3__3724_, data_stage_3__3723_, data_stage_3__3722_, data_stage_3__3721_, data_stage_3__3720_, data_stage_3__3719_, data_stage_3__3718_, data_stage_3__3717_, data_stage_3__3716_, data_stage_3__3715_, data_stage_3__3714_, data_stage_3__3713_, data_stage_3__3712_, data_stage_3__3711_, data_stage_3__3710_, data_stage_3__3709_, data_stage_3__3708_, data_stage_3__3707_, data_stage_3__3706_, data_stage_3__3705_, data_stage_3__3704_, data_stage_3__3703_, data_stage_3__3702_, data_stage_3__3701_, data_stage_3__3700_, data_stage_3__3699_, data_stage_3__3698_, data_stage_3__3697_, data_stage_3__3696_, data_stage_3__3695_, data_stage_3__3694_, data_stage_3__3693_, data_stage_3__3692_, data_stage_3__3691_, data_stage_3__3690_, data_stage_3__3689_, data_stage_3__3688_, data_stage_3__3687_, data_stage_3__3686_, data_stage_3__3685_, data_stage_3__3684_, data_stage_3__3683_, data_stage_3__3682_, data_stage_3__3681_, data_stage_3__3680_, data_stage_3__3679_, data_stage_3__3678_, data_stage_3__3677_, data_stage_3__3676_, data_stage_3__3675_, data_stage_3__3674_, data_stage_3__3673_, data_stage_3__3672_, data_stage_3__3671_, data_stage_3__3670_, data_stage_3__3669_, data_stage_3__3668_, data_stage_3__3667_, data_stage_3__3666_, data_stage_3__3665_, data_stage_3__3664_, data_stage_3__3663_, data_stage_3__3662_, data_stage_3__3661_, data_stage_3__3660_, data_stage_3__3659_, data_stage_3__3658_, data_stage_3__3657_, data_stage_3__3656_, data_stage_3__3655_, data_stage_3__3654_, data_stage_3__3653_, data_stage_3__3652_, data_stage_3__3651_, data_stage_3__3650_, data_stage_3__3649_, data_stage_3__3648_, data_stage_3__3647_, data_stage_3__3646_, data_stage_3__3645_, data_stage_3__3644_, data_stage_3__3643_, data_stage_3__3642_, data_stage_3__3641_, data_stage_3__3640_, data_stage_3__3639_, data_stage_3__3638_, data_stage_3__3637_, data_stage_3__3636_, data_stage_3__3635_, data_stage_3__3634_, data_stage_3__3633_, data_stage_3__3632_, data_stage_3__3631_, data_stage_3__3630_, data_stage_3__3629_, data_stage_3__3628_, data_stage_3__3627_, data_stage_3__3626_, data_stage_3__3625_, data_stage_3__3624_, data_stage_3__3623_, data_stage_3__3622_, data_stage_3__3621_, data_stage_3__3620_, data_stage_3__3619_, data_stage_3__3618_, data_stage_3__3617_, data_stage_3__3616_, data_stage_3__3615_, data_stage_3__3614_, data_stage_3__3613_, data_stage_3__3612_, data_stage_3__3611_, data_stage_3__3610_, data_stage_3__3609_, data_stage_3__3608_, data_stage_3__3607_, data_stage_3__3606_, data_stage_3__3605_, data_stage_3__3604_, data_stage_3__3603_, data_stage_3__3602_, data_stage_3__3601_, data_stage_3__3600_, data_stage_3__3599_, data_stage_3__3598_, data_stage_3__3597_, data_stage_3__3596_, data_stage_3__3595_, data_stage_3__3594_, data_stage_3__3593_, data_stage_3__3592_, data_stage_3__3591_, data_stage_3__3590_, data_stage_3__3589_, data_stage_3__3588_, data_stage_3__3587_, data_stage_3__3586_, data_stage_3__3585_, data_stage_3__3584_, data_stage_3__3583_, data_stage_3__3582_, data_stage_3__3581_, data_stage_3__3580_, data_stage_3__3579_, data_stage_3__3578_, data_stage_3__3577_, data_stage_3__3576_, data_stage_3__3575_, data_stage_3__3574_, data_stage_3__3573_, data_stage_3__3572_, data_stage_3__3571_, data_stage_3__3570_, data_stage_3__3569_, data_stage_3__3568_, data_stage_3__3567_, data_stage_3__3566_, data_stage_3__3565_, data_stage_3__3564_, data_stage_3__3563_, data_stage_3__3562_, data_stage_3__3561_, data_stage_3__3560_, data_stage_3__3559_, data_stage_3__3558_, data_stage_3__3557_, data_stage_3__3556_, data_stage_3__3555_, data_stage_3__3554_, data_stage_3__3553_, data_stage_3__3552_, data_stage_3__3551_, data_stage_3__3550_, data_stage_3__3549_, data_stage_3__3548_, data_stage_3__3547_, data_stage_3__3546_, data_stage_3__3545_, data_stage_3__3544_, data_stage_3__3543_, data_stage_3__3542_, data_stage_3__3541_, data_stage_3__3540_, data_stage_3__3539_, data_stage_3__3538_, data_stage_3__3537_, data_stage_3__3536_, data_stage_3__3535_, data_stage_3__3534_, data_stage_3__3533_, data_stage_3__3532_, data_stage_3__3531_, data_stage_3__3530_, data_stage_3__3529_, data_stage_3__3528_, data_stage_3__3527_, data_stage_3__3526_, data_stage_3__3525_, data_stage_3__3524_, data_stage_3__3523_, data_stage_3__3522_, data_stage_3__3521_, data_stage_3__3520_, data_stage_3__3519_, data_stage_3__3518_, data_stage_3__3517_, data_stage_3__3516_, data_stage_3__3515_, data_stage_3__3514_, data_stage_3__3513_, data_stage_3__3512_, data_stage_3__3511_, data_stage_3__3510_, data_stage_3__3509_, data_stage_3__3508_, data_stage_3__3507_, data_stage_3__3506_, data_stage_3__3505_, data_stage_3__3504_, data_stage_3__3503_, data_stage_3__3502_, data_stage_3__3501_, data_stage_3__3500_, data_stage_3__3499_, data_stage_3__3498_, data_stage_3__3497_, data_stage_3__3496_, data_stage_3__3495_, data_stage_3__3494_, data_stage_3__3493_, data_stage_3__3492_, data_stage_3__3491_, data_stage_3__3490_, data_stage_3__3489_, data_stage_3__3488_, data_stage_3__3487_, data_stage_3__3486_, data_stage_3__3485_, data_stage_3__3484_, data_stage_3__3483_, data_stage_3__3482_, data_stage_3__3481_, data_stage_3__3480_, data_stage_3__3479_, data_stage_3__3478_, data_stage_3__3477_, data_stage_3__3476_, data_stage_3__3475_, data_stage_3__3474_, data_stage_3__3473_, data_stage_3__3472_, data_stage_3__3471_, data_stage_3__3470_, data_stage_3__3469_, data_stage_3__3468_, data_stage_3__3467_, data_stage_3__3466_, data_stage_3__3465_, data_stage_3__3464_, data_stage_3__3463_, data_stage_3__3462_, data_stage_3__3461_, data_stage_3__3460_, data_stage_3__3459_, data_stage_3__3458_, data_stage_3__3457_, data_stage_3__3456_, data_stage_3__3455_, data_stage_3__3454_, data_stage_3__3453_, data_stage_3__3452_, data_stage_3__3451_, data_stage_3__3450_, data_stage_3__3449_, data_stage_3__3448_, data_stage_3__3447_, data_stage_3__3446_, data_stage_3__3445_, data_stage_3__3444_, data_stage_3__3443_, data_stage_3__3442_, data_stage_3__3441_, data_stage_3__3440_, data_stage_3__3439_, data_stage_3__3438_, data_stage_3__3437_, data_stage_3__3436_, data_stage_3__3435_, data_stage_3__3434_, data_stage_3__3433_, data_stage_3__3432_, data_stage_3__3431_, data_stage_3__3430_, data_stage_3__3429_, data_stage_3__3428_, data_stage_3__3427_, data_stage_3__3426_, data_stage_3__3425_, data_stage_3__3424_, data_stage_3__3423_, data_stage_3__3422_, data_stage_3__3421_, data_stage_3__3420_, data_stage_3__3419_, data_stage_3__3418_, data_stage_3__3417_, data_stage_3__3416_, data_stage_3__3415_, data_stage_3__3414_, data_stage_3__3413_, data_stage_3__3412_, data_stage_3__3411_, data_stage_3__3410_, data_stage_3__3409_, data_stage_3__3408_, data_stage_3__3407_, data_stage_3__3406_, data_stage_3__3405_, data_stage_3__3404_, data_stage_3__3403_, data_stage_3__3402_, data_stage_3__3401_, data_stage_3__3400_, data_stage_3__3399_, data_stage_3__3398_, data_stage_3__3397_, data_stage_3__3396_, data_stage_3__3395_, data_stage_3__3394_, data_stage_3__3393_, data_stage_3__3392_, data_stage_3__3391_, data_stage_3__3390_, data_stage_3__3389_, data_stage_3__3388_, data_stage_3__3387_, data_stage_3__3386_, data_stage_3__3385_, data_stage_3__3384_, data_stage_3__3383_, data_stage_3__3382_, data_stage_3__3381_, data_stage_3__3380_, data_stage_3__3379_, data_stage_3__3378_, data_stage_3__3377_, data_stage_3__3376_, data_stage_3__3375_, data_stage_3__3374_, data_stage_3__3373_, data_stage_3__3372_, data_stage_3__3371_, data_stage_3__3370_, data_stage_3__3369_, data_stage_3__3368_, data_stage_3__3367_, data_stage_3__3366_, data_stage_3__3365_, data_stage_3__3364_, data_stage_3__3363_, data_stage_3__3362_, data_stage_3__3361_, data_stage_3__3360_, data_stage_3__3359_, data_stage_3__3358_, data_stage_3__3357_, data_stage_3__3356_, data_stage_3__3355_, data_stage_3__3354_, data_stage_3__3353_, data_stage_3__3352_, data_stage_3__3351_, data_stage_3__3350_, data_stage_3__3349_, data_stage_3__3348_, data_stage_3__3347_, data_stage_3__3346_, data_stage_3__3345_, data_stage_3__3344_, data_stage_3__3343_, data_stage_3__3342_, data_stage_3__3341_, data_stage_3__3340_, data_stage_3__3339_, data_stage_3__3338_, data_stage_3__3337_, data_stage_3__3336_, data_stage_3__3335_, data_stage_3__3334_, data_stage_3__3333_, data_stage_3__3332_, data_stage_3__3331_, data_stage_3__3330_, data_stage_3__3329_, data_stage_3__3328_, data_stage_3__3327_, data_stage_3__3326_, data_stage_3__3325_, data_stage_3__3324_, data_stage_3__3323_, data_stage_3__3322_, data_stage_3__3321_, data_stage_3__3320_, data_stage_3__3319_, data_stage_3__3318_, data_stage_3__3317_, data_stage_3__3316_, data_stage_3__3315_, data_stage_3__3314_, data_stage_3__3313_, data_stage_3__3312_, data_stage_3__3311_, data_stage_3__3310_, data_stage_3__3309_, data_stage_3__3308_, data_stage_3__3307_, data_stage_3__3306_, data_stage_3__3305_, data_stage_3__3304_, data_stage_3__3303_, data_stage_3__3302_, data_stage_3__3301_, data_stage_3__3300_, data_stage_3__3299_, data_stage_3__3298_, data_stage_3__3297_, data_stage_3__3296_, data_stage_3__3295_, data_stage_3__3294_, data_stage_3__3293_, data_stage_3__3292_, data_stage_3__3291_, data_stage_3__3290_, data_stage_3__3289_, data_stage_3__3288_, data_stage_3__3287_, data_stage_3__3286_, data_stage_3__3285_, data_stage_3__3284_, data_stage_3__3283_, data_stage_3__3282_, data_stage_3__3281_, data_stage_3__3280_, data_stage_3__3279_, data_stage_3__3278_, data_stage_3__3277_, data_stage_3__3276_, data_stage_3__3275_, data_stage_3__3274_, data_stage_3__3273_, data_stage_3__3272_, data_stage_3__3271_, data_stage_3__3270_, data_stage_3__3269_, data_stage_3__3268_, data_stage_3__3267_, data_stage_3__3266_, data_stage_3__3265_, data_stage_3__3264_, data_stage_3__3263_, data_stage_3__3262_, data_stage_3__3261_, data_stage_3__3260_, data_stage_3__3259_, data_stage_3__3258_, data_stage_3__3257_, data_stage_3__3256_, data_stage_3__3255_, data_stage_3__3254_, data_stage_3__3253_, data_stage_3__3252_, data_stage_3__3251_, data_stage_3__3250_, data_stage_3__3249_, data_stage_3__3248_, data_stage_3__3247_, data_stage_3__3246_, data_stage_3__3245_, data_stage_3__3244_, data_stage_3__3243_, data_stage_3__3242_, data_stage_3__3241_, data_stage_3__3240_, data_stage_3__3239_, data_stage_3__3238_, data_stage_3__3237_, data_stage_3__3236_, data_stage_3__3235_, data_stage_3__3234_, data_stage_3__3233_, data_stage_3__3232_, data_stage_3__3231_, data_stage_3__3230_, data_stage_3__3229_, data_stage_3__3228_, data_stage_3__3227_, data_stage_3__3226_, data_stage_3__3225_, data_stage_3__3224_, data_stage_3__3223_, data_stage_3__3222_, data_stage_3__3221_, data_stage_3__3220_, data_stage_3__3219_, data_stage_3__3218_, data_stage_3__3217_, data_stage_3__3216_, data_stage_3__3215_, data_stage_3__3214_, data_stage_3__3213_, data_stage_3__3212_, data_stage_3__3211_, data_stage_3__3210_, data_stage_3__3209_, data_stage_3__3208_, data_stage_3__3207_, data_stage_3__3206_, data_stage_3__3205_, data_stage_3__3204_, data_stage_3__3203_, data_stage_3__3202_, data_stage_3__3201_, data_stage_3__3200_, data_stage_3__3199_, data_stage_3__3198_, data_stage_3__3197_, data_stage_3__3196_, data_stage_3__3195_, data_stage_3__3194_, data_stage_3__3193_, data_stage_3__3192_, data_stage_3__3191_, data_stage_3__3190_, data_stage_3__3189_, data_stage_3__3188_, data_stage_3__3187_, data_stage_3__3186_, data_stage_3__3185_, data_stage_3__3184_, data_stage_3__3183_, data_stage_3__3182_, data_stage_3__3181_, data_stage_3__3180_, data_stage_3__3179_, data_stage_3__3178_, data_stage_3__3177_, data_stage_3__3176_, data_stage_3__3175_, data_stage_3__3174_, data_stage_3__3173_, data_stage_3__3172_, data_stage_3__3171_, data_stage_3__3170_, data_stage_3__3169_, data_stage_3__3168_, data_stage_3__3167_, data_stage_3__3166_, data_stage_3__3165_, data_stage_3__3164_, data_stage_3__3163_, data_stage_3__3162_, data_stage_3__3161_, data_stage_3__3160_, data_stage_3__3159_, data_stage_3__3158_, data_stage_3__3157_, data_stage_3__3156_, data_stage_3__3155_, data_stage_3__3154_, data_stage_3__3153_, data_stage_3__3152_, data_stage_3__3151_, data_stage_3__3150_, data_stage_3__3149_, data_stage_3__3148_, data_stage_3__3147_, data_stage_3__3146_, data_stage_3__3145_, data_stage_3__3144_, data_stage_3__3143_, data_stage_3__3142_, data_stage_3__3141_, data_stage_3__3140_, data_stage_3__3139_, data_stage_3__3138_, data_stage_3__3137_, data_stage_3__3136_, data_stage_3__3135_, data_stage_3__3134_, data_stage_3__3133_, data_stage_3__3132_, data_stage_3__3131_, data_stage_3__3130_, data_stage_3__3129_, data_stage_3__3128_, data_stage_3__3127_, data_stage_3__3126_, data_stage_3__3125_, data_stage_3__3124_, data_stage_3__3123_, data_stage_3__3122_, data_stage_3__3121_, data_stage_3__3120_, data_stage_3__3119_, data_stage_3__3118_, data_stage_3__3117_, data_stage_3__3116_, data_stage_3__3115_, data_stage_3__3114_, data_stage_3__3113_, data_stage_3__3112_, data_stage_3__3111_, data_stage_3__3110_, data_stage_3__3109_, data_stage_3__3108_, data_stage_3__3107_, data_stage_3__3106_, data_stage_3__3105_, data_stage_3__3104_, data_stage_3__3103_, data_stage_3__3102_, data_stage_3__3101_, data_stage_3__3100_, data_stage_3__3099_, data_stage_3__3098_, data_stage_3__3097_, data_stage_3__3096_, data_stage_3__3095_, data_stage_3__3094_, data_stage_3__3093_, data_stage_3__3092_, data_stage_3__3091_, data_stage_3__3090_, data_stage_3__3089_, data_stage_3__3088_, data_stage_3__3087_, data_stage_3__3086_, data_stage_3__3085_, data_stage_3__3084_, data_stage_3__3083_, data_stage_3__3082_, data_stage_3__3081_, data_stage_3__3080_, data_stage_3__3079_, data_stage_3__3078_, data_stage_3__3077_, data_stage_3__3076_, data_stage_3__3075_, data_stage_3__3074_, data_stage_3__3073_, data_stage_3__3072_ }),
    .swap_i(sel_i[3]),
    .data_o({ data_stage_4__4095_, data_stage_4__4094_, data_stage_4__4093_, data_stage_4__4092_, data_stage_4__4091_, data_stage_4__4090_, data_stage_4__4089_, data_stage_4__4088_, data_stage_4__4087_, data_stage_4__4086_, data_stage_4__4085_, data_stage_4__4084_, data_stage_4__4083_, data_stage_4__4082_, data_stage_4__4081_, data_stage_4__4080_, data_stage_4__4079_, data_stage_4__4078_, data_stage_4__4077_, data_stage_4__4076_, data_stage_4__4075_, data_stage_4__4074_, data_stage_4__4073_, data_stage_4__4072_, data_stage_4__4071_, data_stage_4__4070_, data_stage_4__4069_, data_stage_4__4068_, data_stage_4__4067_, data_stage_4__4066_, data_stage_4__4065_, data_stage_4__4064_, data_stage_4__4063_, data_stage_4__4062_, data_stage_4__4061_, data_stage_4__4060_, data_stage_4__4059_, data_stage_4__4058_, data_stage_4__4057_, data_stage_4__4056_, data_stage_4__4055_, data_stage_4__4054_, data_stage_4__4053_, data_stage_4__4052_, data_stage_4__4051_, data_stage_4__4050_, data_stage_4__4049_, data_stage_4__4048_, data_stage_4__4047_, data_stage_4__4046_, data_stage_4__4045_, data_stage_4__4044_, data_stage_4__4043_, data_stage_4__4042_, data_stage_4__4041_, data_stage_4__4040_, data_stage_4__4039_, data_stage_4__4038_, data_stage_4__4037_, data_stage_4__4036_, data_stage_4__4035_, data_stage_4__4034_, data_stage_4__4033_, data_stage_4__4032_, data_stage_4__4031_, data_stage_4__4030_, data_stage_4__4029_, data_stage_4__4028_, data_stage_4__4027_, data_stage_4__4026_, data_stage_4__4025_, data_stage_4__4024_, data_stage_4__4023_, data_stage_4__4022_, data_stage_4__4021_, data_stage_4__4020_, data_stage_4__4019_, data_stage_4__4018_, data_stage_4__4017_, data_stage_4__4016_, data_stage_4__4015_, data_stage_4__4014_, data_stage_4__4013_, data_stage_4__4012_, data_stage_4__4011_, data_stage_4__4010_, data_stage_4__4009_, data_stage_4__4008_, data_stage_4__4007_, data_stage_4__4006_, data_stage_4__4005_, data_stage_4__4004_, data_stage_4__4003_, data_stage_4__4002_, data_stage_4__4001_, data_stage_4__4000_, data_stage_4__3999_, data_stage_4__3998_, data_stage_4__3997_, data_stage_4__3996_, data_stage_4__3995_, data_stage_4__3994_, data_stage_4__3993_, data_stage_4__3992_, data_stage_4__3991_, data_stage_4__3990_, data_stage_4__3989_, data_stage_4__3988_, data_stage_4__3987_, data_stage_4__3986_, data_stage_4__3985_, data_stage_4__3984_, data_stage_4__3983_, data_stage_4__3982_, data_stage_4__3981_, data_stage_4__3980_, data_stage_4__3979_, data_stage_4__3978_, data_stage_4__3977_, data_stage_4__3976_, data_stage_4__3975_, data_stage_4__3974_, data_stage_4__3973_, data_stage_4__3972_, data_stage_4__3971_, data_stage_4__3970_, data_stage_4__3969_, data_stage_4__3968_, data_stage_4__3967_, data_stage_4__3966_, data_stage_4__3965_, data_stage_4__3964_, data_stage_4__3963_, data_stage_4__3962_, data_stage_4__3961_, data_stage_4__3960_, data_stage_4__3959_, data_stage_4__3958_, data_stage_4__3957_, data_stage_4__3956_, data_stage_4__3955_, data_stage_4__3954_, data_stage_4__3953_, data_stage_4__3952_, data_stage_4__3951_, data_stage_4__3950_, data_stage_4__3949_, data_stage_4__3948_, data_stage_4__3947_, data_stage_4__3946_, data_stage_4__3945_, data_stage_4__3944_, data_stage_4__3943_, data_stage_4__3942_, data_stage_4__3941_, data_stage_4__3940_, data_stage_4__3939_, data_stage_4__3938_, data_stage_4__3937_, data_stage_4__3936_, data_stage_4__3935_, data_stage_4__3934_, data_stage_4__3933_, data_stage_4__3932_, data_stage_4__3931_, data_stage_4__3930_, data_stage_4__3929_, data_stage_4__3928_, data_stage_4__3927_, data_stage_4__3926_, data_stage_4__3925_, data_stage_4__3924_, data_stage_4__3923_, data_stage_4__3922_, data_stage_4__3921_, data_stage_4__3920_, data_stage_4__3919_, data_stage_4__3918_, data_stage_4__3917_, data_stage_4__3916_, data_stage_4__3915_, data_stage_4__3914_, data_stage_4__3913_, data_stage_4__3912_, data_stage_4__3911_, data_stage_4__3910_, data_stage_4__3909_, data_stage_4__3908_, data_stage_4__3907_, data_stage_4__3906_, data_stage_4__3905_, data_stage_4__3904_, data_stage_4__3903_, data_stage_4__3902_, data_stage_4__3901_, data_stage_4__3900_, data_stage_4__3899_, data_stage_4__3898_, data_stage_4__3897_, data_stage_4__3896_, data_stage_4__3895_, data_stage_4__3894_, data_stage_4__3893_, data_stage_4__3892_, data_stage_4__3891_, data_stage_4__3890_, data_stage_4__3889_, data_stage_4__3888_, data_stage_4__3887_, data_stage_4__3886_, data_stage_4__3885_, data_stage_4__3884_, data_stage_4__3883_, data_stage_4__3882_, data_stage_4__3881_, data_stage_4__3880_, data_stage_4__3879_, data_stage_4__3878_, data_stage_4__3877_, data_stage_4__3876_, data_stage_4__3875_, data_stage_4__3874_, data_stage_4__3873_, data_stage_4__3872_, data_stage_4__3871_, data_stage_4__3870_, data_stage_4__3869_, data_stage_4__3868_, data_stage_4__3867_, data_stage_4__3866_, data_stage_4__3865_, data_stage_4__3864_, data_stage_4__3863_, data_stage_4__3862_, data_stage_4__3861_, data_stage_4__3860_, data_stage_4__3859_, data_stage_4__3858_, data_stage_4__3857_, data_stage_4__3856_, data_stage_4__3855_, data_stage_4__3854_, data_stage_4__3853_, data_stage_4__3852_, data_stage_4__3851_, data_stage_4__3850_, data_stage_4__3849_, data_stage_4__3848_, data_stage_4__3847_, data_stage_4__3846_, data_stage_4__3845_, data_stage_4__3844_, data_stage_4__3843_, data_stage_4__3842_, data_stage_4__3841_, data_stage_4__3840_, data_stage_4__3839_, data_stage_4__3838_, data_stage_4__3837_, data_stage_4__3836_, data_stage_4__3835_, data_stage_4__3834_, data_stage_4__3833_, data_stage_4__3832_, data_stage_4__3831_, data_stage_4__3830_, data_stage_4__3829_, data_stage_4__3828_, data_stage_4__3827_, data_stage_4__3826_, data_stage_4__3825_, data_stage_4__3824_, data_stage_4__3823_, data_stage_4__3822_, data_stage_4__3821_, data_stage_4__3820_, data_stage_4__3819_, data_stage_4__3818_, data_stage_4__3817_, data_stage_4__3816_, data_stage_4__3815_, data_stage_4__3814_, data_stage_4__3813_, data_stage_4__3812_, data_stage_4__3811_, data_stage_4__3810_, data_stage_4__3809_, data_stage_4__3808_, data_stage_4__3807_, data_stage_4__3806_, data_stage_4__3805_, data_stage_4__3804_, data_stage_4__3803_, data_stage_4__3802_, data_stage_4__3801_, data_stage_4__3800_, data_stage_4__3799_, data_stage_4__3798_, data_stage_4__3797_, data_stage_4__3796_, data_stage_4__3795_, data_stage_4__3794_, data_stage_4__3793_, data_stage_4__3792_, data_stage_4__3791_, data_stage_4__3790_, data_stage_4__3789_, data_stage_4__3788_, data_stage_4__3787_, data_stage_4__3786_, data_stage_4__3785_, data_stage_4__3784_, data_stage_4__3783_, data_stage_4__3782_, data_stage_4__3781_, data_stage_4__3780_, data_stage_4__3779_, data_stage_4__3778_, data_stage_4__3777_, data_stage_4__3776_, data_stage_4__3775_, data_stage_4__3774_, data_stage_4__3773_, data_stage_4__3772_, data_stage_4__3771_, data_stage_4__3770_, data_stage_4__3769_, data_stage_4__3768_, data_stage_4__3767_, data_stage_4__3766_, data_stage_4__3765_, data_stage_4__3764_, data_stage_4__3763_, data_stage_4__3762_, data_stage_4__3761_, data_stage_4__3760_, data_stage_4__3759_, data_stage_4__3758_, data_stage_4__3757_, data_stage_4__3756_, data_stage_4__3755_, data_stage_4__3754_, data_stage_4__3753_, data_stage_4__3752_, data_stage_4__3751_, data_stage_4__3750_, data_stage_4__3749_, data_stage_4__3748_, data_stage_4__3747_, data_stage_4__3746_, data_stage_4__3745_, data_stage_4__3744_, data_stage_4__3743_, data_stage_4__3742_, data_stage_4__3741_, data_stage_4__3740_, data_stage_4__3739_, data_stage_4__3738_, data_stage_4__3737_, data_stage_4__3736_, data_stage_4__3735_, data_stage_4__3734_, data_stage_4__3733_, data_stage_4__3732_, data_stage_4__3731_, data_stage_4__3730_, data_stage_4__3729_, data_stage_4__3728_, data_stage_4__3727_, data_stage_4__3726_, data_stage_4__3725_, data_stage_4__3724_, data_stage_4__3723_, data_stage_4__3722_, data_stage_4__3721_, data_stage_4__3720_, data_stage_4__3719_, data_stage_4__3718_, data_stage_4__3717_, data_stage_4__3716_, data_stage_4__3715_, data_stage_4__3714_, data_stage_4__3713_, data_stage_4__3712_, data_stage_4__3711_, data_stage_4__3710_, data_stage_4__3709_, data_stage_4__3708_, data_stage_4__3707_, data_stage_4__3706_, data_stage_4__3705_, data_stage_4__3704_, data_stage_4__3703_, data_stage_4__3702_, data_stage_4__3701_, data_stage_4__3700_, data_stage_4__3699_, data_stage_4__3698_, data_stage_4__3697_, data_stage_4__3696_, data_stage_4__3695_, data_stage_4__3694_, data_stage_4__3693_, data_stage_4__3692_, data_stage_4__3691_, data_stage_4__3690_, data_stage_4__3689_, data_stage_4__3688_, data_stage_4__3687_, data_stage_4__3686_, data_stage_4__3685_, data_stage_4__3684_, data_stage_4__3683_, data_stage_4__3682_, data_stage_4__3681_, data_stage_4__3680_, data_stage_4__3679_, data_stage_4__3678_, data_stage_4__3677_, data_stage_4__3676_, data_stage_4__3675_, data_stage_4__3674_, data_stage_4__3673_, data_stage_4__3672_, data_stage_4__3671_, data_stage_4__3670_, data_stage_4__3669_, data_stage_4__3668_, data_stage_4__3667_, data_stage_4__3666_, data_stage_4__3665_, data_stage_4__3664_, data_stage_4__3663_, data_stage_4__3662_, data_stage_4__3661_, data_stage_4__3660_, data_stage_4__3659_, data_stage_4__3658_, data_stage_4__3657_, data_stage_4__3656_, data_stage_4__3655_, data_stage_4__3654_, data_stage_4__3653_, data_stage_4__3652_, data_stage_4__3651_, data_stage_4__3650_, data_stage_4__3649_, data_stage_4__3648_, data_stage_4__3647_, data_stage_4__3646_, data_stage_4__3645_, data_stage_4__3644_, data_stage_4__3643_, data_stage_4__3642_, data_stage_4__3641_, data_stage_4__3640_, data_stage_4__3639_, data_stage_4__3638_, data_stage_4__3637_, data_stage_4__3636_, data_stage_4__3635_, data_stage_4__3634_, data_stage_4__3633_, data_stage_4__3632_, data_stage_4__3631_, data_stage_4__3630_, data_stage_4__3629_, data_stage_4__3628_, data_stage_4__3627_, data_stage_4__3626_, data_stage_4__3625_, data_stage_4__3624_, data_stage_4__3623_, data_stage_4__3622_, data_stage_4__3621_, data_stage_4__3620_, data_stage_4__3619_, data_stage_4__3618_, data_stage_4__3617_, data_stage_4__3616_, data_stage_4__3615_, data_stage_4__3614_, data_stage_4__3613_, data_stage_4__3612_, data_stage_4__3611_, data_stage_4__3610_, data_stage_4__3609_, data_stage_4__3608_, data_stage_4__3607_, data_stage_4__3606_, data_stage_4__3605_, data_stage_4__3604_, data_stage_4__3603_, data_stage_4__3602_, data_stage_4__3601_, data_stage_4__3600_, data_stage_4__3599_, data_stage_4__3598_, data_stage_4__3597_, data_stage_4__3596_, data_stage_4__3595_, data_stage_4__3594_, data_stage_4__3593_, data_stage_4__3592_, data_stage_4__3591_, data_stage_4__3590_, data_stage_4__3589_, data_stage_4__3588_, data_stage_4__3587_, data_stage_4__3586_, data_stage_4__3585_, data_stage_4__3584_, data_stage_4__3583_, data_stage_4__3582_, data_stage_4__3581_, data_stage_4__3580_, data_stage_4__3579_, data_stage_4__3578_, data_stage_4__3577_, data_stage_4__3576_, data_stage_4__3575_, data_stage_4__3574_, data_stage_4__3573_, data_stage_4__3572_, data_stage_4__3571_, data_stage_4__3570_, data_stage_4__3569_, data_stage_4__3568_, data_stage_4__3567_, data_stage_4__3566_, data_stage_4__3565_, data_stage_4__3564_, data_stage_4__3563_, data_stage_4__3562_, data_stage_4__3561_, data_stage_4__3560_, data_stage_4__3559_, data_stage_4__3558_, data_stage_4__3557_, data_stage_4__3556_, data_stage_4__3555_, data_stage_4__3554_, data_stage_4__3553_, data_stage_4__3552_, data_stage_4__3551_, data_stage_4__3550_, data_stage_4__3549_, data_stage_4__3548_, data_stage_4__3547_, data_stage_4__3546_, data_stage_4__3545_, data_stage_4__3544_, data_stage_4__3543_, data_stage_4__3542_, data_stage_4__3541_, data_stage_4__3540_, data_stage_4__3539_, data_stage_4__3538_, data_stage_4__3537_, data_stage_4__3536_, data_stage_4__3535_, data_stage_4__3534_, data_stage_4__3533_, data_stage_4__3532_, data_stage_4__3531_, data_stage_4__3530_, data_stage_4__3529_, data_stage_4__3528_, data_stage_4__3527_, data_stage_4__3526_, data_stage_4__3525_, data_stage_4__3524_, data_stage_4__3523_, data_stage_4__3522_, data_stage_4__3521_, data_stage_4__3520_, data_stage_4__3519_, data_stage_4__3518_, data_stage_4__3517_, data_stage_4__3516_, data_stage_4__3515_, data_stage_4__3514_, data_stage_4__3513_, data_stage_4__3512_, data_stage_4__3511_, data_stage_4__3510_, data_stage_4__3509_, data_stage_4__3508_, data_stage_4__3507_, data_stage_4__3506_, data_stage_4__3505_, data_stage_4__3504_, data_stage_4__3503_, data_stage_4__3502_, data_stage_4__3501_, data_stage_4__3500_, data_stage_4__3499_, data_stage_4__3498_, data_stage_4__3497_, data_stage_4__3496_, data_stage_4__3495_, data_stage_4__3494_, data_stage_4__3493_, data_stage_4__3492_, data_stage_4__3491_, data_stage_4__3490_, data_stage_4__3489_, data_stage_4__3488_, data_stage_4__3487_, data_stage_4__3486_, data_stage_4__3485_, data_stage_4__3484_, data_stage_4__3483_, data_stage_4__3482_, data_stage_4__3481_, data_stage_4__3480_, data_stage_4__3479_, data_stage_4__3478_, data_stage_4__3477_, data_stage_4__3476_, data_stage_4__3475_, data_stage_4__3474_, data_stage_4__3473_, data_stage_4__3472_, data_stage_4__3471_, data_stage_4__3470_, data_stage_4__3469_, data_stage_4__3468_, data_stage_4__3467_, data_stage_4__3466_, data_stage_4__3465_, data_stage_4__3464_, data_stage_4__3463_, data_stage_4__3462_, data_stage_4__3461_, data_stage_4__3460_, data_stage_4__3459_, data_stage_4__3458_, data_stage_4__3457_, data_stage_4__3456_, data_stage_4__3455_, data_stage_4__3454_, data_stage_4__3453_, data_stage_4__3452_, data_stage_4__3451_, data_stage_4__3450_, data_stage_4__3449_, data_stage_4__3448_, data_stage_4__3447_, data_stage_4__3446_, data_stage_4__3445_, data_stage_4__3444_, data_stage_4__3443_, data_stage_4__3442_, data_stage_4__3441_, data_stage_4__3440_, data_stage_4__3439_, data_stage_4__3438_, data_stage_4__3437_, data_stage_4__3436_, data_stage_4__3435_, data_stage_4__3434_, data_stage_4__3433_, data_stage_4__3432_, data_stage_4__3431_, data_stage_4__3430_, data_stage_4__3429_, data_stage_4__3428_, data_stage_4__3427_, data_stage_4__3426_, data_stage_4__3425_, data_stage_4__3424_, data_stage_4__3423_, data_stage_4__3422_, data_stage_4__3421_, data_stage_4__3420_, data_stage_4__3419_, data_stage_4__3418_, data_stage_4__3417_, data_stage_4__3416_, data_stage_4__3415_, data_stage_4__3414_, data_stage_4__3413_, data_stage_4__3412_, data_stage_4__3411_, data_stage_4__3410_, data_stage_4__3409_, data_stage_4__3408_, data_stage_4__3407_, data_stage_4__3406_, data_stage_4__3405_, data_stage_4__3404_, data_stage_4__3403_, data_stage_4__3402_, data_stage_4__3401_, data_stage_4__3400_, data_stage_4__3399_, data_stage_4__3398_, data_stage_4__3397_, data_stage_4__3396_, data_stage_4__3395_, data_stage_4__3394_, data_stage_4__3393_, data_stage_4__3392_, data_stage_4__3391_, data_stage_4__3390_, data_stage_4__3389_, data_stage_4__3388_, data_stage_4__3387_, data_stage_4__3386_, data_stage_4__3385_, data_stage_4__3384_, data_stage_4__3383_, data_stage_4__3382_, data_stage_4__3381_, data_stage_4__3380_, data_stage_4__3379_, data_stage_4__3378_, data_stage_4__3377_, data_stage_4__3376_, data_stage_4__3375_, data_stage_4__3374_, data_stage_4__3373_, data_stage_4__3372_, data_stage_4__3371_, data_stage_4__3370_, data_stage_4__3369_, data_stage_4__3368_, data_stage_4__3367_, data_stage_4__3366_, data_stage_4__3365_, data_stage_4__3364_, data_stage_4__3363_, data_stage_4__3362_, data_stage_4__3361_, data_stage_4__3360_, data_stage_4__3359_, data_stage_4__3358_, data_stage_4__3357_, data_stage_4__3356_, data_stage_4__3355_, data_stage_4__3354_, data_stage_4__3353_, data_stage_4__3352_, data_stage_4__3351_, data_stage_4__3350_, data_stage_4__3349_, data_stage_4__3348_, data_stage_4__3347_, data_stage_4__3346_, data_stage_4__3345_, data_stage_4__3344_, data_stage_4__3343_, data_stage_4__3342_, data_stage_4__3341_, data_stage_4__3340_, data_stage_4__3339_, data_stage_4__3338_, data_stage_4__3337_, data_stage_4__3336_, data_stage_4__3335_, data_stage_4__3334_, data_stage_4__3333_, data_stage_4__3332_, data_stage_4__3331_, data_stage_4__3330_, data_stage_4__3329_, data_stage_4__3328_, data_stage_4__3327_, data_stage_4__3326_, data_stage_4__3325_, data_stage_4__3324_, data_stage_4__3323_, data_stage_4__3322_, data_stage_4__3321_, data_stage_4__3320_, data_stage_4__3319_, data_stage_4__3318_, data_stage_4__3317_, data_stage_4__3316_, data_stage_4__3315_, data_stage_4__3314_, data_stage_4__3313_, data_stage_4__3312_, data_stage_4__3311_, data_stage_4__3310_, data_stage_4__3309_, data_stage_4__3308_, data_stage_4__3307_, data_stage_4__3306_, data_stage_4__3305_, data_stage_4__3304_, data_stage_4__3303_, data_stage_4__3302_, data_stage_4__3301_, data_stage_4__3300_, data_stage_4__3299_, data_stage_4__3298_, data_stage_4__3297_, data_stage_4__3296_, data_stage_4__3295_, data_stage_4__3294_, data_stage_4__3293_, data_stage_4__3292_, data_stage_4__3291_, data_stage_4__3290_, data_stage_4__3289_, data_stage_4__3288_, data_stage_4__3287_, data_stage_4__3286_, data_stage_4__3285_, data_stage_4__3284_, data_stage_4__3283_, data_stage_4__3282_, data_stage_4__3281_, data_stage_4__3280_, data_stage_4__3279_, data_stage_4__3278_, data_stage_4__3277_, data_stage_4__3276_, data_stage_4__3275_, data_stage_4__3274_, data_stage_4__3273_, data_stage_4__3272_, data_stage_4__3271_, data_stage_4__3270_, data_stage_4__3269_, data_stage_4__3268_, data_stage_4__3267_, data_stage_4__3266_, data_stage_4__3265_, data_stage_4__3264_, data_stage_4__3263_, data_stage_4__3262_, data_stage_4__3261_, data_stage_4__3260_, data_stage_4__3259_, data_stage_4__3258_, data_stage_4__3257_, data_stage_4__3256_, data_stage_4__3255_, data_stage_4__3254_, data_stage_4__3253_, data_stage_4__3252_, data_stage_4__3251_, data_stage_4__3250_, data_stage_4__3249_, data_stage_4__3248_, data_stage_4__3247_, data_stage_4__3246_, data_stage_4__3245_, data_stage_4__3244_, data_stage_4__3243_, data_stage_4__3242_, data_stage_4__3241_, data_stage_4__3240_, data_stage_4__3239_, data_stage_4__3238_, data_stage_4__3237_, data_stage_4__3236_, data_stage_4__3235_, data_stage_4__3234_, data_stage_4__3233_, data_stage_4__3232_, data_stage_4__3231_, data_stage_4__3230_, data_stage_4__3229_, data_stage_4__3228_, data_stage_4__3227_, data_stage_4__3226_, data_stage_4__3225_, data_stage_4__3224_, data_stage_4__3223_, data_stage_4__3222_, data_stage_4__3221_, data_stage_4__3220_, data_stage_4__3219_, data_stage_4__3218_, data_stage_4__3217_, data_stage_4__3216_, data_stage_4__3215_, data_stage_4__3214_, data_stage_4__3213_, data_stage_4__3212_, data_stage_4__3211_, data_stage_4__3210_, data_stage_4__3209_, data_stage_4__3208_, data_stage_4__3207_, data_stage_4__3206_, data_stage_4__3205_, data_stage_4__3204_, data_stage_4__3203_, data_stage_4__3202_, data_stage_4__3201_, data_stage_4__3200_, data_stage_4__3199_, data_stage_4__3198_, data_stage_4__3197_, data_stage_4__3196_, data_stage_4__3195_, data_stage_4__3194_, data_stage_4__3193_, data_stage_4__3192_, data_stage_4__3191_, data_stage_4__3190_, data_stage_4__3189_, data_stage_4__3188_, data_stage_4__3187_, data_stage_4__3186_, data_stage_4__3185_, data_stage_4__3184_, data_stage_4__3183_, data_stage_4__3182_, data_stage_4__3181_, data_stage_4__3180_, data_stage_4__3179_, data_stage_4__3178_, data_stage_4__3177_, data_stage_4__3176_, data_stage_4__3175_, data_stage_4__3174_, data_stage_4__3173_, data_stage_4__3172_, data_stage_4__3171_, data_stage_4__3170_, data_stage_4__3169_, data_stage_4__3168_, data_stage_4__3167_, data_stage_4__3166_, data_stage_4__3165_, data_stage_4__3164_, data_stage_4__3163_, data_stage_4__3162_, data_stage_4__3161_, data_stage_4__3160_, data_stage_4__3159_, data_stage_4__3158_, data_stage_4__3157_, data_stage_4__3156_, data_stage_4__3155_, data_stage_4__3154_, data_stage_4__3153_, data_stage_4__3152_, data_stage_4__3151_, data_stage_4__3150_, data_stage_4__3149_, data_stage_4__3148_, data_stage_4__3147_, data_stage_4__3146_, data_stage_4__3145_, data_stage_4__3144_, data_stage_4__3143_, data_stage_4__3142_, data_stage_4__3141_, data_stage_4__3140_, data_stage_4__3139_, data_stage_4__3138_, data_stage_4__3137_, data_stage_4__3136_, data_stage_4__3135_, data_stage_4__3134_, data_stage_4__3133_, data_stage_4__3132_, data_stage_4__3131_, data_stage_4__3130_, data_stage_4__3129_, data_stage_4__3128_, data_stage_4__3127_, data_stage_4__3126_, data_stage_4__3125_, data_stage_4__3124_, data_stage_4__3123_, data_stage_4__3122_, data_stage_4__3121_, data_stage_4__3120_, data_stage_4__3119_, data_stage_4__3118_, data_stage_4__3117_, data_stage_4__3116_, data_stage_4__3115_, data_stage_4__3114_, data_stage_4__3113_, data_stage_4__3112_, data_stage_4__3111_, data_stage_4__3110_, data_stage_4__3109_, data_stage_4__3108_, data_stage_4__3107_, data_stage_4__3106_, data_stage_4__3105_, data_stage_4__3104_, data_stage_4__3103_, data_stage_4__3102_, data_stage_4__3101_, data_stage_4__3100_, data_stage_4__3099_, data_stage_4__3098_, data_stage_4__3097_, data_stage_4__3096_, data_stage_4__3095_, data_stage_4__3094_, data_stage_4__3093_, data_stage_4__3092_, data_stage_4__3091_, data_stage_4__3090_, data_stage_4__3089_, data_stage_4__3088_, data_stage_4__3087_, data_stage_4__3086_, data_stage_4__3085_, data_stage_4__3084_, data_stage_4__3083_, data_stage_4__3082_, data_stage_4__3081_, data_stage_4__3080_, data_stage_4__3079_, data_stage_4__3078_, data_stage_4__3077_, data_stage_4__3076_, data_stage_4__3075_, data_stage_4__3074_, data_stage_4__3073_, data_stage_4__3072_ })
  );


  bsg_swap_width_p1024
  mux_stage_4__mux_swap_0__swap_inst
  (
    .data_i({ data_stage_4__2047_, data_stage_4__2046_, data_stage_4__2045_, data_stage_4__2044_, data_stage_4__2043_, data_stage_4__2042_, data_stage_4__2041_, data_stage_4__2040_, data_stage_4__2039_, data_stage_4__2038_, data_stage_4__2037_, data_stage_4__2036_, data_stage_4__2035_, data_stage_4__2034_, data_stage_4__2033_, data_stage_4__2032_, data_stage_4__2031_, data_stage_4__2030_, data_stage_4__2029_, data_stage_4__2028_, data_stage_4__2027_, data_stage_4__2026_, data_stage_4__2025_, data_stage_4__2024_, data_stage_4__2023_, data_stage_4__2022_, data_stage_4__2021_, data_stage_4__2020_, data_stage_4__2019_, data_stage_4__2018_, data_stage_4__2017_, data_stage_4__2016_, data_stage_4__2015_, data_stage_4__2014_, data_stage_4__2013_, data_stage_4__2012_, data_stage_4__2011_, data_stage_4__2010_, data_stage_4__2009_, data_stage_4__2008_, data_stage_4__2007_, data_stage_4__2006_, data_stage_4__2005_, data_stage_4__2004_, data_stage_4__2003_, data_stage_4__2002_, data_stage_4__2001_, data_stage_4__2000_, data_stage_4__1999_, data_stage_4__1998_, data_stage_4__1997_, data_stage_4__1996_, data_stage_4__1995_, data_stage_4__1994_, data_stage_4__1993_, data_stage_4__1992_, data_stage_4__1991_, data_stage_4__1990_, data_stage_4__1989_, data_stage_4__1988_, data_stage_4__1987_, data_stage_4__1986_, data_stage_4__1985_, data_stage_4__1984_, data_stage_4__1983_, data_stage_4__1982_, data_stage_4__1981_, data_stage_4__1980_, data_stage_4__1979_, data_stage_4__1978_, data_stage_4__1977_, data_stage_4__1976_, data_stage_4__1975_, data_stage_4__1974_, data_stage_4__1973_, data_stage_4__1972_, data_stage_4__1971_, data_stage_4__1970_, data_stage_4__1969_, data_stage_4__1968_, data_stage_4__1967_, data_stage_4__1966_, data_stage_4__1965_, data_stage_4__1964_, data_stage_4__1963_, data_stage_4__1962_, data_stage_4__1961_, data_stage_4__1960_, data_stage_4__1959_, data_stage_4__1958_, data_stage_4__1957_, data_stage_4__1956_, data_stage_4__1955_, data_stage_4__1954_, data_stage_4__1953_, data_stage_4__1952_, data_stage_4__1951_, data_stage_4__1950_, data_stage_4__1949_, data_stage_4__1948_, data_stage_4__1947_, data_stage_4__1946_, data_stage_4__1945_, data_stage_4__1944_, data_stage_4__1943_, data_stage_4__1942_, data_stage_4__1941_, data_stage_4__1940_, data_stage_4__1939_, data_stage_4__1938_, data_stage_4__1937_, data_stage_4__1936_, data_stage_4__1935_, data_stage_4__1934_, data_stage_4__1933_, data_stage_4__1932_, data_stage_4__1931_, data_stage_4__1930_, data_stage_4__1929_, data_stage_4__1928_, data_stage_4__1927_, data_stage_4__1926_, data_stage_4__1925_, data_stage_4__1924_, data_stage_4__1923_, data_stage_4__1922_, data_stage_4__1921_, data_stage_4__1920_, data_stage_4__1919_, data_stage_4__1918_, data_stage_4__1917_, data_stage_4__1916_, data_stage_4__1915_, data_stage_4__1914_, data_stage_4__1913_, data_stage_4__1912_, data_stage_4__1911_, data_stage_4__1910_, data_stage_4__1909_, data_stage_4__1908_, data_stage_4__1907_, data_stage_4__1906_, data_stage_4__1905_, data_stage_4__1904_, data_stage_4__1903_, data_stage_4__1902_, data_stage_4__1901_, data_stage_4__1900_, data_stage_4__1899_, data_stage_4__1898_, data_stage_4__1897_, data_stage_4__1896_, data_stage_4__1895_, data_stage_4__1894_, data_stage_4__1893_, data_stage_4__1892_, data_stage_4__1891_, data_stage_4__1890_, data_stage_4__1889_, data_stage_4__1888_, data_stage_4__1887_, data_stage_4__1886_, data_stage_4__1885_, data_stage_4__1884_, data_stage_4__1883_, data_stage_4__1882_, data_stage_4__1881_, data_stage_4__1880_, data_stage_4__1879_, data_stage_4__1878_, data_stage_4__1877_, data_stage_4__1876_, data_stage_4__1875_, data_stage_4__1874_, data_stage_4__1873_, data_stage_4__1872_, data_stage_4__1871_, data_stage_4__1870_, data_stage_4__1869_, data_stage_4__1868_, data_stage_4__1867_, data_stage_4__1866_, data_stage_4__1865_, data_stage_4__1864_, data_stage_4__1863_, data_stage_4__1862_, data_stage_4__1861_, data_stage_4__1860_, data_stage_4__1859_, data_stage_4__1858_, data_stage_4__1857_, data_stage_4__1856_, data_stage_4__1855_, data_stage_4__1854_, data_stage_4__1853_, data_stage_4__1852_, data_stage_4__1851_, data_stage_4__1850_, data_stage_4__1849_, data_stage_4__1848_, data_stage_4__1847_, data_stage_4__1846_, data_stage_4__1845_, data_stage_4__1844_, data_stage_4__1843_, data_stage_4__1842_, data_stage_4__1841_, data_stage_4__1840_, data_stage_4__1839_, data_stage_4__1838_, data_stage_4__1837_, data_stage_4__1836_, data_stage_4__1835_, data_stage_4__1834_, data_stage_4__1833_, data_stage_4__1832_, data_stage_4__1831_, data_stage_4__1830_, data_stage_4__1829_, data_stage_4__1828_, data_stage_4__1827_, data_stage_4__1826_, data_stage_4__1825_, data_stage_4__1824_, data_stage_4__1823_, data_stage_4__1822_, data_stage_4__1821_, data_stage_4__1820_, data_stage_4__1819_, data_stage_4__1818_, data_stage_4__1817_, data_stage_4__1816_, data_stage_4__1815_, data_stage_4__1814_, data_stage_4__1813_, data_stage_4__1812_, data_stage_4__1811_, data_stage_4__1810_, data_stage_4__1809_, data_stage_4__1808_, data_stage_4__1807_, data_stage_4__1806_, data_stage_4__1805_, data_stage_4__1804_, data_stage_4__1803_, data_stage_4__1802_, data_stage_4__1801_, data_stage_4__1800_, data_stage_4__1799_, data_stage_4__1798_, data_stage_4__1797_, data_stage_4__1796_, data_stage_4__1795_, data_stage_4__1794_, data_stage_4__1793_, data_stage_4__1792_, data_stage_4__1791_, data_stage_4__1790_, data_stage_4__1789_, data_stage_4__1788_, data_stage_4__1787_, data_stage_4__1786_, data_stage_4__1785_, data_stage_4__1784_, data_stage_4__1783_, data_stage_4__1782_, data_stage_4__1781_, data_stage_4__1780_, data_stage_4__1779_, data_stage_4__1778_, data_stage_4__1777_, data_stage_4__1776_, data_stage_4__1775_, data_stage_4__1774_, data_stage_4__1773_, data_stage_4__1772_, data_stage_4__1771_, data_stage_4__1770_, data_stage_4__1769_, data_stage_4__1768_, data_stage_4__1767_, data_stage_4__1766_, data_stage_4__1765_, data_stage_4__1764_, data_stage_4__1763_, data_stage_4__1762_, data_stage_4__1761_, data_stage_4__1760_, data_stage_4__1759_, data_stage_4__1758_, data_stage_4__1757_, data_stage_4__1756_, data_stage_4__1755_, data_stage_4__1754_, data_stage_4__1753_, data_stage_4__1752_, data_stage_4__1751_, data_stage_4__1750_, data_stage_4__1749_, data_stage_4__1748_, data_stage_4__1747_, data_stage_4__1746_, data_stage_4__1745_, data_stage_4__1744_, data_stage_4__1743_, data_stage_4__1742_, data_stage_4__1741_, data_stage_4__1740_, data_stage_4__1739_, data_stage_4__1738_, data_stage_4__1737_, data_stage_4__1736_, data_stage_4__1735_, data_stage_4__1734_, data_stage_4__1733_, data_stage_4__1732_, data_stage_4__1731_, data_stage_4__1730_, data_stage_4__1729_, data_stage_4__1728_, data_stage_4__1727_, data_stage_4__1726_, data_stage_4__1725_, data_stage_4__1724_, data_stage_4__1723_, data_stage_4__1722_, data_stage_4__1721_, data_stage_4__1720_, data_stage_4__1719_, data_stage_4__1718_, data_stage_4__1717_, data_stage_4__1716_, data_stage_4__1715_, data_stage_4__1714_, data_stage_4__1713_, data_stage_4__1712_, data_stage_4__1711_, data_stage_4__1710_, data_stage_4__1709_, data_stage_4__1708_, data_stage_4__1707_, data_stage_4__1706_, data_stage_4__1705_, data_stage_4__1704_, data_stage_4__1703_, data_stage_4__1702_, data_stage_4__1701_, data_stage_4__1700_, data_stage_4__1699_, data_stage_4__1698_, data_stage_4__1697_, data_stage_4__1696_, data_stage_4__1695_, data_stage_4__1694_, data_stage_4__1693_, data_stage_4__1692_, data_stage_4__1691_, data_stage_4__1690_, data_stage_4__1689_, data_stage_4__1688_, data_stage_4__1687_, data_stage_4__1686_, data_stage_4__1685_, data_stage_4__1684_, data_stage_4__1683_, data_stage_4__1682_, data_stage_4__1681_, data_stage_4__1680_, data_stage_4__1679_, data_stage_4__1678_, data_stage_4__1677_, data_stage_4__1676_, data_stage_4__1675_, data_stage_4__1674_, data_stage_4__1673_, data_stage_4__1672_, data_stage_4__1671_, data_stage_4__1670_, data_stage_4__1669_, data_stage_4__1668_, data_stage_4__1667_, data_stage_4__1666_, data_stage_4__1665_, data_stage_4__1664_, data_stage_4__1663_, data_stage_4__1662_, data_stage_4__1661_, data_stage_4__1660_, data_stage_4__1659_, data_stage_4__1658_, data_stage_4__1657_, data_stage_4__1656_, data_stage_4__1655_, data_stage_4__1654_, data_stage_4__1653_, data_stage_4__1652_, data_stage_4__1651_, data_stage_4__1650_, data_stage_4__1649_, data_stage_4__1648_, data_stage_4__1647_, data_stage_4__1646_, data_stage_4__1645_, data_stage_4__1644_, data_stage_4__1643_, data_stage_4__1642_, data_stage_4__1641_, data_stage_4__1640_, data_stage_4__1639_, data_stage_4__1638_, data_stage_4__1637_, data_stage_4__1636_, data_stage_4__1635_, data_stage_4__1634_, data_stage_4__1633_, data_stage_4__1632_, data_stage_4__1631_, data_stage_4__1630_, data_stage_4__1629_, data_stage_4__1628_, data_stage_4__1627_, data_stage_4__1626_, data_stage_4__1625_, data_stage_4__1624_, data_stage_4__1623_, data_stage_4__1622_, data_stage_4__1621_, data_stage_4__1620_, data_stage_4__1619_, data_stage_4__1618_, data_stage_4__1617_, data_stage_4__1616_, data_stage_4__1615_, data_stage_4__1614_, data_stage_4__1613_, data_stage_4__1612_, data_stage_4__1611_, data_stage_4__1610_, data_stage_4__1609_, data_stage_4__1608_, data_stage_4__1607_, data_stage_4__1606_, data_stage_4__1605_, data_stage_4__1604_, data_stage_4__1603_, data_stage_4__1602_, data_stage_4__1601_, data_stage_4__1600_, data_stage_4__1599_, data_stage_4__1598_, data_stage_4__1597_, data_stage_4__1596_, data_stage_4__1595_, data_stage_4__1594_, data_stage_4__1593_, data_stage_4__1592_, data_stage_4__1591_, data_stage_4__1590_, data_stage_4__1589_, data_stage_4__1588_, data_stage_4__1587_, data_stage_4__1586_, data_stage_4__1585_, data_stage_4__1584_, data_stage_4__1583_, data_stage_4__1582_, data_stage_4__1581_, data_stage_4__1580_, data_stage_4__1579_, data_stage_4__1578_, data_stage_4__1577_, data_stage_4__1576_, data_stage_4__1575_, data_stage_4__1574_, data_stage_4__1573_, data_stage_4__1572_, data_stage_4__1571_, data_stage_4__1570_, data_stage_4__1569_, data_stage_4__1568_, data_stage_4__1567_, data_stage_4__1566_, data_stage_4__1565_, data_stage_4__1564_, data_stage_4__1563_, data_stage_4__1562_, data_stage_4__1561_, data_stage_4__1560_, data_stage_4__1559_, data_stage_4__1558_, data_stage_4__1557_, data_stage_4__1556_, data_stage_4__1555_, data_stage_4__1554_, data_stage_4__1553_, data_stage_4__1552_, data_stage_4__1551_, data_stage_4__1550_, data_stage_4__1549_, data_stage_4__1548_, data_stage_4__1547_, data_stage_4__1546_, data_stage_4__1545_, data_stage_4__1544_, data_stage_4__1543_, data_stage_4__1542_, data_stage_4__1541_, data_stage_4__1540_, data_stage_4__1539_, data_stage_4__1538_, data_stage_4__1537_, data_stage_4__1536_, data_stage_4__1535_, data_stage_4__1534_, data_stage_4__1533_, data_stage_4__1532_, data_stage_4__1531_, data_stage_4__1530_, data_stage_4__1529_, data_stage_4__1528_, data_stage_4__1527_, data_stage_4__1526_, data_stage_4__1525_, data_stage_4__1524_, data_stage_4__1523_, data_stage_4__1522_, data_stage_4__1521_, data_stage_4__1520_, data_stage_4__1519_, data_stage_4__1518_, data_stage_4__1517_, data_stage_4__1516_, data_stage_4__1515_, data_stage_4__1514_, data_stage_4__1513_, data_stage_4__1512_, data_stage_4__1511_, data_stage_4__1510_, data_stage_4__1509_, data_stage_4__1508_, data_stage_4__1507_, data_stage_4__1506_, data_stage_4__1505_, data_stage_4__1504_, data_stage_4__1503_, data_stage_4__1502_, data_stage_4__1501_, data_stage_4__1500_, data_stage_4__1499_, data_stage_4__1498_, data_stage_4__1497_, data_stage_4__1496_, data_stage_4__1495_, data_stage_4__1494_, data_stage_4__1493_, data_stage_4__1492_, data_stage_4__1491_, data_stage_4__1490_, data_stage_4__1489_, data_stage_4__1488_, data_stage_4__1487_, data_stage_4__1486_, data_stage_4__1485_, data_stage_4__1484_, data_stage_4__1483_, data_stage_4__1482_, data_stage_4__1481_, data_stage_4__1480_, data_stage_4__1479_, data_stage_4__1478_, data_stage_4__1477_, data_stage_4__1476_, data_stage_4__1475_, data_stage_4__1474_, data_stage_4__1473_, data_stage_4__1472_, data_stage_4__1471_, data_stage_4__1470_, data_stage_4__1469_, data_stage_4__1468_, data_stage_4__1467_, data_stage_4__1466_, data_stage_4__1465_, data_stage_4__1464_, data_stage_4__1463_, data_stage_4__1462_, data_stage_4__1461_, data_stage_4__1460_, data_stage_4__1459_, data_stage_4__1458_, data_stage_4__1457_, data_stage_4__1456_, data_stage_4__1455_, data_stage_4__1454_, data_stage_4__1453_, data_stage_4__1452_, data_stage_4__1451_, data_stage_4__1450_, data_stage_4__1449_, data_stage_4__1448_, data_stage_4__1447_, data_stage_4__1446_, data_stage_4__1445_, data_stage_4__1444_, data_stage_4__1443_, data_stage_4__1442_, data_stage_4__1441_, data_stage_4__1440_, data_stage_4__1439_, data_stage_4__1438_, data_stage_4__1437_, data_stage_4__1436_, data_stage_4__1435_, data_stage_4__1434_, data_stage_4__1433_, data_stage_4__1432_, data_stage_4__1431_, data_stage_4__1430_, data_stage_4__1429_, data_stage_4__1428_, data_stage_4__1427_, data_stage_4__1426_, data_stage_4__1425_, data_stage_4__1424_, data_stage_4__1423_, data_stage_4__1422_, data_stage_4__1421_, data_stage_4__1420_, data_stage_4__1419_, data_stage_4__1418_, data_stage_4__1417_, data_stage_4__1416_, data_stage_4__1415_, data_stage_4__1414_, data_stage_4__1413_, data_stage_4__1412_, data_stage_4__1411_, data_stage_4__1410_, data_stage_4__1409_, data_stage_4__1408_, data_stage_4__1407_, data_stage_4__1406_, data_stage_4__1405_, data_stage_4__1404_, data_stage_4__1403_, data_stage_4__1402_, data_stage_4__1401_, data_stage_4__1400_, data_stage_4__1399_, data_stage_4__1398_, data_stage_4__1397_, data_stage_4__1396_, data_stage_4__1395_, data_stage_4__1394_, data_stage_4__1393_, data_stage_4__1392_, data_stage_4__1391_, data_stage_4__1390_, data_stage_4__1389_, data_stage_4__1388_, data_stage_4__1387_, data_stage_4__1386_, data_stage_4__1385_, data_stage_4__1384_, data_stage_4__1383_, data_stage_4__1382_, data_stage_4__1381_, data_stage_4__1380_, data_stage_4__1379_, data_stage_4__1378_, data_stage_4__1377_, data_stage_4__1376_, data_stage_4__1375_, data_stage_4__1374_, data_stage_4__1373_, data_stage_4__1372_, data_stage_4__1371_, data_stage_4__1370_, data_stage_4__1369_, data_stage_4__1368_, data_stage_4__1367_, data_stage_4__1366_, data_stage_4__1365_, data_stage_4__1364_, data_stage_4__1363_, data_stage_4__1362_, data_stage_4__1361_, data_stage_4__1360_, data_stage_4__1359_, data_stage_4__1358_, data_stage_4__1357_, data_stage_4__1356_, data_stage_4__1355_, data_stage_4__1354_, data_stage_4__1353_, data_stage_4__1352_, data_stage_4__1351_, data_stage_4__1350_, data_stage_4__1349_, data_stage_4__1348_, data_stage_4__1347_, data_stage_4__1346_, data_stage_4__1345_, data_stage_4__1344_, data_stage_4__1343_, data_stage_4__1342_, data_stage_4__1341_, data_stage_4__1340_, data_stage_4__1339_, data_stage_4__1338_, data_stage_4__1337_, data_stage_4__1336_, data_stage_4__1335_, data_stage_4__1334_, data_stage_4__1333_, data_stage_4__1332_, data_stage_4__1331_, data_stage_4__1330_, data_stage_4__1329_, data_stage_4__1328_, data_stage_4__1327_, data_stage_4__1326_, data_stage_4__1325_, data_stage_4__1324_, data_stage_4__1323_, data_stage_4__1322_, data_stage_4__1321_, data_stage_4__1320_, data_stage_4__1319_, data_stage_4__1318_, data_stage_4__1317_, data_stage_4__1316_, data_stage_4__1315_, data_stage_4__1314_, data_stage_4__1313_, data_stage_4__1312_, data_stage_4__1311_, data_stage_4__1310_, data_stage_4__1309_, data_stage_4__1308_, data_stage_4__1307_, data_stage_4__1306_, data_stage_4__1305_, data_stage_4__1304_, data_stage_4__1303_, data_stage_4__1302_, data_stage_4__1301_, data_stage_4__1300_, data_stage_4__1299_, data_stage_4__1298_, data_stage_4__1297_, data_stage_4__1296_, data_stage_4__1295_, data_stage_4__1294_, data_stage_4__1293_, data_stage_4__1292_, data_stage_4__1291_, data_stage_4__1290_, data_stage_4__1289_, data_stage_4__1288_, data_stage_4__1287_, data_stage_4__1286_, data_stage_4__1285_, data_stage_4__1284_, data_stage_4__1283_, data_stage_4__1282_, data_stage_4__1281_, data_stage_4__1280_, data_stage_4__1279_, data_stage_4__1278_, data_stage_4__1277_, data_stage_4__1276_, data_stage_4__1275_, data_stage_4__1274_, data_stage_4__1273_, data_stage_4__1272_, data_stage_4__1271_, data_stage_4__1270_, data_stage_4__1269_, data_stage_4__1268_, data_stage_4__1267_, data_stage_4__1266_, data_stage_4__1265_, data_stage_4__1264_, data_stage_4__1263_, data_stage_4__1262_, data_stage_4__1261_, data_stage_4__1260_, data_stage_4__1259_, data_stage_4__1258_, data_stage_4__1257_, data_stage_4__1256_, data_stage_4__1255_, data_stage_4__1254_, data_stage_4__1253_, data_stage_4__1252_, data_stage_4__1251_, data_stage_4__1250_, data_stage_4__1249_, data_stage_4__1248_, data_stage_4__1247_, data_stage_4__1246_, data_stage_4__1245_, data_stage_4__1244_, data_stage_4__1243_, data_stage_4__1242_, data_stage_4__1241_, data_stage_4__1240_, data_stage_4__1239_, data_stage_4__1238_, data_stage_4__1237_, data_stage_4__1236_, data_stage_4__1235_, data_stage_4__1234_, data_stage_4__1233_, data_stage_4__1232_, data_stage_4__1231_, data_stage_4__1230_, data_stage_4__1229_, data_stage_4__1228_, data_stage_4__1227_, data_stage_4__1226_, data_stage_4__1225_, data_stage_4__1224_, data_stage_4__1223_, data_stage_4__1222_, data_stage_4__1221_, data_stage_4__1220_, data_stage_4__1219_, data_stage_4__1218_, data_stage_4__1217_, data_stage_4__1216_, data_stage_4__1215_, data_stage_4__1214_, data_stage_4__1213_, data_stage_4__1212_, data_stage_4__1211_, data_stage_4__1210_, data_stage_4__1209_, data_stage_4__1208_, data_stage_4__1207_, data_stage_4__1206_, data_stage_4__1205_, data_stage_4__1204_, data_stage_4__1203_, data_stage_4__1202_, data_stage_4__1201_, data_stage_4__1200_, data_stage_4__1199_, data_stage_4__1198_, data_stage_4__1197_, data_stage_4__1196_, data_stage_4__1195_, data_stage_4__1194_, data_stage_4__1193_, data_stage_4__1192_, data_stage_4__1191_, data_stage_4__1190_, data_stage_4__1189_, data_stage_4__1188_, data_stage_4__1187_, data_stage_4__1186_, data_stage_4__1185_, data_stage_4__1184_, data_stage_4__1183_, data_stage_4__1182_, data_stage_4__1181_, data_stage_4__1180_, data_stage_4__1179_, data_stage_4__1178_, data_stage_4__1177_, data_stage_4__1176_, data_stage_4__1175_, data_stage_4__1174_, data_stage_4__1173_, data_stage_4__1172_, data_stage_4__1171_, data_stage_4__1170_, data_stage_4__1169_, data_stage_4__1168_, data_stage_4__1167_, data_stage_4__1166_, data_stage_4__1165_, data_stage_4__1164_, data_stage_4__1163_, data_stage_4__1162_, data_stage_4__1161_, data_stage_4__1160_, data_stage_4__1159_, data_stage_4__1158_, data_stage_4__1157_, data_stage_4__1156_, data_stage_4__1155_, data_stage_4__1154_, data_stage_4__1153_, data_stage_4__1152_, data_stage_4__1151_, data_stage_4__1150_, data_stage_4__1149_, data_stage_4__1148_, data_stage_4__1147_, data_stage_4__1146_, data_stage_4__1145_, data_stage_4__1144_, data_stage_4__1143_, data_stage_4__1142_, data_stage_4__1141_, data_stage_4__1140_, data_stage_4__1139_, data_stage_4__1138_, data_stage_4__1137_, data_stage_4__1136_, data_stage_4__1135_, data_stage_4__1134_, data_stage_4__1133_, data_stage_4__1132_, data_stage_4__1131_, data_stage_4__1130_, data_stage_4__1129_, data_stage_4__1128_, data_stage_4__1127_, data_stage_4__1126_, data_stage_4__1125_, data_stage_4__1124_, data_stage_4__1123_, data_stage_4__1122_, data_stage_4__1121_, data_stage_4__1120_, data_stage_4__1119_, data_stage_4__1118_, data_stage_4__1117_, data_stage_4__1116_, data_stage_4__1115_, data_stage_4__1114_, data_stage_4__1113_, data_stage_4__1112_, data_stage_4__1111_, data_stage_4__1110_, data_stage_4__1109_, data_stage_4__1108_, data_stage_4__1107_, data_stage_4__1106_, data_stage_4__1105_, data_stage_4__1104_, data_stage_4__1103_, data_stage_4__1102_, data_stage_4__1101_, data_stage_4__1100_, data_stage_4__1099_, data_stage_4__1098_, data_stage_4__1097_, data_stage_4__1096_, data_stage_4__1095_, data_stage_4__1094_, data_stage_4__1093_, data_stage_4__1092_, data_stage_4__1091_, data_stage_4__1090_, data_stage_4__1089_, data_stage_4__1088_, data_stage_4__1087_, data_stage_4__1086_, data_stage_4__1085_, data_stage_4__1084_, data_stage_4__1083_, data_stage_4__1082_, data_stage_4__1081_, data_stage_4__1080_, data_stage_4__1079_, data_stage_4__1078_, data_stage_4__1077_, data_stage_4__1076_, data_stage_4__1075_, data_stage_4__1074_, data_stage_4__1073_, data_stage_4__1072_, data_stage_4__1071_, data_stage_4__1070_, data_stage_4__1069_, data_stage_4__1068_, data_stage_4__1067_, data_stage_4__1066_, data_stage_4__1065_, data_stage_4__1064_, data_stage_4__1063_, data_stage_4__1062_, data_stage_4__1061_, data_stage_4__1060_, data_stage_4__1059_, data_stage_4__1058_, data_stage_4__1057_, data_stage_4__1056_, data_stage_4__1055_, data_stage_4__1054_, data_stage_4__1053_, data_stage_4__1052_, data_stage_4__1051_, data_stage_4__1050_, data_stage_4__1049_, data_stage_4__1048_, data_stage_4__1047_, data_stage_4__1046_, data_stage_4__1045_, data_stage_4__1044_, data_stage_4__1043_, data_stage_4__1042_, data_stage_4__1041_, data_stage_4__1040_, data_stage_4__1039_, data_stage_4__1038_, data_stage_4__1037_, data_stage_4__1036_, data_stage_4__1035_, data_stage_4__1034_, data_stage_4__1033_, data_stage_4__1032_, data_stage_4__1031_, data_stage_4__1030_, data_stage_4__1029_, data_stage_4__1028_, data_stage_4__1027_, data_stage_4__1026_, data_stage_4__1025_, data_stage_4__1024_, data_stage_4__1023_, data_stage_4__1022_, data_stage_4__1021_, data_stage_4__1020_, data_stage_4__1019_, data_stage_4__1018_, data_stage_4__1017_, data_stage_4__1016_, data_stage_4__1015_, data_stage_4__1014_, data_stage_4__1013_, data_stage_4__1012_, data_stage_4__1011_, data_stage_4__1010_, data_stage_4__1009_, data_stage_4__1008_, data_stage_4__1007_, data_stage_4__1006_, data_stage_4__1005_, data_stage_4__1004_, data_stage_4__1003_, data_stage_4__1002_, data_stage_4__1001_, data_stage_4__1000_, data_stage_4__999_, data_stage_4__998_, data_stage_4__997_, data_stage_4__996_, data_stage_4__995_, data_stage_4__994_, data_stage_4__993_, data_stage_4__992_, data_stage_4__991_, data_stage_4__990_, data_stage_4__989_, data_stage_4__988_, data_stage_4__987_, data_stage_4__986_, data_stage_4__985_, data_stage_4__984_, data_stage_4__983_, data_stage_4__982_, data_stage_4__981_, data_stage_4__980_, data_stage_4__979_, data_stage_4__978_, data_stage_4__977_, data_stage_4__976_, data_stage_4__975_, data_stage_4__974_, data_stage_4__973_, data_stage_4__972_, data_stage_4__971_, data_stage_4__970_, data_stage_4__969_, data_stage_4__968_, data_stage_4__967_, data_stage_4__966_, data_stage_4__965_, data_stage_4__964_, data_stage_4__963_, data_stage_4__962_, data_stage_4__961_, data_stage_4__960_, data_stage_4__959_, data_stage_4__958_, data_stage_4__957_, data_stage_4__956_, data_stage_4__955_, data_stage_4__954_, data_stage_4__953_, data_stage_4__952_, data_stage_4__951_, data_stage_4__950_, data_stage_4__949_, data_stage_4__948_, data_stage_4__947_, data_stage_4__946_, data_stage_4__945_, data_stage_4__944_, data_stage_4__943_, data_stage_4__942_, data_stage_4__941_, data_stage_4__940_, data_stage_4__939_, data_stage_4__938_, data_stage_4__937_, data_stage_4__936_, data_stage_4__935_, data_stage_4__934_, data_stage_4__933_, data_stage_4__932_, data_stage_4__931_, data_stage_4__930_, data_stage_4__929_, data_stage_4__928_, data_stage_4__927_, data_stage_4__926_, data_stage_4__925_, data_stage_4__924_, data_stage_4__923_, data_stage_4__922_, data_stage_4__921_, data_stage_4__920_, data_stage_4__919_, data_stage_4__918_, data_stage_4__917_, data_stage_4__916_, data_stage_4__915_, data_stage_4__914_, data_stage_4__913_, data_stage_4__912_, data_stage_4__911_, data_stage_4__910_, data_stage_4__909_, data_stage_4__908_, data_stage_4__907_, data_stage_4__906_, data_stage_4__905_, data_stage_4__904_, data_stage_4__903_, data_stage_4__902_, data_stage_4__901_, data_stage_4__900_, data_stage_4__899_, data_stage_4__898_, data_stage_4__897_, data_stage_4__896_, data_stage_4__895_, data_stage_4__894_, data_stage_4__893_, data_stage_4__892_, data_stage_4__891_, data_stage_4__890_, data_stage_4__889_, data_stage_4__888_, data_stage_4__887_, data_stage_4__886_, data_stage_4__885_, data_stage_4__884_, data_stage_4__883_, data_stage_4__882_, data_stage_4__881_, data_stage_4__880_, data_stage_4__879_, data_stage_4__878_, data_stage_4__877_, data_stage_4__876_, data_stage_4__875_, data_stage_4__874_, data_stage_4__873_, data_stage_4__872_, data_stage_4__871_, data_stage_4__870_, data_stage_4__869_, data_stage_4__868_, data_stage_4__867_, data_stage_4__866_, data_stage_4__865_, data_stage_4__864_, data_stage_4__863_, data_stage_4__862_, data_stage_4__861_, data_stage_4__860_, data_stage_4__859_, data_stage_4__858_, data_stage_4__857_, data_stage_4__856_, data_stage_4__855_, data_stage_4__854_, data_stage_4__853_, data_stage_4__852_, data_stage_4__851_, data_stage_4__850_, data_stage_4__849_, data_stage_4__848_, data_stage_4__847_, data_stage_4__846_, data_stage_4__845_, data_stage_4__844_, data_stage_4__843_, data_stage_4__842_, data_stage_4__841_, data_stage_4__840_, data_stage_4__839_, data_stage_4__838_, data_stage_4__837_, data_stage_4__836_, data_stage_4__835_, data_stage_4__834_, data_stage_4__833_, data_stage_4__832_, data_stage_4__831_, data_stage_4__830_, data_stage_4__829_, data_stage_4__828_, data_stage_4__827_, data_stage_4__826_, data_stage_4__825_, data_stage_4__824_, data_stage_4__823_, data_stage_4__822_, data_stage_4__821_, data_stage_4__820_, data_stage_4__819_, data_stage_4__818_, data_stage_4__817_, data_stage_4__816_, data_stage_4__815_, data_stage_4__814_, data_stage_4__813_, data_stage_4__812_, data_stage_4__811_, data_stage_4__810_, data_stage_4__809_, data_stage_4__808_, data_stage_4__807_, data_stage_4__806_, data_stage_4__805_, data_stage_4__804_, data_stage_4__803_, data_stage_4__802_, data_stage_4__801_, data_stage_4__800_, data_stage_4__799_, data_stage_4__798_, data_stage_4__797_, data_stage_4__796_, data_stage_4__795_, data_stage_4__794_, data_stage_4__793_, data_stage_4__792_, data_stage_4__791_, data_stage_4__790_, data_stage_4__789_, data_stage_4__788_, data_stage_4__787_, data_stage_4__786_, data_stage_4__785_, data_stage_4__784_, data_stage_4__783_, data_stage_4__782_, data_stage_4__781_, data_stage_4__780_, data_stage_4__779_, data_stage_4__778_, data_stage_4__777_, data_stage_4__776_, data_stage_4__775_, data_stage_4__774_, data_stage_4__773_, data_stage_4__772_, data_stage_4__771_, data_stage_4__770_, data_stage_4__769_, data_stage_4__768_, data_stage_4__767_, data_stage_4__766_, data_stage_4__765_, data_stage_4__764_, data_stage_4__763_, data_stage_4__762_, data_stage_4__761_, data_stage_4__760_, data_stage_4__759_, data_stage_4__758_, data_stage_4__757_, data_stage_4__756_, data_stage_4__755_, data_stage_4__754_, data_stage_4__753_, data_stage_4__752_, data_stage_4__751_, data_stage_4__750_, data_stage_4__749_, data_stage_4__748_, data_stage_4__747_, data_stage_4__746_, data_stage_4__745_, data_stage_4__744_, data_stage_4__743_, data_stage_4__742_, data_stage_4__741_, data_stage_4__740_, data_stage_4__739_, data_stage_4__738_, data_stage_4__737_, data_stage_4__736_, data_stage_4__735_, data_stage_4__734_, data_stage_4__733_, data_stage_4__732_, data_stage_4__731_, data_stage_4__730_, data_stage_4__729_, data_stage_4__728_, data_stage_4__727_, data_stage_4__726_, data_stage_4__725_, data_stage_4__724_, data_stage_4__723_, data_stage_4__722_, data_stage_4__721_, data_stage_4__720_, data_stage_4__719_, data_stage_4__718_, data_stage_4__717_, data_stage_4__716_, data_stage_4__715_, data_stage_4__714_, data_stage_4__713_, data_stage_4__712_, data_stage_4__711_, data_stage_4__710_, data_stage_4__709_, data_stage_4__708_, data_stage_4__707_, data_stage_4__706_, data_stage_4__705_, data_stage_4__704_, data_stage_4__703_, data_stage_4__702_, data_stage_4__701_, data_stage_4__700_, data_stage_4__699_, data_stage_4__698_, data_stage_4__697_, data_stage_4__696_, data_stage_4__695_, data_stage_4__694_, data_stage_4__693_, data_stage_4__692_, data_stage_4__691_, data_stage_4__690_, data_stage_4__689_, data_stage_4__688_, data_stage_4__687_, data_stage_4__686_, data_stage_4__685_, data_stage_4__684_, data_stage_4__683_, data_stage_4__682_, data_stage_4__681_, data_stage_4__680_, data_stage_4__679_, data_stage_4__678_, data_stage_4__677_, data_stage_4__676_, data_stage_4__675_, data_stage_4__674_, data_stage_4__673_, data_stage_4__672_, data_stage_4__671_, data_stage_4__670_, data_stage_4__669_, data_stage_4__668_, data_stage_4__667_, data_stage_4__666_, data_stage_4__665_, data_stage_4__664_, data_stage_4__663_, data_stage_4__662_, data_stage_4__661_, data_stage_4__660_, data_stage_4__659_, data_stage_4__658_, data_stage_4__657_, data_stage_4__656_, data_stage_4__655_, data_stage_4__654_, data_stage_4__653_, data_stage_4__652_, data_stage_4__651_, data_stage_4__650_, data_stage_4__649_, data_stage_4__648_, data_stage_4__647_, data_stage_4__646_, data_stage_4__645_, data_stage_4__644_, data_stage_4__643_, data_stage_4__642_, data_stage_4__641_, data_stage_4__640_, data_stage_4__639_, data_stage_4__638_, data_stage_4__637_, data_stage_4__636_, data_stage_4__635_, data_stage_4__634_, data_stage_4__633_, data_stage_4__632_, data_stage_4__631_, data_stage_4__630_, data_stage_4__629_, data_stage_4__628_, data_stage_4__627_, data_stage_4__626_, data_stage_4__625_, data_stage_4__624_, data_stage_4__623_, data_stage_4__622_, data_stage_4__621_, data_stage_4__620_, data_stage_4__619_, data_stage_4__618_, data_stage_4__617_, data_stage_4__616_, data_stage_4__615_, data_stage_4__614_, data_stage_4__613_, data_stage_4__612_, data_stage_4__611_, data_stage_4__610_, data_stage_4__609_, data_stage_4__608_, data_stage_4__607_, data_stage_4__606_, data_stage_4__605_, data_stage_4__604_, data_stage_4__603_, data_stage_4__602_, data_stage_4__601_, data_stage_4__600_, data_stage_4__599_, data_stage_4__598_, data_stage_4__597_, data_stage_4__596_, data_stage_4__595_, data_stage_4__594_, data_stage_4__593_, data_stage_4__592_, data_stage_4__591_, data_stage_4__590_, data_stage_4__589_, data_stage_4__588_, data_stage_4__587_, data_stage_4__586_, data_stage_4__585_, data_stage_4__584_, data_stage_4__583_, data_stage_4__582_, data_stage_4__581_, data_stage_4__580_, data_stage_4__579_, data_stage_4__578_, data_stage_4__577_, data_stage_4__576_, data_stage_4__575_, data_stage_4__574_, data_stage_4__573_, data_stage_4__572_, data_stage_4__571_, data_stage_4__570_, data_stage_4__569_, data_stage_4__568_, data_stage_4__567_, data_stage_4__566_, data_stage_4__565_, data_stage_4__564_, data_stage_4__563_, data_stage_4__562_, data_stage_4__561_, data_stage_4__560_, data_stage_4__559_, data_stage_4__558_, data_stage_4__557_, data_stage_4__556_, data_stage_4__555_, data_stage_4__554_, data_stage_4__553_, data_stage_4__552_, data_stage_4__551_, data_stage_4__550_, data_stage_4__549_, data_stage_4__548_, data_stage_4__547_, data_stage_4__546_, data_stage_4__545_, data_stage_4__544_, data_stage_4__543_, data_stage_4__542_, data_stage_4__541_, data_stage_4__540_, data_stage_4__539_, data_stage_4__538_, data_stage_4__537_, data_stage_4__536_, data_stage_4__535_, data_stage_4__534_, data_stage_4__533_, data_stage_4__532_, data_stage_4__531_, data_stage_4__530_, data_stage_4__529_, data_stage_4__528_, data_stage_4__527_, data_stage_4__526_, data_stage_4__525_, data_stage_4__524_, data_stage_4__523_, data_stage_4__522_, data_stage_4__521_, data_stage_4__520_, data_stage_4__519_, data_stage_4__518_, data_stage_4__517_, data_stage_4__516_, data_stage_4__515_, data_stage_4__514_, data_stage_4__513_, data_stage_4__512_, data_stage_4__511_, data_stage_4__510_, data_stage_4__509_, data_stage_4__508_, data_stage_4__507_, data_stage_4__506_, data_stage_4__505_, data_stage_4__504_, data_stage_4__503_, data_stage_4__502_, data_stage_4__501_, data_stage_4__500_, data_stage_4__499_, data_stage_4__498_, data_stage_4__497_, data_stage_4__496_, data_stage_4__495_, data_stage_4__494_, data_stage_4__493_, data_stage_4__492_, data_stage_4__491_, data_stage_4__490_, data_stage_4__489_, data_stage_4__488_, data_stage_4__487_, data_stage_4__486_, data_stage_4__485_, data_stage_4__484_, data_stage_4__483_, data_stage_4__482_, data_stage_4__481_, data_stage_4__480_, data_stage_4__479_, data_stage_4__478_, data_stage_4__477_, data_stage_4__476_, data_stage_4__475_, data_stage_4__474_, data_stage_4__473_, data_stage_4__472_, data_stage_4__471_, data_stage_4__470_, data_stage_4__469_, data_stage_4__468_, data_stage_4__467_, data_stage_4__466_, data_stage_4__465_, data_stage_4__464_, data_stage_4__463_, data_stage_4__462_, data_stage_4__461_, data_stage_4__460_, data_stage_4__459_, data_stage_4__458_, data_stage_4__457_, data_stage_4__456_, data_stage_4__455_, data_stage_4__454_, data_stage_4__453_, data_stage_4__452_, data_stage_4__451_, data_stage_4__450_, data_stage_4__449_, data_stage_4__448_, data_stage_4__447_, data_stage_4__446_, data_stage_4__445_, data_stage_4__444_, data_stage_4__443_, data_stage_4__442_, data_stage_4__441_, data_stage_4__440_, data_stage_4__439_, data_stage_4__438_, data_stage_4__437_, data_stage_4__436_, data_stage_4__435_, data_stage_4__434_, data_stage_4__433_, data_stage_4__432_, data_stage_4__431_, data_stage_4__430_, data_stage_4__429_, data_stage_4__428_, data_stage_4__427_, data_stage_4__426_, data_stage_4__425_, data_stage_4__424_, data_stage_4__423_, data_stage_4__422_, data_stage_4__421_, data_stage_4__420_, data_stage_4__419_, data_stage_4__418_, data_stage_4__417_, data_stage_4__416_, data_stage_4__415_, data_stage_4__414_, data_stage_4__413_, data_stage_4__412_, data_stage_4__411_, data_stage_4__410_, data_stage_4__409_, data_stage_4__408_, data_stage_4__407_, data_stage_4__406_, data_stage_4__405_, data_stage_4__404_, data_stage_4__403_, data_stage_4__402_, data_stage_4__401_, data_stage_4__400_, data_stage_4__399_, data_stage_4__398_, data_stage_4__397_, data_stage_4__396_, data_stage_4__395_, data_stage_4__394_, data_stage_4__393_, data_stage_4__392_, data_stage_4__391_, data_stage_4__390_, data_stage_4__389_, data_stage_4__388_, data_stage_4__387_, data_stage_4__386_, data_stage_4__385_, data_stage_4__384_, data_stage_4__383_, data_stage_4__382_, data_stage_4__381_, data_stage_4__380_, data_stage_4__379_, data_stage_4__378_, data_stage_4__377_, data_stage_4__376_, data_stage_4__375_, data_stage_4__374_, data_stage_4__373_, data_stage_4__372_, data_stage_4__371_, data_stage_4__370_, data_stage_4__369_, data_stage_4__368_, data_stage_4__367_, data_stage_4__366_, data_stage_4__365_, data_stage_4__364_, data_stage_4__363_, data_stage_4__362_, data_stage_4__361_, data_stage_4__360_, data_stage_4__359_, data_stage_4__358_, data_stage_4__357_, data_stage_4__356_, data_stage_4__355_, data_stage_4__354_, data_stage_4__353_, data_stage_4__352_, data_stage_4__351_, data_stage_4__350_, data_stage_4__349_, data_stage_4__348_, data_stage_4__347_, data_stage_4__346_, data_stage_4__345_, data_stage_4__344_, data_stage_4__343_, data_stage_4__342_, data_stage_4__341_, data_stage_4__340_, data_stage_4__339_, data_stage_4__338_, data_stage_4__337_, data_stage_4__336_, data_stage_4__335_, data_stage_4__334_, data_stage_4__333_, data_stage_4__332_, data_stage_4__331_, data_stage_4__330_, data_stage_4__329_, data_stage_4__328_, data_stage_4__327_, data_stage_4__326_, data_stage_4__325_, data_stage_4__324_, data_stage_4__323_, data_stage_4__322_, data_stage_4__321_, data_stage_4__320_, data_stage_4__319_, data_stage_4__318_, data_stage_4__317_, data_stage_4__316_, data_stage_4__315_, data_stage_4__314_, data_stage_4__313_, data_stage_4__312_, data_stage_4__311_, data_stage_4__310_, data_stage_4__309_, data_stage_4__308_, data_stage_4__307_, data_stage_4__306_, data_stage_4__305_, data_stage_4__304_, data_stage_4__303_, data_stage_4__302_, data_stage_4__301_, data_stage_4__300_, data_stage_4__299_, data_stage_4__298_, data_stage_4__297_, data_stage_4__296_, data_stage_4__295_, data_stage_4__294_, data_stage_4__293_, data_stage_4__292_, data_stage_4__291_, data_stage_4__290_, data_stage_4__289_, data_stage_4__288_, data_stage_4__287_, data_stage_4__286_, data_stage_4__285_, data_stage_4__284_, data_stage_4__283_, data_stage_4__282_, data_stage_4__281_, data_stage_4__280_, data_stage_4__279_, data_stage_4__278_, data_stage_4__277_, data_stage_4__276_, data_stage_4__275_, data_stage_4__274_, data_stage_4__273_, data_stage_4__272_, data_stage_4__271_, data_stage_4__270_, data_stage_4__269_, data_stage_4__268_, data_stage_4__267_, data_stage_4__266_, data_stage_4__265_, data_stage_4__264_, data_stage_4__263_, data_stage_4__262_, data_stage_4__261_, data_stage_4__260_, data_stage_4__259_, data_stage_4__258_, data_stage_4__257_, data_stage_4__256_, data_stage_4__255_, data_stage_4__254_, data_stage_4__253_, data_stage_4__252_, data_stage_4__251_, data_stage_4__250_, data_stage_4__249_, data_stage_4__248_, data_stage_4__247_, data_stage_4__246_, data_stage_4__245_, data_stage_4__244_, data_stage_4__243_, data_stage_4__242_, data_stage_4__241_, data_stage_4__240_, data_stage_4__239_, data_stage_4__238_, data_stage_4__237_, data_stage_4__236_, data_stage_4__235_, data_stage_4__234_, data_stage_4__233_, data_stage_4__232_, data_stage_4__231_, data_stage_4__230_, data_stage_4__229_, data_stage_4__228_, data_stage_4__227_, data_stage_4__226_, data_stage_4__225_, data_stage_4__224_, data_stage_4__223_, data_stage_4__222_, data_stage_4__221_, data_stage_4__220_, data_stage_4__219_, data_stage_4__218_, data_stage_4__217_, data_stage_4__216_, data_stage_4__215_, data_stage_4__214_, data_stage_4__213_, data_stage_4__212_, data_stage_4__211_, data_stage_4__210_, data_stage_4__209_, data_stage_4__208_, data_stage_4__207_, data_stage_4__206_, data_stage_4__205_, data_stage_4__204_, data_stage_4__203_, data_stage_4__202_, data_stage_4__201_, data_stage_4__200_, data_stage_4__199_, data_stage_4__198_, data_stage_4__197_, data_stage_4__196_, data_stage_4__195_, data_stage_4__194_, data_stage_4__193_, data_stage_4__192_, data_stage_4__191_, data_stage_4__190_, data_stage_4__189_, data_stage_4__188_, data_stage_4__187_, data_stage_4__186_, data_stage_4__185_, data_stage_4__184_, data_stage_4__183_, data_stage_4__182_, data_stage_4__181_, data_stage_4__180_, data_stage_4__179_, data_stage_4__178_, data_stage_4__177_, data_stage_4__176_, data_stage_4__175_, data_stage_4__174_, data_stage_4__173_, data_stage_4__172_, data_stage_4__171_, data_stage_4__170_, data_stage_4__169_, data_stage_4__168_, data_stage_4__167_, data_stage_4__166_, data_stage_4__165_, data_stage_4__164_, data_stage_4__163_, data_stage_4__162_, data_stage_4__161_, data_stage_4__160_, data_stage_4__159_, data_stage_4__158_, data_stage_4__157_, data_stage_4__156_, data_stage_4__155_, data_stage_4__154_, data_stage_4__153_, data_stage_4__152_, data_stage_4__151_, data_stage_4__150_, data_stage_4__149_, data_stage_4__148_, data_stage_4__147_, data_stage_4__146_, data_stage_4__145_, data_stage_4__144_, data_stage_4__143_, data_stage_4__142_, data_stage_4__141_, data_stage_4__140_, data_stage_4__139_, data_stage_4__138_, data_stage_4__137_, data_stage_4__136_, data_stage_4__135_, data_stage_4__134_, data_stage_4__133_, data_stage_4__132_, data_stage_4__131_, data_stage_4__130_, data_stage_4__129_, data_stage_4__128_, data_stage_4__127_, data_stage_4__126_, data_stage_4__125_, data_stage_4__124_, data_stage_4__123_, data_stage_4__122_, data_stage_4__121_, data_stage_4__120_, data_stage_4__119_, data_stage_4__118_, data_stage_4__117_, data_stage_4__116_, data_stage_4__115_, data_stage_4__114_, data_stage_4__113_, data_stage_4__112_, data_stage_4__111_, data_stage_4__110_, data_stage_4__109_, data_stage_4__108_, data_stage_4__107_, data_stage_4__106_, data_stage_4__105_, data_stage_4__104_, data_stage_4__103_, data_stage_4__102_, data_stage_4__101_, data_stage_4__100_, data_stage_4__99_, data_stage_4__98_, data_stage_4__97_, data_stage_4__96_, data_stage_4__95_, data_stage_4__94_, data_stage_4__93_, data_stage_4__92_, data_stage_4__91_, data_stage_4__90_, data_stage_4__89_, data_stage_4__88_, data_stage_4__87_, data_stage_4__86_, data_stage_4__85_, data_stage_4__84_, data_stage_4__83_, data_stage_4__82_, data_stage_4__81_, data_stage_4__80_, data_stage_4__79_, data_stage_4__78_, data_stage_4__77_, data_stage_4__76_, data_stage_4__75_, data_stage_4__74_, data_stage_4__73_, data_stage_4__72_, data_stage_4__71_, data_stage_4__70_, data_stage_4__69_, data_stage_4__68_, data_stage_4__67_, data_stage_4__66_, data_stage_4__65_, data_stage_4__64_, data_stage_4__63_, data_stage_4__62_, data_stage_4__61_, data_stage_4__60_, data_stage_4__59_, data_stage_4__58_, data_stage_4__57_, data_stage_4__56_, data_stage_4__55_, data_stage_4__54_, data_stage_4__53_, data_stage_4__52_, data_stage_4__51_, data_stage_4__50_, data_stage_4__49_, data_stage_4__48_, data_stage_4__47_, data_stage_4__46_, data_stage_4__45_, data_stage_4__44_, data_stage_4__43_, data_stage_4__42_, data_stage_4__41_, data_stage_4__40_, data_stage_4__39_, data_stage_4__38_, data_stage_4__37_, data_stage_4__36_, data_stage_4__35_, data_stage_4__34_, data_stage_4__33_, data_stage_4__32_, data_stage_4__31_, data_stage_4__30_, data_stage_4__29_, data_stage_4__28_, data_stage_4__27_, data_stage_4__26_, data_stage_4__25_, data_stage_4__24_, data_stage_4__23_, data_stage_4__22_, data_stage_4__21_, data_stage_4__20_, data_stage_4__19_, data_stage_4__18_, data_stage_4__17_, data_stage_4__16_, data_stage_4__15_, data_stage_4__14_, data_stage_4__13_, data_stage_4__12_, data_stage_4__11_, data_stage_4__10_, data_stage_4__9_, data_stage_4__8_, data_stage_4__7_, data_stage_4__6_, data_stage_4__5_, data_stage_4__4_, data_stage_4__3_, data_stage_4__2_, data_stage_4__1_, data_stage_4__0_ }),
    .swap_i(sel_i[4]),
    .data_o({ data_stage_5__2047_, data_stage_5__2046_, data_stage_5__2045_, data_stage_5__2044_, data_stage_5__2043_, data_stage_5__2042_, data_stage_5__2041_, data_stage_5__2040_, data_stage_5__2039_, data_stage_5__2038_, data_stage_5__2037_, data_stage_5__2036_, data_stage_5__2035_, data_stage_5__2034_, data_stage_5__2033_, data_stage_5__2032_, data_stage_5__2031_, data_stage_5__2030_, data_stage_5__2029_, data_stage_5__2028_, data_stage_5__2027_, data_stage_5__2026_, data_stage_5__2025_, data_stage_5__2024_, data_stage_5__2023_, data_stage_5__2022_, data_stage_5__2021_, data_stage_5__2020_, data_stage_5__2019_, data_stage_5__2018_, data_stage_5__2017_, data_stage_5__2016_, data_stage_5__2015_, data_stage_5__2014_, data_stage_5__2013_, data_stage_5__2012_, data_stage_5__2011_, data_stage_5__2010_, data_stage_5__2009_, data_stage_5__2008_, data_stage_5__2007_, data_stage_5__2006_, data_stage_5__2005_, data_stage_5__2004_, data_stage_5__2003_, data_stage_5__2002_, data_stage_5__2001_, data_stage_5__2000_, data_stage_5__1999_, data_stage_5__1998_, data_stage_5__1997_, data_stage_5__1996_, data_stage_5__1995_, data_stage_5__1994_, data_stage_5__1993_, data_stage_5__1992_, data_stage_5__1991_, data_stage_5__1990_, data_stage_5__1989_, data_stage_5__1988_, data_stage_5__1987_, data_stage_5__1986_, data_stage_5__1985_, data_stage_5__1984_, data_stage_5__1983_, data_stage_5__1982_, data_stage_5__1981_, data_stage_5__1980_, data_stage_5__1979_, data_stage_5__1978_, data_stage_5__1977_, data_stage_5__1976_, data_stage_5__1975_, data_stage_5__1974_, data_stage_5__1973_, data_stage_5__1972_, data_stage_5__1971_, data_stage_5__1970_, data_stage_5__1969_, data_stage_5__1968_, data_stage_5__1967_, data_stage_5__1966_, data_stage_5__1965_, data_stage_5__1964_, data_stage_5__1963_, data_stage_5__1962_, data_stage_5__1961_, data_stage_5__1960_, data_stage_5__1959_, data_stage_5__1958_, data_stage_5__1957_, data_stage_5__1956_, data_stage_5__1955_, data_stage_5__1954_, data_stage_5__1953_, data_stage_5__1952_, data_stage_5__1951_, data_stage_5__1950_, data_stage_5__1949_, data_stage_5__1948_, data_stage_5__1947_, data_stage_5__1946_, data_stage_5__1945_, data_stage_5__1944_, data_stage_5__1943_, data_stage_5__1942_, data_stage_5__1941_, data_stage_5__1940_, data_stage_5__1939_, data_stage_5__1938_, data_stage_5__1937_, data_stage_5__1936_, data_stage_5__1935_, data_stage_5__1934_, data_stage_5__1933_, data_stage_5__1932_, data_stage_5__1931_, data_stage_5__1930_, data_stage_5__1929_, data_stage_5__1928_, data_stage_5__1927_, data_stage_5__1926_, data_stage_5__1925_, data_stage_5__1924_, data_stage_5__1923_, data_stage_5__1922_, data_stage_5__1921_, data_stage_5__1920_, data_stage_5__1919_, data_stage_5__1918_, data_stage_5__1917_, data_stage_5__1916_, data_stage_5__1915_, data_stage_5__1914_, data_stage_5__1913_, data_stage_5__1912_, data_stage_5__1911_, data_stage_5__1910_, data_stage_5__1909_, data_stage_5__1908_, data_stage_5__1907_, data_stage_5__1906_, data_stage_5__1905_, data_stage_5__1904_, data_stage_5__1903_, data_stage_5__1902_, data_stage_5__1901_, data_stage_5__1900_, data_stage_5__1899_, data_stage_5__1898_, data_stage_5__1897_, data_stage_5__1896_, data_stage_5__1895_, data_stage_5__1894_, data_stage_5__1893_, data_stage_5__1892_, data_stage_5__1891_, data_stage_5__1890_, data_stage_5__1889_, data_stage_5__1888_, data_stage_5__1887_, data_stage_5__1886_, data_stage_5__1885_, data_stage_5__1884_, data_stage_5__1883_, data_stage_5__1882_, data_stage_5__1881_, data_stage_5__1880_, data_stage_5__1879_, data_stage_5__1878_, data_stage_5__1877_, data_stage_5__1876_, data_stage_5__1875_, data_stage_5__1874_, data_stage_5__1873_, data_stage_5__1872_, data_stage_5__1871_, data_stage_5__1870_, data_stage_5__1869_, data_stage_5__1868_, data_stage_5__1867_, data_stage_5__1866_, data_stage_5__1865_, data_stage_5__1864_, data_stage_5__1863_, data_stage_5__1862_, data_stage_5__1861_, data_stage_5__1860_, data_stage_5__1859_, data_stage_5__1858_, data_stage_5__1857_, data_stage_5__1856_, data_stage_5__1855_, data_stage_5__1854_, data_stage_5__1853_, data_stage_5__1852_, data_stage_5__1851_, data_stage_5__1850_, data_stage_5__1849_, data_stage_5__1848_, data_stage_5__1847_, data_stage_5__1846_, data_stage_5__1845_, data_stage_5__1844_, data_stage_5__1843_, data_stage_5__1842_, data_stage_5__1841_, data_stage_5__1840_, data_stage_5__1839_, data_stage_5__1838_, data_stage_5__1837_, data_stage_5__1836_, data_stage_5__1835_, data_stage_5__1834_, data_stage_5__1833_, data_stage_5__1832_, data_stage_5__1831_, data_stage_5__1830_, data_stage_5__1829_, data_stage_5__1828_, data_stage_5__1827_, data_stage_5__1826_, data_stage_5__1825_, data_stage_5__1824_, data_stage_5__1823_, data_stage_5__1822_, data_stage_5__1821_, data_stage_5__1820_, data_stage_5__1819_, data_stage_5__1818_, data_stage_5__1817_, data_stage_5__1816_, data_stage_5__1815_, data_stage_5__1814_, data_stage_5__1813_, data_stage_5__1812_, data_stage_5__1811_, data_stage_5__1810_, data_stage_5__1809_, data_stage_5__1808_, data_stage_5__1807_, data_stage_5__1806_, data_stage_5__1805_, data_stage_5__1804_, data_stage_5__1803_, data_stage_5__1802_, data_stage_5__1801_, data_stage_5__1800_, data_stage_5__1799_, data_stage_5__1798_, data_stage_5__1797_, data_stage_5__1796_, data_stage_5__1795_, data_stage_5__1794_, data_stage_5__1793_, data_stage_5__1792_, data_stage_5__1791_, data_stage_5__1790_, data_stage_5__1789_, data_stage_5__1788_, data_stage_5__1787_, data_stage_5__1786_, data_stage_5__1785_, data_stage_5__1784_, data_stage_5__1783_, data_stage_5__1782_, data_stage_5__1781_, data_stage_5__1780_, data_stage_5__1779_, data_stage_5__1778_, data_stage_5__1777_, data_stage_5__1776_, data_stage_5__1775_, data_stage_5__1774_, data_stage_5__1773_, data_stage_5__1772_, data_stage_5__1771_, data_stage_5__1770_, data_stage_5__1769_, data_stage_5__1768_, data_stage_5__1767_, data_stage_5__1766_, data_stage_5__1765_, data_stage_5__1764_, data_stage_5__1763_, data_stage_5__1762_, data_stage_5__1761_, data_stage_5__1760_, data_stage_5__1759_, data_stage_5__1758_, data_stage_5__1757_, data_stage_5__1756_, data_stage_5__1755_, data_stage_5__1754_, data_stage_5__1753_, data_stage_5__1752_, data_stage_5__1751_, data_stage_5__1750_, data_stage_5__1749_, data_stage_5__1748_, data_stage_5__1747_, data_stage_5__1746_, data_stage_5__1745_, data_stage_5__1744_, data_stage_5__1743_, data_stage_5__1742_, data_stage_5__1741_, data_stage_5__1740_, data_stage_5__1739_, data_stage_5__1738_, data_stage_5__1737_, data_stage_5__1736_, data_stage_5__1735_, data_stage_5__1734_, data_stage_5__1733_, data_stage_5__1732_, data_stage_5__1731_, data_stage_5__1730_, data_stage_5__1729_, data_stage_5__1728_, data_stage_5__1727_, data_stage_5__1726_, data_stage_5__1725_, data_stage_5__1724_, data_stage_5__1723_, data_stage_5__1722_, data_stage_5__1721_, data_stage_5__1720_, data_stage_5__1719_, data_stage_5__1718_, data_stage_5__1717_, data_stage_5__1716_, data_stage_5__1715_, data_stage_5__1714_, data_stage_5__1713_, data_stage_5__1712_, data_stage_5__1711_, data_stage_5__1710_, data_stage_5__1709_, data_stage_5__1708_, data_stage_5__1707_, data_stage_5__1706_, data_stage_5__1705_, data_stage_5__1704_, data_stage_5__1703_, data_stage_5__1702_, data_stage_5__1701_, data_stage_5__1700_, data_stage_5__1699_, data_stage_5__1698_, data_stage_5__1697_, data_stage_5__1696_, data_stage_5__1695_, data_stage_5__1694_, data_stage_5__1693_, data_stage_5__1692_, data_stage_5__1691_, data_stage_5__1690_, data_stage_5__1689_, data_stage_5__1688_, data_stage_5__1687_, data_stage_5__1686_, data_stage_5__1685_, data_stage_5__1684_, data_stage_5__1683_, data_stage_5__1682_, data_stage_5__1681_, data_stage_5__1680_, data_stage_5__1679_, data_stage_5__1678_, data_stage_5__1677_, data_stage_5__1676_, data_stage_5__1675_, data_stage_5__1674_, data_stage_5__1673_, data_stage_5__1672_, data_stage_5__1671_, data_stage_5__1670_, data_stage_5__1669_, data_stage_5__1668_, data_stage_5__1667_, data_stage_5__1666_, data_stage_5__1665_, data_stage_5__1664_, data_stage_5__1663_, data_stage_5__1662_, data_stage_5__1661_, data_stage_5__1660_, data_stage_5__1659_, data_stage_5__1658_, data_stage_5__1657_, data_stage_5__1656_, data_stage_5__1655_, data_stage_5__1654_, data_stage_5__1653_, data_stage_5__1652_, data_stage_5__1651_, data_stage_5__1650_, data_stage_5__1649_, data_stage_5__1648_, data_stage_5__1647_, data_stage_5__1646_, data_stage_5__1645_, data_stage_5__1644_, data_stage_5__1643_, data_stage_5__1642_, data_stage_5__1641_, data_stage_5__1640_, data_stage_5__1639_, data_stage_5__1638_, data_stage_5__1637_, data_stage_5__1636_, data_stage_5__1635_, data_stage_5__1634_, data_stage_5__1633_, data_stage_5__1632_, data_stage_5__1631_, data_stage_5__1630_, data_stage_5__1629_, data_stage_5__1628_, data_stage_5__1627_, data_stage_5__1626_, data_stage_5__1625_, data_stage_5__1624_, data_stage_5__1623_, data_stage_5__1622_, data_stage_5__1621_, data_stage_5__1620_, data_stage_5__1619_, data_stage_5__1618_, data_stage_5__1617_, data_stage_5__1616_, data_stage_5__1615_, data_stage_5__1614_, data_stage_5__1613_, data_stage_5__1612_, data_stage_5__1611_, data_stage_5__1610_, data_stage_5__1609_, data_stage_5__1608_, data_stage_5__1607_, data_stage_5__1606_, data_stage_5__1605_, data_stage_5__1604_, data_stage_5__1603_, data_stage_5__1602_, data_stage_5__1601_, data_stage_5__1600_, data_stage_5__1599_, data_stage_5__1598_, data_stage_5__1597_, data_stage_5__1596_, data_stage_5__1595_, data_stage_5__1594_, data_stage_5__1593_, data_stage_5__1592_, data_stage_5__1591_, data_stage_5__1590_, data_stage_5__1589_, data_stage_5__1588_, data_stage_5__1587_, data_stage_5__1586_, data_stage_5__1585_, data_stage_5__1584_, data_stage_5__1583_, data_stage_5__1582_, data_stage_5__1581_, data_stage_5__1580_, data_stage_5__1579_, data_stage_5__1578_, data_stage_5__1577_, data_stage_5__1576_, data_stage_5__1575_, data_stage_5__1574_, data_stage_5__1573_, data_stage_5__1572_, data_stage_5__1571_, data_stage_5__1570_, data_stage_5__1569_, data_stage_5__1568_, data_stage_5__1567_, data_stage_5__1566_, data_stage_5__1565_, data_stage_5__1564_, data_stage_5__1563_, data_stage_5__1562_, data_stage_5__1561_, data_stage_5__1560_, data_stage_5__1559_, data_stage_5__1558_, data_stage_5__1557_, data_stage_5__1556_, data_stage_5__1555_, data_stage_5__1554_, data_stage_5__1553_, data_stage_5__1552_, data_stage_5__1551_, data_stage_5__1550_, data_stage_5__1549_, data_stage_5__1548_, data_stage_5__1547_, data_stage_5__1546_, data_stage_5__1545_, data_stage_5__1544_, data_stage_5__1543_, data_stage_5__1542_, data_stage_5__1541_, data_stage_5__1540_, data_stage_5__1539_, data_stage_5__1538_, data_stage_5__1537_, data_stage_5__1536_, data_stage_5__1535_, data_stage_5__1534_, data_stage_5__1533_, data_stage_5__1532_, data_stage_5__1531_, data_stage_5__1530_, data_stage_5__1529_, data_stage_5__1528_, data_stage_5__1527_, data_stage_5__1526_, data_stage_5__1525_, data_stage_5__1524_, data_stage_5__1523_, data_stage_5__1522_, data_stage_5__1521_, data_stage_5__1520_, data_stage_5__1519_, data_stage_5__1518_, data_stage_5__1517_, data_stage_5__1516_, data_stage_5__1515_, data_stage_5__1514_, data_stage_5__1513_, data_stage_5__1512_, data_stage_5__1511_, data_stage_5__1510_, data_stage_5__1509_, data_stage_5__1508_, data_stage_5__1507_, data_stage_5__1506_, data_stage_5__1505_, data_stage_5__1504_, data_stage_5__1503_, data_stage_5__1502_, data_stage_5__1501_, data_stage_5__1500_, data_stage_5__1499_, data_stage_5__1498_, data_stage_5__1497_, data_stage_5__1496_, data_stage_5__1495_, data_stage_5__1494_, data_stage_5__1493_, data_stage_5__1492_, data_stage_5__1491_, data_stage_5__1490_, data_stage_5__1489_, data_stage_5__1488_, data_stage_5__1487_, data_stage_5__1486_, data_stage_5__1485_, data_stage_5__1484_, data_stage_5__1483_, data_stage_5__1482_, data_stage_5__1481_, data_stage_5__1480_, data_stage_5__1479_, data_stage_5__1478_, data_stage_5__1477_, data_stage_5__1476_, data_stage_5__1475_, data_stage_5__1474_, data_stage_5__1473_, data_stage_5__1472_, data_stage_5__1471_, data_stage_5__1470_, data_stage_5__1469_, data_stage_5__1468_, data_stage_5__1467_, data_stage_5__1466_, data_stage_5__1465_, data_stage_5__1464_, data_stage_5__1463_, data_stage_5__1462_, data_stage_5__1461_, data_stage_5__1460_, data_stage_5__1459_, data_stage_5__1458_, data_stage_5__1457_, data_stage_5__1456_, data_stage_5__1455_, data_stage_5__1454_, data_stage_5__1453_, data_stage_5__1452_, data_stage_5__1451_, data_stage_5__1450_, data_stage_5__1449_, data_stage_5__1448_, data_stage_5__1447_, data_stage_5__1446_, data_stage_5__1445_, data_stage_5__1444_, data_stage_5__1443_, data_stage_5__1442_, data_stage_5__1441_, data_stage_5__1440_, data_stage_5__1439_, data_stage_5__1438_, data_stage_5__1437_, data_stage_5__1436_, data_stage_5__1435_, data_stage_5__1434_, data_stage_5__1433_, data_stage_5__1432_, data_stage_5__1431_, data_stage_5__1430_, data_stage_5__1429_, data_stage_5__1428_, data_stage_5__1427_, data_stage_5__1426_, data_stage_5__1425_, data_stage_5__1424_, data_stage_5__1423_, data_stage_5__1422_, data_stage_5__1421_, data_stage_5__1420_, data_stage_5__1419_, data_stage_5__1418_, data_stage_5__1417_, data_stage_5__1416_, data_stage_5__1415_, data_stage_5__1414_, data_stage_5__1413_, data_stage_5__1412_, data_stage_5__1411_, data_stage_5__1410_, data_stage_5__1409_, data_stage_5__1408_, data_stage_5__1407_, data_stage_5__1406_, data_stage_5__1405_, data_stage_5__1404_, data_stage_5__1403_, data_stage_5__1402_, data_stage_5__1401_, data_stage_5__1400_, data_stage_5__1399_, data_stage_5__1398_, data_stage_5__1397_, data_stage_5__1396_, data_stage_5__1395_, data_stage_5__1394_, data_stage_5__1393_, data_stage_5__1392_, data_stage_5__1391_, data_stage_5__1390_, data_stage_5__1389_, data_stage_5__1388_, data_stage_5__1387_, data_stage_5__1386_, data_stage_5__1385_, data_stage_5__1384_, data_stage_5__1383_, data_stage_5__1382_, data_stage_5__1381_, data_stage_5__1380_, data_stage_5__1379_, data_stage_5__1378_, data_stage_5__1377_, data_stage_5__1376_, data_stage_5__1375_, data_stage_5__1374_, data_stage_5__1373_, data_stage_5__1372_, data_stage_5__1371_, data_stage_5__1370_, data_stage_5__1369_, data_stage_5__1368_, data_stage_5__1367_, data_stage_5__1366_, data_stage_5__1365_, data_stage_5__1364_, data_stage_5__1363_, data_stage_5__1362_, data_stage_5__1361_, data_stage_5__1360_, data_stage_5__1359_, data_stage_5__1358_, data_stage_5__1357_, data_stage_5__1356_, data_stage_5__1355_, data_stage_5__1354_, data_stage_5__1353_, data_stage_5__1352_, data_stage_5__1351_, data_stage_5__1350_, data_stage_5__1349_, data_stage_5__1348_, data_stage_5__1347_, data_stage_5__1346_, data_stage_5__1345_, data_stage_5__1344_, data_stage_5__1343_, data_stage_5__1342_, data_stage_5__1341_, data_stage_5__1340_, data_stage_5__1339_, data_stage_5__1338_, data_stage_5__1337_, data_stage_5__1336_, data_stage_5__1335_, data_stage_5__1334_, data_stage_5__1333_, data_stage_5__1332_, data_stage_5__1331_, data_stage_5__1330_, data_stage_5__1329_, data_stage_5__1328_, data_stage_5__1327_, data_stage_5__1326_, data_stage_5__1325_, data_stage_5__1324_, data_stage_5__1323_, data_stage_5__1322_, data_stage_5__1321_, data_stage_5__1320_, data_stage_5__1319_, data_stage_5__1318_, data_stage_5__1317_, data_stage_5__1316_, data_stage_5__1315_, data_stage_5__1314_, data_stage_5__1313_, data_stage_5__1312_, data_stage_5__1311_, data_stage_5__1310_, data_stage_5__1309_, data_stage_5__1308_, data_stage_5__1307_, data_stage_5__1306_, data_stage_5__1305_, data_stage_5__1304_, data_stage_5__1303_, data_stage_5__1302_, data_stage_5__1301_, data_stage_5__1300_, data_stage_5__1299_, data_stage_5__1298_, data_stage_5__1297_, data_stage_5__1296_, data_stage_5__1295_, data_stage_5__1294_, data_stage_5__1293_, data_stage_5__1292_, data_stage_5__1291_, data_stage_5__1290_, data_stage_5__1289_, data_stage_5__1288_, data_stage_5__1287_, data_stage_5__1286_, data_stage_5__1285_, data_stage_5__1284_, data_stage_5__1283_, data_stage_5__1282_, data_stage_5__1281_, data_stage_5__1280_, data_stage_5__1279_, data_stage_5__1278_, data_stage_5__1277_, data_stage_5__1276_, data_stage_5__1275_, data_stage_5__1274_, data_stage_5__1273_, data_stage_5__1272_, data_stage_5__1271_, data_stage_5__1270_, data_stage_5__1269_, data_stage_5__1268_, data_stage_5__1267_, data_stage_5__1266_, data_stage_5__1265_, data_stage_5__1264_, data_stage_5__1263_, data_stage_5__1262_, data_stage_5__1261_, data_stage_5__1260_, data_stage_5__1259_, data_stage_5__1258_, data_stage_5__1257_, data_stage_5__1256_, data_stage_5__1255_, data_stage_5__1254_, data_stage_5__1253_, data_stage_5__1252_, data_stage_5__1251_, data_stage_5__1250_, data_stage_5__1249_, data_stage_5__1248_, data_stage_5__1247_, data_stage_5__1246_, data_stage_5__1245_, data_stage_5__1244_, data_stage_5__1243_, data_stage_5__1242_, data_stage_5__1241_, data_stage_5__1240_, data_stage_5__1239_, data_stage_5__1238_, data_stage_5__1237_, data_stage_5__1236_, data_stage_5__1235_, data_stage_5__1234_, data_stage_5__1233_, data_stage_5__1232_, data_stage_5__1231_, data_stage_5__1230_, data_stage_5__1229_, data_stage_5__1228_, data_stage_5__1227_, data_stage_5__1226_, data_stage_5__1225_, data_stage_5__1224_, data_stage_5__1223_, data_stage_5__1222_, data_stage_5__1221_, data_stage_5__1220_, data_stage_5__1219_, data_stage_5__1218_, data_stage_5__1217_, data_stage_5__1216_, data_stage_5__1215_, data_stage_5__1214_, data_stage_5__1213_, data_stage_5__1212_, data_stage_5__1211_, data_stage_5__1210_, data_stage_5__1209_, data_stage_5__1208_, data_stage_5__1207_, data_stage_5__1206_, data_stage_5__1205_, data_stage_5__1204_, data_stage_5__1203_, data_stage_5__1202_, data_stage_5__1201_, data_stage_5__1200_, data_stage_5__1199_, data_stage_5__1198_, data_stage_5__1197_, data_stage_5__1196_, data_stage_5__1195_, data_stage_5__1194_, data_stage_5__1193_, data_stage_5__1192_, data_stage_5__1191_, data_stage_5__1190_, data_stage_5__1189_, data_stage_5__1188_, data_stage_5__1187_, data_stage_5__1186_, data_stage_5__1185_, data_stage_5__1184_, data_stage_5__1183_, data_stage_5__1182_, data_stage_5__1181_, data_stage_5__1180_, data_stage_5__1179_, data_stage_5__1178_, data_stage_5__1177_, data_stage_5__1176_, data_stage_5__1175_, data_stage_5__1174_, data_stage_5__1173_, data_stage_5__1172_, data_stage_5__1171_, data_stage_5__1170_, data_stage_5__1169_, data_stage_5__1168_, data_stage_5__1167_, data_stage_5__1166_, data_stage_5__1165_, data_stage_5__1164_, data_stage_5__1163_, data_stage_5__1162_, data_stage_5__1161_, data_stage_5__1160_, data_stage_5__1159_, data_stage_5__1158_, data_stage_5__1157_, data_stage_5__1156_, data_stage_5__1155_, data_stage_5__1154_, data_stage_5__1153_, data_stage_5__1152_, data_stage_5__1151_, data_stage_5__1150_, data_stage_5__1149_, data_stage_5__1148_, data_stage_5__1147_, data_stage_5__1146_, data_stage_5__1145_, data_stage_5__1144_, data_stage_5__1143_, data_stage_5__1142_, data_stage_5__1141_, data_stage_5__1140_, data_stage_5__1139_, data_stage_5__1138_, data_stage_5__1137_, data_stage_5__1136_, data_stage_5__1135_, data_stage_5__1134_, data_stage_5__1133_, data_stage_5__1132_, data_stage_5__1131_, data_stage_5__1130_, data_stage_5__1129_, data_stage_5__1128_, data_stage_5__1127_, data_stage_5__1126_, data_stage_5__1125_, data_stage_5__1124_, data_stage_5__1123_, data_stage_5__1122_, data_stage_5__1121_, data_stage_5__1120_, data_stage_5__1119_, data_stage_5__1118_, data_stage_5__1117_, data_stage_5__1116_, data_stage_5__1115_, data_stage_5__1114_, data_stage_5__1113_, data_stage_5__1112_, data_stage_5__1111_, data_stage_5__1110_, data_stage_5__1109_, data_stage_5__1108_, data_stage_5__1107_, data_stage_5__1106_, data_stage_5__1105_, data_stage_5__1104_, data_stage_5__1103_, data_stage_5__1102_, data_stage_5__1101_, data_stage_5__1100_, data_stage_5__1099_, data_stage_5__1098_, data_stage_5__1097_, data_stage_5__1096_, data_stage_5__1095_, data_stage_5__1094_, data_stage_5__1093_, data_stage_5__1092_, data_stage_5__1091_, data_stage_5__1090_, data_stage_5__1089_, data_stage_5__1088_, data_stage_5__1087_, data_stage_5__1086_, data_stage_5__1085_, data_stage_5__1084_, data_stage_5__1083_, data_stage_5__1082_, data_stage_5__1081_, data_stage_5__1080_, data_stage_5__1079_, data_stage_5__1078_, data_stage_5__1077_, data_stage_5__1076_, data_stage_5__1075_, data_stage_5__1074_, data_stage_5__1073_, data_stage_5__1072_, data_stage_5__1071_, data_stage_5__1070_, data_stage_5__1069_, data_stage_5__1068_, data_stage_5__1067_, data_stage_5__1066_, data_stage_5__1065_, data_stage_5__1064_, data_stage_5__1063_, data_stage_5__1062_, data_stage_5__1061_, data_stage_5__1060_, data_stage_5__1059_, data_stage_5__1058_, data_stage_5__1057_, data_stage_5__1056_, data_stage_5__1055_, data_stage_5__1054_, data_stage_5__1053_, data_stage_5__1052_, data_stage_5__1051_, data_stage_5__1050_, data_stage_5__1049_, data_stage_5__1048_, data_stage_5__1047_, data_stage_5__1046_, data_stage_5__1045_, data_stage_5__1044_, data_stage_5__1043_, data_stage_5__1042_, data_stage_5__1041_, data_stage_5__1040_, data_stage_5__1039_, data_stage_5__1038_, data_stage_5__1037_, data_stage_5__1036_, data_stage_5__1035_, data_stage_5__1034_, data_stage_5__1033_, data_stage_5__1032_, data_stage_5__1031_, data_stage_5__1030_, data_stage_5__1029_, data_stage_5__1028_, data_stage_5__1027_, data_stage_5__1026_, data_stage_5__1025_, data_stage_5__1024_, data_stage_5__1023_, data_stage_5__1022_, data_stage_5__1021_, data_stage_5__1020_, data_stage_5__1019_, data_stage_5__1018_, data_stage_5__1017_, data_stage_5__1016_, data_stage_5__1015_, data_stage_5__1014_, data_stage_5__1013_, data_stage_5__1012_, data_stage_5__1011_, data_stage_5__1010_, data_stage_5__1009_, data_stage_5__1008_, data_stage_5__1007_, data_stage_5__1006_, data_stage_5__1005_, data_stage_5__1004_, data_stage_5__1003_, data_stage_5__1002_, data_stage_5__1001_, data_stage_5__1000_, data_stage_5__999_, data_stage_5__998_, data_stage_5__997_, data_stage_5__996_, data_stage_5__995_, data_stage_5__994_, data_stage_5__993_, data_stage_5__992_, data_stage_5__991_, data_stage_5__990_, data_stage_5__989_, data_stage_5__988_, data_stage_5__987_, data_stage_5__986_, data_stage_5__985_, data_stage_5__984_, data_stage_5__983_, data_stage_5__982_, data_stage_5__981_, data_stage_5__980_, data_stage_5__979_, data_stage_5__978_, data_stage_5__977_, data_stage_5__976_, data_stage_5__975_, data_stage_5__974_, data_stage_5__973_, data_stage_5__972_, data_stage_5__971_, data_stage_5__970_, data_stage_5__969_, data_stage_5__968_, data_stage_5__967_, data_stage_5__966_, data_stage_5__965_, data_stage_5__964_, data_stage_5__963_, data_stage_5__962_, data_stage_5__961_, data_stage_5__960_, data_stage_5__959_, data_stage_5__958_, data_stage_5__957_, data_stage_5__956_, data_stage_5__955_, data_stage_5__954_, data_stage_5__953_, data_stage_5__952_, data_stage_5__951_, data_stage_5__950_, data_stage_5__949_, data_stage_5__948_, data_stage_5__947_, data_stage_5__946_, data_stage_5__945_, data_stage_5__944_, data_stage_5__943_, data_stage_5__942_, data_stage_5__941_, data_stage_5__940_, data_stage_5__939_, data_stage_5__938_, data_stage_5__937_, data_stage_5__936_, data_stage_5__935_, data_stage_5__934_, data_stage_5__933_, data_stage_5__932_, data_stage_5__931_, data_stage_5__930_, data_stage_5__929_, data_stage_5__928_, data_stage_5__927_, data_stage_5__926_, data_stage_5__925_, data_stage_5__924_, data_stage_5__923_, data_stage_5__922_, data_stage_5__921_, data_stage_5__920_, data_stage_5__919_, data_stage_5__918_, data_stage_5__917_, data_stage_5__916_, data_stage_5__915_, data_stage_5__914_, data_stage_5__913_, data_stage_5__912_, data_stage_5__911_, data_stage_5__910_, data_stage_5__909_, data_stage_5__908_, data_stage_5__907_, data_stage_5__906_, data_stage_5__905_, data_stage_5__904_, data_stage_5__903_, data_stage_5__902_, data_stage_5__901_, data_stage_5__900_, data_stage_5__899_, data_stage_5__898_, data_stage_5__897_, data_stage_5__896_, data_stage_5__895_, data_stage_5__894_, data_stage_5__893_, data_stage_5__892_, data_stage_5__891_, data_stage_5__890_, data_stage_5__889_, data_stage_5__888_, data_stage_5__887_, data_stage_5__886_, data_stage_5__885_, data_stage_5__884_, data_stage_5__883_, data_stage_5__882_, data_stage_5__881_, data_stage_5__880_, data_stage_5__879_, data_stage_5__878_, data_stage_5__877_, data_stage_5__876_, data_stage_5__875_, data_stage_5__874_, data_stage_5__873_, data_stage_5__872_, data_stage_5__871_, data_stage_5__870_, data_stage_5__869_, data_stage_5__868_, data_stage_5__867_, data_stage_5__866_, data_stage_5__865_, data_stage_5__864_, data_stage_5__863_, data_stage_5__862_, data_stage_5__861_, data_stage_5__860_, data_stage_5__859_, data_stage_5__858_, data_stage_5__857_, data_stage_5__856_, data_stage_5__855_, data_stage_5__854_, data_stage_5__853_, data_stage_5__852_, data_stage_5__851_, data_stage_5__850_, data_stage_5__849_, data_stage_5__848_, data_stage_5__847_, data_stage_5__846_, data_stage_5__845_, data_stage_5__844_, data_stage_5__843_, data_stage_5__842_, data_stage_5__841_, data_stage_5__840_, data_stage_5__839_, data_stage_5__838_, data_stage_5__837_, data_stage_5__836_, data_stage_5__835_, data_stage_5__834_, data_stage_5__833_, data_stage_5__832_, data_stage_5__831_, data_stage_5__830_, data_stage_5__829_, data_stage_5__828_, data_stage_5__827_, data_stage_5__826_, data_stage_5__825_, data_stage_5__824_, data_stage_5__823_, data_stage_5__822_, data_stage_5__821_, data_stage_5__820_, data_stage_5__819_, data_stage_5__818_, data_stage_5__817_, data_stage_5__816_, data_stage_5__815_, data_stage_5__814_, data_stage_5__813_, data_stage_5__812_, data_stage_5__811_, data_stage_5__810_, data_stage_5__809_, data_stage_5__808_, data_stage_5__807_, data_stage_5__806_, data_stage_5__805_, data_stage_5__804_, data_stage_5__803_, data_stage_5__802_, data_stage_5__801_, data_stage_5__800_, data_stage_5__799_, data_stage_5__798_, data_stage_5__797_, data_stage_5__796_, data_stage_5__795_, data_stage_5__794_, data_stage_5__793_, data_stage_5__792_, data_stage_5__791_, data_stage_5__790_, data_stage_5__789_, data_stage_5__788_, data_stage_5__787_, data_stage_5__786_, data_stage_5__785_, data_stage_5__784_, data_stage_5__783_, data_stage_5__782_, data_stage_5__781_, data_stage_5__780_, data_stage_5__779_, data_stage_5__778_, data_stage_5__777_, data_stage_5__776_, data_stage_5__775_, data_stage_5__774_, data_stage_5__773_, data_stage_5__772_, data_stage_5__771_, data_stage_5__770_, data_stage_5__769_, data_stage_5__768_, data_stage_5__767_, data_stage_5__766_, data_stage_5__765_, data_stage_5__764_, data_stage_5__763_, data_stage_5__762_, data_stage_5__761_, data_stage_5__760_, data_stage_5__759_, data_stage_5__758_, data_stage_5__757_, data_stage_5__756_, data_stage_5__755_, data_stage_5__754_, data_stage_5__753_, data_stage_5__752_, data_stage_5__751_, data_stage_5__750_, data_stage_5__749_, data_stage_5__748_, data_stage_5__747_, data_stage_5__746_, data_stage_5__745_, data_stage_5__744_, data_stage_5__743_, data_stage_5__742_, data_stage_5__741_, data_stage_5__740_, data_stage_5__739_, data_stage_5__738_, data_stage_5__737_, data_stage_5__736_, data_stage_5__735_, data_stage_5__734_, data_stage_5__733_, data_stage_5__732_, data_stage_5__731_, data_stage_5__730_, data_stage_5__729_, data_stage_5__728_, data_stage_5__727_, data_stage_5__726_, data_stage_5__725_, data_stage_5__724_, data_stage_5__723_, data_stage_5__722_, data_stage_5__721_, data_stage_5__720_, data_stage_5__719_, data_stage_5__718_, data_stage_5__717_, data_stage_5__716_, data_stage_5__715_, data_stage_5__714_, data_stage_5__713_, data_stage_5__712_, data_stage_5__711_, data_stage_5__710_, data_stage_5__709_, data_stage_5__708_, data_stage_5__707_, data_stage_5__706_, data_stage_5__705_, data_stage_5__704_, data_stage_5__703_, data_stage_5__702_, data_stage_5__701_, data_stage_5__700_, data_stage_5__699_, data_stage_5__698_, data_stage_5__697_, data_stage_5__696_, data_stage_5__695_, data_stage_5__694_, data_stage_5__693_, data_stage_5__692_, data_stage_5__691_, data_stage_5__690_, data_stage_5__689_, data_stage_5__688_, data_stage_5__687_, data_stage_5__686_, data_stage_5__685_, data_stage_5__684_, data_stage_5__683_, data_stage_5__682_, data_stage_5__681_, data_stage_5__680_, data_stage_5__679_, data_stage_5__678_, data_stage_5__677_, data_stage_5__676_, data_stage_5__675_, data_stage_5__674_, data_stage_5__673_, data_stage_5__672_, data_stage_5__671_, data_stage_5__670_, data_stage_5__669_, data_stage_5__668_, data_stage_5__667_, data_stage_5__666_, data_stage_5__665_, data_stage_5__664_, data_stage_5__663_, data_stage_5__662_, data_stage_5__661_, data_stage_5__660_, data_stage_5__659_, data_stage_5__658_, data_stage_5__657_, data_stage_5__656_, data_stage_5__655_, data_stage_5__654_, data_stage_5__653_, data_stage_5__652_, data_stage_5__651_, data_stage_5__650_, data_stage_5__649_, data_stage_5__648_, data_stage_5__647_, data_stage_5__646_, data_stage_5__645_, data_stage_5__644_, data_stage_5__643_, data_stage_5__642_, data_stage_5__641_, data_stage_5__640_, data_stage_5__639_, data_stage_5__638_, data_stage_5__637_, data_stage_5__636_, data_stage_5__635_, data_stage_5__634_, data_stage_5__633_, data_stage_5__632_, data_stage_5__631_, data_stage_5__630_, data_stage_5__629_, data_stage_5__628_, data_stage_5__627_, data_stage_5__626_, data_stage_5__625_, data_stage_5__624_, data_stage_5__623_, data_stage_5__622_, data_stage_5__621_, data_stage_5__620_, data_stage_5__619_, data_stage_5__618_, data_stage_5__617_, data_stage_5__616_, data_stage_5__615_, data_stage_5__614_, data_stage_5__613_, data_stage_5__612_, data_stage_5__611_, data_stage_5__610_, data_stage_5__609_, data_stage_5__608_, data_stage_5__607_, data_stage_5__606_, data_stage_5__605_, data_stage_5__604_, data_stage_5__603_, data_stage_5__602_, data_stage_5__601_, data_stage_5__600_, data_stage_5__599_, data_stage_5__598_, data_stage_5__597_, data_stage_5__596_, data_stage_5__595_, data_stage_5__594_, data_stage_5__593_, data_stage_5__592_, data_stage_5__591_, data_stage_5__590_, data_stage_5__589_, data_stage_5__588_, data_stage_5__587_, data_stage_5__586_, data_stage_5__585_, data_stage_5__584_, data_stage_5__583_, data_stage_5__582_, data_stage_5__581_, data_stage_5__580_, data_stage_5__579_, data_stage_5__578_, data_stage_5__577_, data_stage_5__576_, data_stage_5__575_, data_stage_5__574_, data_stage_5__573_, data_stage_5__572_, data_stage_5__571_, data_stage_5__570_, data_stage_5__569_, data_stage_5__568_, data_stage_5__567_, data_stage_5__566_, data_stage_5__565_, data_stage_5__564_, data_stage_5__563_, data_stage_5__562_, data_stage_5__561_, data_stage_5__560_, data_stage_5__559_, data_stage_5__558_, data_stage_5__557_, data_stage_5__556_, data_stage_5__555_, data_stage_5__554_, data_stage_5__553_, data_stage_5__552_, data_stage_5__551_, data_stage_5__550_, data_stage_5__549_, data_stage_5__548_, data_stage_5__547_, data_stage_5__546_, data_stage_5__545_, data_stage_5__544_, data_stage_5__543_, data_stage_5__542_, data_stage_5__541_, data_stage_5__540_, data_stage_5__539_, data_stage_5__538_, data_stage_5__537_, data_stage_5__536_, data_stage_5__535_, data_stage_5__534_, data_stage_5__533_, data_stage_5__532_, data_stage_5__531_, data_stage_5__530_, data_stage_5__529_, data_stage_5__528_, data_stage_5__527_, data_stage_5__526_, data_stage_5__525_, data_stage_5__524_, data_stage_5__523_, data_stage_5__522_, data_stage_5__521_, data_stage_5__520_, data_stage_5__519_, data_stage_5__518_, data_stage_5__517_, data_stage_5__516_, data_stage_5__515_, data_stage_5__514_, data_stage_5__513_, data_stage_5__512_, data_stage_5__511_, data_stage_5__510_, data_stage_5__509_, data_stage_5__508_, data_stage_5__507_, data_stage_5__506_, data_stage_5__505_, data_stage_5__504_, data_stage_5__503_, data_stage_5__502_, data_stage_5__501_, data_stage_5__500_, data_stage_5__499_, data_stage_5__498_, data_stage_5__497_, data_stage_5__496_, data_stage_5__495_, data_stage_5__494_, data_stage_5__493_, data_stage_5__492_, data_stage_5__491_, data_stage_5__490_, data_stage_5__489_, data_stage_5__488_, data_stage_5__487_, data_stage_5__486_, data_stage_5__485_, data_stage_5__484_, data_stage_5__483_, data_stage_5__482_, data_stage_5__481_, data_stage_5__480_, data_stage_5__479_, data_stage_5__478_, data_stage_5__477_, data_stage_5__476_, data_stage_5__475_, data_stage_5__474_, data_stage_5__473_, data_stage_5__472_, data_stage_5__471_, data_stage_5__470_, data_stage_5__469_, data_stage_5__468_, data_stage_5__467_, data_stage_5__466_, data_stage_5__465_, data_stage_5__464_, data_stage_5__463_, data_stage_5__462_, data_stage_5__461_, data_stage_5__460_, data_stage_5__459_, data_stage_5__458_, data_stage_5__457_, data_stage_5__456_, data_stage_5__455_, data_stage_5__454_, data_stage_5__453_, data_stage_5__452_, data_stage_5__451_, data_stage_5__450_, data_stage_5__449_, data_stage_5__448_, data_stage_5__447_, data_stage_5__446_, data_stage_5__445_, data_stage_5__444_, data_stage_5__443_, data_stage_5__442_, data_stage_5__441_, data_stage_5__440_, data_stage_5__439_, data_stage_5__438_, data_stage_5__437_, data_stage_5__436_, data_stage_5__435_, data_stage_5__434_, data_stage_5__433_, data_stage_5__432_, data_stage_5__431_, data_stage_5__430_, data_stage_5__429_, data_stage_5__428_, data_stage_5__427_, data_stage_5__426_, data_stage_5__425_, data_stage_5__424_, data_stage_5__423_, data_stage_5__422_, data_stage_5__421_, data_stage_5__420_, data_stage_5__419_, data_stage_5__418_, data_stage_5__417_, data_stage_5__416_, data_stage_5__415_, data_stage_5__414_, data_stage_5__413_, data_stage_5__412_, data_stage_5__411_, data_stage_5__410_, data_stage_5__409_, data_stage_5__408_, data_stage_5__407_, data_stage_5__406_, data_stage_5__405_, data_stage_5__404_, data_stage_5__403_, data_stage_5__402_, data_stage_5__401_, data_stage_5__400_, data_stage_5__399_, data_stage_5__398_, data_stage_5__397_, data_stage_5__396_, data_stage_5__395_, data_stage_5__394_, data_stage_5__393_, data_stage_5__392_, data_stage_5__391_, data_stage_5__390_, data_stage_5__389_, data_stage_5__388_, data_stage_5__387_, data_stage_5__386_, data_stage_5__385_, data_stage_5__384_, data_stage_5__383_, data_stage_5__382_, data_stage_5__381_, data_stage_5__380_, data_stage_5__379_, data_stage_5__378_, data_stage_5__377_, data_stage_5__376_, data_stage_5__375_, data_stage_5__374_, data_stage_5__373_, data_stage_5__372_, data_stage_5__371_, data_stage_5__370_, data_stage_5__369_, data_stage_5__368_, data_stage_5__367_, data_stage_5__366_, data_stage_5__365_, data_stage_5__364_, data_stage_5__363_, data_stage_5__362_, data_stage_5__361_, data_stage_5__360_, data_stage_5__359_, data_stage_5__358_, data_stage_5__357_, data_stage_5__356_, data_stage_5__355_, data_stage_5__354_, data_stage_5__353_, data_stage_5__352_, data_stage_5__351_, data_stage_5__350_, data_stage_5__349_, data_stage_5__348_, data_stage_5__347_, data_stage_5__346_, data_stage_5__345_, data_stage_5__344_, data_stage_5__343_, data_stage_5__342_, data_stage_5__341_, data_stage_5__340_, data_stage_5__339_, data_stage_5__338_, data_stage_5__337_, data_stage_5__336_, data_stage_5__335_, data_stage_5__334_, data_stage_5__333_, data_stage_5__332_, data_stage_5__331_, data_stage_5__330_, data_stage_5__329_, data_stage_5__328_, data_stage_5__327_, data_stage_5__326_, data_stage_5__325_, data_stage_5__324_, data_stage_5__323_, data_stage_5__322_, data_stage_5__321_, data_stage_5__320_, data_stage_5__319_, data_stage_5__318_, data_stage_5__317_, data_stage_5__316_, data_stage_5__315_, data_stage_5__314_, data_stage_5__313_, data_stage_5__312_, data_stage_5__311_, data_stage_5__310_, data_stage_5__309_, data_stage_5__308_, data_stage_5__307_, data_stage_5__306_, data_stage_5__305_, data_stage_5__304_, data_stage_5__303_, data_stage_5__302_, data_stage_5__301_, data_stage_5__300_, data_stage_5__299_, data_stage_5__298_, data_stage_5__297_, data_stage_5__296_, data_stage_5__295_, data_stage_5__294_, data_stage_5__293_, data_stage_5__292_, data_stage_5__291_, data_stage_5__290_, data_stage_5__289_, data_stage_5__288_, data_stage_5__287_, data_stage_5__286_, data_stage_5__285_, data_stage_5__284_, data_stage_5__283_, data_stage_5__282_, data_stage_5__281_, data_stage_5__280_, data_stage_5__279_, data_stage_5__278_, data_stage_5__277_, data_stage_5__276_, data_stage_5__275_, data_stage_5__274_, data_stage_5__273_, data_stage_5__272_, data_stage_5__271_, data_stage_5__270_, data_stage_5__269_, data_stage_5__268_, data_stage_5__267_, data_stage_5__266_, data_stage_5__265_, data_stage_5__264_, data_stage_5__263_, data_stage_5__262_, data_stage_5__261_, data_stage_5__260_, data_stage_5__259_, data_stage_5__258_, data_stage_5__257_, data_stage_5__256_, data_stage_5__255_, data_stage_5__254_, data_stage_5__253_, data_stage_5__252_, data_stage_5__251_, data_stage_5__250_, data_stage_5__249_, data_stage_5__248_, data_stage_5__247_, data_stage_5__246_, data_stage_5__245_, data_stage_5__244_, data_stage_5__243_, data_stage_5__242_, data_stage_5__241_, data_stage_5__240_, data_stage_5__239_, data_stage_5__238_, data_stage_5__237_, data_stage_5__236_, data_stage_5__235_, data_stage_5__234_, data_stage_5__233_, data_stage_5__232_, data_stage_5__231_, data_stage_5__230_, data_stage_5__229_, data_stage_5__228_, data_stage_5__227_, data_stage_5__226_, data_stage_5__225_, data_stage_5__224_, data_stage_5__223_, data_stage_5__222_, data_stage_5__221_, data_stage_5__220_, data_stage_5__219_, data_stage_5__218_, data_stage_5__217_, data_stage_5__216_, data_stage_5__215_, data_stage_5__214_, data_stage_5__213_, data_stage_5__212_, data_stage_5__211_, data_stage_5__210_, data_stage_5__209_, data_stage_5__208_, data_stage_5__207_, data_stage_5__206_, data_stage_5__205_, data_stage_5__204_, data_stage_5__203_, data_stage_5__202_, data_stage_5__201_, data_stage_5__200_, data_stage_5__199_, data_stage_5__198_, data_stage_5__197_, data_stage_5__196_, data_stage_5__195_, data_stage_5__194_, data_stage_5__193_, data_stage_5__192_, data_stage_5__191_, data_stage_5__190_, data_stage_5__189_, data_stage_5__188_, data_stage_5__187_, data_stage_5__186_, data_stage_5__185_, data_stage_5__184_, data_stage_5__183_, data_stage_5__182_, data_stage_5__181_, data_stage_5__180_, data_stage_5__179_, data_stage_5__178_, data_stage_5__177_, data_stage_5__176_, data_stage_5__175_, data_stage_5__174_, data_stage_5__173_, data_stage_5__172_, data_stage_5__171_, data_stage_5__170_, data_stage_5__169_, data_stage_5__168_, data_stage_5__167_, data_stage_5__166_, data_stage_5__165_, data_stage_5__164_, data_stage_5__163_, data_stage_5__162_, data_stage_5__161_, data_stage_5__160_, data_stage_5__159_, data_stage_5__158_, data_stage_5__157_, data_stage_5__156_, data_stage_5__155_, data_stage_5__154_, data_stage_5__153_, data_stage_5__152_, data_stage_5__151_, data_stage_5__150_, data_stage_5__149_, data_stage_5__148_, data_stage_5__147_, data_stage_5__146_, data_stage_5__145_, data_stage_5__144_, data_stage_5__143_, data_stage_5__142_, data_stage_5__141_, data_stage_5__140_, data_stage_5__139_, data_stage_5__138_, data_stage_5__137_, data_stage_5__136_, data_stage_5__135_, data_stage_5__134_, data_stage_5__133_, data_stage_5__132_, data_stage_5__131_, data_stage_5__130_, data_stage_5__129_, data_stage_5__128_, data_stage_5__127_, data_stage_5__126_, data_stage_5__125_, data_stage_5__124_, data_stage_5__123_, data_stage_5__122_, data_stage_5__121_, data_stage_5__120_, data_stage_5__119_, data_stage_5__118_, data_stage_5__117_, data_stage_5__116_, data_stage_5__115_, data_stage_5__114_, data_stage_5__113_, data_stage_5__112_, data_stage_5__111_, data_stage_5__110_, data_stage_5__109_, data_stage_5__108_, data_stage_5__107_, data_stage_5__106_, data_stage_5__105_, data_stage_5__104_, data_stage_5__103_, data_stage_5__102_, data_stage_5__101_, data_stage_5__100_, data_stage_5__99_, data_stage_5__98_, data_stage_5__97_, data_stage_5__96_, data_stage_5__95_, data_stage_5__94_, data_stage_5__93_, data_stage_5__92_, data_stage_5__91_, data_stage_5__90_, data_stage_5__89_, data_stage_5__88_, data_stage_5__87_, data_stage_5__86_, data_stage_5__85_, data_stage_5__84_, data_stage_5__83_, data_stage_5__82_, data_stage_5__81_, data_stage_5__80_, data_stage_5__79_, data_stage_5__78_, data_stage_5__77_, data_stage_5__76_, data_stage_5__75_, data_stage_5__74_, data_stage_5__73_, data_stage_5__72_, data_stage_5__71_, data_stage_5__70_, data_stage_5__69_, data_stage_5__68_, data_stage_5__67_, data_stage_5__66_, data_stage_5__65_, data_stage_5__64_, data_stage_5__63_, data_stage_5__62_, data_stage_5__61_, data_stage_5__60_, data_stage_5__59_, data_stage_5__58_, data_stage_5__57_, data_stage_5__56_, data_stage_5__55_, data_stage_5__54_, data_stage_5__53_, data_stage_5__52_, data_stage_5__51_, data_stage_5__50_, data_stage_5__49_, data_stage_5__48_, data_stage_5__47_, data_stage_5__46_, data_stage_5__45_, data_stage_5__44_, data_stage_5__43_, data_stage_5__42_, data_stage_5__41_, data_stage_5__40_, data_stage_5__39_, data_stage_5__38_, data_stage_5__37_, data_stage_5__36_, data_stage_5__35_, data_stage_5__34_, data_stage_5__33_, data_stage_5__32_, data_stage_5__31_, data_stage_5__30_, data_stage_5__29_, data_stage_5__28_, data_stage_5__27_, data_stage_5__26_, data_stage_5__25_, data_stage_5__24_, data_stage_5__23_, data_stage_5__22_, data_stage_5__21_, data_stage_5__20_, data_stage_5__19_, data_stage_5__18_, data_stage_5__17_, data_stage_5__16_, data_stage_5__15_, data_stage_5__14_, data_stage_5__13_, data_stage_5__12_, data_stage_5__11_, data_stage_5__10_, data_stage_5__9_, data_stage_5__8_, data_stage_5__7_, data_stage_5__6_, data_stage_5__5_, data_stage_5__4_, data_stage_5__3_, data_stage_5__2_, data_stage_5__1_, data_stage_5__0_ })
  );


  bsg_swap_width_p1024
  mux_stage_4__mux_swap_1__swap_inst
  (
    .data_i({ data_stage_4__4095_, data_stage_4__4094_, data_stage_4__4093_, data_stage_4__4092_, data_stage_4__4091_, data_stage_4__4090_, data_stage_4__4089_, data_stage_4__4088_, data_stage_4__4087_, data_stage_4__4086_, data_stage_4__4085_, data_stage_4__4084_, data_stage_4__4083_, data_stage_4__4082_, data_stage_4__4081_, data_stage_4__4080_, data_stage_4__4079_, data_stage_4__4078_, data_stage_4__4077_, data_stage_4__4076_, data_stage_4__4075_, data_stage_4__4074_, data_stage_4__4073_, data_stage_4__4072_, data_stage_4__4071_, data_stage_4__4070_, data_stage_4__4069_, data_stage_4__4068_, data_stage_4__4067_, data_stage_4__4066_, data_stage_4__4065_, data_stage_4__4064_, data_stage_4__4063_, data_stage_4__4062_, data_stage_4__4061_, data_stage_4__4060_, data_stage_4__4059_, data_stage_4__4058_, data_stage_4__4057_, data_stage_4__4056_, data_stage_4__4055_, data_stage_4__4054_, data_stage_4__4053_, data_stage_4__4052_, data_stage_4__4051_, data_stage_4__4050_, data_stage_4__4049_, data_stage_4__4048_, data_stage_4__4047_, data_stage_4__4046_, data_stage_4__4045_, data_stage_4__4044_, data_stage_4__4043_, data_stage_4__4042_, data_stage_4__4041_, data_stage_4__4040_, data_stage_4__4039_, data_stage_4__4038_, data_stage_4__4037_, data_stage_4__4036_, data_stage_4__4035_, data_stage_4__4034_, data_stage_4__4033_, data_stage_4__4032_, data_stage_4__4031_, data_stage_4__4030_, data_stage_4__4029_, data_stage_4__4028_, data_stage_4__4027_, data_stage_4__4026_, data_stage_4__4025_, data_stage_4__4024_, data_stage_4__4023_, data_stage_4__4022_, data_stage_4__4021_, data_stage_4__4020_, data_stage_4__4019_, data_stage_4__4018_, data_stage_4__4017_, data_stage_4__4016_, data_stage_4__4015_, data_stage_4__4014_, data_stage_4__4013_, data_stage_4__4012_, data_stage_4__4011_, data_stage_4__4010_, data_stage_4__4009_, data_stage_4__4008_, data_stage_4__4007_, data_stage_4__4006_, data_stage_4__4005_, data_stage_4__4004_, data_stage_4__4003_, data_stage_4__4002_, data_stage_4__4001_, data_stage_4__4000_, data_stage_4__3999_, data_stage_4__3998_, data_stage_4__3997_, data_stage_4__3996_, data_stage_4__3995_, data_stage_4__3994_, data_stage_4__3993_, data_stage_4__3992_, data_stage_4__3991_, data_stage_4__3990_, data_stage_4__3989_, data_stage_4__3988_, data_stage_4__3987_, data_stage_4__3986_, data_stage_4__3985_, data_stage_4__3984_, data_stage_4__3983_, data_stage_4__3982_, data_stage_4__3981_, data_stage_4__3980_, data_stage_4__3979_, data_stage_4__3978_, data_stage_4__3977_, data_stage_4__3976_, data_stage_4__3975_, data_stage_4__3974_, data_stage_4__3973_, data_stage_4__3972_, data_stage_4__3971_, data_stage_4__3970_, data_stage_4__3969_, data_stage_4__3968_, data_stage_4__3967_, data_stage_4__3966_, data_stage_4__3965_, data_stage_4__3964_, data_stage_4__3963_, data_stage_4__3962_, data_stage_4__3961_, data_stage_4__3960_, data_stage_4__3959_, data_stage_4__3958_, data_stage_4__3957_, data_stage_4__3956_, data_stage_4__3955_, data_stage_4__3954_, data_stage_4__3953_, data_stage_4__3952_, data_stage_4__3951_, data_stage_4__3950_, data_stage_4__3949_, data_stage_4__3948_, data_stage_4__3947_, data_stage_4__3946_, data_stage_4__3945_, data_stage_4__3944_, data_stage_4__3943_, data_stage_4__3942_, data_stage_4__3941_, data_stage_4__3940_, data_stage_4__3939_, data_stage_4__3938_, data_stage_4__3937_, data_stage_4__3936_, data_stage_4__3935_, data_stage_4__3934_, data_stage_4__3933_, data_stage_4__3932_, data_stage_4__3931_, data_stage_4__3930_, data_stage_4__3929_, data_stage_4__3928_, data_stage_4__3927_, data_stage_4__3926_, data_stage_4__3925_, data_stage_4__3924_, data_stage_4__3923_, data_stage_4__3922_, data_stage_4__3921_, data_stage_4__3920_, data_stage_4__3919_, data_stage_4__3918_, data_stage_4__3917_, data_stage_4__3916_, data_stage_4__3915_, data_stage_4__3914_, data_stage_4__3913_, data_stage_4__3912_, data_stage_4__3911_, data_stage_4__3910_, data_stage_4__3909_, data_stage_4__3908_, data_stage_4__3907_, data_stage_4__3906_, data_stage_4__3905_, data_stage_4__3904_, data_stage_4__3903_, data_stage_4__3902_, data_stage_4__3901_, data_stage_4__3900_, data_stage_4__3899_, data_stage_4__3898_, data_stage_4__3897_, data_stage_4__3896_, data_stage_4__3895_, data_stage_4__3894_, data_stage_4__3893_, data_stage_4__3892_, data_stage_4__3891_, data_stage_4__3890_, data_stage_4__3889_, data_stage_4__3888_, data_stage_4__3887_, data_stage_4__3886_, data_stage_4__3885_, data_stage_4__3884_, data_stage_4__3883_, data_stage_4__3882_, data_stage_4__3881_, data_stage_4__3880_, data_stage_4__3879_, data_stage_4__3878_, data_stage_4__3877_, data_stage_4__3876_, data_stage_4__3875_, data_stage_4__3874_, data_stage_4__3873_, data_stage_4__3872_, data_stage_4__3871_, data_stage_4__3870_, data_stage_4__3869_, data_stage_4__3868_, data_stage_4__3867_, data_stage_4__3866_, data_stage_4__3865_, data_stage_4__3864_, data_stage_4__3863_, data_stage_4__3862_, data_stage_4__3861_, data_stage_4__3860_, data_stage_4__3859_, data_stage_4__3858_, data_stage_4__3857_, data_stage_4__3856_, data_stage_4__3855_, data_stage_4__3854_, data_stage_4__3853_, data_stage_4__3852_, data_stage_4__3851_, data_stage_4__3850_, data_stage_4__3849_, data_stage_4__3848_, data_stage_4__3847_, data_stage_4__3846_, data_stage_4__3845_, data_stage_4__3844_, data_stage_4__3843_, data_stage_4__3842_, data_stage_4__3841_, data_stage_4__3840_, data_stage_4__3839_, data_stage_4__3838_, data_stage_4__3837_, data_stage_4__3836_, data_stage_4__3835_, data_stage_4__3834_, data_stage_4__3833_, data_stage_4__3832_, data_stage_4__3831_, data_stage_4__3830_, data_stage_4__3829_, data_stage_4__3828_, data_stage_4__3827_, data_stage_4__3826_, data_stage_4__3825_, data_stage_4__3824_, data_stage_4__3823_, data_stage_4__3822_, data_stage_4__3821_, data_stage_4__3820_, data_stage_4__3819_, data_stage_4__3818_, data_stage_4__3817_, data_stage_4__3816_, data_stage_4__3815_, data_stage_4__3814_, data_stage_4__3813_, data_stage_4__3812_, data_stage_4__3811_, data_stage_4__3810_, data_stage_4__3809_, data_stage_4__3808_, data_stage_4__3807_, data_stage_4__3806_, data_stage_4__3805_, data_stage_4__3804_, data_stage_4__3803_, data_stage_4__3802_, data_stage_4__3801_, data_stage_4__3800_, data_stage_4__3799_, data_stage_4__3798_, data_stage_4__3797_, data_stage_4__3796_, data_stage_4__3795_, data_stage_4__3794_, data_stage_4__3793_, data_stage_4__3792_, data_stage_4__3791_, data_stage_4__3790_, data_stage_4__3789_, data_stage_4__3788_, data_stage_4__3787_, data_stage_4__3786_, data_stage_4__3785_, data_stage_4__3784_, data_stage_4__3783_, data_stage_4__3782_, data_stage_4__3781_, data_stage_4__3780_, data_stage_4__3779_, data_stage_4__3778_, data_stage_4__3777_, data_stage_4__3776_, data_stage_4__3775_, data_stage_4__3774_, data_stage_4__3773_, data_stage_4__3772_, data_stage_4__3771_, data_stage_4__3770_, data_stage_4__3769_, data_stage_4__3768_, data_stage_4__3767_, data_stage_4__3766_, data_stage_4__3765_, data_stage_4__3764_, data_stage_4__3763_, data_stage_4__3762_, data_stage_4__3761_, data_stage_4__3760_, data_stage_4__3759_, data_stage_4__3758_, data_stage_4__3757_, data_stage_4__3756_, data_stage_4__3755_, data_stage_4__3754_, data_stage_4__3753_, data_stage_4__3752_, data_stage_4__3751_, data_stage_4__3750_, data_stage_4__3749_, data_stage_4__3748_, data_stage_4__3747_, data_stage_4__3746_, data_stage_4__3745_, data_stage_4__3744_, data_stage_4__3743_, data_stage_4__3742_, data_stage_4__3741_, data_stage_4__3740_, data_stage_4__3739_, data_stage_4__3738_, data_stage_4__3737_, data_stage_4__3736_, data_stage_4__3735_, data_stage_4__3734_, data_stage_4__3733_, data_stage_4__3732_, data_stage_4__3731_, data_stage_4__3730_, data_stage_4__3729_, data_stage_4__3728_, data_stage_4__3727_, data_stage_4__3726_, data_stage_4__3725_, data_stage_4__3724_, data_stage_4__3723_, data_stage_4__3722_, data_stage_4__3721_, data_stage_4__3720_, data_stage_4__3719_, data_stage_4__3718_, data_stage_4__3717_, data_stage_4__3716_, data_stage_4__3715_, data_stage_4__3714_, data_stage_4__3713_, data_stage_4__3712_, data_stage_4__3711_, data_stage_4__3710_, data_stage_4__3709_, data_stage_4__3708_, data_stage_4__3707_, data_stage_4__3706_, data_stage_4__3705_, data_stage_4__3704_, data_stage_4__3703_, data_stage_4__3702_, data_stage_4__3701_, data_stage_4__3700_, data_stage_4__3699_, data_stage_4__3698_, data_stage_4__3697_, data_stage_4__3696_, data_stage_4__3695_, data_stage_4__3694_, data_stage_4__3693_, data_stage_4__3692_, data_stage_4__3691_, data_stage_4__3690_, data_stage_4__3689_, data_stage_4__3688_, data_stage_4__3687_, data_stage_4__3686_, data_stage_4__3685_, data_stage_4__3684_, data_stage_4__3683_, data_stage_4__3682_, data_stage_4__3681_, data_stage_4__3680_, data_stage_4__3679_, data_stage_4__3678_, data_stage_4__3677_, data_stage_4__3676_, data_stage_4__3675_, data_stage_4__3674_, data_stage_4__3673_, data_stage_4__3672_, data_stage_4__3671_, data_stage_4__3670_, data_stage_4__3669_, data_stage_4__3668_, data_stage_4__3667_, data_stage_4__3666_, data_stage_4__3665_, data_stage_4__3664_, data_stage_4__3663_, data_stage_4__3662_, data_stage_4__3661_, data_stage_4__3660_, data_stage_4__3659_, data_stage_4__3658_, data_stage_4__3657_, data_stage_4__3656_, data_stage_4__3655_, data_stage_4__3654_, data_stage_4__3653_, data_stage_4__3652_, data_stage_4__3651_, data_stage_4__3650_, data_stage_4__3649_, data_stage_4__3648_, data_stage_4__3647_, data_stage_4__3646_, data_stage_4__3645_, data_stage_4__3644_, data_stage_4__3643_, data_stage_4__3642_, data_stage_4__3641_, data_stage_4__3640_, data_stage_4__3639_, data_stage_4__3638_, data_stage_4__3637_, data_stage_4__3636_, data_stage_4__3635_, data_stage_4__3634_, data_stage_4__3633_, data_stage_4__3632_, data_stage_4__3631_, data_stage_4__3630_, data_stage_4__3629_, data_stage_4__3628_, data_stage_4__3627_, data_stage_4__3626_, data_stage_4__3625_, data_stage_4__3624_, data_stage_4__3623_, data_stage_4__3622_, data_stage_4__3621_, data_stage_4__3620_, data_stage_4__3619_, data_stage_4__3618_, data_stage_4__3617_, data_stage_4__3616_, data_stage_4__3615_, data_stage_4__3614_, data_stage_4__3613_, data_stage_4__3612_, data_stage_4__3611_, data_stage_4__3610_, data_stage_4__3609_, data_stage_4__3608_, data_stage_4__3607_, data_stage_4__3606_, data_stage_4__3605_, data_stage_4__3604_, data_stage_4__3603_, data_stage_4__3602_, data_stage_4__3601_, data_stage_4__3600_, data_stage_4__3599_, data_stage_4__3598_, data_stage_4__3597_, data_stage_4__3596_, data_stage_4__3595_, data_stage_4__3594_, data_stage_4__3593_, data_stage_4__3592_, data_stage_4__3591_, data_stage_4__3590_, data_stage_4__3589_, data_stage_4__3588_, data_stage_4__3587_, data_stage_4__3586_, data_stage_4__3585_, data_stage_4__3584_, data_stage_4__3583_, data_stage_4__3582_, data_stage_4__3581_, data_stage_4__3580_, data_stage_4__3579_, data_stage_4__3578_, data_stage_4__3577_, data_stage_4__3576_, data_stage_4__3575_, data_stage_4__3574_, data_stage_4__3573_, data_stage_4__3572_, data_stage_4__3571_, data_stage_4__3570_, data_stage_4__3569_, data_stage_4__3568_, data_stage_4__3567_, data_stage_4__3566_, data_stage_4__3565_, data_stage_4__3564_, data_stage_4__3563_, data_stage_4__3562_, data_stage_4__3561_, data_stage_4__3560_, data_stage_4__3559_, data_stage_4__3558_, data_stage_4__3557_, data_stage_4__3556_, data_stage_4__3555_, data_stage_4__3554_, data_stage_4__3553_, data_stage_4__3552_, data_stage_4__3551_, data_stage_4__3550_, data_stage_4__3549_, data_stage_4__3548_, data_stage_4__3547_, data_stage_4__3546_, data_stage_4__3545_, data_stage_4__3544_, data_stage_4__3543_, data_stage_4__3542_, data_stage_4__3541_, data_stage_4__3540_, data_stage_4__3539_, data_stage_4__3538_, data_stage_4__3537_, data_stage_4__3536_, data_stage_4__3535_, data_stage_4__3534_, data_stage_4__3533_, data_stage_4__3532_, data_stage_4__3531_, data_stage_4__3530_, data_stage_4__3529_, data_stage_4__3528_, data_stage_4__3527_, data_stage_4__3526_, data_stage_4__3525_, data_stage_4__3524_, data_stage_4__3523_, data_stage_4__3522_, data_stage_4__3521_, data_stage_4__3520_, data_stage_4__3519_, data_stage_4__3518_, data_stage_4__3517_, data_stage_4__3516_, data_stage_4__3515_, data_stage_4__3514_, data_stage_4__3513_, data_stage_4__3512_, data_stage_4__3511_, data_stage_4__3510_, data_stage_4__3509_, data_stage_4__3508_, data_stage_4__3507_, data_stage_4__3506_, data_stage_4__3505_, data_stage_4__3504_, data_stage_4__3503_, data_stage_4__3502_, data_stage_4__3501_, data_stage_4__3500_, data_stage_4__3499_, data_stage_4__3498_, data_stage_4__3497_, data_stage_4__3496_, data_stage_4__3495_, data_stage_4__3494_, data_stage_4__3493_, data_stage_4__3492_, data_stage_4__3491_, data_stage_4__3490_, data_stage_4__3489_, data_stage_4__3488_, data_stage_4__3487_, data_stage_4__3486_, data_stage_4__3485_, data_stage_4__3484_, data_stage_4__3483_, data_stage_4__3482_, data_stage_4__3481_, data_stage_4__3480_, data_stage_4__3479_, data_stage_4__3478_, data_stage_4__3477_, data_stage_4__3476_, data_stage_4__3475_, data_stage_4__3474_, data_stage_4__3473_, data_stage_4__3472_, data_stage_4__3471_, data_stage_4__3470_, data_stage_4__3469_, data_stage_4__3468_, data_stage_4__3467_, data_stage_4__3466_, data_stage_4__3465_, data_stage_4__3464_, data_stage_4__3463_, data_stage_4__3462_, data_stage_4__3461_, data_stage_4__3460_, data_stage_4__3459_, data_stage_4__3458_, data_stage_4__3457_, data_stage_4__3456_, data_stage_4__3455_, data_stage_4__3454_, data_stage_4__3453_, data_stage_4__3452_, data_stage_4__3451_, data_stage_4__3450_, data_stage_4__3449_, data_stage_4__3448_, data_stage_4__3447_, data_stage_4__3446_, data_stage_4__3445_, data_stage_4__3444_, data_stage_4__3443_, data_stage_4__3442_, data_stage_4__3441_, data_stage_4__3440_, data_stage_4__3439_, data_stage_4__3438_, data_stage_4__3437_, data_stage_4__3436_, data_stage_4__3435_, data_stage_4__3434_, data_stage_4__3433_, data_stage_4__3432_, data_stage_4__3431_, data_stage_4__3430_, data_stage_4__3429_, data_stage_4__3428_, data_stage_4__3427_, data_stage_4__3426_, data_stage_4__3425_, data_stage_4__3424_, data_stage_4__3423_, data_stage_4__3422_, data_stage_4__3421_, data_stage_4__3420_, data_stage_4__3419_, data_stage_4__3418_, data_stage_4__3417_, data_stage_4__3416_, data_stage_4__3415_, data_stage_4__3414_, data_stage_4__3413_, data_stage_4__3412_, data_stage_4__3411_, data_stage_4__3410_, data_stage_4__3409_, data_stage_4__3408_, data_stage_4__3407_, data_stage_4__3406_, data_stage_4__3405_, data_stage_4__3404_, data_stage_4__3403_, data_stage_4__3402_, data_stage_4__3401_, data_stage_4__3400_, data_stage_4__3399_, data_stage_4__3398_, data_stage_4__3397_, data_stage_4__3396_, data_stage_4__3395_, data_stage_4__3394_, data_stage_4__3393_, data_stage_4__3392_, data_stage_4__3391_, data_stage_4__3390_, data_stage_4__3389_, data_stage_4__3388_, data_stage_4__3387_, data_stage_4__3386_, data_stage_4__3385_, data_stage_4__3384_, data_stage_4__3383_, data_stage_4__3382_, data_stage_4__3381_, data_stage_4__3380_, data_stage_4__3379_, data_stage_4__3378_, data_stage_4__3377_, data_stage_4__3376_, data_stage_4__3375_, data_stage_4__3374_, data_stage_4__3373_, data_stage_4__3372_, data_stage_4__3371_, data_stage_4__3370_, data_stage_4__3369_, data_stage_4__3368_, data_stage_4__3367_, data_stage_4__3366_, data_stage_4__3365_, data_stage_4__3364_, data_stage_4__3363_, data_stage_4__3362_, data_stage_4__3361_, data_stage_4__3360_, data_stage_4__3359_, data_stage_4__3358_, data_stage_4__3357_, data_stage_4__3356_, data_stage_4__3355_, data_stage_4__3354_, data_stage_4__3353_, data_stage_4__3352_, data_stage_4__3351_, data_stage_4__3350_, data_stage_4__3349_, data_stage_4__3348_, data_stage_4__3347_, data_stage_4__3346_, data_stage_4__3345_, data_stage_4__3344_, data_stage_4__3343_, data_stage_4__3342_, data_stage_4__3341_, data_stage_4__3340_, data_stage_4__3339_, data_stage_4__3338_, data_stage_4__3337_, data_stage_4__3336_, data_stage_4__3335_, data_stage_4__3334_, data_stage_4__3333_, data_stage_4__3332_, data_stage_4__3331_, data_stage_4__3330_, data_stage_4__3329_, data_stage_4__3328_, data_stage_4__3327_, data_stage_4__3326_, data_stage_4__3325_, data_stage_4__3324_, data_stage_4__3323_, data_stage_4__3322_, data_stage_4__3321_, data_stage_4__3320_, data_stage_4__3319_, data_stage_4__3318_, data_stage_4__3317_, data_stage_4__3316_, data_stage_4__3315_, data_stage_4__3314_, data_stage_4__3313_, data_stage_4__3312_, data_stage_4__3311_, data_stage_4__3310_, data_stage_4__3309_, data_stage_4__3308_, data_stage_4__3307_, data_stage_4__3306_, data_stage_4__3305_, data_stage_4__3304_, data_stage_4__3303_, data_stage_4__3302_, data_stage_4__3301_, data_stage_4__3300_, data_stage_4__3299_, data_stage_4__3298_, data_stage_4__3297_, data_stage_4__3296_, data_stage_4__3295_, data_stage_4__3294_, data_stage_4__3293_, data_stage_4__3292_, data_stage_4__3291_, data_stage_4__3290_, data_stage_4__3289_, data_stage_4__3288_, data_stage_4__3287_, data_stage_4__3286_, data_stage_4__3285_, data_stage_4__3284_, data_stage_4__3283_, data_stage_4__3282_, data_stage_4__3281_, data_stage_4__3280_, data_stage_4__3279_, data_stage_4__3278_, data_stage_4__3277_, data_stage_4__3276_, data_stage_4__3275_, data_stage_4__3274_, data_stage_4__3273_, data_stage_4__3272_, data_stage_4__3271_, data_stage_4__3270_, data_stage_4__3269_, data_stage_4__3268_, data_stage_4__3267_, data_stage_4__3266_, data_stage_4__3265_, data_stage_4__3264_, data_stage_4__3263_, data_stage_4__3262_, data_stage_4__3261_, data_stage_4__3260_, data_stage_4__3259_, data_stage_4__3258_, data_stage_4__3257_, data_stage_4__3256_, data_stage_4__3255_, data_stage_4__3254_, data_stage_4__3253_, data_stage_4__3252_, data_stage_4__3251_, data_stage_4__3250_, data_stage_4__3249_, data_stage_4__3248_, data_stage_4__3247_, data_stage_4__3246_, data_stage_4__3245_, data_stage_4__3244_, data_stage_4__3243_, data_stage_4__3242_, data_stage_4__3241_, data_stage_4__3240_, data_stage_4__3239_, data_stage_4__3238_, data_stage_4__3237_, data_stage_4__3236_, data_stage_4__3235_, data_stage_4__3234_, data_stage_4__3233_, data_stage_4__3232_, data_stage_4__3231_, data_stage_4__3230_, data_stage_4__3229_, data_stage_4__3228_, data_stage_4__3227_, data_stage_4__3226_, data_stage_4__3225_, data_stage_4__3224_, data_stage_4__3223_, data_stage_4__3222_, data_stage_4__3221_, data_stage_4__3220_, data_stage_4__3219_, data_stage_4__3218_, data_stage_4__3217_, data_stage_4__3216_, data_stage_4__3215_, data_stage_4__3214_, data_stage_4__3213_, data_stage_4__3212_, data_stage_4__3211_, data_stage_4__3210_, data_stage_4__3209_, data_stage_4__3208_, data_stage_4__3207_, data_stage_4__3206_, data_stage_4__3205_, data_stage_4__3204_, data_stage_4__3203_, data_stage_4__3202_, data_stage_4__3201_, data_stage_4__3200_, data_stage_4__3199_, data_stage_4__3198_, data_stage_4__3197_, data_stage_4__3196_, data_stage_4__3195_, data_stage_4__3194_, data_stage_4__3193_, data_stage_4__3192_, data_stage_4__3191_, data_stage_4__3190_, data_stage_4__3189_, data_stage_4__3188_, data_stage_4__3187_, data_stage_4__3186_, data_stage_4__3185_, data_stage_4__3184_, data_stage_4__3183_, data_stage_4__3182_, data_stage_4__3181_, data_stage_4__3180_, data_stage_4__3179_, data_stage_4__3178_, data_stage_4__3177_, data_stage_4__3176_, data_stage_4__3175_, data_stage_4__3174_, data_stage_4__3173_, data_stage_4__3172_, data_stage_4__3171_, data_stage_4__3170_, data_stage_4__3169_, data_stage_4__3168_, data_stage_4__3167_, data_stage_4__3166_, data_stage_4__3165_, data_stage_4__3164_, data_stage_4__3163_, data_stage_4__3162_, data_stage_4__3161_, data_stage_4__3160_, data_stage_4__3159_, data_stage_4__3158_, data_stage_4__3157_, data_stage_4__3156_, data_stage_4__3155_, data_stage_4__3154_, data_stage_4__3153_, data_stage_4__3152_, data_stage_4__3151_, data_stage_4__3150_, data_stage_4__3149_, data_stage_4__3148_, data_stage_4__3147_, data_stage_4__3146_, data_stage_4__3145_, data_stage_4__3144_, data_stage_4__3143_, data_stage_4__3142_, data_stage_4__3141_, data_stage_4__3140_, data_stage_4__3139_, data_stage_4__3138_, data_stage_4__3137_, data_stage_4__3136_, data_stage_4__3135_, data_stage_4__3134_, data_stage_4__3133_, data_stage_4__3132_, data_stage_4__3131_, data_stage_4__3130_, data_stage_4__3129_, data_stage_4__3128_, data_stage_4__3127_, data_stage_4__3126_, data_stage_4__3125_, data_stage_4__3124_, data_stage_4__3123_, data_stage_4__3122_, data_stage_4__3121_, data_stage_4__3120_, data_stage_4__3119_, data_stage_4__3118_, data_stage_4__3117_, data_stage_4__3116_, data_stage_4__3115_, data_stage_4__3114_, data_stage_4__3113_, data_stage_4__3112_, data_stage_4__3111_, data_stage_4__3110_, data_stage_4__3109_, data_stage_4__3108_, data_stage_4__3107_, data_stage_4__3106_, data_stage_4__3105_, data_stage_4__3104_, data_stage_4__3103_, data_stage_4__3102_, data_stage_4__3101_, data_stage_4__3100_, data_stage_4__3099_, data_stage_4__3098_, data_stage_4__3097_, data_stage_4__3096_, data_stage_4__3095_, data_stage_4__3094_, data_stage_4__3093_, data_stage_4__3092_, data_stage_4__3091_, data_stage_4__3090_, data_stage_4__3089_, data_stage_4__3088_, data_stage_4__3087_, data_stage_4__3086_, data_stage_4__3085_, data_stage_4__3084_, data_stage_4__3083_, data_stage_4__3082_, data_stage_4__3081_, data_stage_4__3080_, data_stage_4__3079_, data_stage_4__3078_, data_stage_4__3077_, data_stage_4__3076_, data_stage_4__3075_, data_stage_4__3074_, data_stage_4__3073_, data_stage_4__3072_, data_stage_4__3071_, data_stage_4__3070_, data_stage_4__3069_, data_stage_4__3068_, data_stage_4__3067_, data_stage_4__3066_, data_stage_4__3065_, data_stage_4__3064_, data_stage_4__3063_, data_stage_4__3062_, data_stage_4__3061_, data_stage_4__3060_, data_stage_4__3059_, data_stage_4__3058_, data_stage_4__3057_, data_stage_4__3056_, data_stage_4__3055_, data_stage_4__3054_, data_stage_4__3053_, data_stage_4__3052_, data_stage_4__3051_, data_stage_4__3050_, data_stage_4__3049_, data_stage_4__3048_, data_stage_4__3047_, data_stage_4__3046_, data_stage_4__3045_, data_stage_4__3044_, data_stage_4__3043_, data_stage_4__3042_, data_stage_4__3041_, data_stage_4__3040_, data_stage_4__3039_, data_stage_4__3038_, data_stage_4__3037_, data_stage_4__3036_, data_stage_4__3035_, data_stage_4__3034_, data_stage_4__3033_, data_stage_4__3032_, data_stage_4__3031_, data_stage_4__3030_, data_stage_4__3029_, data_stage_4__3028_, data_stage_4__3027_, data_stage_4__3026_, data_stage_4__3025_, data_stage_4__3024_, data_stage_4__3023_, data_stage_4__3022_, data_stage_4__3021_, data_stage_4__3020_, data_stage_4__3019_, data_stage_4__3018_, data_stage_4__3017_, data_stage_4__3016_, data_stage_4__3015_, data_stage_4__3014_, data_stage_4__3013_, data_stage_4__3012_, data_stage_4__3011_, data_stage_4__3010_, data_stage_4__3009_, data_stage_4__3008_, data_stage_4__3007_, data_stage_4__3006_, data_stage_4__3005_, data_stage_4__3004_, data_stage_4__3003_, data_stage_4__3002_, data_stage_4__3001_, data_stage_4__3000_, data_stage_4__2999_, data_stage_4__2998_, data_stage_4__2997_, data_stage_4__2996_, data_stage_4__2995_, data_stage_4__2994_, data_stage_4__2993_, data_stage_4__2992_, data_stage_4__2991_, data_stage_4__2990_, data_stage_4__2989_, data_stage_4__2988_, data_stage_4__2987_, data_stage_4__2986_, data_stage_4__2985_, data_stage_4__2984_, data_stage_4__2983_, data_stage_4__2982_, data_stage_4__2981_, data_stage_4__2980_, data_stage_4__2979_, data_stage_4__2978_, data_stage_4__2977_, data_stage_4__2976_, data_stage_4__2975_, data_stage_4__2974_, data_stage_4__2973_, data_stage_4__2972_, data_stage_4__2971_, data_stage_4__2970_, data_stage_4__2969_, data_stage_4__2968_, data_stage_4__2967_, data_stage_4__2966_, data_stage_4__2965_, data_stage_4__2964_, data_stage_4__2963_, data_stage_4__2962_, data_stage_4__2961_, data_stage_4__2960_, data_stage_4__2959_, data_stage_4__2958_, data_stage_4__2957_, data_stage_4__2956_, data_stage_4__2955_, data_stage_4__2954_, data_stage_4__2953_, data_stage_4__2952_, data_stage_4__2951_, data_stage_4__2950_, data_stage_4__2949_, data_stage_4__2948_, data_stage_4__2947_, data_stage_4__2946_, data_stage_4__2945_, data_stage_4__2944_, data_stage_4__2943_, data_stage_4__2942_, data_stage_4__2941_, data_stage_4__2940_, data_stage_4__2939_, data_stage_4__2938_, data_stage_4__2937_, data_stage_4__2936_, data_stage_4__2935_, data_stage_4__2934_, data_stage_4__2933_, data_stage_4__2932_, data_stage_4__2931_, data_stage_4__2930_, data_stage_4__2929_, data_stage_4__2928_, data_stage_4__2927_, data_stage_4__2926_, data_stage_4__2925_, data_stage_4__2924_, data_stage_4__2923_, data_stage_4__2922_, data_stage_4__2921_, data_stage_4__2920_, data_stage_4__2919_, data_stage_4__2918_, data_stage_4__2917_, data_stage_4__2916_, data_stage_4__2915_, data_stage_4__2914_, data_stage_4__2913_, data_stage_4__2912_, data_stage_4__2911_, data_stage_4__2910_, data_stage_4__2909_, data_stage_4__2908_, data_stage_4__2907_, data_stage_4__2906_, data_stage_4__2905_, data_stage_4__2904_, data_stage_4__2903_, data_stage_4__2902_, data_stage_4__2901_, data_stage_4__2900_, data_stage_4__2899_, data_stage_4__2898_, data_stage_4__2897_, data_stage_4__2896_, data_stage_4__2895_, data_stage_4__2894_, data_stage_4__2893_, data_stage_4__2892_, data_stage_4__2891_, data_stage_4__2890_, data_stage_4__2889_, data_stage_4__2888_, data_stage_4__2887_, data_stage_4__2886_, data_stage_4__2885_, data_stage_4__2884_, data_stage_4__2883_, data_stage_4__2882_, data_stage_4__2881_, data_stage_4__2880_, data_stage_4__2879_, data_stage_4__2878_, data_stage_4__2877_, data_stage_4__2876_, data_stage_4__2875_, data_stage_4__2874_, data_stage_4__2873_, data_stage_4__2872_, data_stage_4__2871_, data_stage_4__2870_, data_stage_4__2869_, data_stage_4__2868_, data_stage_4__2867_, data_stage_4__2866_, data_stage_4__2865_, data_stage_4__2864_, data_stage_4__2863_, data_stage_4__2862_, data_stage_4__2861_, data_stage_4__2860_, data_stage_4__2859_, data_stage_4__2858_, data_stage_4__2857_, data_stage_4__2856_, data_stage_4__2855_, data_stage_4__2854_, data_stage_4__2853_, data_stage_4__2852_, data_stage_4__2851_, data_stage_4__2850_, data_stage_4__2849_, data_stage_4__2848_, data_stage_4__2847_, data_stage_4__2846_, data_stage_4__2845_, data_stage_4__2844_, data_stage_4__2843_, data_stage_4__2842_, data_stage_4__2841_, data_stage_4__2840_, data_stage_4__2839_, data_stage_4__2838_, data_stage_4__2837_, data_stage_4__2836_, data_stage_4__2835_, data_stage_4__2834_, data_stage_4__2833_, data_stage_4__2832_, data_stage_4__2831_, data_stage_4__2830_, data_stage_4__2829_, data_stage_4__2828_, data_stage_4__2827_, data_stage_4__2826_, data_stage_4__2825_, data_stage_4__2824_, data_stage_4__2823_, data_stage_4__2822_, data_stage_4__2821_, data_stage_4__2820_, data_stage_4__2819_, data_stage_4__2818_, data_stage_4__2817_, data_stage_4__2816_, data_stage_4__2815_, data_stage_4__2814_, data_stage_4__2813_, data_stage_4__2812_, data_stage_4__2811_, data_stage_4__2810_, data_stage_4__2809_, data_stage_4__2808_, data_stage_4__2807_, data_stage_4__2806_, data_stage_4__2805_, data_stage_4__2804_, data_stage_4__2803_, data_stage_4__2802_, data_stage_4__2801_, data_stage_4__2800_, data_stage_4__2799_, data_stage_4__2798_, data_stage_4__2797_, data_stage_4__2796_, data_stage_4__2795_, data_stage_4__2794_, data_stage_4__2793_, data_stage_4__2792_, data_stage_4__2791_, data_stage_4__2790_, data_stage_4__2789_, data_stage_4__2788_, data_stage_4__2787_, data_stage_4__2786_, data_stage_4__2785_, data_stage_4__2784_, data_stage_4__2783_, data_stage_4__2782_, data_stage_4__2781_, data_stage_4__2780_, data_stage_4__2779_, data_stage_4__2778_, data_stage_4__2777_, data_stage_4__2776_, data_stage_4__2775_, data_stage_4__2774_, data_stage_4__2773_, data_stage_4__2772_, data_stage_4__2771_, data_stage_4__2770_, data_stage_4__2769_, data_stage_4__2768_, data_stage_4__2767_, data_stage_4__2766_, data_stage_4__2765_, data_stage_4__2764_, data_stage_4__2763_, data_stage_4__2762_, data_stage_4__2761_, data_stage_4__2760_, data_stage_4__2759_, data_stage_4__2758_, data_stage_4__2757_, data_stage_4__2756_, data_stage_4__2755_, data_stage_4__2754_, data_stage_4__2753_, data_stage_4__2752_, data_stage_4__2751_, data_stage_4__2750_, data_stage_4__2749_, data_stage_4__2748_, data_stage_4__2747_, data_stage_4__2746_, data_stage_4__2745_, data_stage_4__2744_, data_stage_4__2743_, data_stage_4__2742_, data_stage_4__2741_, data_stage_4__2740_, data_stage_4__2739_, data_stage_4__2738_, data_stage_4__2737_, data_stage_4__2736_, data_stage_4__2735_, data_stage_4__2734_, data_stage_4__2733_, data_stage_4__2732_, data_stage_4__2731_, data_stage_4__2730_, data_stage_4__2729_, data_stage_4__2728_, data_stage_4__2727_, data_stage_4__2726_, data_stage_4__2725_, data_stage_4__2724_, data_stage_4__2723_, data_stage_4__2722_, data_stage_4__2721_, data_stage_4__2720_, data_stage_4__2719_, data_stage_4__2718_, data_stage_4__2717_, data_stage_4__2716_, data_stage_4__2715_, data_stage_4__2714_, data_stage_4__2713_, data_stage_4__2712_, data_stage_4__2711_, data_stage_4__2710_, data_stage_4__2709_, data_stage_4__2708_, data_stage_4__2707_, data_stage_4__2706_, data_stage_4__2705_, data_stage_4__2704_, data_stage_4__2703_, data_stage_4__2702_, data_stage_4__2701_, data_stage_4__2700_, data_stage_4__2699_, data_stage_4__2698_, data_stage_4__2697_, data_stage_4__2696_, data_stage_4__2695_, data_stage_4__2694_, data_stage_4__2693_, data_stage_4__2692_, data_stage_4__2691_, data_stage_4__2690_, data_stage_4__2689_, data_stage_4__2688_, data_stage_4__2687_, data_stage_4__2686_, data_stage_4__2685_, data_stage_4__2684_, data_stage_4__2683_, data_stage_4__2682_, data_stage_4__2681_, data_stage_4__2680_, data_stage_4__2679_, data_stage_4__2678_, data_stage_4__2677_, data_stage_4__2676_, data_stage_4__2675_, data_stage_4__2674_, data_stage_4__2673_, data_stage_4__2672_, data_stage_4__2671_, data_stage_4__2670_, data_stage_4__2669_, data_stage_4__2668_, data_stage_4__2667_, data_stage_4__2666_, data_stage_4__2665_, data_stage_4__2664_, data_stage_4__2663_, data_stage_4__2662_, data_stage_4__2661_, data_stage_4__2660_, data_stage_4__2659_, data_stage_4__2658_, data_stage_4__2657_, data_stage_4__2656_, data_stage_4__2655_, data_stage_4__2654_, data_stage_4__2653_, data_stage_4__2652_, data_stage_4__2651_, data_stage_4__2650_, data_stage_4__2649_, data_stage_4__2648_, data_stage_4__2647_, data_stage_4__2646_, data_stage_4__2645_, data_stage_4__2644_, data_stage_4__2643_, data_stage_4__2642_, data_stage_4__2641_, data_stage_4__2640_, data_stage_4__2639_, data_stage_4__2638_, data_stage_4__2637_, data_stage_4__2636_, data_stage_4__2635_, data_stage_4__2634_, data_stage_4__2633_, data_stage_4__2632_, data_stage_4__2631_, data_stage_4__2630_, data_stage_4__2629_, data_stage_4__2628_, data_stage_4__2627_, data_stage_4__2626_, data_stage_4__2625_, data_stage_4__2624_, data_stage_4__2623_, data_stage_4__2622_, data_stage_4__2621_, data_stage_4__2620_, data_stage_4__2619_, data_stage_4__2618_, data_stage_4__2617_, data_stage_4__2616_, data_stage_4__2615_, data_stage_4__2614_, data_stage_4__2613_, data_stage_4__2612_, data_stage_4__2611_, data_stage_4__2610_, data_stage_4__2609_, data_stage_4__2608_, data_stage_4__2607_, data_stage_4__2606_, data_stage_4__2605_, data_stage_4__2604_, data_stage_4__2603_, data_stage_4__2602_, data_stage_4__2601_, data_stage_4__2600_, data_stage_4__2599_, data_stage_4__2598_, data_stage_4__2597_, data_stage_4__2596_, data_stage_4__2595_, data_stage_4__2594_, data_stage_4__2593_, data_stage_4__2592_, data_stage_4__2591_, data_stage_4__2590_, data_stage_4__2589_, data_stage_4__2588_, data_stage_4__2587_, data_stage_4__2586_, data_stage_4__2585_, data_stage_4__2584_, data_stage_4__2583_, data_stage_4__2582_, data_stage_4__2581_, data_stage_4__2580_, data_stage_4__2579_, data_stage_4__2578_, data_stage_4__2577_, data_stage_4__2576_, data_stage_4__2575_, data_stage_4__2574_, data_stage_4__2573_, data_stage_4__2572_, data_stage_4__2571_, data_stage_4__2570_, data_stage_4__2569_, data_stage_4__2568_, data_stage_4__2567_, data_stage_4__2566_, data_stage_4__2565_, data_stage_4__2564_, data_stage_4__2563_, data_stage_4__2562_, data_stage_4__2561_, data_stage_4__2560_, data_stage_4__2559_, data_stage_4__2558_, data_stage_4__2557_, data_stage_4__2556_, data_stage_4__2555_, data_stage_4__2554_, data_stage_4__2553_, data_stage_4__2552_, data_stage_4__2551_, data_stage_4__2550_, data_stage_4__2549_, data_stage_4__2548_, data_stage_4__2547_, data_stage_4__2546_, data_stage_4__2545_, data_stage_4__2544_, data_stage_4__2543_, data_stage_4__2542_, data_stage_4__2541_, data_stage_4__2540_, data_stage_4__2539_, data_stage_4__2538_, data_stage_4__2537_, data_stage_4__2536_, data_stage_4__2535_, data_stage_4__2534_, data_stage_4__2533_, data_stage_4__2532_, data_stage_4__2531_, data_stage_4__2530_, data_stage_4__2529_, data_stage_4__2528_, data_stage_4__2527_, data_stage_4__2526_, data_stage_4__2525_, data_stage_4__2524_, data_stage_4__2523_, data_stage_4__2522_, data_stage_4__2521_, data_stage_4__2520_, data_stage_4__2519_, data_stage_4__2518_, data_stage_4__2517_, data_stage_4__2516_, data_stage_4__2515_, data_stage_4__2514_, data_stage_4__2513_, data_stage_4__2512_, data_stage_4__2511_, data_stage_4__2510_, data_stage_4__2509_, data_stage_4__2508_, data_stage_4__2507_, data_stage_4__2506_, data_stage_4__2505_, data_stage_4__2504_, data_stage_4__2503_, data_stage_4__2502_, data_stage_4__2501_, data_stage_4__2500_, data_stage_4__2499_, data_stage_4__2498_, data_stage_4__2497_, data_stage_4__2496_, data_stage_4__2495_, data_stage_4__2494_, data_stage_4__2493_, data_stage_4__2492_, data_stage_4__2491_, data_stage_4__2490_, data_stage_4__2489_, data_stage_4__2488_, data_stage_4__2487_, data_stage_4__2486_, data_stage_4__2485_, data_stage_4__2484_, data_stage_4__2483_, data_stage_4__2482_, data_stage_4__2481_, data_stage_4__2480_, data_stage_4__2479_, data_stage_4__2478_, data_stage_4__2477_, data_stage_4__2476_, data_stage_4__2475_, data_stage_4__2474_, data_stage_4__2473_, data_stage_4__2472_, data_stage_4__2471_, data_stage_4__2470_, data_stage_4__2469_, data_stage_4__2468_, data_stage_4__2467_, data_stage_4__2466_, data_stage_4__2465_, data_stage_4__2464_, data_stage_4__2463_, data_stage_4__2462_, data_stage_4__2461_, data_stage_4__2460_, data_stage_4__2459_, data_stage_4__2458_, data_stage_4__2457_, data_stage_4__2456_, data_stage_4__2455_, data_stage_4__2454_, data_stage_4__2453_, data_stage_4__2452_, data_stage_4__2451_, data_stage_4__2450_, data_stage_4__2449_, data_stage_4__2448_, data_stage_4__2447_, data_stage_4__2446_, data_stage_4__2445_, data_stage_4__2444_, data_stage_4__2443_, data_stage_4__2442_, data_stage_4__2441_, data_stage_4__2440_, data_stage_4__2439_, data_stage_4__2438_, data_stage_4__2437_, data_stage_4__2436_, data_stage_4__2435_, data_stage_4__2434_, data_stage_4__2433_, data_stage_4__2432_, data_stage_4__2431_, data_stage_4__2430_, data_stage_4__2429_, data_stage_4__2428_, data_stage_4__2427_, data_stage_4__2426_, data_stage_4__2425_, data_stage_4__2424_, data_stage_4__2423_, data_stage_4__2422_, data_stage_4__2421_, data_stage_4__2420_, data_stage_4__2419_, data_stage_4__2418_, data_stage_4__2417_, data_stage_4__2416_, data_stage_4__2415_, data_stage_4__2414_, data_stage_4__2413_, data_stage_4__2412_, data_stage_4__2411_, data_stage_4__2410_, data_stage_4__2409_, data_stage_4__2408_, data_stage_4__2407_, data_stage_4__2406_, data_stage_4__2405_, data_stage_4__2404_, data_stage_4__2403_, data_stage_4__2402_, data_stage_4__2401_, data_stage_4__2400_, data_stage_4__2399_, data_stage_4__2398_, data_stage_4__2397_, data_stage_4__2396_, data_stage_4__2395_, data_stage_4__2394_, data_stage_4__2393_, data_stage_4__2392_, data_stage_4__2391_, data_stage_4__2390_, data_stage_4__2389_, data_stage_4__2388_, data_stage_4__2387_, data_stage_4__2386_, data_stage_4__2385_, data_stage_4__2384_, data_stage_4__2383_, data_stage_4__2382_, data_stage_4__2381_, data_stage_4__2380_, data_stage_4__2379_, data_stage_4__2378_, data_stage_4__2377_, data_stage_4__2376_, data_stage_4__2375_, data_stage_4__2374_, data_stage_4__2373_, data_stage_4__2372_, data_stage_4__2371_, data_stage_4__2370_, data_stage_4__2369_, data_stage_4__2368_, data_stage_4__2367_, data_stage_4__2366_, data_stage_4__2365_, data_stage_4__2364_, data_stage_4__2363_, data_stage_4__2362_, data_stage_4__2361_, data_stage_4__2360_, data_stage_4__2359_, data_stage_4__2358_, data_stage_4__2357_, data_stage_4__2356_, data_stage_4__2355_, data_stage_4__2354_, data_stage_4__2353_, data_stage_4__2352_, data_stage_4__2351_, data_stage_4__2350_, data_stage_4__2349_, data_stage_4__2348_, data_stage_4__2347_, data_stage_4__2346_, data_stage_4__2345_, data_stage_4__2344_, data_stage_4__2343_, data_stage_4__2342_, data_stage_4__2341_, data_stage_4__2340_, data_stage_4__2339_, data_stage_4__2338_, data_stage_4__2337_, data_stage_4__2336_, data_stage_4__2335_, data_stage_4__2334_, data_stage_4__2333_, data_stage_4__2332_, data_stage_4__2331_, data_stage_4__2330_, data_stage_4__2329_, data_stage_4__2328_, data_stage_4__2327_, data_stage_4__2326_, data_stage_4__2325_, data_stage_4__2324_, data_stage_4__2323_, data_stage_4__2322_, data_stage_4__2321_, data_stage_4__2320_, data_stage_4__2319_, data_stage_4__2318_, data_stage_4__2317_, data_stage_4__2316_, data_stage_4__2315_, data_stage_4__2314_, data_stage_4__2313_, data_stage_4__2312_, data_stage_4__2311_, data_stage_4__2310_, data_stage_4__2309_, data_stage_4__2308_, data_stage_4__2307_, data_stage_4__2306_, data_stage_4__2305_, data_stage_4__2304_, data_stage_4__2303_, data_stage_4__2302_, data_stage_4__2301_, data_stage_4__2300_, data_stage_4__2299_, data_stage_4__2298_, data_stage_4__2297_, data_stage_4__2296_, data_stage_4__2295_, data_stage_4__2294_, data_stage_4__2293_, data_stage_4__2292_, data_stage_4__2291_, data_stage_4__2290_, data_stage_4__2289_, data_stage_4__2288_, data_stage_4__2287_, data_stage_4__2286_, data_stage_4__2285_, data_stage_4__2284_, data_stage_4__2283_, data_stage_4__2282_, data_stage_4__2281_, data_stage_4__2280_, data_stage_4__2279_, data_stage_4__2278_, data_stage_4__2277_, data_stage_4__2276_, data_stage_4__2275_, data_stage_4__2274_, data_stage_4__2273_, data_stage_4__2272_, data_stage_4__2271_, data_stage_4__2270_, data_stage_4__2269_, data_stage_4__2268_, data_stage_4__2267_, data_stage_4__2266_, data_stage_4__2265_, data_stage_4__2264_, data_stage_4__2263_, data_stage_4__2262_, data_stage_4__2261_, data_stage_4__2260_, data_stage_4__2259_, data_stage_4__2258_, data_stage_4__2257_, data_stage_4__2256_, data_stage_4__2255_, data_stage_4__2254_, data_stage_4__2253_, data_stage_4__2252_, data_stage_4__2251_, data_stage_4__2250_, data_stage_4__2249_, data_stage_4__2248_, data_stage_4__2247_, data_stage_4__2246_, data_stage_4__2245_, data_stage_4__2244_, data_stage_4__2243_, data_stage_4__2242_, data_stage_4__2241_, data_stage_4__2240_, data_stage_4__2239_, data_stage_4__2238_, data_stage_4__2237_, data_stage_4__2236_, data_stage_4__2235_, data_stage_4__2234_, data_stage_4__2233_, data_stage_4__2232_, data_stage_4__2231_, data_stage_4__2230_, data_stage_4__2229_, data_stage_4__2228_, data_stage_4__2227_, data_stage_4__2226_, data_stage_4__2225_, data_stage_4__2224_, data_stage_4__2223_, data_stage_4__2222_, data_stage_4__2221_, data_stage_4__2220_, data_stage_4__2219_, data_stage_4__2218_, data_stage_4__2217_, data_stage_4__2216_, data_stage_4__2215_, data_stage_4__2214_, data_stage_4__2213_, data_stage_4__2212_, data_stage_4__2211_, data_stage_4__2210_, data_stage_4__2209_, data_stage_4__2208_, data_stage_4__2207_, data_stage_4__2206_, data_stage_4__2205_, data_stage_4__2204_, data_stage_4__2203_, data_stage_4__2202_, data_stage_4__2201_, data_stage_4__2200_, data_stage_4__2199_, data_stage_4__2198_, data_stage_4__2197_, data_stage_4__2196_, data_stage_4__2195_, data_stage_4__2194_, data_stage_4__2193_, data_stage_4__2192_, data_stage_4__2191_, data_stage_4__2190_, data_stage_4__2189_, data_stage_4__2188_, data_stage_4__2187_, data_stage_4__2186_, data_stage_4__2185_, data_stage_4__2184_, data_stage_4__2183_, data_stage_4__2182_, data_stage_4__2181_, data_stage_4__2180_, data_stage_4__2179_, data_stage_4__2178_, data_stage_4__2177_, data_stage_4__2176_, data_stage_4__2175_, data_stage_4__2174_, data_stage_4__2173_, data_stage_4__2172_, data_stage_4__2171_, data_stage_4__2170_, data_stage_4__2169_, data_stage_4__2168_, data_stage_4__2167_, data_stage_4__2166_, data_stage_4__2165_, data_stage_4__2164_, data_stage_4__2163_, data_stage_4__2162_, data_stage_4__2161_, data_stage_4__2160_, data_stage_4__2159_, data_stage_4__2158_, data_stage_4__2157_, data_stage_4__2156_, data_stage_4__2155_, data_stage_4__2154_, data_stage_4__2153_, data_stage_4__2152_, data_stage_4__2151_, data_stage_4__2150_, data_stage_4__2149_, data_stage_4__2148_, data_stage_4__2147_, data_stage_4__2146_, data_stage_4__2145_, data_stage_4__2144_, data_stage_4__2143_, data_stage_4__2142_, data_stage_4__2141_, data_stage_4__2140_, data_stage_4__2139_, data_stage_4__2138_, data_stage_4__2137_, data_stage_4__2136_, data_stage_4__2135_, data_stage_4__2134_, data_stage_4__2133_, data_stage_4__2132_, data_stage_4__2131_, data_stage_4__2130_, data_stage_4__2129_, data_stage_4__2128_, data_stage_4__2127_, data_stage_4__2126_, data_stage_4__2125_, data_stage_4__2124_, data_stage_4__2123_, data_stage_4__2122_, data_stage_4__2121_, data_stage_4__2120_, data_stage_4__2119_, data_stage_4__2118_, data_stage_4__2117_, data_stage_4__2116_, data_stage_4__2115_, data_stage_4__2114_, data_stage_4__2113_, data_stage_4__2112_, data_stage_4__2111_, data_stage_4__2110_, data_stage_4__2109_, data_stage_4__2108_, data_stage_4__2107_, data_stage_4__2106_, data_stage_4__2105_, data_stage_4__2104_, data_stage_4__2103_, data_stage_4__2102_, data_stage_4__2101_, data_stage_4__2100_, data_stage_4__2099_, data_stage_4__2098_, data_stage_4__2097_, data_stage_4__2096_, data_stage_4__2095_, data_stage_4__2094_, data_stage_4__2093_, data_stage_4__2092_, data_stage_4__2091_, data_stage_4__2090_, data_stage_4__2089_, data_stage_4__2088_, data_stage_4__2087_, data_stage_4__2086_, data_stage_4__2085_, data_stage_4__2084_, data_stage_4__2083_, data_stage_4__2082_, data_stage_4__2081_, data_stage_4__2080_, data_stage_4__2079_, data_stage_4__2078_, data_stage_4__2077_, data_stage_4__2076_, data_stage_4__2075_, data_stage_4__2074_, data_stage_4__2073_, data_stage_4__2072_, data_stage_4__2071_, data_stage_4__2070_, data_stage_4__2069_, data_stage_4__2068_, data_stage_4__2067_, data_stage_4__2066_, data_stage_4__2065_, data_stage_4__2064_, data_stage_4__2063_, data_stage_4__2062_, data_stage_4__2061_, data_stage_4__2060_, data_stage_4__2059_, data_stage_4__2058_, data_stage_4__2057_, data_stage_4__2056_, data_stage_4__2055_, data_stage_4__2054_, data_stage_4__2053_, data_stage_4__2052_, data_stage_4__2051_, data_stage_4__2050_, data_stage_4__2049_, data_stage_4__2048_ }),
    .swap_i(sel_i[4]),
    .data_o({ data_stage_5__4095_, data_stage_5__4094_, data_stage_5__4093_, data_stage_5__4092_, data_stage_5__4091_, data_stage_5__4090_, data_stage_5__4089_, data_stage_5__4088_, data_stage_5__4087_, data_stage_5__4086_, data_stage_5__4085_, data_stage_5__4084_, data_stage_5__4083_, data_stage_5__4082_, data_stage_5__4081_, data_stage_5__4080_, data_stage_5__4079_, data_stage_5__4078_, data_stage_5__4077_, data_stage_5__4076_, data_stage_5__4075_, data_stage_5__4074_, data_stage_5__4073_, data_stage_5__4072_, data_stage_5__4071_, data_stage_5__4070_, data_stage_5__4069_, data_stage_5__4068_, data_stage_5__4067_, data_stage_5__4066_, data_stage_5__4065_, data_stage_5__4064_, data_stage_5__4063_, data_stage_5__4062_, data_stage_5__4061_, data_stage_5__4060_, data_stage_5__4059_, data_stage_5__4058_, data_stage_5__4057_, data_stage_5__4056_, data_stage_5__4055_, data_stage_5__4054_, data_stage_5__4053_, data_stage_5__4052_, data_stage_5__4051_, data_stage_5__4050_, data_stage_5__4049_, data_stage_5__4048_, data_stage_5__4047_, data_stage_5__4046_, data_stage_5__4045_, data_stage_5__4044_, data_stage_5__4043_, data_stage_5__4042_, data_stage_5__4041_, data_stage_5__4040_, data_stage_5__4039_, data_stage_5__4038_, data_stage_5__4037_, data_stage_5__4036_, data_stage_5__4035_, data_stage_5__4034_, data_stage_5__4033_, data_stage_5__4032_, data_stage_5__4031_, data_stage_5__4030_, data_stage_5__4029_, data_stage_5__4028_, data_stage_5__4027_, data_stage_5__4026_, data_stage_5__4025_, data_stage_5__4024_, data_stage_5__4023_, data_stage_5__4022_, data_stage_5__4021_, data_stage_5__4020_, data_stage_5__4019_, data_stage_5__4018_, data_stage_5__4017_, data_stage_5__4016_, data_stage_5__4015_, data_stage_5__4014_, data_stage_5__4013_, data_stage_5__4012_, data_stage_5__4011_, data_stage_5__4010_, data_stage_5__4009_, data_stage_5__4008_, data_stage_5__4007_, data_stage_5__4006_, data_stage_5__4005_, data_stage_5__4004_, data_stage_5__4003_, data_stage_5__4002_, data_stage_5__4001_, data_stage_5__4000_, data_stage_5__3999_, data_stage_5__3998_, data_stage_5__3997_, data_stage_5__3996_, data_stage_5__3995_, data_stage_5__3994_, data_stage_5__3993_, data_stage_5__3992_, data_stage_5__3991_, data_stage_5__3990_, data_stage_5__3989_, data_stage_5__3988_, data_stage_5__3987_, data_stage_5__3986_, data_stage_5__3985_, data_stage_5__3984_, data_stage_5__3983_, data_stage_5__3982_, data_stage_5__3981_, data_stage_5__3980_, data_stage_5__3979_, data_stage_5__3978_, data_stage_5__3977_, data_stage_5__3976_, data_stage_5__3975_, data_stage_5__3974_, data_stage_5__3973_, data_stage_5__3972_, data_stage_5__3971_, data_stage_5__3970_, data_stage_5__3969_, data_stage_5__3968_, data_stage_5__3967_, data_stage_5__3966_, data_stage_5__3965_, data_stage_5__3964_, data_stage_5__3963_, data_stage_5__3962_, data_stage_5__3961_, data_stage_5__3960_, data_stage_5__3959_, data_stage_5__3958_, data_stage_5__3957_, data_stage_5__3956_, data_stage_5__3955_, data_stage_5__3954_, data_stage_5__3953_, data_stage_5__3952_, data_stage_5__3951_, data_stage_5__3950_, data_stage_5__3949_, data_stage_5__3948_, data_stage_5__3947_, data_stage_5__3946_, data_stage_5__3945_, data_stage_5__3944_, data_stage_5__3943_, data_stage_5__3942_, data_stage_5__3941_, data_stage_5__3940_, data_stage_5__3939_, data_stage_5__3938_, data_stage_5__3937_, data_stage_5__3936_, data_stage_5__3935_, data_stage_5__3934_, data_stage_5__3933_, data_stage_5__3932_, data_stage_5__3931_, data_stage_5__3930_, data_stage_5__3929_, data_stage_5__3928_, data_stage_5__3927_, data_stage_5__3926_, data_stage_5__3925_, data_stage_5__3924_, data_stage_5__3923_, data_stage_5__3922_, data_stage_5__3921_, data_stage_5__3920_, data_stage_5__3919_, data_stage_5__3918_, data_stage_5__3917_, data_stage_5__3916_, data_stage_5__3915_, data_stage_5__3914_, data_stage_5__3913_, data_stage_5__3912_, data_stage_5__3911_, data_stage_5__3910_, data_stage_5__3909_, data_stage_5__3908_, data_stage_5__3907_, data_stage_5__3906_, data_stage_5__3905_, data_stage_5__3904_, data_stage_5__3903_, data_stage_5__3902_, data_stage_5__3901_, data_stage_5__3900_, data_stage_5__3899_, data_stage_5__3898_, data_stage_5__3897_, data_stage_5__3896_, data_stage_5__3895_, data_stage_5__3894_, data_stage_5__3893_, data_stage_5__3892_, data_stage_5__3891_, data_stage_5__3890_, data_stage_5__3889_, data_stage_5__3888_, data_stage_5__3887_, data_stage_5__3886_, data_stage_5__3885_, data_stage_5__3884_, data_stage_5__3883_, data_stage_5__3882_, data_stage_5__3881_, data_stage_5__3880_, data_stage_5__3879_, data_stage_5__3878_, data_stage_5__3877_, data_stage_5__3876_, data_stage_5__3875_, data_stage_5__3874_, data_stage_5__3873_, data_stage_5__3872_, data_stage_5__3871_, data_stage_5__3870_, data_stage_5__3869_, data_stage_5__3868_, data_stage_5__3867_, data_stage_5__3866_, data_stage_5__3865_, data_stage_5__3864_, data_stage_5__3863_, data_stage_5__3862_, data_stage_5__3861_, data_stage_5__3860_, data_stage_5__3859_, data_stage_5__3858_, data_stage_5__3857_, data_stage_5__3856_, data_stage_5__3855_, data_stage_5__3854_, data_stage_5__3853_, data_stage_5__3852_, data_stage_5__3851_, data_stage_5__3850_, data_stage_5__3849_, data_stage_5__3848_, data_stage_5__3847_, data_stage_5__3846_, data_stage_5__3845_, data_stage_5__3844_, data_stage_5__3843_, data_stage_5__3842_, data_stage_5__3841_, data_stage_5__3840_, data_stage_5__3839_, data_stage_5__3838_, data_stage_5__3837_, data_stage_5__3836_, data_stage_5__3835_, data_stage_5__3834_, data_stage_5__3833_, data_stage_5__3832_, data_stage_5__3831_, data_stage_5__3830_, data_stage_5__3829_, data_stage_5__3828_, data_stage_5__3827_, data_stage_5__3826_, data_stage_5__3825_, data_stage_5__3824_, data_stage_5__3823_, data_stage_5__3822_, data_stage_5__3821_, data_stage_5__3820_, data_stage_5__3819_, data_stage_5__3818_, data_stage_5__3817_, data_stage_5__3816_, data_stage_5__3815_, data_stage_5__3814_, data_stage_5__3813_, data_stage_5__3812_, data_stage_5__3811_, data_stage_5__3810_, data_stage_5__3809_, data_stage_5__3808_, data_stage_5__3807_, data_stage_5__3806_, data_stage_5__3805_, data_stage_5__3804_, data_stage_5__3803_, data_stage_5__3802_, data_stage_5__3801_, data_stage_5__3800_, data_stage_5__3799_, data_stage_5__3798_, data_stage_5__3797_, data_stage_5__3796_, data_stage_5__3795_, data_stage_5__3794_, data_stage_5__3793_, data_stage_5__3792_, data_stage_5__3791_, data_stage_5__3790_, data_stage_5__3789_, data_stage_5__3788_, data_stage_5__3787_, data_stage_5__3786_, data_stage_5__3785_, data_stage_5__3784_, data_stage_5__3783_, data_stage_5__3782_, data_stage_5__3781_, data_stage_5__3780_, data_stage_5__3779_, data_stage_5__3778_, data_stage_5__3777_, data_stage_5__3776_, data_stage_5__3775_, data_stage_5__3774_, data_stage_5__3773_, data_stage_5__3772_, data_stage_5__3771_, data_stage_5__3770_, data_stage_5__3769_, data_stage_5__3768_, data_stage_5__3767_, data_stage_5__3766_, data_stage_5__3765_, data_stage_5__3764_, data_stage_5__3763_, data_stage_5__3762_, data_stage_5__3761_, data_stage_5__3760_, data_stage_5__3759_, data_stage_5__3758_, data_stage_5__3757_, data_stage_5__3756_, data_stage_5__3755_, data_stage_5__3754_, data_stage_5__3753_, data_stage_5__3752_, data_stage_5__3751_, data_stage_5__3750_, data_stage_5__3749_, data_stage_5__3748_, data_stage_5__3747_, data_stage_5__3746_, data_stage_5__3745_, data_stage_5__3744_, data_stage_5__3743_, data_stage_5__3742_, data_stage_5__3741_, data_stage_5__3740_, data_stage_5__3739_, data_stage_5__3738_, data_stage_5__3737_, data_stage_5__3736_, data_stage_5__3735_, data_stage_5__3734_, data_stage_5__3733_, data_stage_5__3732_, data_stage_5__3731_, data_stage_5__3730_, data_stage_5__3729_, data_stage_5__3728_, data_stage_5__3727_, data_stage_5__3726_, data_stage_5__3725_, data_stage_5__3724_, data_stage_5__3723_, data_stage_5__3722_, data_stage_5__3721_, data_stage_5__3720_, data_stage_5__3719_, data_stage_5__3718_, data_stage_5__3717_, data_stage_5__3716_, data_stage_5__3715_, data_stage_5__3714_, data_stage_5__3713_, data_stage_5__3712_, data_stage_5__3711_, data_stage_5__3710_, data_stage_5__3709_, data_stage_5__3708_, data_stage_5__3707_, data_stage_5__3706_, data_stage_5__3705_, data_stage_5__3704_, data_stage_5__3703_, data_stage_5__3702_, data_stage_5__3701_, data_stage_5__3700_, data_stage_5__3699_, data_stage_5__3698_, data_stage_5__3697_, data_stage_5__3696_, data_stage_5__3695_, data_stage_5__3694_, data_stage_5__3693_, data_stage_5__3692_, data_stage_5__3691_, data_stage_5__3690_, data_stage_5__3689_, data_stage_5__3688_, data_stage_5__3687_, data_stage_5__3686_, data_stage_5__3685_, data_stage_5__3684_, data_stage_5__3683_, data_stage_5__3682_, data_stage_5__3681_, data_stage_5__3680_, data_stage_5__3679_, data_stage_5__3678_, data_stage_5__3677_, data_stage_5__3676_, data_stage_5__3675_, data_stage_5__3674_, data_stage_5__3673_, data_stage_5__3672_, data_stage_5__3671_, data_stage_5__3670_, data_stage_5__3669_, data_stage_5__3668_, data_stage_5__3667_, data_stage_5__3666_, data_stage_5__3665_, data_stage_5__3664_, data_stage_5__3663_, data_stage_5__3662_, data_stage_5__3661_, data_stage_5__3660_, data_stage_5__3659_, data_stage_5__3658_, data_stage_5__3657_, data_stage_5__3656_, data_stage_5__3655_, data_stage_5__3654_, data_stage_5__3653_, data_stage_5__3652_, data_stage_5__3651_, data_stage_5__3650_, data_stage_5__3649_, data_stage_5__3648_, data_stage_5__3647_, data_stage_5__3646_, data_stage_5__3645_, data_stage_5__3644_, data_stage_5__3643_, data_stage_5__3642_, data_stage_5__3641_, data_stage_5__3640_, data_stage_5__3639_, data_stage_5__3638_, data_stage_5__3637_, data_stage_5__3636_, data_stage_5__3635_, data_stage_5__3634_, data_stage_5__3633_, data_stage_5__3632_, data_stage_5__3631_, data_stage_5__3630_, data_stage_5__3629_, data_stage_5__3628_, data_stage_5__3627_, data_stage_5__3626_, data_stage_5__3625_, data_stage_5__3624_, data_stage_5__3623_, data_stage_5__3622_, data_stage_5__3621_, data_stage_5__3620_, data_stage_5__3619_, data_stage_5__3618_, data_stage_5__3617_, data_stage_5__3616_, data_stage_5__3615_, data_stage_5__3614_, data_stage_5__3613_, data_stage_5__3612_, data_stage_5__3611_, data_stage_5__3610_, data_stage_5__3609_, data_stage_5__3608_, data_stage_5__3607_, data_stage_5__3606_, data_stage_5__3605_, data_stage_5__3604_, data_stage_5__3603_, data_stage_5__3602_, data_stage_5__3601_, data_stage_5__3600_, data_stage_5__3599_, data_stage_5__3598_, data_stage_5__3597_, data_stage_5__3596_, data_stage_5__3595_, data_stage_5__3594_, data_stage_5__3593_, data_stage_5__3592_, data_stage_5__3591_, data_stage_5__3590_, data_stage_5__3589_, data_stage_5__3588_, data_stage_5__3587_, data_stage_5__3586_, data_stage_5__3585_, data_stage_5__3584_, data_stage_5__3583_, data_stage_5__3582_, data_stage_5__3581_, data_stage_5__3580_, data_stage_5__3579_, data_stage_5__3578_, data_stage_5__3577_, data_stage_5__3576_, data_stage_5__3575_, data_stage_5__3574_, data_stage_5__3573_, data_stage_5__3572_, data_stage_5__3571_, data_stage_5__3570_, data_stage_5__3569_, data_stage_5__3568_, data_stage_5__3567_, data_stage_5__3566_, data_stage_5__3565_, data_stage_5__3564_, data_stage_5__3563_, data_stage_5__3562_, data_stage_5__3561_, data_stage_5__3560_, data_stage_5__3559_, data_stage_5__3558_, data_stage_5__3557_, data_stage_5__3556_, data_stage_5__3555_, data_stage_5__3554_, data_stage_5__3553_, data_stage_5__3552_, data_stage_5__3551_, data_stage_5__3550_, data_stage_5__3549_, data_stage_5__3548_, data_stage_5__3547_, data_stage_5__3546_, data_stage_5__3545_, data_stage_5__3544_, data_stage_5__3543_, data_stage_5__3542_, data_stage_5__3541_, data_stage_5__3540_, data_stage_5__3539_, data_stage_5__3538_, data_stage_5__3537_, data_stage_5__3536_, data_stage_5__3535_, data_stage_5__3534_, data_stage_5__3533_, data_stage_5__3532_, data_stage_5__3531_, data_stage_5__3530_, data_stage_5__3529_, data_stage_5__3528_, data_stage_5__3527_, data_stage_5__3526_, data_stage_5__3525_, data_stage_5__3524_, data_stage_5__3523_, data_stage_5__3522_, data_stage_5__3521_, data_stage_5__3520_, data_stage_5__3519_, data_stage_5__3518_, data_stage_5__3517_, data_stage_5__3516_, data_stage_5__3515_, data_stage_5__3514_, data_stage_5__3513_, data_stage_5__3512_, data_stage_5__3511_, data_stage_5__3510_, data_stage_5__3509_, data_stage_5__3508_, data_stage_5__3507_, data_stage_5__3506_, data_stage_5__3505_, data_stage_5__3504_, data_stage_5__3503_, data_stage_5__3502_, data_stage_5__3501_, data_stage_5__3500_, data_stage_5__3499_, data_stage_5__3498_, data_stage_5__3497_, data_stage_5__3496_, data_stage_5__3495_, data_stage_5__3494_, data_stage_5__3493_, data_stage_5__3492_, data_stage_5__3491_, data_stage_5__3490_, data_stage_5__3489_, data_stage_5__3488_, data_stage_5__3487_, data_stage_5__3486_, data_stage_5__3485_, data_stage_5__3484_, data_stage_5__3483_, data_stage_5__3482_, data_stage_5__3481_, data_stage_5__3480_, data_stage_5__3479_, data_stage_5__3478_, data_stage_5__3477_, data_stage_5__3476_, data_stage_5__3475_, data_stage_5__3474_, data_stage_5__3473_, data_stage_5__3472_, data_stage_5__3471_, data_stage_5__3470_, data_stage_5__3469_, data_stage_5__3468_, data_stage_5__3467_, data_stage_5__3466_, data_stage_5__3465_, data_stage_5__3464_, data_stage_5__3463_, data_stage_5__3462_, data_stage_5__3461_, data_stage_5__3460_, data_stage_5__3459_, data_stage_5__3458_, data_stage_5__3457_, data_stage_5__3456_, data_stage_5__3455_, data_stage_5__3454_, data_stage_5__3453_, data_stage_5__3452_, data_stage_5__3451_, data_stage_5__3450_, data_stage_5__3449_, data_stage_5__3448_, data_stage_5__3447_, data_stage_5__3446_, data_stage_5__3445_, data_stage_5__3444_, data_stage_5__3443_, data_stage_5__3442_, data_stage_5__3441_, data_stage_5__3440_, data_stage_5__3439_, data_stage_5__3438_, data_stage_5__3437_, data_stage_5__3436_, data_stage_5__3435_, data_stage_5__3434_, data_stage_5__3433_, data_stage_5__3432_, data_stage_5__3431_, data_stage_5__3430_, data_stage_5__3429_, data_stage_5__3428_, data_stage_5__3427_, data_stage_5__3426_, data_stage_5__3425_, data_stage_5__3424_, data_stage_5__3423_, data_stage_5__3422_, data_stage_5__3421_, data_stage_5__3420_, data_stage_5__3419_, data_stage_5__3418_, data_stage_5__3417_, data_stage_5__3416_, data_stage_5__3415_, data_stage_5__3414_, data_stage_5__3413_, data_stage_5__3412_, data_stage_5__3411_, data_stage_5__3410_, data_stage_5__3409_, data_stage_5__3408_, data_stage_5__3407_, data_stage_5__3406_, data_stage_5__3405_, data_stage_5__3404_, data_stage_5__3403_, data_stage_5__3402_, data_stage_5__3401_, data_stage_5__3400_, data_stage_5__3399_, data_stage_5__3398_, data_stage_5__3397_, data_stage_5__3396_, data_stage_5__3395_, data_stage_5__3394_, data_stage_5__3393_, data_stage_5__3392_, data_stage_5__3391_, data_stage_5__3390_, data_stage_5__3389_, data_stage_5__3388_, data_stage_5__3387_, data_stage_5__3386_, data_stage_5__3385_, data_stage_5__3384_, data_stage_5__3383_, data_stage_5__3382_, data_stage_5__3381_, data_stage_5__3380_, data_stage_5__3379_, data_stage_5__3378_, data_stage_5__3377_, data_stage_5__3376_, data_stage_5__3375_, data_stage_5__3374_, data_stage_5__3373_, data_stage_5__3372_, data_stage_5__3371_, data_stage_5__3370_, data_stage_5__3369_, data_stage_5__3368_, data_stage_5__3367_, data_stage_5__3366_, data_stage_5__3365_, data_stage_5__3364_, data_stage_5__3363_, data_stage_5__3362_, data_stage_5__3361_, data_stage_5__3360_, data_stage_5__3359_, data_stage_5__3358_, data_stage_5__3357_, data_stage_5__3356_, data_stage_5__3355_, data_stage_5__3354_, data_stage_5__3353_, data_stage_5__3352_, data_stage_5__3351_, data_stage_5__3350_, data_stage_5__3349_, data_stage_5__3348_, data_stage_5__3347_, data_stage_5__3346_, data_stage_5__3345_, data_stage_5__3344_, data_stage_5__3343_, data_stage_5__3342_, data_stage_5__3341_, data_stage_5__3340_, data_stage_5__3339_, data_stage_5__3338_, data_stage_5__3337_, data_stage_5__3336_, data_stage_5__3335_, data_stage_5__3334_, data_stage_5__3333_, data_stage_5__3332_, data_stage_5__3331_, data_stage_5__3330_, data_stage_5__3329_, data_stage_5__3328_, data_stage_5__3327_, data_stage_5__3326_, data_stage_5__3325_, data_stage_5__3324_, data_stage_5__3323_, data_stage_5__3322_, data_stage_5__3321_, data_stage_5__3320_, data_stage_5__3319_, data_stage_5__3318_, data_stage_5__3317_, data_stage_5__3316_, data_stage_5__3315_, data_stage_5__3314_, data_stage_5__3313_, data_stage_5__3312_, data_stage_5__3311_, data_stage_5__3310_, data_stage_5__3309_, data_stage_5__3308_, data_stage_5__3307_, data_stage_5__3306_, data_stage_5__3305_, data_stage_5__3304_, data_stage_5__3303_, data_stage_5__3302_, data_stage_5__3301_, data_stage_5__3300_, data_stage_5__3299_, data_stage_5__3298_, data_stage_5__3297_, data_stage_5__3296_, data_stage_5__3295_, data_stage_5__3294_, data_stage_5__3293_, data_stage_5__3292_, data_stage_5__3291_, data_stage_5__3290_, data_stage_5__3289_, data_stage_5__3288_, data_stage_5__3287_, data_stage_5__3286_, data_stage_5__3285_, data_stage_5__3284_, data_stage_5__3283_, data_stage_5__3282_, data_stage_5__3281_, data_stage_5__3280_, data_stage_5__3279_, data_stage_5__3278_, data_stage_5__3277_, data_stage_5__3276_, data_stage_5__3275_, data_stage_5__3274_, data_stage_5__3273_, data_stage_5__3272_, data_stage_5__3271_, data_stage_5__3270_, data_stage_5__3269_, data_stage_5__3268_, data_stage_5__3267_, data_stage_5__3266_, data_stage_5__3265_, data_stage_5__3264_, data_stage_5__3263_, data_stage_5__3262_, data_stage_5__3261_, data_stage_5__3260_, data_stage_5__3259_, data_stage_5__3258_, data_stage_5__3257_, data_stage_5__3256_, data_stage_5__3255_, data_stage_5__3254_, data_stage_5__3253_, data_stage_5__3252_, data_stage_5__3251_, data_stage_5__3250_, data_stage_5__3249_, data_stage_5__3248_, data_stage_5__3247_, data_stage_5__3246_, data_stage_5__3245_, data_stage_5__3244_, data_stage_5__3243_, data_stage_5__3242_, data_stage_5__3241_, data_stage_5__3240_, data_stage_5__3239_, data_stage_5__3238_, data_stage_5__3237_, data_stage_5__3236_, data_stage_5__3235_, data_stage_5__3234_, data_stage_5__3233_, data_stage_5__3232_, data_stage_5__3231_, data_stage_5__3230_, data_stage_5__3229_, data_stage_5__3228_, data_stage_5__3227_, data_stage_5__3226_, data_stage_5__3225_, data_stage_5__3224_, data_stage_5__3223_, data_stage_5__3222_, data_stage_5__3221_, data_stage_5__3220_, data_stage_5__3219_, data_stage_5__3218_, data_stage_5__3217_, data_stage_5__3216_, data_stage_5__3215_, data_stage_5__3214_, data_stage_5__3213_, data_stage_5__3212_, data_stage_5__3211_, data_stage_5__3210_, data_stage_5__3209_, data_stage_5__3208_, data_stage_5__3207_, data_stage_5__3206_, data_stage_5__3205_, data_stage_5__3204_, data_stage_5__3203_, data_stage_5__3202_, data_stage_5__3201_, data_stage_5__3200_, data_stage_5__3199_, data_stage_5__3198_, data_stage_5__3197_, data_stage_5__3196_, data_stage_5__3195_, data_stage_5__3194_, data_stage_5__3193_, data_stage_5__3192_, data_stage_5__3191_, data_stage_5__3190_, data_stage_5__3189_, data_stage_5__3188_, data_stage_5__3187_, data_stage_5__3186_, data_stage_5__3185_, data_stage_5__3184_, data_stage_5__3183_, data_stage_5__3182_, data_stage_5__3181_, data_stage_5__3180_, data_stage_5__3179_, data_stage_5__3178_, data_stage_5__3177_, data_stage_5__3176_, data_stage_5__3175_, data_stage_5__3174_, data_stage_5__3173_, data_stage_5__3172_, data_stage_5__3171_, data_stage_5__3170_, data_stage_5__3169_, data_stage_5__3168_, data_stage_5__3167_, data_stage_5__3166_, data_stage_5__3165_, data_stage_5__3164_, data_stage_5__3163_, data_stage_5__3162_, data_stage_5__3161_, data_stage_5__3160_, data_stage_5__3159_, data_stage_5__3158_, data_stage_5__3157_, data_stage_5__3156_, data_stage_5__3155_, data_stage_5__3154_, data_stage_5__3153_, data_stage_5__3152_, data_stage_5__3151_, data_stage_5__3150_, data_stage_5__3149_, data_stage_5__3148_, data_stage_5__3147_, data_stage_5__3146_, data_stage_5__3145_, data_stage_5__3144_, data_stage_5__3143_, data_stage_5__3142_, data_stage_5__3141_, data_stage_5__3140_, data_stage_5__3139_, data_stage_5__3138_, data_stage_5__3137_, data_stage_5__3136_, data_stage_5__3135_, data_stage_5__3134_, data_stage_5__3133_, data_stage_5__3132_, data_stage_5__3131_, data_stage_5__3130_, data_stage_5__3129_, data_stage_5__3128_, data_stage_5__3127_, data_stage_5__3126_, data_stage_5__3125_, data_stage_5__3124_, data_stage_5__3123_, data_stage_5__3122_, data_stage_5__3121_, data_stage_5__3120_, data_stage_5__3119_, data_stage_5__3118_, data_stage_5__3117_, data_stage_5__3116_, data_stage_5__3115_, data_stage_5__3114_, data_stage_5__3113_, data_stage_5__3112_, data_stage_5__3111_, data_stage_5__3110_, data_stage_5__3109_, data_stage_5__3108_, data_stage_5__3107_, data_stage_5__3106_, data_stage_5__3105_, data_stage_5__3104_, data_stage_5__3103_, data_stage_5__3102_, data_stage_5__3101_, data_stage_5__3100_, data_stage_5__3099_, data_stage_5__3098_, data_stage_5__3097_, data_stage_5__3096_, data_stage_5__3095_, data_stage_5__3094_, data_stage_5__3093_, data_stage_5__3092_, data_stage_5__3091_, data_stage_5__3090_, data_stage_5__3089_, data_stage_5__3088_, data_stage_5__3087_, data_stage_5__3086_, data_stage_5__3085_, data_stage_5__3084_, data_stage_5__3083_, data_stage_5__3082_, data_stage_5__3081_, data_stage_5__3080_, data_stage_5__3079_, data_stage_5__3078_, data_stage_5__3077_, data_stage_5__3076_, data_stage_5__3075_, data_stage_5__3074_, data_stage_5__3073_, data_stage_5__3072_, data_stage_5__3071_, data_stage_5__3070_, data_stage_5__3069_, data_stage_5__3068_, data_stage_5__3067_, data_stage_5__3066_, data_stage_5__3065_, data_stage_5__3064_, data_stage_5__3063_, data_stage_5__3062_, data_stage_5__3061_, data_stage_5__3060_, data_stage_5__3059_, data_stage_5__3058_, data_stage_5__3057_, data_stage_5__3056_, data_stage_5__3055_, data_stage_5__3054_, data_stage_5__3053_, data_stage_5__3052_, data_stage_5__3051_, data_stage_5__3050_, data_stage_5__3049_, data_stage_5__3048_, data_stage_5__3047_, data_stage_5__3046_, data_stage_5__3045_, data_stage_5__3044_, data_stage_5__3043_, data_stage_5__3042_, data_stage_5__3041_, data_stage_5__3040_, data_stage_5__3039_, data_stage_5__3038_, data_stage_5__3037_, data_stage_5__3036_, data_stage_5__3035_, data_stage_5__3034_, data_stage_5__3033_, data_stage_5__3032_, data_stage_5__3031_, data_stage_5__3030_, data_stage_5__3029_, data_stage_5__3028_, data_stage_5__3027_, data_stage_5__3026_, data_stage_5__3025_, data_stage_5__3024_, data_stage_5__3023_, data_stage_5__3022_, data_stage_5__3021_, data_stage_5__3020_, data_stage_5__3019_, data_stage_5__3018_, data_stage_5__3017_, data_stage_5__3016_, data_stage_5__3015_, data_stage_5__3014_, data_stage_5__3013_, data_stage_5__3012_, data_stage_5__3011_, data_stage_5__3010_, data_stage_5__3009_, data_stage_5__3008_, data_stage_5__3007_, data_stage_5__3006_, data_stage_5__3005_, data_stage_5__3004_, data_stage_5__3003_, data_stage_5__3002_, data_stage_5__3001_, data_stage_5__3000_, data_stage_5__2999_, data_stage_5__2998_, data_stage_5__2997_, data_stage_5__2996_, data_stage_5__2995_, data_stage_5__2994_, data_stage_5__2993_, data_stage_5__2992_, data_stage_5__2991_, data_stage_5__2990_, data_stage_5__2989_, data_stage_5__2988_, data_stage_5__2987_, data_stage_5__2986_, data_stage_5__2985_, data_stage_5__2984_, data_stage_5__2983_, data_stage_5__2982_, data_stage_5__2981_, data_stage_5__2980_, data_stage_5__2979_, data_stage_5__2978_, data_stage_5__2977_, data_stage_5__2976_, data_stage_5__2975_, data_stage_5__2974_, data_stage_5__2973_, data_stage_5__2972_, data_stage_5__2971_, data_stage_5__2970_, data_stage_5__2969_, data_stage_5__2968_, data_stage_5__2967_, data_stage_5__2966_, data_stage_5__2965_, data_stage_5__2964_, data_stage_5__2963_, data_stage_5__2962_, data_stage_5__2961_, data_stage_5__2960_, data_stage_5__2959_, data_stage_5__2958_, data_stage_5__2957_, data_stage_5__2956_, data_stage_5__2955_, data_stage_5__2954_, data_stage_5__2953_, data_stage_5__2952_, data_stage_5__2951_, data_stage_5__2950_, data_stage_5__2949_, data_stage_5__2948_, data_stage_5__2947_, data_stage_5__2946_, data_stage_5__2945_, data_stage_5__2944_, data_stage_5__2943_, data_stage_5__2942_, data_stage_5__2941_, data_stage_5__2940_, data_stage_5__2939_, data_stage_5__2938_, data_stage_5__2937_, data_stage_5__2936_, data_stage_5__2935_, data_stage_5__2934_, data_stage_5__2933_, data_stage_5__2932_, data_stage_5__2931_, data_stage_5__2930_, data_stage_5__2929_, data_stage_5__2928_, data_stage_5__2927_, data_stage_5__2926_, data_stage_5__2925_, data_stage_5__2924_, data_stage_5__2923_, data_stage_5__2922_, data_stage_5__2921_, data_stage_5__2920_, data_stage_5__2919_, data_stage_5__2918_, data_stage_5__2917_, data_stage_5__2916_, data_stage_5__2915_, data_stage_5__2914_, data_stage_5__2913_, data_stage_5__2912_, data_stage_5__2911_, data_stage_5__2910_, data_stage_5__2909_, data_stage_5__2908_, data_stage_5__2907_, data_stage_5__2906_, data_stage_5__2905_, data_stage_5__2904_, data_stage_5__2903_, data_stage_5__2902_, data_stage_5__2901_, data_stage_5__2900_, data_stage_5__2899_, data_stage_5__2898_, data_stage_5__2897_, data_stage_5__2896_, data_stage_5__2895_, data_stage_5__2894_, data_stage_5__2893_, data_stage_5__2892_, data_stage_5__2891_, data_stage_5__2890_, data_stage_5__2889_, data_stage_5__2888_, data_stage_5__2887_, data_stage_5__2886_, data_stage_5__2885_, data_stage_5__2884_, data_stage_5__2883_, data_stage_5__2882_, data_stage_5__2881_, data_stage_5__2880_, data_stage_5__2879_, data_stage_5__2878_, data_stage_5__2877_, data_stage_5__2876_, data_stage_5__2875_, data_stage_5__2874_, data_stage_5__2873_, data_stage_5__2872_, data_stage_5__2871_, data_stage_5__2870_, data_stage_5__2869_, data_stage_5__2868_, data_stage_5__2867_, data_stage_5__2866_, data_stage_5__2865_, data_stage_5__2864_, data_stage_5__2863_, data_stage_5__2862_, data_stage_5__2861_, data_stage_5__2860_, data_stage_5__2859_, data_stage_5__2858_, data_stage_5__2857_, data_stage_5__2856_, data_stage_5__2855_, data_stage_5__2854_, data_stage_5__2853_, data_stage_5__2852_, data_stage_5__2851_, data_stage_5__2850_, data_stage_5__2849_, data_stage_5__2848_, data_stage_5__2847_, data_stage_5__2846_, data_stage_5__2845_, data_stage_5__2844_, data_stage_5__2843_, data_stage_5__2842_, data_stage_5__2841_, data_stage_5__2840_, data_stage_5__2839_, data_stage_5__2838_, data_stage_5__2837_, data_stage_5__2836_, data_stage_5__2835_, data_stage_5__2834_, data_stage_5__2833_, data_stage_5__2832_, data_stage_5__2831_, data_stage_5__2830_, data_stage_5__2829_, data_stage_5__2828_, data_stage_5__2827_, data_stage_5__2826_, data_stage_5__2825_, data_stage_5__2824_, data_stage_5__2823_, data_stage_5__2822_, data_stage_5__2821_, data_stage_5__2820_, data_stage_5__2819_, data_stage_5__2818_, data_stage_5__2817_, data_stage_5__2816_, data_stage_5__2815_, data_stage_5__2814_, data_stage_5__2813_, data_stage_5__2812_, data_stage_5__2811_, data_stage_5__2810_, data_stage_5__2809_, data_stage_5__2808_, data_stage_5__2807_, data_stage_5__2806_, data_stage_5__2805_, data_stage_5__2804_, data_stage_5__2803_, data_stage_5__2802_, data_stage_5__2801_, data_stage_5__2800_, data_stage_5__2799_, data_stage_5__2798_, data_stage_5__2797_, data_stage_5__2796_, data_stage_5__2795_, data_stage_5__2794_, data_stage_5__2793_, data_stage_5__2792_, data_stage_5__2791_, data_stage_5__2790_, data_stage_5__2789_, data_stage_5__2788_, data_stage_5__2787_, data_stage_5__2786_, data_stage_5__2785_, data_stage_5__2784_, data_stage_5__2783_, data_stage_5__2782_, data_stage_5__2781_, data_stage_5__2780_, data_stage_5__2779_, data_stage_5__2778_, data_stage_5__2777_, data_stage_5__2776_, data_stage_5__2775_, data_stage_5__2774_, data_stage_5__2773_, data_stage_5__2772_, data_stage_5__2771_, data_stage_5__2770_, data_stage_5__2769_, data_stage_5__2768_, data_stage_5__2767_, data_stage_5__2766_, data_stage_5__2765_, data_stage_5__2764_, data_stage_5__2763_, data_stage_5__2762_, data_stage_5__2761_, data_stage_5__2760_, data_stage_5__2759_, data_stage_5__2758_, data_stage_5__2757_, data_stage_5__2756_, data_stage_5__2755_, data_stage_5__2754_, data_stage_5__2753_, data_stage_5__2752_, data_stage_5__2751_, data_stage_5__2750_, data_stage_5__2749_, data_stage_5__2748_, data_stage_5__2747_, data_stage_5__2746_, data_stage_5__2745_, data_stage_5__2744_, data_stage_5__2743_, data_stage_5__2742_, data_stage_5__2741_, data_stage_5__2740_, data_stage_5__2739_, data_stage_5__2738_, data_stage_5__2737_, data_stage_5__2736_, data_stage_5__2735_, data_stage_5__2734_, data_stage_5__2733_, data_stage_5__2732_, data_stage_5__2731_, data_stage_5__2730_, data_stage_5__2729_, data_stage_5__2728_, data_stage_5__2727_, data_stage_5__2726_, data_stage_5__2725_, data_stage_5__2724_, data_stage_5__2723_, data_stage_5__2722_, data_stage_5__2721_, data_stage_5__2720_, data_stage_5__2719_, data_stage_5__2718_, data_stage_5__2717_, data_stage_5__2716_, data_stage_5__2715_, data_stage_5__2714_, data_stage_5__2713_, data_stage_5__2712_, data_stage_5__2711_, data_stage_5__2710_, data_stage_5__2709_, data_stage_5__2708_, data_stage_5__2707_, data_stage_5__2706_, data_stage_5__2705_, data_stage_5__2704_, data_stage_5__2703_, data_stage_5__2702_, data_stage_5__2701_, data_stage_5__2700_, data_stage_5__2699_, data_stage_5__2698_, data_stage_5__2697_, data_stage_5__2696_, data_stage_5__2695_, data_stage_5__2694_, data_stage_5__2693_, data_stage_5__2692_, data_stage_5__2691_, data_stage_5__2690_, data_stage_5__2689_, data_stage_5__2688_, data_stage_5__2687_, data_stage_5__2686_, data_stage_5__2685_, data_stage_5__2684_, data_stage_5__2683_, data_stage_5__2682_, data_stage_5__2681_, data_stage_5__2680_, data_stage_5__2679_, data_stage_5__2678_, data_stage_5__2677_, data_stage_5__2676_, data_stage_5__2675_, data_stage_5__2674_, data_stage_5__2673_, data_stage_5__2672_, data_stage_5__2671_, data_stage_5__2670_, data_stage_5__2669_, data_stage_5__2668_, data_stage_5__2667_, data_stage_5__2666_, data_stage_5__2665_, data_stage_5__2664_, data_stage_5__2663_, data_stage_5__2662_, data_stage_5__2661_, data_stage_5__2660_, data_stage_5__2659_, data_stage_5__2658_, data_stage_5__2657_, data_stage_5__2656_, data_stage_5__2655_, data_stage_5__2654_, data_stage_5__2653_, data_stage_5__2652_, data_stage_5__2651_, data_stage_5__2650_, data_stage_5__2649_, data_stage_5__2648_, data_stage_5__2647_, data_stage_5__2646_, data_stage_5__2645_, data_stage_5__2644_, data_stage_5__2643_, data_stage_5__2642_, data_stage_5__2641_, data_stage_5__2640_, data_stage_5__2639_, data_stage_5__2638_, data_stage_5__2637_, data_stage_5__2636_, data_stage_5__2635_, data_stage_5__2634_, data_stage_5__2633_, data_stage_5__2632_, data_stage_5__2631_, data_stage_5__2630_, data_stage_5__2629_, data_stage_5__2628_, data_stage_5__2627_, data_stage_5__2626_, data_stage_5__2625_, data_stage_5__2624_, data_stage_5__2623_, data_stage_5__2622_, data_stage_5__2621_, data_stage_5__2620_, data_stage_5__2619_, data_stage_5__2618_, data_stage_5__2617_, data_stage_5__2616_, data_stage_5__2615_, data_stage_5__2614_, data_stage_5__2613_, data_stage_5__2612_, data_stage_5__2611_, data_stage_5__2610_, data_stage_5__2609_, data_stage_5__2608_, data_stage_5__2607_, data_stage_5__2606_, data_stage_5__2605_, data_stage_5__2604_, data_stage_5__2603_, data_stage_5__2602_, data_stage_5__2601_, data_stage_5__2600_, data_stage_5__2599_, data_stage_5__2598_, data_stage_5__2597_, data_stage_5__2596_, data_stage_5__2595_, data_stage_5__2594_, data_stage_5__2593_, data_stage_5__2592_, data_stage_5__2591_, data_stage_5__2590_, data_stage_5__2589_, data_stage_5__2588_, data_stage_5__2587_, data_stage_5__2586_, data_stage_5__2585_, data_stage_5__2584_, data_stage_5__2583_, data_stage_5__2582_, data_stage_5__2581_, data_stage_5__2580_, data_stage_5__2579_, data_stage_5__2578_, data_stage_5__2577_, data_stage_5__2576_, data_stage_5__2575_, data_stage_5__2574_, data_stage_5__2573_, data_stage_5__2572_, data_stage_5__2571_, data_stage_5__2570_, data_stage_5__2569_, data_stage_5__2568_, data_stage_5__2567_, data_stage_5__2566_, data_stage_5__2565_, data_stage_5__2564_, data_stage_5__2563_, data_stage_5__2562_, data_stage_5__2561_, data_stage_5__2560_, data_stage_5__2559_, data_stage_5__2558_, data_stage_5__2557_, data_stage_5__2556_, data_stage_5__2555_, data_stage_5__2554_, data_stage_5__2553_, data_stage_5__2552_, data_stage_5__2551_, data_stage_5__2550_, data_stage_5__2549_, data_stage_5__2548_, data_stage_5__2547_, data_stage_5__2546_, data_stage_5__2545_, data_stage_5__2544_, data_stage_5__2543_, data_stage_5__2542_, data_stage_5__2541_, data_stage_5__2540_, data_stage_5__2539_, data_stage_5__2538_, data_stage_5__2537_, data_stage_5__2536_, data_stage_5__2535_, data_stage_5__2534_, data_stage_5__2533_, data_stage_5__2532_, data_stage_5__2531_, data_stage_5__2530_, data_stage_5__2529_, data_stage_5__2528_, data_stage_5__2527_, data_stage_5__2526_, data_stage_5__2525_, data_stage_5__2524_, data_stage_5__2523_, data_stage_5__2522_, data_stage_5__2521_, data_stage_5__2520_, data_stage_5__2519_, data_stage_5__2518_, data_stage_5__2517_, data_stage_5__2516_, data_stage_5__2515_, data_stage_5__2514_, data_stage_5__2513_, data_stage_5__2512_, data_stage_5__2511_, data_stage_5__2510_, data_stage_5__2509_, data_stage_5__2508_, data_stage_5__2507_, data_stage_5__2506_, data_stage_5__2505_, data_stage_5__2504_, data_stage_5__2503_, data_stage_5__2502_, data_stage_5__2501_, data_stage_5__2500_, data_stage_5__2499_, data_stage_5__2498_, data_stage_5__2497_, data_stage_5__2496_, data_stage_5__2495_, data_stage_5__2494_, data_stage_5__2493_, data_stage_5__2492_, data_stage_5__2491_, data_stage_5__2490_, data_stage_5__2489_, data_stage_5__2488_, data_stage_5__2487_, data_stage_5__2486_, data_stage_5__2485_, data_stage_5__2484_, data_stage_5__2483_, data_stage_5__2482_, data_stage_5__2481_, data_stage_5__2480_, data_stage_5__2479_, data_stage_5__2478_, data_stage_5__2477_, data_stage_5__2476_, data_stage_5__2475_, data_stage_5__2474_, data_stage_5__2473_, data_stage_5__2472_, data_stage_5__2471_, data_stage_5__2470_, data_stage_5__2469_, data_stage_5__2468_, data_stage_5__2467_, data_stage_5__2466_, data_stage_5__2465_, data_stage_5__2464_, data_stage_5__2463_, data_stage_5__2462_, data_stage_5__2461_, data_stage_5__2460_, data_stage_5__2459_, data_stage_5__2458_, data_stage_5__2457_, data_stage_5__2456_, data_stage_5__2455_, data_stage_5__2454_, data_stage_5__2453_, data_stage_5__2452_, data_stage_5__2451_, data_stage_5__2450_, data_stage_5__2449_, data_stage_5__2448_, data_stage_5__2447_, data_stage_5__2446_, data_stage_5__2445_, data_stage_5__2444_, data_stage_5__2443_, data_stage_5__2442_, data_stage_5__2441_, data_stage_5__2440_, data_stage_5__2439_, data_stage_5__2438_, data_stage_5__2437_, data_stage_5__2436_, data_stage_5__2435_, data_stage_5__2434_, data_stage_5__2433_, data_stage_5__2432_, data_stage_5__2431_, data_stage_5__2430_, data_stage_5__2429_, data_stage_5__2428_, data_stage_5__2427_, data_stage_5__2426_, data_stage_5__2425_, data_stage_5__2424_, data_stage_5__2423_, data_stage_5__2422_, data_stage_5__2421_, data_stage_5__2420_, data_stage_5__2419_, data_stage_5__2418_, data_stage_5__2417_, data_stage_5__2416_, data_stage_5__2415_, data_stage_5__2414_, data_stage_5__2413_, data_stage_5__2412_, data_stage_5__2411_, data_stage_5__2410_, data_stage_5__2409_, data_stage_5__2408_, data_stage_5__2407_, data_stage_5__2406_, data_stage_5__2405_, data_stage_5__2404_, data_stage_5__2403_, data_stage_5__2402_, data_stage_5__2401_, data_stage_5__2400_, data_stage_5__2399_, data_stage_5__2398_, data_stage_5__2397_, data_stage_5__2396_, data_stage_5__2395_, data_stage_5__2394_, data_stage_5__2393_, data_stage_5__2392_, data_stage_5__2391_, data_stage_5__2390_, data_stage_5__2389_, data_stage_5__2388_, data_stage_5__2387_, data_stage_5__2386_, data_stage_5__2385_, data_stage_5__2384_, data_stage_5__2383_, data_stage_5__2382_, data_stage_5__2381_, data_stage_5__2380_, data_stage_5__2379_, data_stage_5__2378_, data_stage_5__2377_, data_stage_5__2376_, data_stage_5__2375_, data_stage_5__2374_, data_stage_5__2373_, data_stage_5__2372_, data_stage_5__2371_, data_stage_5__2370_, data_stage_5__2369_, data_stage_5__2368_, data_stage_5__2367_, data_stage_5__2366_, data_stage_5__2365_, data_stage_5__2364_, data_stage_5__2363_, data_stage_5__2362_, data_stage_5__2361_, data_stage_5__2360_, data_stage_5__2359_, data_stage_5__2358_, data_stage_5__2357_, data_stage_5__2356_, data_stage_5__2355_, data_stage_5__2354_, data_stage_5__2353_, data_stage_5__2352_, data_stage_5__2351_, data_stage_5__2350_, data_stage_5__2349_, data_stage_5__2348_, data_stage_5__2347_, data_stage_5__2346_, data_stage_5__2345_, data_stage_5__2344_, data_stage_5__2343_, data_stage_5__2342_, data_stage_5__2341_, data_stage_5__2340_, data_stage_5__2339_, data_stage_5__2338_, data_stage_5__2337_, data_stage_5__2336_, data_stage_5__2335_, data_stage_5__2334_, data_stage_5__2333_, data_stage_5__2332_, data_stage_5__2331_, data_stage_5__2330_, data_stage_5__2329_, data_stage_5__2328_, data_stage_5__2327_, data_stage_5__2326_, data_stage_5__2325_, data_stage_5__2324_, data_stage_5__2323_, data_stage_5__2322_, data_stage_5__2321_, data_stage_5__2320_, data_stage_5__2319_, data_stage_5__2318_, data_stage_5__2317_, data_stage_5__2316_, data_stage_5__2315_, data_stage_5__2314_, data_stage_5__2313_, data_stage_5__2312_, data_stage_5__2311_, data_stage_5__2310_, data_stage_5__2309_, data_stage_5__2308_, data_stage_5__2307_, data_stage_5__2306_, data_stage_5__2305_, data_stage_5__2304_, data_stage_5__2303_, data_stage_5__2302_, data_stage_5__2301_, data_stage_5__2300_, data_stage_5__2299_, data_stage_5__2298_, data_stage_5__2297_, data_stage_5__2296_, data_stage_5__2295_, data_stage_5__2294_, data_stage_5__2293_, data_stage_5__2292_, data_stage_5__2291_, data_stage_5__2290_, data_stage_5__2289_, data_stage_5__2288_, data_stage_5__2287_, data_stage_5__2286_, data_stage_5__2285_, data_stage_5__2284_, data_stage_5__2283_, data_stage_5__2282_, data_stage_5__2281_, data_stage_5__2280_, data_stage_5__2279_, data_stage_5__2278_, data_stage_5__2277_, data_stage_5__2276_, data_stage_5__2275_, data_stage_5__2274_, data_stage_5__2273_, data_stage_5__2272_, data_stage_5__2271_, data_stage_5__2270_, data_stage_5__2269_, data_stage_5__2268_, data_stage_5__2267_, data_stage_5__2266_, data_stage_5__2265_, data_stage_5__2264_, data_stage_5__2263_, data_stage_5__2262_, data_stage_5__2261_, data_stage_5__2260_, data_stage_5__2259_, data_stage_5__2258_, data_stage_5__2257_, data_stage_5__2256_, data_stage_5__2255_, data_stage_5__2254_, data_stage_5__2253_, data_stage_5__2252_, data_stage_5__2251_, data_stage_5__2250_, data_stage_5__2249_, data_stage_5__2248_, data_stage_5__2247_, data_stage_5__2246_, data_stage_5__2245_, data_stage_5__2244_, data_stage_5__2243_, data_stage_5__2242_, data_stage_5__2241_, data_stage_5__2240_, data_stage_5__2239_, data_stage_5__2238_, data_stage_5__2237_, data_stage_5__2236_, data_stage_5__2235_, data_stage_5__2234_, data_stage_5__2233_, data_stage_5__2232_, data_stage_5__2231_, data_stage_5__2230_, data_stage_5__2229_, data_stage_5__2228_, data_stage_5__2227_, data_stage_5__2226_, data_stage_5__2225_, data_stage_5__2224_, data_stage_5__2223_, data_stage_5__2222_, data_stage_5__2221_, data_stage_5__2220_, data_stage_5__2219_, data_stage_5__2218_, data_stage_5__2217_, data_stage_5__2216_, data_stage_5__2215_, data_stage_5__2214_, data_stage_5__2213_, data_stage_5__2212_, data_stage_5__2211_, data_stage_5__2210_, data_stage_5__2209_, data_stage_5__2208_, data_stage_5__2207_, data_stage_5__2206_, data_stage_5__2205_, data_stage_5__2204_, data_stage_5__2203_, data_stage_5__2202_, data_stage_5__2201_, data_stage_5__2200_, data_stage_5__2199_, data_stage_5__2198_, data_stage_5__2197_, data_stage_5__2196_, data_stage_5__2195_, data_stage_5__2194_, data_stage_5__2193_, data_stage_5__2192_, data_stage_5__2191_, data_stage_5__2190_, data_stage_5__2189_, data_stage_5__2188_, data_stage_5__2187_, data_stage_5__2186_, data_stage_5__2185_, data_stage_5__2184_, data_stage_5__2183_, data_stage_5__2182_, data_stage_5__2181_, data_stage_5__2180_, data_stage_5__2179_, data_stage_5__2178_, data_stage_5__2177_, data_stage_5__2176_, data_stage_5__2175_, data_stage_5__2174_, data_stage_5__2173_, data_stage_5__2172_, data_stage_5__2171_, data_stage_5__2170_, data_stage_5__2169_, data_stage_5__2168_, data_stage_5__2167_, data_stage_5__2166_, data_stage_5__2165_, data_stage_5__2164_, data_stage_5__2163_, data_stage_5__2162_, data_stage_5__2161_, data_stage_5__2160_, data_stage_5__2159_, data_stage_5__2158_, data_stage_5__2157_, data_stage_5__2156_, data_stage_5__2155_, data_stage_5__2154_, data_stage_5__2153_, data_stage_5__2152_, data_stage_5__2151_, data_stage_5__2150_, data_stage_5__2149_, data_stage_5__2148_, data_stage_5__2147_, data_stage_5__2146_, data_stage_5__2145_, data_stage_5__2144_, data_stage_5__2143_, data_stage_5__2142_, data_stage_5__2141_, data_stage_5__2140_, data_stage_5__2139_, data_stage_5__2138_, data_stage_5__2137_, data_stage_5__2136_, data_stage_5__2135_, data_stage_5__2134_, data_stage_5__2133_, data_stage_5__2132_, data_stage_5__2131_, data_stage_5__2130_, data_stage_5__2129_, data_stage_5__2128_, data_stage_5__2127_, data_stage_5__2126_, data_stage_5__2125_, data_stage_5__2124_, data_stage_5__2123_, data_stage_5__2122_, data_stage_5__2121_, data_stage_5__2120_, data_stage_5__2119_, data_stage_5__2118_, data_stage_5__2117_, data_stage_5__2116_, data_stage_5__2115_, data_stage_5__2114_, data_stage_5__2113_, data_stage_5__2112_, data_stage_5__2111_, data_stage_5__2110_, data_stage_5__2109_, data_stage_5__2108_, data_stage_5__2107_, data_stage_5__2106_, data_stage_5__2105_, data_stage_5__2104_, data_stage_5__2103_, data_stage_5__2102_, data_stage_5__2101_, data_stage_5__2100_, data_stage_5__2099_, data_stage_5__2098_, data_stage_5__2097_, data_stage_5__2096_, data_stage_5__2095_, data_stage_5__2094_, data_stage_5__2093_, data_stage_5__2092_, data_stage_5__2091_, data_stage_5__2090_, data_stage_5__2089_, data_stage_5__2088_, data_stage_5__2087_, data_stage_5__2086_, data_stage_5__2085_, data_stage_5__2084_, data_stage_5__2083_, data_stage_5__2082_, data_stage_5__2081_, data_stage_5__2080_, data_stage_5__2079_, data_stage_5__2078_, data_stage_5__2077_, data_stage_5__2076_, data_stage_5__2075_, data_stage_5__2074_, data_stage_5__2073_, data_stage_5__2072_, data_stage_5__2071_, data_stage_5__2070_, data_stage_5__2069_, data_stage_5__2068_, data_stage_5__2067_, data_stage_5__2066_, data_stage_5__2065_, data_stage_5__2064_, data_stage_5__2063_, data_stage_5__2062_, data_stage_5__2061_, data_stage_5__2060_, data_stage_5__2059_, data_stage_5__2058_, data_stage_5__2057_, data_stage_5__2056_, data_stage_5__2055_, data_stage_5__2054_, data_stage_5__2053_, data_stage_5__2052_, data_stage_5__2051_, data_stage_5__2050_, data_stage_5__2049_, data_stage_5__2048_ })
  );


  bsg_swap_width_p2048
  mux_stage_5__mux_swap_0__swap_inst
  (
    .data_i({ data_stage_5__4095_, data_stage_5__4094_, data_stage_5__4093_, data_stage_5__4092_, data_stage_5__4091_, data_stage_5__4090_, data_stage_5__4089_, data_stage_5__4088_, data_stage_5__4087_, data_stage_5__4086_, data_stage_5__4085_, data_stage_5__4084_, data_stage_5__4083_, data_stage_5__4082_, data_stage_5__4081_, data_stage_5__4080_, data_stage_5__4079_, data_stage_5__4078_, data_stage_5__4077_, data_stage_5__4076_, data_stage_5__4075_, data_stage_5__4074_, data_stage_5__4073_, data_stage_5__4072_, data_stage_5__4071_, data_stage_5__4070_, data_stage_5__4069_, data_stage_5__4068_, data_stage_5__4067_, data_stage_5__4066_, data_stage_5__4065_, data_stage_5__4064_, data_stage_5__4063_, data_stage_5__4062_, data_stage_5__4061_, data_stage_5__4060_, data_stage_5__4059_, data_stage_5__4058_, data_stage_5__4057_, data_stage_5__4056_, data_stage_5__4055_, data_stage_5__4054_, data_stage_5__4053_, data_stage_5__4052_, data_stage_5__4051_, data_stage_5__4050_, data_stage_5__4049_, data_stage_5__4048_, data_stage_5__4047_, data_stage_5__4046_, data_stage_5__4045_, data_stage_5__4044_, data_stage_5__4043_, data_stage_5__4042_, data_stage_5__4041_, data_stage_5__4040_, data_stage_5__4039_, data_stage_5__4038_, data_stage_5__4037_, data_stage_5__4036_, data_stage_5__4035_, data_stage_5__4034_, data_stage_5__4033_, data_stage_5__4032_, data_stage_5__4031_, data_stage_5__4030_, data_stage_5__4029_, data_stage_5__4028_, data_stage_5__4027_, data_stage_5__4026_, data_stage_5__4025_, data_stage_5__4024_, data_stage_5__4023_, data_stage_5__4022_, data_stage_5__4021_, data_stage_5__4020_, data_stage_5__4019_, data_stage_5__4018_, data_stage_5__4017_, data_stage_5__4016_, data_stage_5__4015_, data_stage_5__4014_, data_stage_5__4013_, data_stage_5__4012_, data_stage_5__4011_, data_stage_5__4010_, data_stage_5__4009_, data_stage_5__4008_, data_stage_5__4007_, data_stage_5__4006_, data_stage_5__4005_, data_stage_5__4004_, data_stage_5__4003_, data_stage_5__4002_, data_stage_5__4001_, data_stage_5__4000_, data_stage_5__3999_, data_stage_5__3998_, data_stage_5__3997_, data_stage_5__3996_, data_stage_5__3995_, data_stage_5__3994_, data_stage_5__3993_, data_stage_5__3992_, data_stage_5__3991_, data_stage_5__3990_, data_stage_5__3989_, data_stage_5__3988_, data_stage_5__3987_, data_stage_5__3986_, data_stage_5__3985_, data_stage_5__3984_, data_stage_5__3983_, data_stage_5__3982_, data_stage_5__3981_, data_stage_5__3980_, data_stage_5__3979_, data_stage_5__3978_, data_stage_5__3977_, data_stage_5__3976_, data_stage_5__3975_, data_stage_5__3974_, data_stage_5__3973_, data_stage_5__3972_, data_stage_5__3971_, data_stage_5__3970_, data_stage_5__3969_, data_stage_5__3968_, data_stage_5__3967_, data_stage_5__3966_, data_stage_5__3965_, data_stage_5__3964_, data_stage_5__3963_, data_stage_5__3962_, data_stage_5__3961_, data_stage_5__3960_, data_stage_5__3959_, data_stage_5__3958_, data_stage_5__3957_, data_stage_5__3956_, data_stage_5__3955_, data_stage_5__3954_, data_stage_5__3953_, data_stage_5__3952_, data_stage_5__3951_, data_stage_5__3950_, data_stage_5__3949_, data_stage_5__3948_, data_stage_5__3947_, data_stage_5__3946_, data_stage_5__3945_, data_stage_5__3944_, data_stage_5__3943_, data_stage_5__3942_, data_stage_5__3941_, data_stage_5__3940_, data_stage_5__3939_, data_stage_5__3938_, data_stage_5__3937_, data_stage_5__3936_, data_stage_5__3935_, data_stage_5__3934_, data_stage_5__3933_, data_stage_5__3932_, data_stage_5__3931_, data_stage_5__3930_, data_stage_5__3929_, data_stage_5__3928_, data_stage_5__3927_, data_stage_5__3926_, data_stage_5__3925_, data_stage_5__3924_, data_stage_5__3923_, data_stage_5__3922_, data_stage_5__3921_, data_stage_5__3920_, data_stage_5__3919_, data_stage_5__3918_, data_stage_5__3917_, data_stage_5__3916_, data_stage_5__3915_, data_stage_5__3914_, data_stage_5__3913_, data_stage_5__3912_, data_stage_5__3911_, data_stage_5__3910_, data_stage_5__3909_, data_stage_5__3908_, data_stage_5__3907_, data_stage_5__3906_, data_stage_5__3905_, data_stage_5__3904_, data_stage_5__3903_, data_stage_5__3902_, data_stage_5__3901_, data_stage_5__3900_, data_stage_5__3899_, data_stage_5__3898_, data_stage_5__3897_, data_stage_5__3896_, data_stage_5__3895_, data_stage_5__3894_, data_stage_5__3893_, data_stage_5__3892_, data_stage_5__3891_, data_stage_5__3890_, data_stage_5__3889_, data_stage_5__3888_, data_stage_5__3887_, data_stage_5__3886_, data_stage_5__3885_, data_stage_5__3884_, data_stage_5__3883_, data_stage_5__3882_, data_stage_5__3881_, data_stage_5__3880_, data_stage_5__3879_, data_stage_5__3878_, data_stage_5__3877_, data_stage_5__3876_, data_stage_5__3875_, data_stage_5__3874_, data_stage_5__3873_, data_stage_5__3872_, data_stage_5__3871_, data_stage_5__3870_, data_stage_5__3869_, data_stage_5__3868_, data_stage_5__3867_, data_stage_5__3866_, data_stage_5__3865_, data_stage_5__3864_, data_stage_5__3863_, data_stage_5__3862_, data_stage_5__3861_, data_stage_5__3860_, data_stage_5__3859_, data_stage_5__3858_, data_stage_5__3857_, data_stage_5__3856_, data_stage_5__3855_, data_stage_5__3854_, data_stage_5__3853_, data_stage_5__3852_, data_stage_5__3851_, data_stage_5__3850_, data_stage_5__3849_, data_stage_5__3848_, data_stage_5__3847_, data_stage_5__3846_, data_stage_5__3845_, data_stage_5__3844_, data_stage_5__3843_, data_stage_5__3842_, data_stage_5__3841_, data_stage_5__3840_, data_stage_5__3839_, data_stage_5__3838_, data_stage_5__3837_, data_stage_5__3836_, data_stage_5__3835_, data_stage_5__3834_, data_stage_5__3833_, data_stage_5__3832_, data_stage_5__3831_, data_stage_5__3830_, data_stage_5__3829_, data_stage_5__3828_, data_stage_5__3827_, data_stage_5__3826_, data_stage_5__3825_, data_stage_5__3824_, data_stage_5__3823_, data_stage_5__3822_, data_stage_5__3821_, data_stage_5__3820_, data_stage_5__3819_, data_stage_5__3818_, data_stage_5__3817_, data_stage_5__3816_, data_stage_5__3815_, data_stage_5__3814_, data_stage_5__3813_, data_stage_5__3812_, data_stage_5__3811_, data_stage_5__3810_, data_stage_5__3809_, data_stage_5__3808_, data_stage_5__3807_, data_stage_5__3806_, data_stage_5__3805_, data_stage_5__3804_, data_stage_5__3803_, data_stage_5__3802_, data_stage_5__3801_, data_stage_5__3800_, data_stage_5__3799_, data_stage_5__3798_, data_stage_5__3797_, data_stage_5__3796_, data_stage_5__3795_, data_stage_5__3794_, data_stage_5__3793_, data_stage_5__3792_, data_stage_5__3791_, data_stage_5__3790_, data_stage_5__3789_, data_stage_5__3788_, data_stage_5__3787_, data_stage_5__3786_, data_stage_5__3785_, data_stage_5__3784_, data_stage_5__3783_, data_stage_5__3782_, data_stage_5__3781_, data_stage_5__3780_, data_stage_5__3779_, data_stage_5__3778_, data_stage_5__3777_, data_stage_5__3776_, data_stage_5__3775_, data_stage_5__3774_, data_stage_5__3773_, data_stage_5__3772_, data_stage_5__3771_, data_stage_5__3770_, data_stage_5__3769_, data_stage_5__3768_, data_stage_5__3767_, data_stage_5__3766_, data_stage_5__3765_, data_stage_5__3764_, data_stage_5__3763_, data_stage_5__3762_, data_stage_5__3761_, data_stage_5__3760_, data_stage_5__3759_, data_stage_5__3758_, data_stage_5__3757_, data_stage_5__3756_, data_stage_5__3755_, data_stage_5__3754_, data_stage_5__3753_, data_stage_5__3752_, data_stage_5__3751_, data_stage_5__3750_, data_stage_5__3749_, data_stage_5__3748_, data_stage_5__3747_, data_stage_5__3746_, data_stage_5__3745_, data_stage_5__3744_, data_stage_5__3743_, data_stage_5__3742_, data_stage_5__3741_, data_stage_5__3740_, data_stage_5__3739_, data_stage_5__3738_, data_stage_5__3737_, data_stage_5__3736_, data_stage_5__3735_, data_stage_5__3734_, data_stage_5__3733_, data_stage_5__3732_, data_stage_5__3731_, data_stage_5__3730_, data_stage_5__3729_, data_stage_5__3728_, data_stage_5__3727_, data_stage_5__3726_, data_stage_5__3725_, data_stage_5__3724_, data_stage_5__3723_, data_stage_5__3722_, data_stage_5__3721_, data_stage_5__3720_, data_stage_5__3719_, data_stage_5__3718_, data_stage_5__3717_, data_stage_5__3716_, data_stage_5__3715_, data_stage_5__3714_, data_stage_5__3713_, data_stage_5__3712_, data_stage_5__3711_, data_stage_5__3710_, data_stage_5__3709_, data_stage_5__3708_, data_stage_5__3707_, data_stage_5__3706_, data_stage_5__3705_, data_stage_5__3704_, data_stage_5__3703_, data_stage_5__3702_, data_stage_5__3701_, data_stage_5__3700_, data_stage_5__3699_, data_stage_5__3698_, data_stage_5__3697_, data_stage_5__3696_, data_stage_5__3695_, data_stage_5__3694_, data_stage_5__3693_, data_stage_5__3692_, data_stage_5__3691_, data_stage_5__3690_, data_stage_5__3689_, data_stage_5__3688_, data_stage_5__3687_, data_stage_5__3686_, data_stage_5__3685_, data_stage_5__3684_, data_stage_5__3683_, data_stage_5__3682_, data_stage_5__3681_, data_stage_5__3680_, data_stage_5__3679_, data_stage_5__3678_, data_stage_5__3677_, data_stage_5__3676_, data_stage_5__3675_, data_stage_5__3674_, data_stage_5__3673_, data_stage_5__3672_, data_stage_5__3671_, data_stage_5__3670_, data_stage_5__3669_, data_stage_5__3668_, data_stage_5__3667_, data_stage_5__3666_, data_stage_5__3665_, data_stage_5__3664_, data_stage_5__3663_, data_stage_5__3662_, data_stage_5__3661_, data_stage_5__3660_, data_stage_5__3659_, data_stage_5__3658_, data_stage_5__3657_, data_stage_5__3656_, data_stage_5__3655_, data_stage_5__3654_, data_stage_5__3653_, data_stage_5__3652_, data_stage_5__3651_, data_stage_5__3650_, data_stage_5__3649_, data_stage_5__3648_, data_stage_5__3647_, data_stage_5__3646_, data_stage_5__3645_, data_stage_5__3644_, data_stage_5__3643_, data_stage_5__3642_, data_stage_5__3641_, data_stage_5__3640_, data_stage_5__3639_, data_stage_5__3638_, data_stage_5__3637_, data_stage_5__3636_, data_stage_5__3635_, data_stage_5__3634_, data_stage_5__3633_, data_stage_5__3632_, data_stage_5__3631_, data_stage_5__3630_, data_stage_5__3629_, data_stage_5__3628_, data_stage_5__3627_, data_stage_5__3626_, data_stage_5__3625_, data_stage_5__3624_, data_stage_5__3623_, data_stage_5__3622_, data_stage_5__3621_, data_stage_5__3620_, data_stage_5__3619_, data_stage_5__3618_, data_stage_5__3617_, data_stage_5__3616_, data_stage_5__3615_, data_stage_5__3614_, data_stage_5__3613_, data_stage_5__3612_, data_stage_5__3611_, data_stage_5__3610_, data_stage_5__3609_, data_stage_5__3608_, data_stage_5__3607_, data_stage_5__3606_, data_stage_5__3605_, data_stage_5__3604_, data_stage_5__3603_, data_stage_5__3602_, data_stage_5__3601_, data_stage_5__3600_, data_stage_5__3599_, data_stage_5__3598_, data_stage_5__3597_, data_stage_5__3596_, data_stage_5__3595_, data_stage_5__3594_, data_stage_5__3593_, data_stage_5__3592_, data_stage_5__3591_, data_stage_5__3590_, data_stage_5__3589_, data_stage_5__3588_, data_stage_5__3587_, data_stage_5__3586_, data_stage_5__3585_, data_stage_5__3584_, data_stage_5__3583_, data_stage_5__3582_, data_stage_5__3581_, data_stage_5__3580_, data_stage_5__3579_, data_stage_5__3578_, data_stage_5__3577_, data_stage_5__3576_, data_stage_5__3575_, data_stage_5__3574_, data_stage_5__3573_, data_stage_5__3572_, data_stage_5__3571_, data_stage_5__3570_, data_stage_5__3569_, data_stage_5__3568_, data_stage_5__3567_, data_stage_5__3566_, data_stage_5__3565_, data_stage_5__3564_, data_stage_5__3563_, data_stage_5__3562_, data_stage_5__3561_, data_stage_5__3560_, data_stage_5__3559_, data_stage_5__3558_, data_stage_5__3557_, data_stage_5__3556_, data_stage_5__3555_, data_stage_5__3554_, data_stage_5__3553_, data_stage_5__3552_, data_stage_5__3551_, data_stage_5__3550_, data_stage_5__3549_, data_stage_5__3548_, data_stage_5__3547_, data_stage_5__3546_, data_stage_5__3545_, data_stage_5__3544_, data_stage_5__3543_, data_stage_5__3542_, data_stage_5__3541_, data_stage_5__3540_, data_stage_5__3539_, data_stage_5__3538_, data_stage_5__3537_, data_stage_5__3536_, data_stage_5__3535_, data_stage_5__3534_, data_stage_5__3533_, data_stage_5__3532_, data_stage_5__3531_, data_stage_5__3530_, data_stage_5__3529_, data_stage_5__3528_, data_stage_5__3527_, data_stage_5__3526_, data_stage_5__3525_, data_stage_5__3524_, data_stage_5__3523_, data_stage_5__3522_, data_stage_5__3521_, data_stage_5__3520_, data_stage_5__3519_, data_stage_5__3518_, data_stage_5__3517_, data_stage_5__3516_, data_stage_5__3515_, data_stage_5__3514_, data_stage_5__3513_, data_stage_5__3512_, data_stage_5__3511_, data_stage_5__3510_, data_stage_5__3509_, data_stage_5__3508_, data_stage_5__3507_, data_stage_5__3506_, data_stage_5__3505_, data_stage_5__3504_, data_stage_5__3503_, data_stage_5__3502_, data_stage_5__3501_, data_stage_5__3500_, data_stage_5__3499_, data_stage_5__3498_, data_stage_5__3497_, data_stage_5__3496_, data_stage_5__3495_, data_stage_5__3494_, data_stage_5__3493_, data_stage_5__3492_, data_stage_5__3491_, data_stage_5__3490_, data_stage_5__3489_, data_stage_5__3488_, data_stage_5__3487_, data_stage_5__3486_, data_stage_5__3485_, data_stage_5__3484_, data_stage_5__3483_, data_stage_5__3482_, data_stage_5__3481_, data_stage_5__3480_, data_stage_5__3479_, data_stage_5__3478_, data_stage_5__3477_, data_stage_5__3476_, data_stage_5__3475_, data_stage_5__3474_, data_stage_5__3473_, data_stage_5__3472_, data_stage_5__3471_, data_stage_5__3470_, data_stage_5__3469_, data_stage_5__3468_, data_stage_5__3467_, data_stage_5__3466_, data_stage_5__3465_, data_stage_5__3464_, data_stage_5__3463_, data_stage_5__3462_, data_stage_5__3461_, data_stage_5__3460_, data_stage_5__3459_, data_stage_5__3458_, data_stage_5__3457_, data_stage_5__3456_, data_stage_5__3455_, data_stage_5__3454_, data_stage_5__3453_, data_stage_5__3452_, data_stage_5__3451_, data_stage_5__3450_, data_stage_5__3449_, data_stage_5__3448_, data_stage_5__3447_, data_stage_5__3446_, data_stage_5__3445_, data_stage_5__3444_, data_stage_5__3443_, data_stage_5__3442_, data_stage_5__3441_, data_stage_5__3440_, data_stage_5__3439_, data_stage_5__3438_, data_stage_5__3437_, data_stage_5__3436_, data_stage_5__3435_, data_stage_5__3434_, data_stage_5__3433_, data_stage_5__3432_, data_stage_5__3431_, data_stage_5__3430_, data_stage_5__3429_, data_stage_5__3428_, data_stage_5__3427_, data_stage_5__3426_, data_stage_5__3425_, data_stage_5__3424_, data_stage_5__3423_, data_stage_5__3422_, data_stage_5__3421_, data_stage_5__3420_, data_stage_5__3419_, data_stage_5__3418_, data_stage_5__3417_, data_stage_5__3416_, data_stage_5__3415_, data_stage_5__3414_, data_stage_5__3413_, data_stage_5__3412_, data_stage_5__3411_, data_stage_5__3410_, data_stage_5__3409_, data_stage_5__3408_, data_stage_5__3407_, data_stage_5__3406_, data_stage_5__3405_, data_stage_5__3404_, data_stage_5__3403_, data_stage_5__3402_, data_stage_5__3401_, data_stage_5__3400_, data_stage_5__3399_, data_stage_5__3398_, data_stage_5__3397_, data_stage_5__3396_, data_stage_5__3395_, data_stage_5__3394_, data_stage_5__3393_, data_stage_5__3392_, data_stage_5__3391_, data_stage_5__3390_, data_stage_5__3389_, data_stage_5__3388_, data_stage_5__3387_, data_stage_5__3386_, data_stage_5__3385_, data_stage_5__3384_, data_stage_5__3383_, data_stage_5__3382_, data_stage_5__3381_, data_stage_5__3380_, data_stage_5__3379_, data_stage_5__3378_, data_stage_5__3377_, data_stage_5__3376_, data_stage_5__3375_, data_stage_5__3374_, data_stage_5__3373_, data_stage_5__3372_, data_stage_5__3371_, data_stage_5__3370_, data_stage_5__3369_, data_stage_5__3368_, data_stage_5__3367_, data_stage_5__3366_, data_stage_5__3365_, data_stage_5__3364_, data_stage_5__3363_, data_stage_5__3362_, data_stage_5__3361_, data_stage_5__3360_, data_stage_5__3359_, data_stage_5__3358_, data_stage_5__3357_, data_stage_5__3356_, data_stage_5__3355_, data_stage_5__3354_, data_stage_5__3353_, data_stage_5__3352_, data_stage_5__3351_, data_stage_5__3350_, data_stage_5__3349_, data_stage_5__3348_, data_stage_5__3347_, data_stage_5__3346_, data_stage_5__3345_, data_stage_5__3344_, data_stage_5__3343_, data_stage_5__3342_, data_stage_5__3341_, data_stage_5__3340_, data_stage_5__3339_, data_stage_5__3338_, data_stage_5__3337_, data_stage_5__3336_, data_stage_5__3335_, data_stage_5__3334_, data_stage_5__3333_, data_stage_5__3332_, data_stage_5__3331_, data_stage_5__3330_, data_stage_5__3329_, data_stage_5__3328_, data_stage_5__3327_, data_stage_5__3326_, data_stage_5__3325_, data_stage_5__3324_, data_stage_5__3323_, data_stage_5__3322_, data_stage_5__3321_, data_stage_5__3320_, data_stage_5__3319_, data_stage_5__3318_, data_stage_5__3317_, data_stage_5__3316_, data_stage_5__3315_, data_stage_5__3314_, data_stage_5__3313_, data_stage_5__3312_, data_stage_5__3311_, data_stage_5__3310_, data_stage_5__3309_, data_stage_5__3308_, data_stage_5__3307_, data_stage_5__3306_, data_stage_5__3305_, data_stage_5__3304_, data_stage_5__3303_, data_stage_5__3302_, data_stage_5__3301_, data_stage_5__3300_, data_stage_5__3299_, data_stage_5__3298_, data_stage_5__3297_, data_stage_5__3296_, data_stage_5__3295_, data_stage_5__3294_, data_stage_5__3293_, data_stage_5__3292_, data_stage_5__3291_, data_stage_5__3290_, data_stage_5__3289_, data_stage_5__3288_, data_stage_5__3287_, data_stage_5__3286_, data_stage_5__3285_, data_stage_5__3284_, data_stage_5__3283_, data_stage_5__3282_, data_stage_5__3281_, data_stage_5__3280_, data_stage_5__3279_, data_stage_5__3278_, data_stage_5__3277_, data_stage_5__3276_, data_stage_5__3275_, data_stage_5__3274_, data_stage_5__3273_, data_stage_5__3272_, data_stage_5__3271_, data_stage_5__3270_, data_stage_5__3269_, data_stage_5__3268_, data_stage_5__3267_, data_stage_5__3266_, data_stage_5__3265_, data_stage_5__3264_, data_stage_5__3263_, data_stage_5__3262_, data_stage_5__3261_, data_stage_5__3260_, data_stage_5__3259_, data_stage_5__3258_, data_stage_5__3257_, data_stage_5__3256_, data_stage_5__3255_, data_stage_5__3254_, data_stage_5__3253_, data_stage_5__3252_, data_stage_5__3251_, data_stage_5__3250_, data_stage_5__3249_, data_stage_5__3248_, data_stage_5__3247_, data_stage_5__3246_, data_stage_5__3245_, data_stage_5__3244_, data_stage_5__3243_, data_stage_5__3242_, data_stage_5__3241_, data_stage_5__3240_, data_stage_5__3239_, data_stage_5__3238_, data_stage_5__3237_, data_stage_5__3236_, data_stage_5__3235_, data_stage_5__3234_, data_stage_5__3233_, data_stage_5__3232_, data_stage_5__3231_, data_stage_5__3230_, data_stage_5__3229_, data_stage_5__3228_, data_stage_5__3227_, data_stage_5__3226_, data_stage_5__3225_, data_stage_5__3224_, data_stage_5__3223_, data_stage_5__3222_, data_stage_5__3221_, data_stage_5__3220_, data_stage_5__3219_, data_stage_5__3218_, data_stage_5__3217_, data_stage_5__3216_, data_stage_5__3215_, data_stage_5__3214_, data_stage_5__3213_, data_stage_5__3212_, data_stage_5__3211_, data_stage_5__3210_, data_stage_5__3209_, data_stage_5__3208_, data_stage_5__3207_, data_stage_5__3206_, data_stage_5__3205_, data_stage_5__3204_, data_stage_5__3203_, data_stage_5__3202_, data_stage_5__3201_, data_stage_5__3200_, data_stage_5__3199_, data_stage_5__3198_, data_stage_5__3197_, data_stage_5__3196_, data_stage_5__3195_, data_stage_5__3194_, data_stage_5__3193_, data_stage_5__3192_, data_stage_5__3191_, data_stage_5__3190_, data_stage_5__3189_, data_stage_5__3188_, data_stage_5__3187_, data_stage_5__3186_, data_stage_5__3185_, data_stage_5__3184_, data_stage_5__3183_, data_stage_5__3182_, data_stage_5__3181_, data_stage_5__3180_, data_stage_5__3179_, data_stage_5__3178_, data_stage_5__3177_, data_stage_5__3176_, data_stage_5__3175_, data_stage_5__3174_, data_stage_5__3173_, data_stage_5__3172_, data_stage_5__3171_, data_stage_5__3170_, data_stage_5__3169_, data_stage_5__3168_, data_stage_5__3167_, data_stage_5__3166_, data_stage_5__3165_, data_stage_5__3164_, data_stage_5__3163_, data_stage_5__3162_, data_stage_5__3161_, data_stage_5__3160_, data_stage_5__3159_, data_stage_5__3158_, data_stage_5__3157_, data_stage_5__3156_, data_stage_5__3155_, data_stage_5__3154_, data_stage_5__3153_, data_stage_5__3152_, data_stage_5__3151_, data_stage_5__3150_, data_stage_5__3149_, data_stage_5__3148_, data_stage_5__3147_, data_stage_5__3146_, data_stage_5__3145_, data_stage_5__3144_, data_stage_5__3143_, data_stage_5__3142_, data_stage_5__3141_, data_stage_5__3140_, data_stage_5__3139_, data_stage_5__3138_, data_stage_5__3137_, data_stage_5__3136_, data_stage_5__3135_, data_stage_5__3134_, data_stage_5__3133_, data_stage_5__3132_, data_stage_5__3131_, data_stage_5__3130_, data_stage_5__3129_, data_stage_5__3128_, data_stage_5__3127_, data_stage_5__3126_, data_stage_5__3125_, data_stage_5__3124_, data_stage_5__3123_, data_stage_5__3122_, data_stage_5__3121_, data_stage_5__3120_, data_stage_5__3119_, data_stage_5__3118_, data_stage_5__3117_, data_stage_5__3116_, data_stage_5__3115_, data_stage_5__3114_, data_stage_5__3113_, data_stage_5__3112_, data_stage_5__3111_, data_stage_5__3110_, data_stage_5__3109_, data_stage_5__3108_, data_stage_5__3107_, data_stage_5__3106_, data_stage_5__3105_, data_stage_5__3104_, data_stage_5__3103_, data_stage_5__3102_, data_stage_5__3101_, data_stage_5__3100_, data_stage_5__3099_, data_stage_5__3098_, data_stage_5__3097_, data_stage_5__3096_, data_stage_5__3095_, data_stage_5__3094_, data_stage_5__3093_, data_stage_5__3092_, data_stage_5__3091_, data_stage_5__3090_, data_stage_5__3089_, data_stage_5__3088_, data_stage_5__3087_, data_stage_5__3086_, data_stage_5__3085_, data_stage_5__3084_, data_stage_5__3083_, data_stage_5__3082_, data_stage_5__3081_, data_stage_5__3080_, data_stage_5__3079_, data_stage_5__3078_, data_stage_5__3077_, data_stage_5__3076_, data_stage_5__3075_, data_stage_5__3074_, data_stage_5__3073_, data_stage_5__3072_, data_stage_5__3071_, data_stage_5__3070_, data_stage_5__3069_, data_stage_5__3068_, data_stage_5__3067_, data_stage_5__3066_, data_stage_5__3065_, data_stage_5__3064_, data_stage_5__3063_, data_stage_5__3062_, data_stage_5__3061_, data_stage_5__3060_, data_stage_5__3059_, data_stage_5__3058_, data_stage_5__3057_, data_stage_5__3056_, data_stage_5__3055_, data_stage_5__3054_, data_stage_5__3053_, data_stage_5__3052_, data_stage_5__3051_, data_stage_5__3050_, data_stage_5__3049_, data_stage_5__3048_, data_stage_5__3047_, data_stage_5__3046_, data_stage_5__3045_, data_stage_5__3044_, data_stage_5__3043_, data_stage_5__3042_, data_stage_5__3041_, data_stage_5__3040_, data_stage_5__3039_, data_stage_5__3038_, data_stage_5__3037_, data_stage_5__3036_, data_stage_5__3035_, data_stage_5__3034_, data_stage_5__3033_, data_stage_5__3032_, data_stage_5__3031_, data_stage_5__3030_, data_stage_5__3029_, data_stage_5__3028_, data_stage_5__3027_, data_stage_5__3026_, data_stage_5__3025_, data_stage_5__3024_, data_stage_5__3023_, data_stage_5__3022_, data_stage_5__3021_, data_stage_5__3020_, data_stage_5__3019_, data_stage_5__3018_, data_stage_5__3017_, data_stage_5__3016_, data_stage_5__3015_, data_stage_5__3014_, data_stage_5__3013_, data_stage_5__3012_, data_stage_5__3011_, data_stage_5__3010_, data_stage_5__3009_, data_stage_5__3008_, data_stage_5__3007_, data_stage_5__3006_, data_stage_5__3005_, data_stage_5__3004_, data_stage_5__3003_, data_stage_5__3002_, data_stage_5__3001_, data_stage_5__3000_, data_stage_5__2999_, data_stage_5__2998_, data_stage_5__2997_, data_stage_5__2996_, data_stage_5__2995_, data_stage_5__2994_, data_stage_5__2993_, data_stage_5__2992_, data_stage_5__2991_, data_stage_5__2990_, data_stage_5__2989_, data_stage_5__2988_, data_stage_5__2987_, data_stage_5__2986_, data_stage_5__2985_, data_stage_5__2984_, data_stage_5__2983_, data_stage_5__2982_, data_stage_5__2981_, data_stage_5__2980_, data_stage_5__2979_, data_stage_5__2978_, data_stage_5__2977_, data_stage_5__2976_, data_stage_5__2975_, data_stage_5__2974_, data_stage_5__2973_, data_stage_5__2972_, data_stage_5__2971_, data_stage_5__2970_, data_stage_5__2969_, data_stage_5__2968_, data_stage_5__2967_, data_stage_5__2966_, data_stage_5__2965_, data_stage_5__2964_, data_stage_5__2963_, data_stage_5__2962_, data_stage_5__2961_, data_stage_5__2960_, data_stage_5__2959_, data_stage_5__2958_, data_stage_5__2957_, data_stage_5__2956_, data_stage_5__2955_, data_stage_5__2954_, data_stage_5__2953_, data_stage_5__2952_, data_stage_5__2951_, data_stage_5__2950_, data_stage_5__2949_, data_stage_5__2948_, data_stage_5__2947_, data_stage_5__2946_, data_stage_5__2945_, data_stage_5__2944_, data_stage_5__2943_, data_stage_5__2942_, data_stage_5__2941_, data_stage_5__2940_, data_stage_5__2939_, data_stage_5__2938_, data_stage_5__2937_, data_stage_5__2936_, data_stage_5__2935_, data_stage_5__2934_, data_stage_5__2933_, data_stage_5__2932_, data_stage_5__2931_, data_stage_5__2930_, data_stage_5__2929_, data_stage_5__2928_, data_stage_5__2927_, data_stage_5__2926_, data_stage_5__2925_, data_stage_5__2924_, data_stage_5__2923_, data_stage_5__2922_, data_stage_5__2921_, data_stage_5__2920_, data_stage_5__2919_, data_stage_5__2918_, data_stage_5__2917_, data_stage_5__2916_, data_stage_5__2915_, data_stage_5__2914_, data_stage_5__2913_, data_stage_5__2912_, data_stage_5__2911_, data_stage_5__2910_, data_stage_5__2909_, data_stage_5__2908_, data_stage_5__2907_, data_stage_5__2906_, data_stage_5__2905_, data_stage_5__2904_, data_stage_5__2903_, data_stage_5__2902_, data_stage_5__2901_, data_stage_5__2900_, data_stage_5__2899_, data_stage_5__2898_, data_stage_5__2897_, data_stage_5__2896_, data_stage_5__2895_, data_stage_5__2894_, data_stage_5__2893_, data_stage_5__2892_, data_stage_5__2891_, data_stage_5__2890_, data_stage_5__2889_, data_stage_5__2888_, data_stage_5__2887_, data_stage_5__2886_, data_stage_5__2885_, data_stage_5__2884_, data_stage_5__2883_, data_stage_5__2882_, data_stage_5__2881_, data_stage_5__2880_, data_stage_5__2879_, data_stage_5__2878_, data_stage_5__2877_, data_stage_5__2876_, data_stage_5__2875_, data_stage_5__2874_, data_stage_5__2873_, data_stage_5__2872_, data_stage_5__2871_, data_stage_5__2870_, data_stage_5__2869_, data_stage_5__2868_, data_stage_5__2867_, data_stage_5__2866_, data_stage_5__2865_, data_stage_5__2864_, data_stage_5__2863_, data_stage_5__2862_, data_stage_5__2861_, data_stage_5__2860_, data_stage_5__2859_, data_stage_5__2858_, data_stage_5__2857_, data_stage_5__2856_, data_stage_5__2855_, data_stage_5__2854_, data_stage_5__2853_, data_stage_5__2852_, data_stage_5__2851_, data_stage_5__2850_, data_stage_5__2849_, data_stage_5__2848_, data_stage_5__2847_, data_stage_5__2846_, data_stage_5__2845_, data_stage_5__2844_, data_stage_5__2843_, data_stage_5__2842_, data_stage_5__2841_, data_stage_5__2840_, data_stage_5__2839_, data_stage_5__2838_, data_stage_5__2837_, data_stage_5__2836_, data_stage_5__2835_, data_stage_5__2834_, data_stage_5__2833_, data_stage_5__2832_, data_stage_5__2831_, data_stage_5__2830_, data_stage_5__2829_, data_stage_5__2828_, data_stage_5__2827_, data_stage_5__2826_, data_stage_5__2825_, data_stage_5__2824_, data_stage_5__2823_, data_stage_5__2822_, data_stage_5__2821_, data_stage_5__2820_, data_stage_5__2819_, data_stage_5__2818_, data_stage_5__2817_, data_stage_5__2816_, data_stage_5__2815_, data_stage_5__2814_, data_stage_5__2813_, data_stage_5__2812_, data_stage_5__2811_, data_stage_5__2810_, data_stage_5__2809_, data_stage_5__2808_, data_stage_5__2807_, data_stage_5__2806_, data_stage_5__2805_, data_stage_5__2804_, data_stage_5__2803_, data_stage_5__2802_, data_stage_5__2801_, data_stage_5__2800_, data_stage_5__2799_, data_stage_5__2798_, data_stage_5__2797_, data_stage_5__2796_, data_stage_5__2795_, data_stage_5__2794_, data_stage_5__2793_, data_stage_5__2792_, data_stage_5__2791_, data_stage_5__2790_, data_stage_5__2789_, data_stage_5__2788_, data_stage_5__2787_, data_stage_5__2786_, data_stage_5__2785_, data_stage_5__2784_, data_stage_5__2783_, data_stage_5__2782_, data_stage_5__2781_, data_stage_5__2780_, data_stage_5__2779_, data_stage_5__2778_, data_stage_5__2777_, data_stage_5__2776_, data_stage_5__2775_, data_stage_5__2774_, data_stage_5__2773_, data_stage_5__2772_, data_stage_5__2771_, data_stage_5__2770_, data_stage_5__2769_, data_stage_5__2768_, data_stage_5__2767_, data_stage_5__2766_, data_stage_5__2765_, data_stage_5__2764_, data_stage_5__2763_, data_stage_5__2762_, data_stage_5__2761_, data_stage_5__2760_, data_stage_5__2759_, data_stage_5__2758_, data_stage_5__2757_, data_stage_5__2756_, data_stage_5__2755_, data_stage_5__2754_, data_stage_5__2753_, data_stage_5__2752_, data_stage_5__2751_, data_stage_5__2750_, data_stage_5__2749_, data_stage_5__2748_, data_stage_5__2747_, data_stage_5__2746_, data_stage_5__2745_, data_stage_5__2744_, data_stage_5__2743_, data_stage_5__2742_, data_stage_5__2741_, data_stage_5__2740_, data_stage_5__2739_, data_stage_5__2738_, data_stage_5__2737_, data_stage_5__2736_, data_stage_5__2735_, data_stage_5__2734_, data_stage_5__2733_, data_stage_5__2732_, data_stage_5__2731_, data_stage_5__2730_, data_stage_5__2729_, data_stage_5__2728_, data_stage_5__2727_, data_stage_5__2726_, data_stage_5__2725_, data_stage_5__2724_, data_stage_5__2723_, data_stage_5__2722_, data_stage_5__2721_, data_stage_5__2720_, data_stage_5__2719_, data_stage_5__2718_, data_stage_5__2717_, data_stage_5__2716_, data_stage_5__2715_, data_stage_5__2714_, data_stage_5__2713_, data_stage_5__2712_, data_stage_5__2711_, data_stage_5__2710_, data_stage_5__2709_, data_stage_5__2708_, data_stage_5__2707_, data_stage_5__2706_, data_stage_5__2705_, data_stage_5__2704_, data_stage_5__2703_, data_stage_5__2702_, data_stage_5__2701_, data_stage_5__2700_, data_stage_5__2699_, data_stage_5__2698_, data_stage_5__2697_, data_stage_5__2696_, data_stage_5__2695_, data_stage_5__2694_, data_stage_5__2693_, data_stage_5__2692_, data_stage_5__2691_, data_stage_5__2690_, data_stage_5__2689_, data_stage_5__2688_, data_stage_5__2687_, data_stage_5__2686_, data_stage_5__2685_, data_stage_5__2684_, data_stage_5__2683_, data_stage_5__2682_, data_stage_5__2681_, data_stage_5__2680_, data_stage_5__2679_, data_stage_5__2678_, data_stage_5__2677_, data_stage_5__2676_, data_stage_5__2675_, data_stage_5__2674_, data_stage_5__2673_, data_stage_5__2672_, data_stage_5__2671_, data_stage_5__2670_, data_stage_5__2669_, data_stage_5__2668_, data_stage_5__2667_, data_stage_5__2666_, data_stage_5__2665_, data_stage_5__2664_, data_stage_5__2663_, data_stage_5__2662_, data_stage_5__2661_, data_stage_5__2660_, data_stage_5__2659_, data_stage_5__2658_, data_stage_5__2657_, data_stage_5__2656_, data_stage_5__2655_, data_stage_5__2654_, data_stage_5__2653_, data_stage_5__2652_, data_stage_5__2651_, data_stage_5__2650_, data_stage_5__2649_, data_stage_5__2648_, data_stage_5__2647_, data_stage_5__2646_, data_stage_5__2645_, data_stage_5__2644_, data_stage_5__2643_, data_stage_5__2642_, data_stage_5__2641_, data_stage_5__2640_, data_stage_5__2639_, data_stage_5__2638_, data_stage_5__2637_, data_stage_5__2636_, data_stage_5__2635_, data_stage_5__2634_, data_stage_5__2633_, data_stage_5__2632_, data_stage_5__2631_, data_stage_5__2630_, data_stage_5__2629_, data_stage_5__2628_, data_stage_5__2627_, data_stage_5__2626_, data_stage_5__2625_, data_stage_5__2624_, data_stage_5__2623_, data_stage_5__2622_, data_stage_5__2621_, data_stage_5__2620_, data_stage_5__2619_, data_stage_5__2618_, data_stage_5__2617_, data_stage_5__2616_, data_stage_5__2615_, data_stage_5__2614_, data_stage_5__2613_, data_stage_5__2612_, data_stage_5__2611_, data_stage_5__2610_, data_stage_5__2609_, data_stage_5__2608_, data_stage_5__2607_, data_stage_5__2606_, data_stage_5__2605_, data_stage_5__2604_, data_stage_5__2603_, data_stage_5__2602_, data_stage_5__2601_, data_stage_5__2600_, data_stage_5__2599_, data_stage_5__2598_, data_stage_5__2597_, data_stage_5__2596_, data_stage_5__2595_, data_stage_5__2594_, data_stage_5__2593_, data_stage_5__2592_, data_stage_5__2591_, data_stage_5__2590_, data_stage_5__2589_, data_stage_5__2588_, data_stage_5__2587_, data_stage_5__2586_, data_stage_5__2585_, data_stage_5__2584_, data_stage_5__2583_, data_stage_5__2582_, data_stage_5__2581_, data_stage_5__2580_, data_stage_5__2579_, data_stage_5__2578_, data_stage_5__2577_, data_stage_5__2576_, data_stage_5__2575_, data_stage_5__2574_, data_stage_5__2573_, data_stage_5__2572_, data_stage_5__2571_, data_stage_5__2570_, data_stage_5__2569_, data_stage_5__2568_, data_stage_5__2567_, data_stage_5__2566_, data_stage_5__2565_, data_stage_5__2564_, data_stage_5__2563_, data_stage_5__2562_, data_stage_5__2561_, data_stage_5__2560_, data_stage_5__2559_, data_stage_5__2558_, data_stage_5__2557_, data_stage_5__2556_, data_stage_5__2555_, data_stage_5__2554_, data_stage_5__2553_, data_stage_5__2552_, data_stage_5__2551_, data_stage_5__2550_, data_stage_5__2549_, data_stage_5__2548_, data_stage_5__2547_, data_stage_5__2546_, data_stage_5__2545_, data_stage_5__2544_, data_stage_5__2543_, data_stage_5__2542_, data_stage_5__2541_, data_stage_5__2540_, data_stage_5__2539_, data_stage_5__2538_, data_stage_5__2537_, data_stage_5__2536_, data_stage_5__2535_, data_stage_5__2534_, data_stage_5__2533_, data_stage_5__2532_, data_stage_5__2531_, data_stage_5__2530_, data_stage_5__2529_, data_stage_5__2528_, data_stage_5__2527_, data_stage_5__2526_, data_stage_5__2525_, data_stage_5__2524_, data_stage_5__2523_, data_stage_5__2522_, data_stage_5__2521_, data_stage_5__2520_, data_stage_5__2519_, data_stage_5__2518_, data_stage_5__2517_, data_stage_5__2516_, data_stage_5__2515_, data_stage_5__2514_, data_stage_5__2513_, data_stage_5__2512_, data_stage_5__2511_, data_stage_5__2510_, data_stage_5__2509_, data_stage_5__2508_, data_stage_5__2507_, data_stage_5__2506_, data_stage_5__2505_, data_stage_5__2504_, data_stage_5__2503_, data_stage_5__2502_, data_stage_5__2501_, data_stage_5__2500_, data_stage_5__2499_, data_stage_5__2498_, data_stage_5__2497_, data_stage_5__2496_, data_stage_5__2495_, data_stage_5__2494_, data_stage_5__2493_, data_stage_5__2492_, data_stage_5__2491_, data_stage_5__2490_, data_stage_5__2489_, data_stage_5__2488_, data_stage_5__2487_, data_stage_5__2486_, data_stage_5__2485_, data_stage_5__2484_, data_stage_5__2483_, data_stage_5__2482_, data_stage_5__2481_, data_stage_5__2480_, data_stage_5__2479_, data_stage_5__2478_, data_stage_5__2477_, data_stage_5__2476_, data_stage_5__2475_, data_stage_5__2474_, data_stage_5__2473_, data_stage_5__2472_, data_stage_5__2471_, data_stage_5__2470_, data_stage_5__2469_, data_stage_5__2468_, data_stage_5__2467_, data_stage_5__2466_, data_stage_5__2465_, data_stage_5__2464_, data_stage_5__2463_, data_stage_5__2462_, data_stage_5__2461_, data_stage_5__2460_, data_stage_5__2459_, data_stage_5__2458_, data_stage_5__2457_, data_stage_5__2456_, data_stage_5__2455_, data_stage_5__2454_, data_stage_5__2453_, data_stage_5__2452_, data_stage_5__2451_, data_stage_5__2450_, data_stage_5__2449_, data_stage_5__2448_, data_stage_5__2447_, data_stage_5__2446_, data_stage_5__2445_, data_stage_5__2444_, data_stage_5__2443_, data_stage_5__2442_, data_stage_5__2441_, data_stage_5__2440_, data_stage_5__2439_, data_stage_5__2438_, data_stage_5__2437_, data_stage_5__2436_, data_stage_5__2435_, data_stage_5__2434_, data_stage_5__2433_, data_stage_5__2432_, data_stage_5__2431_, data_stage_5__2430_, data_stage_5__2429_, data_stage_5__2428_, data_stage_5__2427_, data_stage_5__2426_, data_stage_5__2425_, data_stage_5__2424_, data_stage_5__2423_, data_stage_5__2422_, data_stage_5__2421_, data_stage_5__2420_, data_stage_5__2419_, data_stage_5__2418_, data_stage_5__2417_, data_stage_5__2416_, data_stage_5__2415_, data_stage_5__2414_, data_stage_5__2413_, data_stage_5__2412_, data_stage_5__2411_, data_stage_5__2410_, data_stage_5__2409_, data_stage_5__2408_, data_stage_5__2407_, data_stage_5__2406_, data_stage_5__2405_, data_stage_5__2404_, data_stage_5__2403_, data_stage_5__2402_, data_stage_5__2401_, data_stage_5__2400_, data_stage_5__2399_, data_stage_5__2398_, data_stage_5__2397_, data_stage_5__2396_, data_stage_5__2395_, data_stage_5__2394_, data_stage_5__2393_, data_stage_5__2392_, data_stage_5__2391_, data_stage_5__2390_, data_stage_5__2389_, data_stage_5__2388_, data_stage_5__2387_, data_stage_5__2386_, data_stage_5__2385_, data_stage_5__2384_, data_stage_5__2383_, data_stage_5__2382_, data_stage_5__2381_, data_stage_5__2380_, data_stage_5__2379_, data_stage_5__2378_, data_stage_5__2377_, data_stage_5__2376_, data_stage_5__2375_, data_stage_5__2374_, data_stage_5__2373_, data_stage_5__2372_, data_stage_5__2371_, data_stage_5__2370_, data_stage_5__2369_, data_stage_5__2368_, data_stage_5__2367_, data_stage_5__2366_, data_stage_5__2365_, data_stage_5__2364_, data_stage_5__2363_, data_stage_5__2362_, data_stage_5__2361_, data_stage_5__2360_, data_stage_5__2359_, data_stage_5__2358_, data_stage_5__2357_, data_stage_5__2356_, data_stage_5__2355_, data_stage_5__2354_, data_stage_5__2353_, data_stage_5__2352_, data_stage_5__2351_, data_stage_5__2350_, data_stage_5__2349_, data_stage_5__2348_, data_stage_5__2347_, data_stage_5__2346_, data_stage_5__2345_, data_stage_5__2344_, data_stage_5__2343_, data_stage_5__2342_, data_stage_5__2341_, data_stage_5__2340_, data_stage_5__2339_, data_stage_5__2338_, data_stage_5__2337_, data_stage_5__2336_, data_stage_5__2335_, data_stage_5__2334_, data_stage_5__2333_, data_stage_5__2332_, data_stage_5__2331_, data_stage_5__2330_, data_stage_5__2329_, data_stage_5__2328_, data_stage_5__2327_, data_stage_5__2326_, data_stage_5__2325_, data_stage_5__2324_, data_stage_5__2323_, data_stage_5__2322_, data_stage_5__2321_, data_stage_5__2320_, data_stage_5__2319_, data_stage_5__2318_, data_stage_5__2317_, data_stage_5__2316_, data_stage_5__2315_, data_stage_5__2314_, data_stage_5__2313_, data_stage_5__2312_, data_stage_5__2311_, data_stage_5__2310_, data_stage_5__2309_, data_stage_5__2308_, data_stage_5__2307_, data_stage_5__2306_, data_stage_5__2305_, data_stage_5__2304_, data_stage_5__2303_, data_stage_5__2302_, data_stage_5__2301_, data_stage_5__2300_, data_stage_5__2299_, data_stage_5__2298_, data_stage_5__2297_, data_stage_5__2296_, data_stage_5__2295_, data_stage_5__2294_, data_stage_5__2293_, data_stage_5__2292_, data_stage_5__2291_, data_stage_5__2290_, data_stage_5__2289_, data_stage_5__2288_, data_stage_5__2287_, data_stage_5__2286_, data_stage_5__2285_, data_stage_5__2284_, data_stage_5__2283_, data_stage_5__2282_, data_stage_5__2281_, data_stage_5__2280_, data_stage_5__2279_, data_stage_5__2278_, data_stage_5__2277_, data_stage_5__2276_, data_stage_5__2275_, data_stage_5__2274_, data_stage_5__2273_, data_stage_5__2272_, data_stage_5__2271_, data_stage_5__2270_, data_stage_5__2269_, data_stage_5__2268_, data_stage_5__2267_, data_stage_5__2266_, data_stage_5__2265_, data_stage_5__2264_, data_stage_5__2263_, data_stage_5__2262_, data_stage_5__2261_, data_stage_5__2260_, data_stage_5__2259_, data_stage_5__2258_, data_stage_5__2257_, data_stage_5__2256_, data_stage_5__2255_, data_stage_5__2254_, data_stage_5__2253_, data_stage_5__2252_, data_stage_5__2251_, data_stage_5__2250_, data_stage_5__2249_, data_stage_5__2248_, data_stage_5__2247_, data_stage_5__2246_, data_stage_5__2245_, data_stage_5__2244_, data_stage_5__2243_, data_stage_5__2242_, data_stage_5__2241_, data_stage_5__2240_, data_stage_5__2239_, data_stage_5__2238_, data_stage_5__2237_, data_stage_5__2236_, data_stage_5__2235_, data_stage_5__2234_, data_stage_5__2233_, data_stage_5__2232_, data_stage_5__2231_, data_stage_5__2230_, data_stage_5__2229_, data_stage_5__2228_, data_stage_5__2227_, data_stage_5__2226_, data_stage_5__2225_, data_stage_5__2224_, data_stage_5__2223_, data_stage_5__2222_, data_stage_5__2221_, data_stage_5__2220_, data_stage_5__2219_, data_stage_5__2218_, data_stage_5__2217_, data_stage_5__2216_, data_stage_5__2215_, data_stage_5__2214_, data_stage_5__2213_, data_stage_5__2212_, data_stage_5__2211_, data_stage_5__2210_, data_stage_5__2209_, data_stage_5__2208_, data_stage_5__2207_, data_stage_5__2206_, data_stage_5__2205_, data_stage_5__2204_, data_stage_5__2203_, data_stage_5__2202_, data_stage_5__2201_, data_stage_5__2200_, data_stage_5__2199_, data_stage_5__2198_, data_stage_5__2197_, data_stage_5__2196_, data_stage_5__2195_, data_stage_5__2194_, data_stage_5__2193_, data_stage_5__2192_, data_stage_5__2191_, data_stage_5__2190_, data_stage_5__2189_, data_stage_5__2188_, data_stage_5__2187_, data_stage_5__2186_, data_stage_5__2185_, data_stage_5__2184_, data_stage_5__2183_, data_stage_5__2182_, data_stage_5__2181_, data_stage_5__2180_, data_stage_5__2179_, data_stage_5__2178_, data_stage_5__2177_, data_stage_5__2176_, data_stage_5__2175_, data_stage_5__2174_, data_stage_5__2173_, data_stage_5__2172_, data_stage_5__2171_, data_stage_5__2170_, data_stage_5__2169_, data_stage_5__2168_, data_stage_5__2167_, data_stage_5__2166_, data_stage_5__2165_, data_stage_5__2164_, data_stage_5__2163_, data_stage_5__2162_, data_stage_5__2161_, data_stage_5__2160_, data_stage_5__2159_, data_stage_5__2158_, data_stage_5__2157_, data_stage_5__2156_, data_stage_5__2155_, data_stage_5__2154_, data_stage_5__2153_, data_stage_5__2152_, data_stage_5__2151_, data_stage_5__2150_, data_stage_5__2149_, data_stage_5__2148_, data_stage_5__2147_, data_stage_5__2146_, data_stage_5__2145_, data_stage_5__2144_, data_stage_5__2143_, data_stage_5__2142_, data_stage_5__2141_, data_stage_5__2140_, data_stage_5__2139_, data_stage_5__2138_, data_stage_5__2137_, data_stage_5__2136_, data_stage_5__2135_, data_stage_5__2134_, data_stage_5__2133_, data_stage_5__2132_, data_stage_5__2131_, data_stage_5__2130_, data_stage_5__2129_, data_stage_5__2128_, data_stage_5__2127_, data_stage_5__2126_, data_stage_5__2125_, data_stage_5__2124_, data_stage_5__2123_, data_stage_5__2122_, data_stage_5__2121_, data_stage_5__2120_, data_stage_5__2119_, data_stage_5__2118_, data_stage_5__2117_, data_stage_5__2116_, data_stage_5__2115_, data_stage_5__2114_, data_stage_5__2113_, data_stage_5__2112_, data_stage_5__2111_, data_stage_5__2110_, data_stage_5__2109_, data_stage_5__2108_, data_stage_5__2107_, data_stage_5__2106_, data_stage_5__2105_, data_stage_5__2104_, data_stage_5__2103_, data_stage_5__2102_, data_stage_5__2101_, data_stage_5__2100_, data_stage_5__2099_, data_stage_5__2098_, data_stage_5__2097_, data_stage_5__2096_, data_stage_5__2095_, data_stage_5__2094_, data_stage_5__2093_, data_stage_5__2092_, data_stage_5__2091_, data_stage_5__2090_, data_stage_5__2089_, data_stage_5__2088_, data_stage_5__2087_, data_stage_5__2086_, data_stage_5__2085_, data_stage_5__2084_, data_stage_5__2083_, data_stage_5__2082_, data_stage_5__2081_, data_stage_5__2080_, data_stage_5__2079_, data_stage_5__2078_, data_stage_5__2077_, data_stage_5__2076_, data_stage_5__2075_, data_stage_5__2074_, data_stage_5__2073_, data_stage_5__2072_, data_stage_5__2071_, data_stage_5__2070_, data_stage_5__2069_, data_stage_5__2068_, data_stage_5__2067_, data_stage_5__2066_, data_stage_5__2065_, data_stage_5__2064_, data_stage_5__2063_, data_stage_5__2062_, data_stage_5__2061_, data_stage_5__2060_, data_stage_5__2059_, data_stage_5__2058_, data_stage_5__2057_, data_stage_5__2056_, data_stage_5__2055_, data_stage_5__2054_, data_stage_5__2053_, data_stage_5__2052_, data_stage_5__2051_, data_stage_5__2050_, data_stage_5__2049_, data_stage_5__2048_, data_stage_5__2047_, data_stage_5__2046_, data_stage_5__2045_, data_stage_5__2044_, data_stage_5__2043_, data_stage_5__2042_, data_stage_5__2041_, data_stage_5__2040_, data_stage_5__2039_, data_stage_5__2038_, data_stage_5__2037_, data_stage_5__2036_, data_stage_5__2035_, data_stage_5__2034_, data_stage_5__2033_, data_stage_5__2032_, data_stage_5__2031_, data_stage_5__2030_, data_stage_5__2029_, data_stage_5__2028_, data_stage_5__2027_, data_stage_5__2026_, data_stage_5__2025_, data_stage_5__2024_, data_stage_5__2023_, data_stage_5__2022_, data_stage_5__2021_, data_stage_5__2020_, data_stage_5__2019_, data_stage_5__2018_, data_stage_5__2017_, data_stage_5__2016_, data_stage_5__2015_, data_stage_5__2014_, data_stage_5__2013_, data_stage_5__2012_, data_stage_5__2011_, data_stage_5__2010_, data_stage_5__2009_, data_stage_5__2008_, data_stage_5__2007_, data_stage_5__2006_, data_stage_5__2005_, data_stage_5__2004_, data_stage_5__2003_, data_stage_5__2002_, data_stage_5__2001_, data_stage_5__2000_, data_stage_5__1999_, data_stage_5__1998_, data_stage_5__1997_, data_stage_5__1996_, data_stage_5__1995_, data_stage_5__1994_, data_stage_5__1993_, data_stage_5__1992_, data_stage_5__1991_, data_stage_5__1990_, data_stage_5__1989_, data_stage_5__1988_, data_stage_5__1987_, data_stage_5__1986_, data_stage_5__1985_, data_stage_5__1984_, data_stage_5__1983_, data_stage_5__1982_, data_stage_5__1981_, data_stage_5__1980_, data_stage_5__1979_, data_stage_5__1978_, data_stage_5__1977_, data_stage_5__1976_, data_stage_5__1975_, data_stage_5__1974_, data_stage_5__1973_, data_stage_5__1972_, data_stage_5__1971_, data_stage_5__1970_, data_stage_5__1969_, data_stage_5__1968_, data_stage_5__1967_, data_stage_5__1966_, data_stage_5__1965_, data_stage_5__1964_, data_stage_5__1963_, data_stage_5__1962_, data_stage_5__1961_, data_stage_5__1960_, data_stage_5__1959_, data_stage_5__1958_, data_stage_5__1957_, data_stage_5__1956_, data_stage_5__1955_, data_stage_5__1954_, data_stage_5__1953_, data_stage_5__1952_, data_stage_5__1951_, data_stage_5__1950_, data_stage_5__1949_, data_stage_5__1948_, data_stage_5__1947_, data_stage_5__1946_, data_stage_5__1945_, data_stage_5__1944_, data_stage_5__1943_, data_stage_5__1942_, data_stage_5__1941_, data_stage_5__1940_, data_stage_5__1939_, data_stage_5__1938_, data_stage_5__1937_, data_stage_5__1936_, data_stage_5__1935_, data_stage_5__1934_, data_stage_5__1933_, data_stage_5__1932_, data_stage_5__1931_, data_stage_5__1930_, data_stage_5__1929_, data_stage_5__1928_, data_stage_5__1927_, data_stage_5__1926_, data_stage_5__1925_, data_stage_5__1924_, data_stage_5__1923_, data_stage_5__1922_, data_stage_5__1921_, data_stage_5__1920_, data_stage_5__1919_, data_stage_5__1918_, data_stage_5__1917_, data_stage_5__1916_, data_stage_5__1915_, data_stage_5__1914_, data_stage_5__1913_, data_stage_5__1912_, data_stage_5__1911_, data_stage_5__1910_, data_stage_5__1909_, data_stage_5__1908_, data_stage_5__1907_, data_stage_5__1906_, data_stage_5__1905_, data_stage_5__1904_, data_stage_5__1903_, data_stage_5__1902_, data_stage_5__1901_, data_stage_5__1900_, data_stage_5__1899_, data_stage_5__1898_, data_stage_5__1897_, data_stage_5__1896_, data_stage_5__1895_, data_stage_5__1894_, data_stage_5__1893_, data_stage_5__1892_, data_stage_5__1891_, data_stage_5__1890_, data_stage_5__1889_, data_stage_5__1888_, data_stage_5__1887_, data_stage_5__1886_, data_stage_5__1885_, data_stage_5__1884_, data_stage_5__1883_, data_stage_5__1882_, data_stage_5__1881_, data_stage_5__1880_, data_stage_5__1879_, data_stage_5__1878_, data_stage_5__1877_, data_stage_5__1876_, data_stage_5__1875_, data_stage_5__1874_, data_stage_5__1873_, data_stage_5__1872_, data_stage_5__1871_, data_stage_5__1870_, data_stage_5__1869_, data_stage_5__1868_, data_stage_5__1867_, data_stage_5__1866_, data_stage_5__1865_, data_stage_5__1864_, data_stage_5__1863_, data_stage_5__1862_, data_stage_5__1861_, data_stage_5__1860_, data_stage_5__1859_, data_stage_5__1858_, data_stage_5__1857_, data_stage_5__1856_, data_stage_5__1855_, data_stage_5__1854_, data_stage_5__1853_, data_stage_5__1852_, data_stage_5__1851_, data_stage_5__1850_, data_stage_5__1849_, data_stage_5__1848_, data_stage_5__1847_, data_stage_5__1846_, data_stage_5__1845_, data_stage_5__1844_, data_stage_5__1843_, data_stage_5__1842_, data_stage_5__1841_, data_stage_5__1840_, data_stage_5__1839_, data_stage_5__1838_, data_stage_5__1837_, data_stage_5__1836_, data_stage_5__1835_, data_stage_5__1834_, data_stage_5__1833_, data_stage_5__1832_, data_stage_5__1831_, data_stage_5__1830_, data_stage_5__1829_, data_stage_5__1828_, data_stage_5__1827_, data_stage_5__1826_, data_stage_5__1825_, data_stage_5__1824_, data_stage_5__1823_, data_stage_5__1822_, data_stage_5__1821_, data_stage_5__1820_, data_stage_5__1819_, data_stage_5__1818_, data_stage_5__1817_, data_stage_5__1816_, data_stage_5__1815_, data_stage_5__1814_, data_stage_5__1813_, data_stage_5__1812_, data_stage_5__1811_, data_stage_5__1810_, data_stage_5__1809_, data_stage_5__1808_, data_stage_5__1807_, data_stage_5__1806_, data_stage_5__1805_, data_stage_5__1804_, data_stage_5__1803_, data_stage_5__1802_, data_stage_5__1801_, data_stage_5__1800_, data_stage_5__1799_, data_stage_5__1798_, data_stage_5__1797_, data_stage_5__1796_, data_stage_5__1795_, data_stage_5__1794_, data_stage_5__1793_, data_stage_5__1792_, data_stage_5__1791_, data_stage_5__1790_, data_stage_5__1789_, data_stage_5__1788_, data_stage_5__1787_, data_stage_5__1786_, data_stage_5__1785_, data_stage_5__1784_, data_stage_5__1783_, data_stage_5__1782_, data_stage_5__1781_, data_stage_5__1780_, data_stage_5__1779_, data_stage_5__1778_, data_stage_5__1777_, data_stage_5__1776_, data_stage_5__1775_, data_stage_5__1774_, data_stage_5__1773_, data_stage_5__1772_, data_stage_5__1771_, data_stage_5__1770_, data_stage_5__1769_, data_stage_5__1768_, data_stage_5__1767_, data_stage_5__1766_, data_stage_5__1765_, data_stage_5__1764_, data_stage_5__1763_, data_stage_5__1762_, data_stage_5__1761_, data_stage_5__1760_, data_stage_5__1759_, data_stage_5__1758_, data_stage_5__1757_, data_stage_5__1756_, data_stage_5__1755_, data_stage_5__1754_, data_stage_5__1753_, data_stage_5__1752_, data_stage_5__1751_, data_stage_5__1750_, data_stage_5__1749_, data_stage_5__1748_, data_stage_5__1747_, data_stage_5__1746_, data_stage_5__1745_, data_stage_5__1744_, data_stage_5__1743_, data_stage_5__1742_, data_stage_5__1741_, data_stage_5__1740_, data_stage_5__1739_, data_stage_5__1738_, data_stage_5__1737_, data_stage_5__1736_, data_stage_5__1735_, data_stage_5__1734_, data_stage_5__1733_, data_stage_5__1732_, data_stage_5__1731_, data_stage_5__1730_, data_stage_5__1729_, data_stage_5__1728_, data_stage_5__1727_, data_stage_5__1726_, data_stage_5__1725_, data_stage_5__1724_, data_stage_5__1723_, data_stage_5__1722_, data_stage_5__1721_, data_stage_5__1720_, data_stage_5__1719_, data_stage_5__1718_, data_stage_5__1717_, data_stage_5__1716_, data_stage_5__1715_, data_stage_5__1714_, data_stage_5__1713_, data_stage_5__1712_, data_stage_5__1711_, data_stage_5__1710_, data_stage_5__1709_, data_stage_5__1708_, data_stage_5__1707_, data_stage_5__1706_, data_stage_5__1705_, data_stage_5__1704_, data_stage_5__1703_, data_stage_5__1702_, data_stage_5__1701_, data_stage_5__1700_, data_stage_5__1699_, data_stage_5__1698_, data_stage_5__1697_, data_stage_5__1696_, data_stage_5__1695_, data_stage_5__1694_, data_stage_5__1693_, data_stage_5__1692_, data_stage_5__1691_, data_stage_5__1690_, data_stage_5__1689_, data_stage_5__1688_, data_stage_5__1687_, data_stage_5__1686_, data_stage_5__1685_, data_stage_5__1684_, data_stage_5__1683_, data_stage_5__1682_, data_stage_5__1681_, data_stage_5__1680_, data_stage_5__1679_, data_stage_5__1678_, data_stage_5__1677_, data_stage_5__1676_, data_stage_5__1675_, data_stage_5__1674_, data_stage_5__1673_, data_stage_5__1672_, data_stage_5__1671_, data_stage_5__1670_, data_stage_5__1669_, data_stage_5__1668_, data_stage_5__1667_, data_stage_5__1666_, data_stage_5__1665_, data_stage_5__1664_, data_stage_5__1663_, data_stage_5__1662_, data_stage_5__1661_, data_stage_5__1660_, data_stage_5__1659_, data_stage_5__1658_, data_stage_5__1657_, data_stage_5__1656_, data_stage_5__1655_, data_stage_5__1654_, data_stage_5__1653_, data_stage_5__1652_, data_stage_5__1651_, data_stage_5__1650_, data_stage_5__1649_, data_stage_5__1648_, data_stage_5__1647_, data_stage_5__1646_, data_stage_5__1645_, data_stage_5__1644_, data_stage_5__1643_, data_stage_5__1642_, data_stage_5__1641_, data_stage_5__1640_, data_stage_5__1639_, data_stage_5__1638_, data_stage_5__1637_, data_stage_5__1636_, data_stage_5__1635_, data_stage_5__1634_, data_stage_5__1633_, data_stage_5__1632_, data_stage_5__1631_, data_stage_5__1630_, data_stage_5__1629_, data_stage_5__1628_, data_stage_5__1627_, data_stage_5__1626_, data_stage_5__1625_, data_stage_5__1624_, data_stage_5__1623_, data_stage_5__1622_, data_stage_5__1621_, data_stage_5__1620_, data_stage_5__1619_, data_stage_5__1618_, data_stage_5__1617_, data_stage_5__1616_, data_stage_5__1615_, data_stage_5__1614_, data_stage_5__1613_, data_stage_5__1612_, data_stage_5__1611_, data_stage_5__1610_, data_stage_5__1609_, data_stage_5__1608_, data_stage_5__1607_, data_stage_5__1606_, data_stage_5__1605_, data_stage_5__1604_, data_stage_5__1603_, data_stage_5__1602_, data_stage_5__1601_, data_stage_5__1600_, data_stage_5__1599_, data_stage_5__1598_, data_stage_5__1597_, data_stage_5__1596_, data_stage_5__1595_, data_stage_5__1594_, data_stage_5__1593_, data_stage_5__1592_, data_stage_5__1591_, data_stage_5__1590_, data_stage_5__1589_, data_stage_5__1588_, data_stage_5__1587_, data_stage_5__1586_, data_stage_5__1585_, data_stage_5__1584_, data_stage_5__1583_, data_stage_5__1582_, data_stage_5__1581_, data_stage_5__1580_, data_stage_5__1579_, data_stage_5__1578_, data_stage_5__1577_, data_stage_5__1576_, data_stage_5__1575_, data_stage_5__1574_, data_stage_5__1573_, data_stage_5__1572_, data_stage_5__1571_, data_stage_5__1570_, data_stage_5__1569_, data_stage_5__1568_, data_stage_5__1567_, data_stage_5__1566_, data_stage_5__1565_, data_stage_5__1564_, data_stage_5__1563_, data_stage_5__1562_, data_stage_5__1561_, data_stage_5__1560_, data_stage_5__1559_, data_stage_5__1558_, data_stage_5__1557_, data_stage_5__1556_, data_stage_5__1555_, data_stage_5__1554_, data_stage_5__1553_, data_stage_5__1552_, data_stage_5__1551_, data_stage_5__1550_, data_stage_5__1549_, data_stage_5__1548_, data_stage_5__1547_, data_stage_5__1546_, data_stage_5__1545_, data_stage_5__1544_, data_stage_5__1543_, data_stage_5__1542_, data_stage_5__1541_, data_stage_5__1540_, data_stage_5__1539_, data_stage_5__1538_, data_stage_5__1537_, data_stage_5__1536_, data_stage_5__1535_, data_stage_5__1534_, data_stage_5__1533_, data_stage_5__1532_, data_stage_5__1531_, data_stage_5__1530_, data_stage_5__1529_, data_stage_5__1528_, data_stage_5__1527_, data_stage_5__1526_, data_stage_5__1525_, data_stage_5__1524_, data_stage_5__1523_, data_stage_5__1522_, data_stage_5__1521_, data_stage_5__1520_, data_stage_5__1519_, data_stage_5__1518_, data_stage_5__1517_, data_stage_5__1516_, data_stage_5__1515_, data_stage_5__1514_, data_stage_5__1513_, data_stage_5__1512_, data_stage_5__1511_, data_stage_5__1510_, data_stage_5__1509_, data_stage_5__1508_, data_stage_5__1507_, data_stage_5__1506_, data_stage_5__1505_, data_stage_5__1504_, data_stage_5__1503_, data_stage_5__1502_, data_stage_5__1501_, data_stage_5__1500_, data_stage_5__1499_, data_stage_5__1498_, data_stage_5__1497_, data_stage_5__1496_, data_stage_5__1495_, data_stage_5__1494_, data_stage_5__1493_, data_stage_5__1492_, data_stage_5__1491_, data_stage_5__1490_, data_stage_5__1489_, data_stage_5__1488_, data_stage_5__1487_, data_stage_5__1486_, data_stage_5__1485_, data_stage_5__1484_, data_stage_5__1483_, data_stage_5__1482_, data_stage_5__1481_, data_stage_5__1480_, data_stage_5__1479_, data_stage_5__1478_, data_stage_5__1477_, data_stage_5__1476_, data_stage_5__1475_, data_stage_5__1474_, data_stage_5__1473_, data_stage_5__1472_, data_stage_5__1471_, data_stage_5__1470_, data_stage_5__1469_, data_stage_5__1468_, data_stage_5__1467_, data_stage_5__1466_, data_stage_5__1465_, data_stage_5__1464_, data_stage_5__1463_, data_stage_5__1462_, data_stage_5__1461_, data_stage_5__1460_, data_stage_5__1459_, data_stage_5__1458_, data_stage_5__1457_, data_stage_5__1456_, data_stage_5__1455_, data_stage_5__1454_, data_stage_5__1453_, data_stage_5__1452_, data_stage_5__1451_, data_stage_5__1450_, data_stage_5__1449_, data_stage_5__1448_, data_stage_5__1447_, data_stage_5__1446_, data_stage_5__1445_, data_stage_5__1444_, data_stage_5__1443_, data_stage_5__1442_, data_stage_5__1441_, data_stage_5__1440_, data_stage_5__1439_, data_stage_5__1438_, data_stage_5__1437_, data_stage_5__1436_, data_stage_5__1435_, data_stage_5__1434_, data_stage_5__1433_, data_stage_5__1432_, data_stage_5__1431_, data_stage_5__1430_, data_stage_5__1429_, data_stage_5__1428_, data_stage_5__1427_, data_stage_5__1426_, data_stage_5__1425_, data_stage_5__1424_, data_stage_5__1423_, data_stage_5__1422_, data_stage_5__1421_, data_stage_5__1420_, data_stage_5__1419_, data_stage_5__1418_, data_stage_5__1417_, data_stage_5__1416_, data_stage_5__1415_, data_stage_5__1414_, data_stage_5__1413_, data_stage_5__1412_, data_stage_5__1411_, data_stage_5__1410_, data_stage_5__1409_, data_stage_5__1408_, data_stage_5__1407_, data_stage_5__1406_, data_stage_5__1405_, data_stage_5__1404_, data_stage_5__1403_, data_stage_5__1402_, data_stage_5__1401_, data_stage_5__1400_, data_stage_5__1399_, data_stage_5__1398_, data_stage_5__1397_, data_stage_5__1396_, data_stage_5__1395_, data_stage_5__1394_, data_stage_5__1393_, data_stage_5__1392_, data_stage_5__1391_, data_stage_5__1390_, data_stage_5__1389_, data_stage_5__1388_, data_stage_5__1387_, data_stage_5__1386_, data_stage_5__1385_, data_stage_5__1384_, data_stage_5__1383_, data_stage_5__1382_, data_stage_5__1381_, data_stage_5__1380_, data_stage_5__1379_, data_stage_5__1378_, data_stage_5__1377_, data_stage_5__1376_, data_stage_5__1375_, data_stage_5__1374_, data_stage_5__1373_, data_stage_5__1372_, data_stage_5__1371_, data_stage_5__1370_, data_stage_5__1369_, data_stage_5__1368_, data_stage_5__1367_, data_stage_5__1366_, data_stage_5__1365_, data_stage_5__1364_, data_stage_5__1363_, data_stage_5__1362_, data_stage_5__1361_, data_stage_5__1360_, data_stage_5__1359_, data_stage_5__1358_, data_stage_5__1357_, data_stage_5__1356_, data_stage_5__1355_, data_stage_5__1354_, data_stage_5__1353_, data_stage_5__1352_, data_stage_5__1351_, data_stage_5__1350_, data_stage_5__1349_, data_stage_5__1348_, data_stage_5__1347_, data_stage_5__1346_, data_stage_5__1345_, data_stage_5__1344_, data_stage_5__1343_, data_stage_5__1342_, data_stage_5__1341_, data_stage_5__1340_, data_stage_5__1339_, data_stage_5__1338_, data_stage_5__1337_, data_stage_5__1336_, data_stage_5__1335_, data_stage_5__1334_, data_stage_5__1333_, data_stage_5__1332_, data_stage_5__1331_, data_stage_5__1330_, data_stage_5__1329_, data_stage_5__1328_, data_stage_5__1327_, data_stage_5__1326_, data_stage_5__1325_, data_stage_5__1324_, data_stage_5__1323_, data_stage_5__1322_, data_stage_5__1321_, data_stage_5__1320_, data_stage_5__1319_, data_stage_5__1318_, data_stage_5__1317_, data_stage_5__1316_, data_stage_5__1315_, data_stage_5__1314_, data_stage_5__1313_, data_stage_5__1312_, data_stage_5__1311_, data_stage_5__1310_, data_stage_5__1309_, data_stage_5__1308_, data_stage_5__1307_, data_stage_5__1306_, data_stage_5__1305_, data_stage_5__1304_, data_stage_5__1303_, data_stage_5__1302_, data_stage_5__1301_, data_stage_5__1300_, data_stage_5__1299_, data_stage_5__1298_, data_stage_5__1297_, data_stage_5__1296_, data_stage_5__1295_, data_stage_5__1294_, data_stage_5__1293_, data_stage_5__1292_, data_stage_5__1291_, data_stage_5__1290_, data_stage_5__1289_, data_stage_5__1288_, data_stage_5__1287_, data_stage_5__1286_, data_stage_5__1285_, data_stage_5__1284_, data_stage_5__1283_, data_stage_5__1282_, data_stage_5__1281_, data_stage_5__1280_, data_stage_5__1279_, data_stage_5__1278_, data_stage_5__1277_, data_stage_5__1276_, data_stage_5__1275_, data_stage_5__1274_, data_stage_5__1273_, data_stage_5__1272_, data_stage_5__1271_, data_stage_5__1270_, data_stage_5__1269_, data_stage_5__1268_, data_stage_5__1267_, data_stage_5__1266_, data_stage_5__1265_, data_stage_5__1264_, data_stage_5__1263_, data_stage_5__1262_, data_stage_5__1261_, data_stage_5__1260_, data_stage_5__1259_, data_stage_5__1258_, data_stage_5__1257_, data_stage_5__1256_, data_stage_5__1255_, data_stage_5__1254_, data_stage_5__1253_, data_stage_5__1252_, data_stage_5__1251_, data_stage_5__1250_, data_stage_5__1249_, data_stage_5__1248_, data_stage_5__1247_, data_stage_5__1246_, data_stage_5__1245_, data_stage_5__1244_, data_stage_5__1243_, data_stage_5__1242_, data_stage_5__1241_, data_stage_5__1240_, data_stage_5__1239_, data_stage_5__1238_, data_stage_5__1237_, data_stage_5__1236_, data_stage_5__1235_, data_stage_5__1234_, data_stage_5__1233_, data_stage_5__1232_, data_stage_5__1231_, data_stage_5__1230_, data_stage_5__1229_, data_stage_5__1228_, data_stage_5__1227_, data_stage_5__1226_, data_stage_5__1225_, data_stage_5__1224_, data_stage_5__1223_, data_stage_5__1222_, data_stage_5__1221_, data_stage_5__1220_, data_stage_5__1219_, data_stage_5__1218_, data_stage_5__1217_, data_stage_5__1216_, data_stage_5__1215_, data_stage_5__1214_, data_stage_5__1213_, data_stage_5__1212_, data_stage_5__1211_, data_stage_5__1210_, data_stage_5__1209_, data_stage_5__1208_, data_stage_5__1207_, data_stage_5__1206_, data_stage_5__1205_, data_stage_5__1204_, data_stage_5__1203_, data_stage_5__1202_, data_stage_5__1201_, data_stage_5__1200_, data_stage_5__1199_, data_stage_5__1198_, data_stage_5__1197_, data_stage_5__1196_, data_stage_5__1195_, data_stage_5__1194_, data_stage_5__1193_, data_stage_5__1192_, data_stage_5__1191_, data_stage_5__1190_, data_stage_5__1189_, data_stage_5__1188_, data_stage_5__1187_, data_stage_5__1186_, data_stage_5__1185_, data_stage_5__1184_, data_stage_5__1183_, data_stage_5__1182_, data_stage_5__1181_, data_stage_5__1180_, data_stage_5__1179_, data_stage_5__1178_, data_stage_5__1177_, data_stage_5__1176_, data_stage_5__1175_, data_stage_5__1174_, data_stage_5__1173_, data_stage_5__1172_, data_stage_5__1171_, data_stage_5__1170_, data_stage_5__1169_, data_stage_5__1168_, data_stage_5__1167_, data_stage_5__1166_, data_stage_5__1165_, data_stage_5__1164_, data_stage_5__1163_, data_stage_5__1162_, data_stage_5__1161_, data_stage_5__1160_, data_stage_5__1159_, data_stage_5__1158_, data_stage_5__1157_, data_stage_5__1156_, data_stage_5__1155_, data_stage_5__1154_, data_stage_5__1153_, data_stage_5__1152_, data_stage_5__1151_, data_stage_5__1150_, data_stage_5__1149_, data_stage_5__1148_, data_stage_5__1147_, data_stage_5__1146_, data_stage_5__1145_, data_stage_5__1144_, data_stage_5__1143_, data_stage_5__1142_, data_stage_5__1141_, data_stage_5__1140_, data_stage_5__1139_, data_stage_5__1138_, data_stage_5__1137_, data_stage_5__1136_, data_stage_5__1135_, data_stage_5__1134_, data_stage_5__1133_, data_stage_5__1132_, data_stage_5__1131_, data_stage_5__1130_, data_stage_5__1129_, data_stage_5__1128_, data_stage_5__1127_, data_stage_5__1126_, data_stage_5__1125_, data_stage_5__1124_, data_stage_5__1123_, data_stage_5__1122_, data_stage_5__1121_, data_stage_5__1120_, data_stage_5__1119_, data_stage_5__1118_, data_stage_5__1117_, data_stage_5__1116_, data_stage_5__1115_, data_stage_5__1114_, data_stage_5__1113_, data_stage_5__1112_, data_stage_5__1111_, data_stage_5__1110_, data_stage_5__1109_, data_stage_5__1108_, data_stage_5__1107_, data_stage_5__1106_, data_stage_5__1105_, data_stage_5__1104_, data_stage_5__1103_, data_stage_5__1102_, data_stage_5__1101_, data_stage_5__1100_, data_stage_5__1099_, data_stage_5__1098_, data_stage_5__1097_, data_stage_5__1096_, data_stage_5__1095_, data_stage_5__1094_, data_stage_5__1093_, data_stage_5__1092_, data_stage_5__1091_, data_stage_5__1090_, data_stage_5__1089_, data_stage_5__1088_, data_stage_5__1087_, data_stage_5__1086_, data_stage_5__1085_, data_stage_5__1084_, data_stage_5__1083_, data_stage_5__1082_, data_stage_5__1081_, data_stage_5__1080_, data_stage_5__1079_, data_stage_5__1078_, data_stage_5__1077_, data_stage_5__1076_, data_stage_5__1075_, data_stage_5__1074_, data_stage_5__1073_, data_stage_5__1072_, data_stage_5__1071_, data_stage_5__1070_, data_stage_5__1069_, data_stage_5__1068_, data_stage_5__1067_, data_stage_5__1066_, data_stage_5__1065_, data_stage_5__1064_, data_stage_5__1063_, data_stage_5__1062_, data_stage_5__1061_, data_stage_5__1060_, data_stage_5__1059_, data_stage_5__1058_, data_stage_5__1057_, data_stage_5__1056_, data_stage_5__1055_, data_stage_5__1054_, data_stage_5__1053_, data_stage_5__1052_, data_stage_5__1051_, data_stage_5__1050_, data_stage_5__1049_, data_stage_5__1048_, data_stage_5__1047_, data_stage_5__1046_, data_stage_5__1045_, data_stage_5__1044_, data_stage_5__1043_, data_stage_5__1042_, data_stage_5__1041_, data_stage_5__1040_, data_stage_5__1039_, data_stage_5__1038_, data_stage_5__1037_, data_stage_5__1036_, data_stage_5__1035_, data_stage_5__1034_, data_stage_5__1033_, data_stage_5__1032_, data_stage_5__1031_, data_stage_5__1030_, data_stage_5__1029_, data_stage_5__1028_, data_stage_5__1027_, data_stage_5__1026_, data_stage_5__1025_, data_stage_5__1024_, data_stage_5__1023_, data_stage_5__1022_, data_stage_5__1021_, data_stage_5__1020_, data_stage_5__1019_, data_stage_5__1018_, data_stage_5__1017_, data_stage_5__1016_, data_stage_5__1015_, data_stage_5__1014_, data_stage_5__1013_, data_stage_5__1012_, data_stage_5__1011_, data_stage_5__1010_, data_stage_5__1009_, data_stage_5__1008_, data_stage_5__1007_, data_stage_5__1006_, data_stage_5__1005_, data_stage_5__1004_, data_stage_5__1003_, data_stage_5__1002_, data_stage_5__1001_, data_stage_5__1000_, data_stage_5__999_, data_stage_5__998_, data_stage_5__997_, data_stage_5__996_, data_stage_5__995_, data_stage_5__994_, data_stage_5__993_, data_stage_5__992_, data_stage_5__991_, data_stage_5__990_, data_stage_5__989_, data_stage_5__988_, data_stage_5__987_, data_stage_5__986_, data_stage_5__985_, data_stage_5__984_, data_stage_5__983_, data_stage_5__982_, data_stage_5__981_, data_stage_5__980_, data_stage_5__979_, data_stage_5__978_, data_stage_5__977_, data_stage_5__976_, data_stage_5__975_, data_stage_5__974_, data_stage_5__973_, data_stage_5__972_, data_stage_5__971_, data_stage_5__970_, data_stage_5__969_, data_stage_5__968_, data_stage_5__967_, data_stage_5__966_, data_stage_5__965_, data_stage_5__964_, data_stage_5__963_, data_stage_5__962_, data_stage_5__961_, data_stage_5__960_, data_stage_5__959_, data_stage_5__958_, data_stage_5__957_, data_stage_5__956_, data_stage_5__955_, data_stage_5__954_, data_stage_5__953_, data_stage_5__952_, data_stage_5__951_, data_stage_5__950_, data_stage_5__949_, data_stage_5__948_, data_stage_5__947_, data_stage_5__946_, data_stage_5__945_, data_stage_5__944_, data_stage_5__943_, data_stage_5__942_, data_stage_5__941_, data_stage_5__940_, data_stage_5__939_, data_stage_5__938_, data_stage_5__937_, data_stage_5__936_, data_stage_5__935_, data_stage_5__934_, data_stage_5__933_, data_stage_5__932_, data_stage_5__931_, data_stage_5__930_, data_stage_5__929_, data_stage_5__928_, data_stage_5__927_, data_stage_5__926_, data_stage_5__925_, data_stage_5__924_, data_stage_5__923_, data_stage_5__922_, data_stage_5__921_, data_stage_5__920_, data_stage_5__919_, data_stage_5__918_, data_stage_5__917_, data_stage_5__916_, data_stage_5__915_, data_stage_5__914_, data_stage_5__913_, data_stage_5__912_, data_stage_5__911_, data_stage_5__910_, data_stage_5__909_, data_stage_5__908_, data_stage_5__907_, data_stage_5__906_, data_stage_5__905_, data_stage_5__904_, data_stage_5__903_, data_stage_5__902_, data_stage_5__901_, data_stage_5__900_, data_stage_5__899_, data_stage_5__898_, data_stage_5__897_, data_stage_5__896_, data_stage_5__895_, data_stage_5__894_, data_stage_5__893_, data_stage_5__892_, data_stage_5__891_, data_stage_5__890_, data_stage_5__889_, data_stage_5__888_, data_stage_5__887_, data_stage_5__886_, data_stage_5__885_, data_stage_5__884_, data_stage_5__883_, data_stage_5__882_, data_stage_5__881_, data_stage_5__880_, data_stage_5__879_, data_stage_5__878_, data_stage_5__877_, data_stage_5__876_, data_stage_5__875_, data_stage_5__874_, data_stage_5__873_, data_stage_5__872_, data_stage_5__871_, data_stage_5__870_, data_stage_5__869_, data_stage_5__868_, data_stage_5__867_, data_stage_5__866_, data_stage_5__865_, data_stage_5__864_, data_stage_5__863_, data_stage_5__862_, data_stage_5__861_, data_stage_5__860_, data_stage_5__859_, data_stage_5__858_, data_stage_5__857_, data_stage_5__856_, data_stage_5__855_, data_stage_5__854_, data_stage_5__853_, data_stage_5__852_, data_stage_5__851_, data_stage_5__850_, data_stage_5__849_, data_stage_5__848_, data_stage_5__847_, data_stage_5__846_, data_stage_5__845_, data_stage_5__844_, data_stage_5__843_, data_stage_5__842_, data_stage_5__841_, data_stage_5__840_, data_stage_5__839_, data_stage_5__838_, data_stage_5__837_, data_stage_5__836_, data_stage_5__835_, data_stage_5__834_, data_stage_5__833_, data_stage_5__832_, data_stage_5__831_, data_stage_5__830_, data_stage_5__829_, data_stage_5__828_, data_stage_5__827_, data_stage_5__826_, data_stage_5__825_, data_stage_5__824_, data_stage_5__823_, data_stage_5__822_, data_stage_5__821_, data_stage_5__820_, data_stage_5__819_, data_stage_5__818_, data_stage_5__817_, data_stage_5__816_, data_stage_5__815_, data_stage_5__814_, data_stage_5__813_, data_stage_5__812_, data_stage_5__811_, data_stage_5__810_, data_stage_5__809_, data_stage_5__808_, data_stage_5__807_, data_stage_5__806_, data_stage_5__805_, data_stage_5__804_, data_stage_5__803_, data_stage_5__802_, data_stage_5__801_, data_stage_5__800_, data_stage_5__799_, data_stage_5__798_, data_stage_5__797_, data_stage_5__796_, data_stage_5__795_, data_stage_5__794_, data_stage_5__793_, data_stage_5__792_, data_stage_5__791_, data_stage_5__790_, data_stage_5__789_, data_stage_5__788_, data_stage_5__787_, data_stage_5__786_, data_stage_5__785_, data_stage_5__784_, data_stage_5__783_, data_stage_5__782_, data_stage_5__781_, data_stage_5__780_, data_stage_5__779_, data_stage_5__778_, data_stage_5__777_, data_stage_5__776_, data_stage_5__775_, data_stage_5__774_, data_stage_5__773_, data_stage_5__772_, data_stage_5__771_, data_stage_5__770_, data_stage_5__769_, data_stage_5__768_, data_stage_5__767_, data_stage_5__766_, data_stage_5__765_, data_stage_5__764_, data_stage_5__763_, data_stage_5__762_, data_stage_5__761_, data_stage_5__760_, data_stage_5__759_, data_stage_5__758_, data_stage_5__757_, data_stage_5__756_, data_stage_5__755_, data_stage_5__754_, data_stage_5__753_, data_stage_5__752_, data_stage_5__751_, data_stage_5__750_, data_stage_5__749_, data_stage_5__748_, data_stage_5__747_, data_stage_5__746_, data_stage_5__745_, data_stage_5__744_, data_stage_5__743_, data_stage_5__742_, data_stage_5__741_, data_stage_5__740_, data_stage_5__739_, data_stage_5__738_, data_stage_5__737_, data_stage_5__736_, data_stage_5__735_, data_stage_5__734_, data_stage_5__733_, data_stage_5__732_, data_stage_5__731_, data_stage_5__730_, data_stage_5__729_, data_stage_5__728_, data_stage_5__727_, data_stage_5__726_, data_stage_5__725_, data_stage_5__724_, data_stage_5__723_, data_stage_5__722_, data_stage_5__721_, data_stage_5__720_, data_stage_5__719_, data_stage_5__718_, data_stage_5__717_, data_stage_5__716_, data_stage_5__715_, data_stage_5__714_, data_stage_5__713_, data_stage_5__712_, data_stage_5__711_, data_stage_5__710_, data_stage_5__709_, data_stage_5__708_, data_stage_5__707_, data_stage_5__706_, data_stage_5__705_, data_stage_5__704_, data_stage_5__703_, data_stage_5__702_, data_stage_5__701_, data_stage_5__700_, data_stage_5__699_, data_stage_5__698_, data_stage_5__697_, data_stage_5__696_, data_stage_5__695_, data_stage_5__694_, data_stage_5__693_, data_stage_5__692_, data_stage_5__691_, data_stage_5__690_, data_stage_5__689_, data_stage_5__688_, data_stage_5__687_, data_stage_5__686_, data_stage_5__685_, data_stage_5__684_, data_stage_5__683_, data_stage_5__682_, data_stage_5__681_, data_stage_5__680_, data_stage_5__679_, data_stage_5__678_, data_stage_5__677_, data_stage_5__676_, data_stage_5__675_, data_stage_5__674_, data_stage_5__673_, data_stage_5__672_, data_stage_5__671_, data_stage_5__670_, data_stage_5__669_, data_stage_5__668_, data_stage_5__667_, data_stage_5__666_, data_stage_5__665_, data_stage_5__664_, data_stage_5__663_, data_stage_5__662_, data_stage_5__661_, data_stage_5__660_, data_stage_5__659_, data_stage_5__658_, data_stage_5__657_, data_stage_5__656_, data_stage_5__655_, data_stage_5__654_, data_stage_5__653_, data_stage_5__652_, data_stage_5__651_, data_stage_5__650_, data_stage_5__649_, data_stage_5__648_, data_stage_5__647_, data_stage_5__646_, data_stage_5__645_, data_stage_5__644_, data_stage_5__643_, data_stage_5__642_, data_stage_5__641_, data_stage_5__640_, data_stage_5__639_, data_stage_5__638_, data_stage_5__637_, data_stage_5__636_, data_stage_5__635_, data_stage_5__634_, data_stage_5__633_, data_stage_5__632_, data_stage_5__631_, data_stage_5__630_, data_stage_5__629_, data_stage_5__628_, data_stage_5__627_, data_stage_5__626_, data_stage_5__625_, data_stage_5__624_, data_stage_5__623_, data_stage_5__622_, data_stage_5__621_, data_stage_5__620_, data_stage_5__619_, data_stage_5__618_, data_stage_5__617_, data_stage_5__616_, data_stage_5__615_, data_stage_5__614_, data_stage_5__613_, data_stage_5__612_, data_stage_5__611_, data_stage_5__610_, data_stage_5__609_, data_stage_5__608_, data_stage_5__607_, data_stage_5__606_, data_stage_5__605_, data_stage_5__604_, data_stage_5__603_, data_stage_5__602_, data_stage_5__601_, data_stage_5__600_, data_stage_5__599_, data_stage_5__598_, data_stage_5__597_, data_stage_5__596_, data_stage_5__595_, data_stage_5__594_, data_stage_5__593_, data_stage_5__592_, data_stage_5__591_, data_stage_5__590_, data_stage_5__589_, data_stage_5__588_, data_stage_5__587_, data_stage_5__586_, data_stage_5__585_, data_stage_5__584_, data_stage_5__583_, data_stage_5__582_, data_stage_5__581_, data_stage_5__580_, data_stage_5__579_, data_stage_5__578_, data_stage_5__577_, data_stage_5__576_, data_stage_5__575_, data_stage_5__574_, data_stage_5__573_, data_stage_5__572_, data_stage_5__571_, data_stage_5__570_, data_stage_5__569_, data_stage_5__568_, data_stage_5__567_, data_stage_5__566_, data_stage_5__565_, data_stage_5__564_, data_stage_5__563_, data_stage_5__562_, data_stage_5__561_, data_stage_5__560_, data_stage_5__559_, data_stage_5__558_, data_stage_5__557_, data_stage_5__556_, data_stage_5__555_, data_stage_5__554_, data_stage_5__553_, data_stage_5__552_, data_stage_5__551_, data_stage_5__550_, data_stage_5__549_, data_stage_5__548_, data_stage_5__547_, data_stage_5__546_, data_stage_5__545_, data_stage_5__544_, data_stage_5__543_, data_stage_5__542_, data_stage_5__541_, data_stage_5__540_, data_stage_5__539_, data_stage_5__538_, data_stage_5__537_, data_stage_5__536_, data_stage_5__535_, data_stage_5__534_, data_stage_5__533_, data_stage_5__532_, data_stage_5__531_, data_stage_5__530_, data_stage_5__529_, data_stage_5__528_, data_stage_5__527_, data_stage_5__526_, data_stage_5__525_, data_stage_5__524_, data_stage_5__523_, data_stage_5__522_, data_stage_5__521_, data_stage_5__520_, data_stage_5__519_, data_stage_5__518_, data_stage_5__517_, data_stage_5__516_, data_stage_5__515_, data_stage_5__514_, data_stage_5__513_, data_stage_5__512_, data_stage_5__511_, data_stage_5__510_, data_stage_5__509_, data_stage_5__508_, data_stage_5__507_, data_stage_5__506_, data_stage_5__505_, data_stage_5__504_, data_stage_5__503_, data_stage_5__502_, data_stage_5__501_, data_stage_5__500_, data_stage_5__499_, data_stage_5__498_, data_stage_5__497_, data_stage_5__496_, data_stage_5__495_, data_stage_5__494_, data_stage_5__493_, data_stage_5__492_, data_stage_5__491_, data_stage_5__490_, data_stage_5__489_, data_stage_5__488_, data_stage_5__487_, data_stage_5__486_, data_stage_5__485_, data_stage_5__484_, data_stage_5__483_, data_stage_5__482_, data_stage_5__481_, data_stage_5__480_, data_stage_5__479_, data_stage_5__478_, data_stage_5__477_, data_stage_5__476_, data_stage_5__475_, data_stage_5__474_, data_stage_5__473_, data_stage_5__472_, data_stage_5__471_, data_stage_5__470_, data_stage_5__469_, data_stage_5__468_, data_stage_5__467_, data_stage_5__466_, data_stage_5__465_, data_stage_5__464_, data_stage_5__463_, data_stage_5__462_, data_stage_5__461_, data_stage_5__460_, data_stage_5__459_, data_stage_5__458_, data_stage_5__457_, data_stage_5__456_, data_stage_5__455_, data_stage_5__454_, data_stage_5__453_, data_stage_5__452_, data_stage_5__451_, data_stage_5__450_, data_stage_5__449_, data_stage_5__448_, data_stage_5__447_, data_stage_5__446_, data_stage_5__445_, data_stage_5__444_, data_stage_5__443_, data_stage_5__442_, data_stage_5__441_, data_stage_5__440_, data_stage_5__439_, data_stage_5__438_, data_stage_5__437_, data_stage_5__436_, data_stage_5__435_, data_stage_5__434_, data_stage_5__433_, data_stage_5__432_, data_stage_5__431_, data_stage_5__430_, data_stage_5__429_, data_stage_5__428_, data_stage_5__427_, data_stage_5__426_, data_stage_5__425_, data_stage_5__424_, data_stage_5__423_, data_stage_5__422_, data_stage_5__421_, data_stage_5__420_, data_stage_5__419_, data_stage_5__418_, data_stage_5__417_, data_stage_5__416_, data_stage_5__415_, data_stage_5__414_, data_stage_5__413_, data_stage_5__412_, data_stage_5__411_, data_stage_5__410_, data_stage_5__409_, data_stage_5__408_, data_stage_5__407_, data_stage_5__406_, data_stage_5__405_, data_stage_5__404_, data_stage_5__403_, data_stage_5__402_, data_stage_5__401_, data_stage_5__400_, data_stage_5__399_, data_stage_5__398_, data_stage_5__397_, data_stage_5__396_, data_stage_5__395_, data_stage_5__394_, data_stage_5__393_, data_stage_5__392_, data_stage_5__391_, data_stage_5__390_, data_stage_5__389_, data_stage_5__388_, data_stage_5__387_, data_stage_5__386_, data_stage_5__385_, data_stage_5__384_, data_stage_5__383_, data_stage_5__382_, data_stage_5__381_, data_stage_5__380_, data_stage_5__379_, data_stage_5__378_, data_stage_5__377_, data_stage_5__376_, data_stage_5__375_, data_stage_5__374_, data_stage_5__373_, data_stage_5__372_, data_stage_5__371_, data_stage_5__370_, data_stage_5__369_, data_stage_5__368_, data_stage_5__367_, data_stage_5__366_, data_stage_5__365_, data_stage_5__364_, data_stage_5__363_, data_stage_5__362_, data_stage_5__361_, data_stage_5__360_, data_stage_5__359_, data_stage_5__358_, data_stage_5__357_, data_stage_5__356_, data_stage_5__355_, data_stage_5__354_, data_stage_5__353_, data_stage_5__352_, data_stage_5__351_, data_stage_5__350_, data_stage_5__349_, data_stage_5__348_, data_stage_5__347_, data_stage_5__346_, data_stage_5__345_, data_stage_5__344_, data_stage_5__343_, data_stage_5__342_, data_stage_5__341_, data_stage_5__340_, data_stage_5__339_, data_stage_5__338_, data_stage_5__337_, data_stage_5__336_, data_stage_5__335_, data_stage_5__334_, data_stage_5__333_, data_stage_5__332_, data_stage_5__331_, data_stage_5__330_, data_stage_5__329_, data_stage_5__328_, data_stage_5__327_, data_stage_5__326_, data_stage_5__325_, data_stage_5__324_, data_stage_5__323_, data_stage_5__322_, data_stage_5__321_, data_stage_5__320_, data_stage_5__319_, data_stage_5__318_, data_stage_5__317_, data_stage_5__316_, data_stage_5__315_, data_stage_5__314_, data_stage_5__313_, data_stage_5__312_, data_stage_5__311_, data_stage_5__310_, data_stage_5__309_, data_stage_5__308_, data_stage_5__307_, data_stage_5__306_, data_stage_5__305_, data_stage_5__304_, data_stage_5__303_, data_stage_5__302_, data_stage_5__301_, data_stage_5__300_, data_stage_5__299_, data_stage_5__298_, data_stage_5__297_, data_stage_5__296_, data_stage_5__295_, data_stage_5__294_, data_stage_5__293_, data_stage_5__292_, data_stage_5__291_, data_stage_5__290_, data_stage_5__289_, data_stage_5__288_, data_stage_5__287_, data_stage_5__286_, data_stage_5__285_, data_stage_5__284_, data_stage_5__283_, data_stage_5__282_, data_stage_5__281_, data_stage_5__280_, data_stage_5__279_, data_stage_5__278_, data_stage_5__277_, data_stage_5__276_, data_stage_5__275_, data_stage_5__274_, data_stage_5__273_, data_stage_5__272_, data_stage_5__271_, data_stage_5__270_, data_stage_5__269_, data_stage_5__268_, data_stage_5__267_, data_stage_5__266_, data_stage_5__265_, data_stage_5__264_, data_stage_5__263_, data_stage_5__262_, data_stage_5__261_, data_stage_5__260_, data_stage_5__259_, data_stage_5__258_, data_stage_5__257_, data_stage_5__256_, data_stage_5__255_, data_stage_5__254_, data_stage_5__253_, data_stage_5__252_, data_stage_5__251_, data_stage_5__250_, data_stage_5__249_, data_stage_5__248_, data_stage_5__247_, data_stage_5__246_, data_stage_5__245_, data_stage_5__244_, data_stage_5__243_, data_stage_5__242_, data_stage_5__241_, data_stage_5__240_, data_stage_5__239_, data_stage_5__238_, data_stage_5__237_, data_stage_5__236_, data_stage_5__235_, data_stage_5__234_, data_stage_5__233_, data_stage_5__232_, data_stage_5__231_, data_stage_5__230_, data_stage_5__229_, data_stage_5__228_, data_stage_5__227_, data_stage_5__226_, data_stage_5__225_, data_stage_5__224_, data_stage_5__223_, data_stage_5__222_, data_stage_5__221_, data_stage_5__220_, data_stage_5__219_, data_stage_5__218_, data_stage_5__217_, data_stage_5__216_, data_stage_5__215_, data_stage_5__214_, data_stage_5__213_, data_stage_5__212_, data_stage_5__211_, data_stage_5__210_, data_stage_5__209_, data_stage_5__208_, data_stage_5__207_, data_stage_5__206_, data_stage_5__205_, data_stage_5__204_, data_stage_5__203_, data_stage_5__202_, data_stage_5__201_, data_stage_5__200_, data_stage_5__199_, data_stage_5__198_, data_stage_5__197_, data_stage_5__196_, data_stage_5__195_, data_stage_5__194_, data_stage_5__193_, data_stage_5__192_, data_stage_5__191_, data_stage_5__190_, data_stage_5__189_, data_stage_5__188_, data_stage_5__187_, data_stage_5__186_, data_stage_5__185_, data_stage_5__184_, data_stage_5__183_, data_stage_5__182_, data_stage_5__181_, data_stage_5__180_, data_stage_5__179_, data_stage_5__178_, data_stage_5__177_, data_stage_5__176_, data_stage_5__175_, data_stage_5__174_, data_stage_5__173_, data_stage_5__172_, data_stage_5__171_, data_stage_5__170_, data_stage_5__169_, data_stage_5__168_, data_stage_5__167_, data_stage_5__166_, data_stage_5__165_, data_stage_5__164_, data_stage_5__163_, data_stage_5__162_, data_stage_5__161_, data_stage_5__160_, data_stage_5__159_, data_stage_5__158_, data_stage_5__157_, data_stage_5__156_, data_stage_5__155_, data_stage_5__154_, data_stage_5__153_, data_stage_5__152_, data_stage_5__151_, data_stage_5__150_, data_stage_5__149_, data_stage_5__148_, data_stage_5__147_, data_stage_5__146_, data_stage_5__145_, data_stage_5__144_, data_stage_5__143_, data_stage_5__142_, data_stage_5__141_, data_stage_5__140_, data_stage_5__139_, data_stage_5__138_, data_stage_5__137_, data_stage_5__136_, data_stage_5__135_, data_stage_5__134_, data_stage_5__133_, data_stage_5__132_, data_stage_5__131_, data_stage_5__130_, data_stage_5__129_, data_stage_5__128_, data_stage_5__127_, data_stage_5__126_, data_stage_5__125_, data_stage_5__124_, data_stage_5__123_, data_stage_5__122_, data_stage_5__121_, data_stage_5__120_, data_stage_5__119_, data_stage_5__118_, data_stage_5__117_, data_stage_5__116_, data_stage_5__115_, data_stage_5__114_, data_stage_5__113_, data_stage_5__112_, data_stage_5__111_, data_stage_5__110_, data_stage_5__109_, data_stage_5__108_, data_stage_5__107_, data_stage_5__106_, data_stage_5__105_, data_stage_5__104_, data_stage_5__103_, data_stage_5__102_, data_stage_5__101_, data_stage_5__100_, data_stage_5__99_, data_stage_5__98_, data_stage_5__97_, data_stage_5__96_, data_stage_5__95_, data_stage_5__94_, data_stage_5__93_, data_stage_5__92_, data_stage_5__91_, data_stage_5__90_, data_stage_5__89_, data_stage_5__88_, data_stage_5__87_, data_stage_5__86_, data_stage_5__85_, data_stage_5__84_, data_stage_5__83_, data_stage_5__82_, data_stage_5__81_, data_stage_5__80_, data_stage_5__79_, data_stage_5__78_, data_stage_5__77_, data_stage_5__76_, data_stage_5__75_, data_stage_5__74_, data_stage_5__73_, data_stage_5__72_, data_stage_5__71_, data_stage_5__70_, data_stage_5__69_, data_stage_5__68_, data_stage_5__67_, data_stage_5__66_, data_stage_5__65_, data_stage_5__64_, data_stage_5__63_, data_stage_5__62_, data_stage_5__61_, data_stage_5__60_, data_stage_5__59_, data_stage_5__58_, data_stage_5__57_, data_stage_5__56_, data_stage_5__55_, data_stage_5__54_, data_stage_5__53_, data_stage_5__52_, data_stage_5__51_, data_stage_5__50_, data_stage_5__49_, data_stage_5__48_, data_stage_5__47_, data_stage_5__46_, data_stage_5__45_, data_stage_5__44_, data_stage_5__43_, data_stage_5__42_, data_stage_5__41_, data_stage_5__40_, data_stage_5__39_, data_stage_5__38_, data_stage_5__37_, data_stage_5__36_, data_stage_5__35_, data_stage_5__34_, data_stage_5__33_, data_stage_5__32_, data_stage_5__31_, data_stage_5__30_, data_stage_5__29_, data_stage_5__28_, data_stage_5__27_, data_stage_5__26_, data_stage_5__25_, data_stage_5__24_, data_stage_5__23_, data_stage_5__22_, data_stage_5__21_, data_stage_5__20_, data_stage_5__19_, data_stage_5__18_, data_stage_5__17_, data_stage_5__16_, data_stage_5__15_, data_stage_5__14_, data_stage_5__13_, data_stage_5__12_, data_stage_5__11_, data_stage_5__10_, data_stage_5__9_, data_stage_5__8_, data_stage_5__7_, data_stage_5__6_, data_stage_5__5_, data_stage_5__4_, data_stage_5__3_, data_stage_5__2_, data_stage_5__1_, data_stage_5__0_ }),
    .swap_i(sel_i[5]),
    .data_o(data_o)
  );


endmodule

