

module top
(
  gray_i,
  binary_o
);

  input [63:0] gray_i;
  output [63:0] binary_o;

  bsg_gray_to_binary
  wrapper
  (
    .gray_i(gray_i),
    .binary_o(binary_o)
  );


endmodule



module bsg_scan_width_p64_xor_p1
(
  i,
  o
);

  input [63:0] i;
  output [63:0] o;
  wire [63:0] o;
  wire t_5__63_,t_5__62_,t_5__61_,t_5__60_,t_5__59_,t_5__58_,t_5__57_,t_5__56_,
  t_5__55_,t_5__54_,t_5__53_,t_5__52_,t_5__51_,t_5__50_,t_5__49_,t_5__48_,t_5__47_,
  t_5__46_,t_5__45_,t_5__44_,t_5__43_,t_5__42_,t_5__41_,t_5__40_,t_5__39_,t_5__38_,
  t_5__37_,t_5__36_,t_5__35_,t_5__34_,t_5__33_,t_5__32_,t_5__31_,t_5__30_,t_5__29_,
  t_5__28_,t_5__27_,t_5__26_,t_5__25_,t_5__24_,t_5__23_,t_5__22_,t_5__21_,t_5__20_,
  t_5__19_,t_5__18_,t_5__17_,t_5__16_,t_5__15_,t_5__14_,t_5__13_,t_5__12_,t_5__11_,
  t_5__10_,t_5__9_,t_5__8_,t_5__7_,t_5__6_,t_5__5_,t_5__4_,t_5__3_,t_5__2_,t_5__1_,
  t_5__0_,t_4__63_,t_4__62_,t_4__61_,t_4__60_,t_4__59_,t_4__58_,t_4__57_,t_4__56_,
  t_4__55_,t_4__54_,t_4__53_,t_4__52_,t_4__51_,t_4__50_,t_4__49_,t_4__48_,t_4__47_,
  t_4__46_,t_4__45_,t_4__44_,t_4__43_,t_4__42_,t_4__41_,t_4__40_,t_4__39_,t_4__38_,
  t_4__37_,t_4__36_,t_4__35_,t_4__34_,t_4__33_,t_4__32_,t_4__31_,t_4__30_,
  t_4__29_,t_4__28_,t_4__27_,t_4__26_,t_4__25_,t_4__24_,t_4__23_,t_4__22_,t_4__21_,
  t_4__20_,t_4__19_,t_4__18_,t_4__17_,t_4__16_,t_4__15_,t_4__14_,t_4__13_,t_4__12_,
  t_4__11_,t_4__10_,t_4__9_,t_4__8_,t_4__7_,t_4__6_,t_4__5_,t_4__4_,t_4__3_,t_4__2_,
  t_4__1_,t_4__0_,t_3__63_,t_3__62_,t_3__61_,t_3__60_,t_3__59_,t_3__58_,t_3__57_,
  t_3__56_,t_3__55_,t_3__54_,t_3__53_,t_3__52_,t_3__51_,t_3__50_,t_3__49_,t_3__48_,
  t_3__47_,t_3__46_,t_3__45_,t_3__44_,t_3__43_,t_3__42_,t_3__41_,t_3__40_,t_3__39_,
  t_3__38_,t_3__37_,t_3__36_,t_3__35_,t_3__34_,t_3__33_,t_3__32_,t_3__31_,t_3__30_,
  t_3__29_,t_3__28_,t_3__27_,t_3__26_,t_3__25_,t_3__24_,t_3__23_,t_3__22_,t_3__21_,
  t_3__20_,t_3__19_,t_3__18_,t_3__17_,t_3__16_,t_3__15_,t_3__14_,t_3__13_,t_3__12_,
  t_3__11_,t_3__10_,t_3__9_,t_3__8_,t_3__7_,t_3__6_,t_3__5_,t_3__4_,t_3__3_,
  t_3__2_,t_3__1_,t_3__0_,t_2__63_,t_2__62_,t_2__61_,t_2__60_,t_2__59_,t_2__58_,
  t_2__57_,t_2__56_,t_2__55_,t_2__54_,t_2__53_,t_2__52_,t_2__51_,t_2__50_,t_2__49_,
  t_2__48_,t_2__47_,t_2__46_,t_2__45_,t_2__44_,t_2__43_,t_2__42_,t_2__41_,t_2__40_,
  t_2__39_,t_2__38_,t_2__37_,t_2__36_,t_2__35_,t_2__34_,t_2__33_,t_2__32_,t_2__31_,
  t_2__30_,t_2__29_,t_2__28_,t_2__27_,t_2__26_,t_2__25_,t_2__24_,t_2__23_,t_2__22_,
  t_2__21_,t_2__20_,t_2__19_,t_2__18_,t_2__17_,t_2__16_,t_2__15_,t_2__14_,t_2__13_,
  t_2__12_,t_2__11_,t_2__10_,t_2__9_,t_2__8_,t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,
  t_2__2_,t_2__1_,t_2__0_,t_1__63_,t_1__62_,t_1__61_,t_1__60_,t_1__59_,t_1__58_,
  t_1__57_,t_1__56_,t_1__55_,t_1__54_,t_1__53_,t_1__52_,t_1__51_,t_1__50_,t_1__49_,
  t_1__48_,t_1__47_,t_1__46_,t_1__45_,t_1__44_,t_1__43_,t_1__42_,t_1__41_,t_1__40_,
  t_1__39_,t_1__38_,t_1__37_,t_1__36_,t_1__35_,t_1__34_,t_1__33_,t_1__32_,
  t_1__31_,t_1__30_,t_1__29_,t_1__28_,t_1__27_,t_1__26_,t_1__25_,t_1__24_,t_1__23_,
  t_1__22_,t_1__21_,t_1__20_,t_1__19_,t_1__18_,t_1__17_,t_1__16_,t_1__15_,t_1__14_,
  t_1__13_,t_1__12_,t_1__11_,t_1__10_,t_1__9_,t_1__8_,t_1__7_,t_1__6_,t_1__5_,t_1__4_,
  t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__63_ = i[63] ^ 1'b0;
  assign t_1__62_ = i[62] ^ i[63];
  assign t_1__61_ = i[61] ^ i[62];
  assign t_1__60_ = i[60] ^ i[61];
  assign t_1__59_ = i[59] ^ i[60];
  assign t_1__58_ = i[58] ^ i[59];
  assign t_1__57_ = i[57] ^ i[58];
  assign t_1__56_ = i[56] ^ i[57];
  assign t_1__55_ = i[55] ^ i[56];
  assign t_1__54_ = i[54] ^ i[55];
  assign t_1__53_ = i[53] ^ i[54];
  assign t_1__52_ = i[52] ^ i[53];
  assign t_1__51_ = i[51] ^ i[52];
  assign t_1__50_ = i[50] ^ i[51];
  assign t_1__49_ = i[49] ^ i[50];
  assign t_1__48_ = i[48] ^ i[49];
  assign t_1__47_ = i[47] ^ i[48];
  assign t_1__46_ = i[46] ^ i[47];
  assign t_1__45_ = i[45] ^ i[46];
  assign t_1__44_ = i[44] ^ i[45];
  assign t_1__43_ = i[43] ^ i[44];
  assign t_1__42_ = i[42] ^ i[43];
  assign t_1__41_ = i[41] ^ i[42];
  assign t_1__40_ = i[40] ^ i[41];
  assign t_1__39_ = i[39] ^ i[40];
  assign t_1__38_ = i[38] ^ i[39];
  assign t_1__37_ = i[37] ^ i[38];
  assign t_1__36_ = i[36] ^ i[37];
  assign t_1__35_ = i[35] ^ i[36];
  assign t_1__34_ = i[34] ^ i[35];
  assign t_1__33_ = i[33] ^ i[34];
  assign t_1__32_ = i[32] ^ i[33];
  assign t_1__31_ = i[31] ^ i[32];
  assign t_1__30_ = i[30] ^ i[31];
  assign t_1__29_ = i[29] ^ i[30];
  assign t_1__28_ = i[28] ^ i[29];
  assign t_1__27_ = i[27] ^ i[28];
  assign t_1__26_ = i[26] ^ i[27];
  assign t_1__25_ = i[25] ^ i[26];
  assign t_1__24_ = i[24] ^ i[25];
  assign t_1__23_ = i[23] ^ i[24];
  assign t_1__22_ = i[22] ^ i[23];
  assign t_1__21_ = i[21] ^ i[22];
  assign t_1__20_ = i[20] ^ i[21];
  assign t_1__19_ = i[19] ^ i[20];
  assign t_1__18_ = i[18] ^ i[19];
  assign t_1__17_ = i[17] ^ i[18];
  assign t_1__16_ = i[16] ^ i[17];
  assign t_1__15_ = i[15] ^ i[16];
  assign t_1__14_ = i[14] ^ i[15];
  assign t_1__13_ = i[13] ^ i[14];
  assign t_1__12_ = i[12] ^ i[13];
  assign t_1__11_ = i[11] ^ i[12];
  assign t_1__10_ = i[10] ^ i[11];
  assign t_1__9_ = i[9] ^ i[10];
  assign t_1__8_ = i[8] ^ i[9];
  assign t_1__7_ = i[7] ^ i[8];
  assign t_1__6_ = i[6] ^ i[7];
  assign t_1__5_ = i[5] ^ i[6];
  assign t_1__4_ = i[4] ^ i[5];
  assign t_1__3_ = i[3] ^ i[4];
  assign t_1__2_ = i[2] ^ i[3];
  assign t_1__1_ = i[1] ^ i[2];
  assign t_1__0_ = i[0] ^ i[1];
  assign t_2__63_ = t_1__63_ ^ 1'b0;
  assign t_2__62_ = t_1__62_ ^ 1'b0;
  assign t_2__61_ = t_1__61_ ^ t_1__63_;
  assign t_2__60_ = t_1__60_ ^ t_1__62_;
  assign t_2__59_ = t_1__59_ ^ t_1__61_;
  assign t_2__58_ = t_1__58_ ^ t_1__60_;
  assign t_2__57_ = t_1__57_ ^ t_1__59_;
  assign t_2__56_ = t_1__56_ ^ t_1__58_;
  assign t_2__55_ = t_1__55_ ^ t_1__57_;
  assign t_2__54_ = t_1__54_ ^ t_1__56_;
  assign t_2__53_ = t_1__53_ ^ t_1__55_;
  assign t_2__52_ = t_1__52_ ^ t_1__54_;
  assign t_2__51_ = t_1__51_ ^ t_1__53_;
  assign t_2__50_ = t_1__50_ ^ t_1__52_;
  assign t_2__49_ = t_1__49_ ^ t_1__51_;
  assign t_2__48_ = t_1__48_ ^ t_1__50_;
  assign t_2__47_ = t_1__47_ ^ t_1__49_;
  assign t_2__46_ = t_1__46_ ^ t_1__48_;
  assign t_2__45_ = t_1__45_ ^ t_1__47_;
  assign t_2__44_ = t_1__44_ ^ t_1__46_;
  assign t_2__43_ = t_1__43_ ^ t_1__45_;
  assign t_2__42_ = t_1__42_ ^ t_1__44_;
  assign t_2__41_ = t_1__41_ ^ t_1__43_;
  assign t_2__40_ = t_1__40_ ^ t_1__42_;
  assign t_2__39_ = t_1__39_ ^ t_1__41_;
  assign t_2__38_ = t_1__38_ ^ t_1__40_;
  assign t_2__37_ = t_1__37_ ^ t_1__39_;
  assign t_2__36_ = t_1__36_ ^ t_1__38_;
  assign t_2__35_ = t_1__35_ ^ t_1__37_;
  assign t_2__34_ = t_1__34_ ^ t_1__36_;
  assign t_2__33_ = t_1__33_ ^ t_1__35_;
  assign t_2__32_ = t_1__32_ ^ t_1__34_;
  assign t_2__31_ = t_1__31_ ^ t_1__33_;
  assign t_2__30_ = t_1__30_ ^ t_1__32_;
  assign t_2__29_ = t_1__29_ ^ t_1__31_;
  assign t_2__28_ = t_1__28_ ^ t_1__30_;
  assign t_2__27_ = t_1__27_ ^ t_1__29_;
  assign t_2__26_ = t_1__26_ ^ t_1__28_;
  assign t_2__25_ = t_1__25_ ^ t_1__27_;
  assign t_2__24_ = t_1__24_ ^ t_1__26_;
  assign t_2__23_ = t_1__23_ ^ t_1__25_;
  assign t_2__22_ = t_1__22_ ^ t_1__24_;
  assign t_2__21_ = t_1__21_ ^ t_1__23_;
  assign t_2__20_ = t_1__20_ ^ t_1__22_;
  assign t_2__19_ = t_1__19_ ^ t_1__21_;
  assign t_2__18_ = t_1__18_ ^ t_1__20_;
  assign t_2__17_ = t_1__17_ ^ t_1__19_;
  assign t_2__16_ = t_1__16_ ^ t_1__18_;
  assign t_2__15_ = t_1__15_ ^ t_1__17_;
  assign t_2__14_ = t_1__14_ ^ t_1__16_;
  assign t_2__13_ = t_1__13_ ^ t_1__15_;
  assign t_2__12_ = t_1__12_ ^ t_1__14_;
  assign t_2__11_ = t_1__11_ ^ t_1__13_;
  assign t_2__10_ = t_1__10_ ^ t_1__12_;
  assign t_2__9_ = t_1__9_ ^ t_1__11_;
  assign t_2__8_ = t_1__8_ ^ t_1__10_;
  assign t_2__7_ = t_1__7_ ^ t_1__9_;
  assign t_2__6_ = t_1__6_ ^ t_1__8_;
  assign t_2__5_ = t_1__5_ ^ t_1__7_;
  assign t_2__4_ = t_1__4_ ^ t_1__6_;
  assign t_2__3_ = t_1__3_ ^ t_1__5_;
  assign t_2__2_ = t_1__2_ ^ t_1__4_;
  assign t_2__1_ = t_1__1_ ^ t_1__3_;
  assign t_2__0_ = t_1__0_ ^ t_1__2_;
  assign t_3__63_ = t_2__63_ ^ 1'b0;
  assign t_3__62_ = t_2__62_ ^ 1'b0;
  assign t_3__61_ = t_2__61_ ^ 1'b0;
  assign t_3__60_ = t_2__60_ ^ 1'b0;
  assign t_3__59_ = t_2__59_ ^ t_2__63_;
  assign t_3__58_ = t_2__58_ ^ t_2__62_;
  assign t_3__57_ = t_2__57_ ^ t_2__61_;
  assign t_3__56_ = t_2__56_ ^ t_2__60_;
  assign t_3__55_ = t_2__55_ ^ t_2__59_;
  assign t_3__54_ = t_2__54_ ^ t_2__58_;
  assign t_3__53_ = t_2__53_ ^ t_2__57_;
  assign t_3__52_ = t_2__52_ ^ t_2__56_;
  assign t_3__51_ = t_2__51_ ^ t_2__55_;
  assign t_3__50_ = t_2__50_ ^ t_2__54_;
  assign t_3__49_ = t_2__49_ ^ t_2__53_;
  assign t_3__48_ = t_2__48_ ^ t_2__52_;
  assign t_3__47_ = t_2__47_ ^ t_2__51_;
  assign t_3__46_ = t_2__46_ ^ t_2__50_;
  assign t_3__45_ = t_2__45_ ^ t_2__49_;
  assign t_3__44_ = t_2__44_ ^ t_2__48_;
  assign t_3__43_ = t_2__43_ ^ t_2__47_;
  assign t_3__42_ = t_2__42_ ^ t_2__46_;
  assign t_3__41_ = t_2__41_ ^ t_2__45_;
  assign t_3__40_ = t_2__40_ ^ t_2__44_;
  assign t_3__39_ = t_2__39_ ^ t_2__43_;
  assign t_3__38_ = t_2__38_ ^ t_2__42_;
  assign t_3__37_ = t_2__37_ ^ t_2__41_;
  assign t_3__36_ = t_2__36_ ^ t_2__40_;
  assign t_3__35_ = t_2__35_ ^ t_2__39_;
  assign t_3__34_ = t_2__34_ ^ t_2__38_;
  assign t_3__33_ = t_2__33_ ^ t_2__37_;
  assign t_3__32_ = t_2__32_ ^ t_2__36_;
  assign t_3__31_ = t_2__31_ ^ t_2__35_;
  assign t_3__30_ = t_2__30_ ^ t_2__34_;
  assign t_3__29_ = t_2__29_ ^ t_2__33_;
  assign t_3__28_ = t_2__28_ ^ t_2__32_;
  assign t_3__27_ = t_2__27_ ^ t_2__31_;
  assign t_3__26_ = t_2__26_ ^ t_2__30_;
  assign t_3__25_ = t_2__25_ ^ t_2__29_;
  assign t_3__24_ = t_2__24_ ^ t_2__28_;
  assign t_3__23_ = t_2__23_ ^ t_2__27_;
  assign t_3__22_ = t_2__22_ ^ t_2__26_;
  assign t_3__21_ = t_2__21_ ^ t_2__25_;
  assign t_3__20_ = t_2__20_ ^ t_2__24_;
  assign t_3__19_ = t_2__19_ ^ t_2__23_;
  assign t_3__18_ = t_2__18_ ^ t_2__22_;
  assign t_3__17_ = t_2__17_ ^ t_2__21_;
  assign t_3__16_ = t_2__16_ ^ t_2__20_;
  assign t_3__15_ = t_2__15_ ^ t_2__19_;
  assign t_3__14_ = t_2__14_ ^ t_2__18_;
  assign t_3__13_ = t_2__13_ ^ t_2__17_;
  assign t_3__12_ = t_2__12_ ^ t_2__16_;
  assign t_3__11_ = t_2__11_ ^ t_2__15_;
  assign t_3__10_ = t_2__10_ ^ t_2__14_;
  assign t_3__9_ = t_2__9_ ^ t_2__13_;
  assign t_3__8_ = t_2__8_ ^ t_2__12_;
  assign t_3__7_ = t_2__7_ ^ t_2__11_;
  assign t_3__6_ = t_2__6_ ^ t_2__10_;
  assign t_3__5_ = t_2__5_ ^ t_2__9_;
  assign t_3__4_ = t_2__4_ ^ t_2__8_;
  assign t_3__3_ = t_2__3_ ^ t_2__7_;
  assign t_3__2_ = t_2__2_ ^ t_2__6_;
  assign t_3__1_ = t_2__1_ ^ t_2__5_;
  assign t_3__0_ = t_2__0_ ^ t_2__4_;
  assign t_4__63_ = t_3__63_ ^ 1'b0;
  assign t_4__62_ = t_3__62_ ^ 1'b0;
  assign t_4__61_ = t_3__61_ ^ 1'b0;
  assign t_4__60_ = t_3__60_ ^ 1'b0;
  assign t_4__59_ = t_3__59_ ^ 1'b0;
  assign t_4__58_ = t_3__58_ ^ 1'b0;
  assign t_4__57_ = t_3__57_ ^ 1'b0;
  assign t_4__56_ = t_3__56_ ^ 1'b0;
  assign t_4__55_ = t_3__55_ ^ t_3__63_;
  assign t_4__54_ = t_3__54_ ^ t_3__62_;
  assign t_4__53_ = t_3__53_ ^ t_3__61_;
  assign t_4__52_ = t_3__52_ ^ t_3__60_;
  assign t_4__51_ = t_3__51_ ^ t_3__59_;
  assign t_4__50_ = t_3__50_ ^ t_3__58_;
  assign t_4__49_ = t_3__49_ ^ t_3__57_;
  assign t_4__48_ = t_3__48_ ^ t_3__56_;
  assign t_4__47_ = t_3__47_ ^ t_3__55_;
  assign t_4__46_ = t_3__46_ ^ t_3__54_;
  assign t_4__45_ = t_3__45_ ^ t_3__53_;
  assign t_4__44_ = t_3__44_ ^ t_3__52_;
  assign t_4__43_ = t_3__43_ ^ t_3__51_;
  assign t_4__42_ = t_3__42_ ^ t_3__50_;
  assign t_4__41_ = t_3__41_ ^ t_3__49_;
  assign t_4__40_ = t_3__40_ ^ t_3__48_;
  assign t_4__39_ = t_3__39_ ^ t_3__47_;
  assign t_4__38_ = t_3__38_ ^ t_3__46_;
  assign t_4__37_ = t_3__37_ ^ t_3__45_;
  assign t_4__36_ = t_3__36_ ^ t_3__44_;
  assign t_4__35_ = t_3__35_ ^ t_3__43_;
  assign t_4__34_ = t_3__34_ ^ t_3__42_;
  assign t_4__33_ = t_3__33_ ^ t_3__41_;
  assign t_4__32_ = t_3__32_ ^ t_3__40_;
  assign t_4__31_ = t_3__31_ ^ t_3__39_;
  assign t_4__30_ = t_3__30_ ^ t_3__38_;
  assign t_4__29_ = t_3__29_ ^ t_3__37_;
  assign t_4__28_ = t_3__28_ ^ t_3__36_;
  assign t_4__27_ = t_3__27_ ^ t_3__35_;
  assign t_4__26_ = t_3__26_ ^ t_3__34_;
  assign t_4__25_ = t_3__25_ ^ t_3__33_;
  assign t_4__24_ = t_3__24_ ^ t_3__32_;
  assign t_4__23_ = t_3__23_ ^ t_3__31_;
  assign t_4__22_ = t_3__22_ ^ t_3__30_;
  assign t_4__21_ = t_3__21_ ^ t_3__29_;
  assign t_4__20_ = t_3__20_ ^ t_3__28_;
  assign t_4__19_ = t_3__19_ ^ t_3__27_;
  assign t_4__18_ = t_3__18_ ^ t_3__26_;
  assign t_4__17_ = t_3__17_ ^ t_3__25_;
  assign t_4__16_ = t_3__16_ ^ t_3__24_;
  assign t_4__15_ = t_3__15_ ^ t_3__23_;
  assign t_4__14_ = t_3__14_ ^ t_3__22_;
  assign t_4__13_ = t_3__13_ ^ t_3__21_;
  assign t_4__12_ = t_3__12_ ^ t_3__20_;
  assign t_4__11_ = t_3__11_ ^ t_3__19_;
  assign t_4__10_ = t_3__10_ ^ t_3__18_;
  assign t_4__9_ = t_3__9_ ^ t_3__17_;
  assign t_4__8_ = t_3__8_ ^ t_3__16_;
  assign t_4__7_ = t_3__7_ ^ t_3__15_;
  assign t_4__6_ = t_3__6_ ^ t_3__14_;
  assign t_4__5_ = t_3__5_ ^ t_3__13_;
  assign t_4__4_ = t_3__4_ ^ t_3__12_;
  assign t_4__3_ = t_3__3_ ^ t_3__11_;
  assign t_4__2_ = t_3__2_ ^ t_3__10_;
  assign t_4__1_ = t_3__1_ ^ t_3__9_;
  assign t_4__0_ = t_3__0_ ^ t_3__8_;
  assign t_5__63_ = t_4__63_ ^ 1'b0;
  assign t_5__62_ = t_4__62_ ^ 1'b0;
  assign t_5__61_ = t_4__61_ ^ 1'b0;
  assign t_5__60_ = t_4__60_ ^ 1'b0;
  assign t_5__59_ = t_4__59_ ^ 1'b0;
  assign t_5__58_ = t_4__58_ ^ 1'b0;
  assign t_5__57_ = t_4__57_ ^ 1'b0;
  assign t_5__56_ = t_4__56_ ^ 1'b0;
  assign t_5__55_ = t_4__55_ ^ 1'b0;
  assign t_5__54_ = t_4__54_ ^ 1'b0;
  assign t_5__53_ = t_4__53_ ^ 1'b0;
  assign t_5__52_ = t_4__52_ ^ 1'b0;
  assign t_5__51_ = t_4__51_ ^ 1'b0;
  assign t_5__50_ = t_4__50_ ^ 1'b0;
  assign t_5__49_ = t_4__49_ ^ 1'b0;
  assign t_5__48_ = t_4__48_ ^ 1'b0;
  assign t_5__47_ = t_4__47_ ^ t_4__63_;
  assign t_5__46_ = t_4__46_ ^ t_4__62_;
  assign t_5__45_ = t_4__45_ ^ t_4__61_;
  assign t_5__44_ = t_4__44_ ^ t_4__60_;
  assign t_5__43_ = t_4__43_ ^ t_4__59_;
  assign t_5__42_ = t_4__42_ ^ t_4__58_;
  assign t_5__41_ = t_4__41_ ^ t_4__57_;
  assign t_5__40_ = t_4__40_ ^ t_4__56_;
  assign t_5__39_ = t_4__39_ ^ t_4__55_;
  assign t_5__38_ = t_4__38_ ^ t_4__54_;
  assign t_5__37_ = t_4__37_ ^ t_4__53_;
  assign t_5__36_ = t_4__36_ ^ t_4__52_;
  assign t_5__35_ = t_4__35_ ^ t_4__51_;
  assign t_5__34_ = t_4__34_ ^ t_4__50_;
  assign t_5__33_ = t_4__33_ ^ t_4__49_;
  assign t_5__32_ = t_4__32_ ^ t_4__48_;
  assign t_5__31_ = t_4__31_ ^ t_4__47_;
  assign t_5__30_ = t_4__30_ ^ t_4__46_;
  assign t_5__29_ = t_4__29_ ^ t_4__45_;
  assign t_5__28_ = t_4__28_ ^ t_4__44_;
  assign t_5__27_ = t_4__27_ ^ t_4__43_;
  assign t_5__26_ = t_4__26_ ^ t_4__42_;
  assign t_5__25_ = t_4__25_ ^ t_4__41_;
  assign t_5__24_ = t_4__24_ ^ t_4__40_;
  assign t_5__23_ = t_4__23_ ^ t_4__39_;
  assign t_5__22_ = t_4__22_ ^ t_4__38_;
  assign t_5__21_ = t_4__21_ ^ t_4__37_;
  assign t_5__20_ = t_4__20_ ^ t_4__36_;
  assign t_5__19_ = t_4__19_ ^ t_4__35_;
  assign t_5__18_ = t_4__18_ ^ t_4__34_;
  assign t_5__17_ = t_4__17_ ^ t_4__33_;
  assign t_5__16_ = t_4__16_ ^ t_4__32_;
  assign t_5__15_ = t_4__15_ ^ t_4__31_;
  assign t_5__14_ = t_4__14_ ^ t_4__30_;
  assign t_5__13_ = t_4__13_ ^ t_4__29_;
  assign t_5__12_ = t_4__12_ ^ t_4__28_;
  assign t_5__11_ = t_4__11_ ^ t_4__27_;
  assign t_5__10_ = t_4__10_ ^ t_4__26_;
  assign t_5__9_ = t_4__9_ ^ t_4__25_;
  assign t_5__8_ = t_4__8_ ^ t_4__24_;
  assign t_5__7_ = t_4__7_ ^ t_4__23_;
  assign t_5__6_ = t_4__6_ ^ t_4__22_;
  assign t_5__5_ = t_4__5_ ^ t_4__21_;
  assign t_5__4_ = t_4__4_ ^ t_4__20_;
  assign t_5__3_ = t_4__3_ ^ t_4__19_;
  assign t_5__2_ = t_4__2_ ^ t_4__18_;
  assign t_5__1_ = t_4__1_ ^ t_4__17_;
  assign t_5__0_ = t_4__0_ ^ t_4__16_;
  assign o[63] = t_5__63_ ^ 1'b0;
  assign o[62] = t_5__62_ ^ 1'b0;
  assign o[61] = t_5__61_ ^ 1'b0;
  assign o[60] = t_5__60_ ^ 1'b0;
  assign o[59] = t_5__59_ ^ 1'b0;
  assign o[58] = t_5__58_ ^ 1'b0;
  assign o[57] = t_5__57_ ^ 1'b0;
  assign o[56] = t_5__56_ ^ 1'b0;
  assign o[55] = t_5__55_ ^ 1'b0;
  assign o[54] = t_5__54_ ^ 1'b0;
  assign o[53] = t_5__53_ ^ 1'b0;
  assign o[52] = t_5__52_ ^ 1'b0;
  assign o[51] = t_5__51_ ^ 1'b0;
  assign o[50] = t_5__50_ ^ 1'b0;
  assign o[49] = t_5__49_ ^ 1'b0;
  assign o[48] = t_5__48_ ^ 1'b0;
  assign o[47] = t_5__47_ ^ 1'b0;
  assign o[46] = t_5__46_ ^ 1'b0;
  assign o[45] = t_5__45_ ^ 1'b0;
  assign o[44] = t_5__44_ ^ 1'b0;
  assign o[43] = t_5__43_ ^ 1'b0;
  assign o[42] = t_5__42_ ^ 1'b0;
  assign o[41] = t_5__41_ ^ 1'b0;
  assign o[40] = t_5__40_ ^ 1'b0;
  assign o[39] = t_5__39_ ^ 1'b0;
  assign o[38] = t_5__38_ ^ 1'b0;
  assign o[37] = t_5__37_ ^ 1'b0;
  assign o[36] = t_5__36_ ^ 1'b0;
  assign o[35] = t_5__35_ ^ 1'b0;
  assign o[34] = t_5__34_ ^ 1'b0;
  assign o[33] = t_5__33_ ^ 1'b0;
  assign o[32] = t_5__32_ ^ 1'b0;
  assign o[31] = t_5__31_ ^ t_5__63_;
  assign o[30] = t_5__30_ ^ t_5__62_;
  assign o[29] = t_5__29_ ^ t_5__61_;
  assign o[28] = t_5__28_ ^ t_5__60_;
  assign o[27] = t_5__27_ ^ t_5__59_;
  assign o[26] = t_5__26_ ^ t_5__58_;
  assign o[25] = t_5__25_ ^ t_5__57_;
  assign o[24] = t_5__24_ ^ t_5__56_;
  assign o[23] = t_5__23_ ^ t_5__55_;
  assign o[22] = t_5__22_ ^ t_5__54_;
  assign o[21] = t_5__21_ ^ t_5__53_;
  assign o[20] = t_5__20_ ^ t_5__52_;
  assign o[19] = t_5__19_ ^ t_5__51_;
  assign o[18] = t_5__18_ ^ t_5__50_;
  assign o[17] = t_5__17_ ^ t_5__49_;
  assign o[16] = t_5__16_ ^ t_5__48_;
  assign o[15] = t_5__15_ ^ t_5__47_;
  assign o[14] = t_5__14_ ^ t_5__46_;
  assign o[13] = t_5__13_ ^ t_5__45_;
  assign o[12] = t_5__12_ ^ t_5__44_;
  assign o[11] = t_5__11_ ^ t_5__43_;
  assign o[10] = t_5__10_ ^ t_5__42_;
  assign o[9] = t_5__9_ ^ t_5__41_;
  assign o[8] = t_5__8_ ^ t_5__40_;
  assign o[7] = t_5__7_ ^ t_5__39_;
  assign o[6] = t_5__6_ ^ t_5__38_;
  assign o[5] = t_5__5_ ^ t_5__37_;
  assign o[4] = t_5__4_ ^ t_5__36_;
  assign o[3] = t_5__3_ ^ t_5__35_;
  assign o[2] = t_5__2_ ^ t_5__34_;
  assign o[1] = t_5__1_ ^ t_5__33_;
  assign o[0] = t_5__0_ ^ t_5__32_;

endmodule



module bsg_gray_to_binary
(
  gray_i,
  binary_o
);

  input [63:0] gray_i;
  output [63:0] binary_o;
  wire [63:0] binary_o;

  bsg_scan_width_p64_xor_p1
  scan_xor
  (
    .i(gray_i),
    .o(binary_o)
  );


endmodule

