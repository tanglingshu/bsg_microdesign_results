

module top
(
  data_i,
  select_i,
  data_o
);

  input [1023:0] data_i;
  input [255:0] select_i;
  output [1023:0] data_o;

  bsg_permute_box
  wrapper
  (
    .data_i(data_i),
    .select_i(select_i),
    .data_o(data_o)
  );


endmodule



module bsg_permute_box
(
  data_i,
  select_i,
  data_o
);

  input [1023:0] data_i;
  input [255:0] select_i;
  output [1023:0] data_o;
  wire [1023:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119;
  assign data_o[127] = (N7)? data_i[127] : 
                       (N9)? data_i[255] : 
                       (N11)? data_i[383] : 
                       (N13)? data_i[511] : 
                       (N8)? data_i[639] : 
                       (N10)? data_i[767] : 
                       (N12)? data_i[895] : 
                       (N14)? data_i[1023] : 1'b0;
  assign data_o[126] = (N7)? data_i[126] : 
                       (N9)? data_i[254] : 
                       (N11)? data_i[382] : 
                       (N13)? data_i[510] : 
                       (N8)? data_i[638] : 
                       (N10)? data_i[766] : 
                       (N12)? data_i[894] : 
                       (N14)? data_i[1022] : 1'b0;
  assign data_o[125] = (N7)? data_i[125] : 
                       (N9)? data_i[253] : 
                       (N11)? data_i[381] : 
                       (N13)? data_i[509] : 
                       (N8)? data_i[637] : 
                       (N10)? data_i[765] : 
                       (N12)? data_i[893] : 
                       (N14)? data_i[1021] : 1'b0;
  assign data_o[124] = (N7)? data_i[124] : 
                       (N9)? data_i[252] : 
                       (N11)? data_i[380] : 
                       (N13)? data_i[508] : 
                       (N8)? data_i[636] : 
                       (N10)? data_i[764] : 
                       (N12)? data_i[892] : 
                       (N14)? data_i[1020] : 1'b0;
  assign data_o[123] = (N7)? data_i[123] : 
                       (N9)? data_i[251] : 
                       (N11)? data_i[379] : 
                       (N13)? data_i[507] : 
                       (N8)? data_i[635] : 
                       (N10)? data_i[763] : 
                       (N12)? data_i[891] : 
                       (N14)? data_i[1019] : 1'b0;
  assign data_o[122] = (N7)? data_i[122] : 
                       (N9)? data_i[250] : 
                       (N11)? data_i[378] : 
                       (N13)? data_i[506] : 
                       (N8)? data_i[634] : 
                       (N10)? data_i[762] : 
                       (N12)? data_i[890] : 
                       (N14)? data_i[1018] : 1'b0;
  assign data_o[121] = (N7)? data_i[121] : 
                       (N9)? data_i[249] : 
                       (N11)? data_i[377] : 
                       (N13)? data_i[505] : 
                       (N8)? data_i[633] : 
                       (N10)? data_i[761] : 
                       (N12)? data_i[889] : 
                       (N14)? data_i[1017] : 1'b0;
  assign data_o[120] = (N7)? data_i[120] : 
                       (N9)? data_i[248] : 
                       (N11)? data_i[376] : 
                       (N13)? data_i[504] : 
                       (N8)? data_i[632] : 
                       (N10)? data_i[760] : 
                       (N12)? data_i[888] : 
                       (N14)? data_i[1016] : 1'b0;
  assign data_o[119] = (N7)? data_i[119] : 
                       (N9)? data_i[247] : 
                       (N11)? data_i[375] : 
                       (N13)? data_i[503] : 
                       (N8)? data_i[631] : 
                       (N10)? data_i[759] : 
                       (N12)? data_i[887] : 
                       (N14)? data_i[1015] : 1'b0;
  assign data_o[118] = (N7)? data_i[118] : 
                       (N9)? data_i[246] : 
                       (N11)? data_i[374] : 
                       (N13)? data_i[502] : 
                       (N8)? data_i[630] : 
                       (N10)? data_i[758] : 
                       (N12)? data_i[886] : 
                       (N14)? data_i[1014] : 1'b0;
  assign data_o[117] = (N7)? data_i[117] : 
                       (N9)? data_i[245] : 
                       (N11)? data_i[373] : 
                       (N13)? data_i[501] : 
                       (N8)? data_i[629] : 
                       (N10)? data_i[757] : 
                       (N12)? data_i[885] : 
                       (N14)? data_i[1013] : 1'b0;
  assign data_o[116] = (N7)? data_i[116] : 
                       (N9)? data_i[244] : 
                       (N11)? data_i[372] : 
                       (N13)? data_i[500] : 
                       (N8)? data_i[628] : 
                       (N10)? data_i[756] : 
                       (N12)? data_i[884] : 
                       (N14)? data_i[1012] : 1'b0;
  assign data_o[115] = (N7)? data_i[115] : 
                       (N9)? data_i[243] : 
                       (N11)? data_i[371] : 
                       (N13)? data_i[499] : 
                       (N8)? data_i[627] : 
                       (N10)? data_i[755] : 
                       (N12)? data_i[883] : 
                       (N14)? data_i[1011] : 1'b0;
  assign data_o[114] = (N7)? data_i[114] : 
                       (N9)? data_i[242] : 
                       (N11)? data_i[370] : 
                       (N13)? data_i[498] : 
                       (N8)? data_i[626] : 
                       (N10)? data_i[754] : 
                       (N12)? data_i[882] : 
                       (N14)? data_i[1010] : 1'b0;
  assign data_o[113] = (N7)? data_i[113] : 
                       (N9)? data_i[241] : 
                       (N11)? data_i[369] : 
                       (N13)? data_i[497] : 
                       (N8)? data_i[625] : 
                       (N10)? data_i[753] : 
                       (N12)? data_i[881] : 
                       (N14)? data_i[1009] : 1'b0;
  assign data_o[112] = (N7)? data_i[112] : 
                       (N9)? data_i[240] : 
                       (N11)? data_i[368] : 
                       (N13)? data_i[496] : 
                       (N8)? data_i[624] : 
                       (N10)? data_i[752] : 
                       (N12)? data_i[880] : 
                       (N14)? data_i[1008] : 1'b0;
  assign data_o[111] = (N7)? data_i[111] : 
                       (N9)? data_i[239] : 
                       (N11)? data_i[367] : 
                       (N13)? data_i[495] : 
                       (N8)? data_i[623] : 
                       (N10)? data_i[751] : 
                       (N12)? data_i[879] : 
                       (N14)? data_i[1007] : 1'b0;
  assign data_o[110] = (N7)? data_i[110] : 
                       (N9)? data_i[238] : 
                       (N11)? data_i[366] : 
                       (N13)? data_i[494] : 
                       (N8)? data_i[622] : 
                       (N10)? data_i[750] : 
                       (N12)? data_i[878] : 
                       (N14)? data_i[1006] : 1'b0;
  assign data_o[109] = (N7)? data_i[109] : 
                       (N9)? data_i[237] : 
                       (N11)? data_i[365] : 
                       (N13)? data_i[493] : 
                       (N8)? data_i[621] : 
                       (N10)? data_i[749] : 
                       (N12)? data_i[877] : 
                       (N14)? data_i[1005] : 1'b0;
  assign data_o[108] = (N7)? data_i[108] : 
                       (N9)? data_i[236] : 
                       (N11)? data_i[364] : 
                       (N13)? data_i[492] : 
                       (N8)? data_i[620] : 
                       (N10)? data_i[748] : 
                       (N12)? data_i[876] : 
                       (N14)? data_i[1004] : 1'b0;
  assign data_o[107] = (N7)? data_i[107] : 
                       (N9)? data_i[235] : 
                       (N11)? data_i[363] : 
                       (N13)? data_i[491] : 
                       (N8)? data_i[619] : 
                       (N10)? data_i[747] : 
                       (N12)? data_i[875] : 
                       (N14)? data_i[1003] : 1'b0;
  assign data_o[106] = (N7)? data_i[106] : 
                       (N9)? data_i[234] : 
                       (N11)? data_i[362] : 
                       (N13)? data_i[490] : 
                       (N8)? data_i[618] : 
                       (N10)? data_i[746] : 
                       (N12)? data_i[874] : 
                       (N14)? data_i[1002] : 1'b0;
  assign data_o[105] = (N7)? data_i[105] : 
                       (N9)? data_i[233] : 
                       (N11)? data_i[361] : 
                       (N13)? data_i[489] : 
                       (N8)? data_i[617] : 
                       (N10)? data_i[745] : 
                       (N12)? data_i[873] : 
                       (N14)? data_i[1001] : 1'b0;
  assign data_o[104] = (N7)? data_i[104] : 
                       (N9)? data_i[232] : 
                       (N11)? data_i[360] : 
                       (N13)? data_i[488] : 
                       (N8)? data_i[616] : 
                       (N10)? data_i[744] : 
                       (N12)? data_i[872] : 
                       (N14)? data_i[1000] : 1'b0;
  assign data_o[103] = (N7)? data_i[103] : 
                       (N9)? data_i[231] : 
                       (N11)? data_i[359] : 
                       (N13)? data_i[487] : 
                       (N8)? data_i[615] : 
                       (N10)? data_i[743] : 
                       (N12)? data_i[871] : 
                       (N14)? data_i[999] : 1'b0;
  assign data_o[102] = (N7)? data_i[102] : 
                       (N9)? data_i[230] : 
                       (N11)? data_i[358] : 
                       (N13)? data_i[486] : 
                       (N8)? data_i[614] : 
                       (N10)? data_i[742] : 
                       (N12)? data_i[870] : 
                       (N14)? data_i[998] : 1'b0;
  assign data_o[101] = (N7)? data_i[101] : 
                       (N9)? data_i[229] : 
                       (N11)? data_i[357] : 
                       (N13)? data_i[485] : 
                       (N8)? data_i[613] : 
                       (N10)? data_i[741] : 
                       (N12)? data_i[869] : 
                       (N14)? data_i[997] : 1'b0;
  assign data_o[100] = (N7)? data_i[100] : 
                       (N9)? data_i[228] : 
                       (N11)? data_i[356] : 
                       (N13)? data_i[484] : 
                       (N8)? data_i[612] : 
                       (N10)? data_i[740] : 
                       (N12)? data_i[868] : 
                       (N14)? data_i[996] : 1'b0;
  assign data_o[99] = (N7)? data_i[99] : 
                      (N9)? data_i[227] : 
                      (N11)? data_i[355] : 
                      (N13)? data_i[483] : 
                      (N8)? data_i[611] : 
                      (N10)? data_i[739] : 
                      (N12)? data_i[867] : 
                      (N14)? data_i[995] : 1'b0;
  assign data_o[98] = (N7)? data_i[98] : 
                      (N9)? data_i[226] : 
                      (N11)? data_i[354] : 
                      (N13)? data_i[482] : 
                      (N8)? data_i[610] : 
                      (N10)? data_i[738] : 
                      (N12)? data_i[866] : 
                      (N14)? data_i[994] : 1'b0;
  assign data_o[97] = (N7)? data_i[97] : 
                      (N9)? data_i[225] : 
                      (N11)? data_i[353] : 
                      (N13)? data_i[481] : 
                      (N8)? data_i[609] : 
                      (N10)? data_i[737] : 
                      (N12)? data_i[865] : 
                      (N14)? data_i[993] : 1'b0;
  assign data_o[96] = (N7)? data_i[96] : 
                      (N9)? data_i[224] : 
                      (N11)? data_i[352] : 
                      (N13)? data_i[480] : 
                      (N8)? data_i[608] : 
                      (N10)? data_i[736] : 
                      (N12)? data_i[864] : 
                      (N14)? data_i[992] : 1'b0;
  assign data_o[95] = (N7)? data_i[95] : 
                      (N9)? data_i[223] : 
                      (N11)? data_i[351] : 
                      (N13)? data_i[479] : 
                      (N8)? data_i[607] : 
                      (N10)? data_i[735] : 
                      (N12)? data_i[863] : 
                      (N14)? data_i[991] : 1'b0;
  assign data_o[94] = (N7)? data_i[94] : 
                      (N9)? data_i[222] : 
                      (N11)? data_i[350] : 
                      (N13)? data_i[478] : 
                      (N8)? data_i[606] : 
                      (N10)? data_i[734] : 
                      (N12)? data_i[862] : 
                      (N14)? data_i[990] : 1'b0;
  assign data_o[93] = (N7)? data_i[93] : 
                      (N9)? data_i[221] : 
                      (N11)? data_i[349] : 
                      (N13)? data_i[477] : 
                      (N8)? data_i[605] : 
                      (N10)? data_i[733] : 
                      (N12)? data_i[861] : 
                      (N14)? data_i[989] : 1'b0;
  assign data_o[92] = (N7)? data_i[92] : 
                      (N9)? data_i[220] : 
                      (N11)? data_i[348] : 
                      (N13)? data_i[476] : 
                      (N8)? data_i[604] : 
                      (N10)? data_i[732] : 
                      (N12)? data_i[860] : 
                      (N14)? data_i[988] : 1'b0;
  assign data_o[91] = (N7)? data_i[91] : 
                      (N9)? data_i[219] : 
                      (N11)? data_i[347] : 
                      (N13)? data_i[475] : 
                      (N8)? data_i[603] : 
                      (N10)? data_i[731] : 
                      (N12)? data_i[859] : 
                      (N14)? data_i[987] : 1'b0;
  assign data_o[90] = (N7)? data_i[90] : 
                      (N9)? data_i[218] : 
                      (N11)? data_i[346] : 
                      (N13)? data_i[474] : 
                      (N8)? data_i[602] : 
                      (N10)? data_i[730] : 
                      (N12)? data_i[858] : 
                      (N14)? data_i[986] : 1'b0;
  assign data_o[89] = (N7)? data_i[89] : 
                      (N9)? data_i[217] : 
                      (N11)? data_i[345] : 
                      (N13)? data_i[473] : 
                      (N8)? data_i[601] : 
                      (N10)? data_i[729] : 
                      (N12)? data_i[857] : 
                      (N14)? data_i[985] : 1'b0;
  assign data_o[88] = (N7)? data_i[88] : 
                      (N9)? data_i[216] : 
                      (N11)? data_i[344] : 
                      (N13)? data_i[472] : 
                      (N8)? data_i[600] : 
                      (N10)? data_i[728] : 
                      (N12)? data_i[856] : 
                      (N14)? data_i[984] : 1'b0;
  assign data_o[87] = (N7)? data_i[87] : 
                      (N9)? data_i[215] : 
                      (N11)? data_i[343] : 
                      (N13)? data_i[471] : 
                      (N8)? data_i[599] : 
                      (N10)? data_i[727] : 
                      (N12)? data_i[855] : 
                      (N14)? data_i[983] : 1'b0;
  assign data_o[86] = (N7)? data_i[86] : 
                      (N9)? data_i[214] : 
                      (N11)? data_i[342] : 
                      (N13)? data_i[470] : 
                      (N8)? data_i[598] : 
                      (N10)? data_i[726] : 
                      (N12)? data_i[854] : 
                      (N14)? data_i[982] : 1'b0;
  assign data_o[85] = (N7)? data_i[85] : 
                      (N9)? data_i[213] : 
                      (N11)? data_i[341] : 
                      (N13)? data_i[469] : 
                      (N8)? data_i[597] : 
                      (N10)? data_i[725] : 
                      (N12)? data_i[853] : 
                      (N14)? data_i[981] : 1'b0;
  assign data_o[84] = (N7)? data_i[84] : 
                      (N9)? data_i[212] : 
                      (N11)? data_i[340] : 
                      (N13)? data_i[468] : 
                      (N8)? data_i[596] : 
                      (N10)? data_i[724] : 
                      (N12)? data_i[852] : 
                      (N14)? data_i[980] : 1'b0;
  assign data_o[83] = (N7)? data_i[83] : 
                      (N9)? data_i[211] : 
                      (N11)? data_i[339] : 
                      (N13)? data_i[467] : 
                      (N8)? data_i[595] : 
                      (N10)? data_i[723] : 
                      (N12)? data_i[851] : 
                      (N14)? data_i[979] : 1'b0;
  assign data_o[82] = (N7)? data_i[82] : 
                      (N9)? data_i[210] : 
                      (N11)? data_i[338] : 
                      (N13)? data_i[466] : 
                      (N8)? data_i[594] : 
                      (N10)? data_i[722] : 
                      (N12)? data_i[850] : 
                      (N14)? data_i[978] : 1'b0;
  assign data_o[81] = (N7)? data_i[81] : 
                      (N9)? data_i[209] : 
                      (N11)? data_i[337] : 
                      (N13)? data_i[465] : 
                      (N8)? data_i[593] : 
                      (N10)? data_i[721] : 
                      (N12)? data_i[849] : 
                      (N14)? data_i[977] : 1'b0;
  assign data_o[80] = (N7)? data_i[80] : 
                      (N9)? data_i[208] : 
                      (N11)? data_i[336] : 
                      (N13)? data_i[464] : 
                      (N8)? data_i[592] : 
                      (N10)? data_i[720] : 
                      (N12)? data_i[848] : 
                      (N14)? data_i[976] : 1'b0;
  assign data_o[79] = (N7)? data_i[79] : 
                      (N9)? data_i[207] : 
                      (N11)? data_i[335] : 
                      (N13)? data_i[463] : 
                      (N8)? data_i[591] : 
                      (N10)? data_i[719] : 
                      (N12)? data_i[847] : 
                      (N14)? data_i[975] : 1'b0;
  assign data_o[78] = (N7)? data_i[78] : 
                      (N9)? data_i[206] : 
                      (N11)? data_i[334] : 
                      (N13)? data_i[462] : 
                      (N8)? data_i[590] : 
                      (N10)? data_i[718] : 
                      (N12)? data_i[846] : 
                      (N14)? data_i[974] : 1'b0;
  assign data_o[77] = (N7)? data_i[77] : 
                      (N9)? data_i[205] : 
                      (N11)? data_i[333] : 
                      (N13)? data_i[461] : 
                      (N8)? data_i[589] : 
                      (N10)? data_i[717] : 
                      (N12)? data_i[845] : 
                      (N14)? data_i[973] : 1'b0;
  assign data_o[76] = (N7)? data_i[76] : 
                      (N9)? data_i[204] : 
                      (N11)? data_i[332] : 
                      (N13)? data_i[460] : 
                      (N8)? data_i[588] : 
                      (N10)? data_i[716] : 
                      (N12)? data_i[844] : 
                      (N14)? data_i[972] : 1'b0;
  assign data_o[75] = (N7)? data_i[75] : 
                      (N9)? data_i[203] : 
                      (N11)? data_i[331] : 
                      (N13)? data_i[459] : 
                      (N8)? data_i[587] : 
                      (N10)? data_i[715] : 
                      (N12)? data_i[843] : 
                      (N14)? data_i[971] : 1'b0;
  assign data_o[74] = (N7)? data_i[74] : 
                      (N9)? data_i[202] : 
                      (N11)? data_i[330] : 
                      (N13)? data_i[458] : 
                      (N8)? data_i[586] : 
                      (N10)? data_i[714] : 
                      (N12)? data_i[842] : 
                      (N14)? data_i[970] : 1'b0;
  assign data_o[73] = (N7)? data_i[73] : 
                      (N9)? data_i[201] : 
                      (N11)? data_i[329] : 
                      (N13)? data_i[457] : 
                      (N8)? data_i[585] : 
                      (N10)? data_i[713] : 
                      (N12)? data_i[841] : 
                      (N14)? data_i[969] : 1'b0;
  assign data_o[72] = (N7)? data_i[72] : 
                      (N9)? data_i[200] : 
                      (N11)? data_i[328] : 
                      (N13)? data_i[456] : 
                      (N8)? data_i[584] : 
                      (N10)? data_i[712] : 
                      (N12)? data_i[840] : 
                      (N14)? data_i[968] : 1'b0;
  assign data_o[71] = (N7)? data_i[71] : 
                      (N9)? data_i[199] : 
                      (N11)? data_i[327] : 
                      (N13)? data_i[455] : 
                      (N8)? data_i[583] : 
                      (N10)? data_i[711] : 
                      (N12)? data_i[839] : 
                      (N14)? data_i[967] : 1'b0;
  assign data_o[70] = (N7)? data_i[70] : 
                      (N9)? data_i[198] : 
                      (N11)? data_i[326] : 
                      (N13)? data_i[454] : 
                      (N8)? data_i[582] : 
                      (N10)? data_i[710] : 
                      (N12)? data_i[838] : 
                      (N14)? data_i[966] : 1'b0;
  assign data_o[69] = (N7)? data_i[69] : 
                      (N9)? data_i[197] : 
                      (N11)? data_i[325] : 
                      (N13)? data_i[453] : 
                      (N8)? data_i[581] : 
                      (N10)? data_i[709] : 
                      (N12)? data_i[837] : 
                      (N14)? data_i[965] : 1'b0;
  assign data_o[68] = (N7)? data_i[68] : 
                      (N9)? data_i[196] : 
                      (N11)? data_i[324] : 
                      (N13)? data_i[452] : 
                      (N8)? data_i[580] : 
                      (N10)? data_i[708] : 
                      (N12)? data_i[836] : 
                      (N14)? data_i[964] : 1'b0;
  assign data_o[67] = (N7)? data_i[67] : 
                      (N9)? data_i[195] : 
                      (N11)? data_i[323] : 
                      (N13)? data_i[451] : 
                      (N8)? data_i[579] : 
                      (N10)? data_i[707] : 
                      (N12)? data_i[835] : 
                      (N14)? data_i[963] : 1'b0;
  assign data_o[66] = (N7)? data_i[66] : 
                      (N9)? data_i[194] : 
                      (N11)? data_i[322] : 
                      (N13)? data_i[450] : 
                      (N8)? data_i[578] : 
                      (N10)? data_i[706] : 
                      (N12)? data_i[834] : 
                      (N14)? data_i[962] : 1'b0;
  assign data_o[65] = (N7)? data_i[65] : 
                      (N9)? data_i[193] : 
                      (N11)? data_i[321] : 
                      (N13)? data_i[449] : 
                      (N8)? data_i[577] : 
                      (N10)? data_i[705] : 
                      (N12)? data_i[833] : 
                      (N14)? data_i[961] : 1'b0;
  assign data_o[64] = (N7)? data_i[64] : 
                      (N9)? data_i[192] : 
                      (N11)? data_i[320] : 
                      (N13)? data_i[448] : 
                      (N8)? data_i[576] : 
                      (N10)? data_i[704] : 
                      (N12)? data_i[832] : 
                      (N14)? data_i[960] : 1'b0;
  assign data_o[63] = (N7)? data_i[63] : 
                      (N9)? data_i[191] : 
                      (N11)? data_i[319] : 
                      (N13)? data_i[447] : 
                      (N8)? data_i[575] : 
                      (N10)? data_i[703] : 
                      (N12)? data_i[831] : 
                      (N14)? data_i[959] : 1'b0;
  assign data_o[62] = (N7)? data_i[62] : 
                      (N9)? data_i[190] : 
                      (N11)? data_i[318] : 
                      (N13)? data_i[446] : 
                      (N8)? data_i[574] : 
                      (N10)? data_i[702] : 
                      (N12)? data_i[830] : 
                      (N14)? data_i[958] : 1'b0;
  assign data_o[61] = (N7)? data_i[61] : 
                      (N9)? data_i[189] : 
                      (N11)? data_i[317] : 
                      (N13)? data_i[445] : 
                      (N8)? data_i[573] : 
                      (N10)? data_i[701] : 
                      (N12)? data_i[829] : 
                      (N14)? data_i[957] : 1'b0;
  assign data_o[60] = (N7)? data_i[60] : 
                      (N9)? data_i[188] : 
                      (N11)? data_i[316] : 
                      (N13)? data_i[444] : 
                      (N8)? data_i[572] : 
                      (N10)? data_i[700] : 
                      (N12)? data_i[828] : 
                      (N14)? data_i[956] : 1'b0;
  assign data_o[59] = (N7)? data_i[59] : 
                      (N9)? data_i[187] : 
                      (N11)? data_i[315] : 
                      (N13)? data_i[443] : 
                      (N8)? data_i[571] : 
                      (N10)? data_i[699] : 
                      (N12)? data_i[827] : 
                      (N14)? data_i[955] : 1'b0;
  assign data_o[58] = (N7)? data_i[58] : 
                      (N9)? data_i[186] : 
                      (N11)? data_i[314] : 
                      (N13)? data_i[442] : 
                      (N8)? data_i[570] : 
                      (N10)? data_i[698] : 
                      (N12)? data_i[826] : 
                      (N14)? data_i[954] : 1'b0;
  assign data_o[57] = (N7)? data_i[57] : 
                      (N9)? data_i[185] : 
                      (N11)? data_i[313] : 
                      (N13)? data_i[441] : 
                      (N8)? data_i[569] : 
                      (N10)? data_i[697] : 
                      (N12)? data_i[825] : 
                      (N14)? data_i[953] : 1'b0;
  assign data_o[56] = (N7)? data_i[56] : 
                      (N9)? data_i[184] : 
                      (N11)? data_i[312] : 
                      (N13)? data_i[440] : 
                      (N8)? data_i[568] : 
                      (N10)? data_i[696] : 
                      (N12)? data_i[824] : 
                      (N14)? data_i[952] : 1'b0;
  assign data_o[55] = (N7)? data_i[55] : 
                      (N9)? data_i[183] : 
                      (N11)? data_i[311] : 
                      (N13)? data_i[439] : 
                      (N8)? data_i[567] : 
                      (N10)? data_i[695] : 
                      (N12)? data_i[823] : 
                      (N14)? data_i[951] : 1'b0;
  assign data_o[54] = (N7)? data_i[54] : 
                      (N9)? data_i[182] : 
                      (N11)? data_i[310] : 
                      (N13)? data_i[438] : 
                      (N8)? data_i[566] : 
                      (N10)? data_i[694] : 
                      (N12)? data_i[822] : 
                      (N14)? data_i[950] : 1'b0;
  assign data_o[53] = (N7)? data_i[53] : 
                      (N9)? data_i[181] : 
                      (N11)? data_i[309] : 
                      (N13)? data_i[437] : 
                      (N8)? data_i[565] : 
                      (N10)? data_i[693] : 
                      (N12)? data_i[821] : 
                      (N14)? data_i[949] : 1'b0;
  assign data_o[52] = (N7)? data_i[52] : 
                      (N9)? data_i[180] : 
                      (N11)? data_i[308] : 
                      (N13)? data_i[436] : 
                      (N8)? data_i[564] : 
                      (N10)? data_i[692] : 
                      (N12)? data_i[820] : 
                      (N14)? data_i[948] : 1'b0;
  assign data_o[51] = (N7)? data_i[51] : 
                      (N9)? data_i[179] : 
                      (N11)? data_i[307] : 
                      (N13)? data_i[435] : 
                      (N8)? data_i[563] : 
                      (N10)? data_i[691] : 
                      (N12)? data_i[819] : 
                      (N14)? data_i[947] : 1'b0;
  assign data_o[50] = (N7)? data_i[50] : 
                      (N9)? data_i[178] : 
                      (N11)? data_i[306] : 
                      (N13)? data_i[434] : 
                      (N8)? data_i[562] : 
                      (N10)? data_i[690] : 
                      (N12)? data_i[818] : 
                      (N14)? data_i[946] : 1'b0;
  assign data_o[49] = (N7)? data_i[49] : 
                      (N9)? data_i[177] : 
                      (N11)? data_i[305] : 
                      (N13)? data_i[433] : 
                      (N8)? data_i[561] : 
                      (N10)? data_i[689] : 
                      (N12)? data_i[817] : 
                      (N14)? data_i[945] : 1'b0;
  assign data_o[48] = (N7)? data_i[48] : 
                      (N9)? data_i[176] : 
                      (N11)? data_i[304] : 
                      (N13)? data_i[432] : 
                      (N8)? data_i[560] : 
                      (N10)? data_i[688] : 
                      (N12)? data_i[816] : 
                      (N14)? data_i[944] : 1'b0;
  assign data_o[47] = (N7)? data_i[47] : 
                      (N9)? data_i[175] : 
                      (N11)? data_i[303] : 
                      (N13)? data_i[431] : 
                      (N8)? data_i[559] : 
                      (N10)? data_i[687] : 
                      (N12)? data_i[815] : 
                      (N14)? data_i[943] : 1'b0;
  assign data_o[46] = (N7)? data_i[46] : 
                      (N9)? data_i[174] : 
                      (N11)? data_i[302] : 
                      (N13)? data_i[430] : 
                      (N8)? data_i[558] : 
                      (N10)? data_i[686] : 
                      (N12)? data_i[814] : 
                      (N14)? data_i[942] : 1'b0;
  assign data_o[45] = (N7)? data_i[45] : 
                      (N9)? data_i[173] : 
                      (N11)? data_i[301] : 
                      (N13)? data_i[429] : 
                      (N8)? data_i[557] : 
                      (N10)? data_i[685] : 
                      (N12)? data_i[813] : 
                      (N14)? data_i[941] : 1'b0;
  assign data_o[44] = (N7)? data_i[44] : 
                      (N9)? data_i[172] : 
                      (N11)? data_i[300] : 
                      (N13)? data_i[428] : 
                      (N8)? data_i[556] : 
                      (N10)? data_i[684] : 
                      (N12)? data_i[812] : 
                      (N14)? data_i[940] : 1'b0;
  assign data_o[43] = (N7)? data_i[43] : 
                      (N9)? data_i[171] : 
                      (N11)? data_i[299] : 
                      (N13)? data_i[427] : 
                      (N8)? data_i[555] : 
                      (N10)? data_i[683] : 
                      (N12)? data_i[811] : 
                      (N14)? data_i[939] : 1'b0;
  assign data_o[42] = (N7)? data_i[42] : 
                      (N9)? data_i[170] : 
                      (N11)? data_i[298] : 
                      (N13)? data_i[426] : 
                      (N8)? data_i[554] : 
                      (N10)? data_i[682] : 
                      (N12)? data_i[810] : 
                      (N14)? data_i[938] : 1'b0;
  assign data_o[41] = (N7)? data_i[41] : 
                      (N9)? data_i[169] : 
                      (N11)? data_i[297] : 
                      (N13)? data_i[425] : 
                      (N8)? data_i[553] : 
                      (N10)? data_i[681] : 
                      (N12)? data_i[809] : 
                      (N14)? data_i[937] : 1'b0;
  assign data_o[40] = (N7)? data_i[40] : 
                      (N9)? data_i[168] : 
                      (N11)? data_i[296] : 
                      (N13)? data_i[424] : 
                      (N8)? data_i[552] : 
                      (N10)? data_i[680] : 
                      (N12)? data_i[808] : 
                      (N14)? data_i[936] : 1'b0;
  assign data_o[39] = (N7)? data_i[39] : 
                      (N9)? data_i[167] : 
                      (N11)? data_i[295] : 
                      (N13)? data_i[423] : 
                      (N8)? data_i[551] : 
                      (N10)? data_i[679] : 
                      (N12)? data_i[807] : 
                      (N14)? data_i[935] : 1'b0;
  assign data_o[38] = (N7)? data_i[38] : 
                      (N9)? data_i[166] : 
                      (N11)? data_i[294] : 
                      (N13)? data_i[422] : 
                      (N8)? data_i[550] : 
                      (N10)? data_i[678] : 
                      (N12)? data_i[806] : 
                      (N14)? data_i[934] : 1'b0;
  assign data_o[37] = (N7)? data_i[37] : 
                      (N9)? data_i[165] : 
                      (N11)? data_i[293] : 
                      (N13)? data_i[421] : 
                      (N8)? data_i[549] : 
                      (N10)? data_i[677] : 
                      (N12)? data_i[805] : 
                      (N14)? data_i[933] : 1'b0;
  assign data_o[36] = (N7)? data_i[36] : 
                      (N9)? data_i[164] : 
                      (N11)? data_i[292] : 
                      (N13)? data_i[420] : 
                      (N8)? data_i[548] : 
                      (N10)? data_i[676] : 
                      (N12)? data_i[804] : 
                      (N14)? data_i[932] : 1'b0;
  assign data_o[35] = (N7)? data_i[35] : 
                      (N9)? data_i[163] : 
                      (N11)? data_i[291] : 
                      (N13)? data_i[419] : 
                      (N8)? data_i[547] : 
                      (N10)? data_i[675] : 
                      (N12)? data_i[803] : 
                      (N14)? data_i[931] : 1'b0;
  assign data_o[34] = (N7)? data_i[34] : 
                      (N9)? data_i[162] : 
                      (N11)? data_i[290] : 
                      (N13)? data_i[418] : 
                      (N8)? data_i[546] : 
                      (N10)? data_i[674] : 
                      (N12)? data_i[802] : 
                      (N14)? data_i[930] : 1'b0;
  assign data_o[33] = (N7)? data_i[33] : 
                      (N9)? data_i[161] : 
                      (N11)? data_i[289] : 
                      (N13)? data_i[417] : 
                      (N8)? data_i[545] : 
                      (N10)? data_i[673] : 
                      (N12)? data_i[801] : 
                      (N14)? data_i[929] : 1'b0;
  assign data_o[32] = (N7)? data_i[32] : 
                      (N9)? data_i[160] : 
                      (N11)? data_i[288] : 
                      (N13)? data_i[416] : 
                      (N8)? data_i[544] : 
                      (N10)? data_i[672] : 
                      (N12)? data_i[800] : 
                      (N14)? data_i[928] : 1'b0;
  assign data_o[31] = (N7)? data_i[31] : 
                      (N9)? data_i[159] : 
                      (N11)? data_i[287] : 
                      (N13)? data_i[415] : 
                      (N8)? data_i[543] : 
                      (N10)? data_i[671] : 
                      (N12)? data_i[799] : 
                      (N14)? data_i[927] : 1'b0;
  assign data_o[30] = (N7)? data_i[30] : 
                      (N9)? data_i[158] : 
                      (N11)? data_i[286] : 
                      (N13)? data_i[414] : 
                      (N8)? data_i[542] : 
                      (N10)? data_i[670] : 
                      (N12)? data_i[798] : 
                      (N14)? data_i[926] : 1'b0;
  assign data_o[29] = (N7)? data_i[29] : 
                      (N9)? data_i[157] : 
                      (N11)? data_i[285] : 
                      (N13)? data_i[413] : 
                      (N8)? data_i[541] : 
                      (N10)? data_i[669] : 
                      (N12)? data_i[797] : 
                      (N14)? data_i[925] : 1'b0;
  assign data_o[28] = (N7)? data_i[28] : 
                      (N9)? data_i[156] : 
                      (N11)? data_i[284] : 
                      (N13)? data_i[412] : 
                      (N8)? data_i[540] : 
                      (N10)? data_i[668] : 
                      (N12)? data_i[796] : 
                      (N14)? data_i[924] : 1'b0;
  assign data_o[27] = (N7)? data_i[27] : 
                      (N9)? data_i[155] : 
                      (N11)? data_i[283] : 
                      (N13)? data_i[411] : 
                      (N8)? data_i[539] : 
                      (N10)? data_i[667] : 
                      (N12)? data_i[795] : 
                      (N14)? data_i[923] : 1'b0;
  assign data_o[26] = (N7)? data_i[26] : 
                      (N9)? data_i[154] : 
                      (N11)? data_i[282] : 
                      (N13)? data_i[410] : 
                      (N8)? data_i[538] : 
                      (N10)? data_i[666] : 
                      (N12)? data_i[794] : 
                      (N14)? data_i[922] : 1'b0;
  assign data_o[25] = (N7)? data_i[25] : 
                      (N9)? data_i[153] : 
                      (N11)? data_i[281] : 
                      (N13)? data_i[409] : 
                      (N8)? data_i[537] : 
                      (N10)? data_i[665] : 
                      (N12)? data_i[793] : 
                      (N14)? data_i[921] : 1'b0;
  assign data_o[24] = (N7)? data_i[24] : 
                      (N9)? data_i[152] : 
                      (N11)? data_i[280] : 
                      (N13)? data_i[408] : 
                      (N8)? data_i[536] : 
                      (N10)? data_i[664] : 
                      (N12)? data_i[792] : 
                      (N14)? data_i[920] : 1'b0;
  assign data_o[23] = (N7)? data_i[23] : 
                      (N9)? data_i[151] : 
                      (N11)? data_i[279] : 
                      (N13)? data_i[407] : 
                      (N8)? data_i[535] : 
                      (N10)? data_i[663] : 
                      (N12)? data_i[791] : 
                      (N14)? data_i[919] : 1'b0;
  assign data_o[22] = (N7)? data_i[22] : 
                      (N9)? data_i[150] : 
                      (N11)? data_i[278] : 
                      (N13)? data_i[406] : 
                      (N8)? data_i[534] : 
                      (N10)? data_i[662] : 
                      (N12)? data_i[790] : 
                      (N14)? data_i[918] : 1'b0;
  assign data_o[21] = (N7)? data_i[21] : 
                      (N9)? data_i[149] : 
                      (N11)? data_i[277] : 
                      (N13)? data_i[405] : 
                      (N8)? data_i[533] : 
                      (N10)? data_i[661] : 
                      (N12)? data_i[789] : 
                      (N14)? data_i[917] : 1'b0;
  assign data_o[20] = (N7)? data_i[20] : 
                      (N9)? data_i[148] : 
                      (N11)? data_i[276] : 
                      (N13)? data_i[404] : 
                      (N8)? data_i[532] : 
                      (N10)? data_i[660] : 
                      (N12)? data_i[788] : 
                      (N14)? data_i[916] : 1'b0;
  assign data_o[19] = (N7)? data_i[19] : 
                      (N9)? data_i[147] : 
                      (N11)? data_i[275] : 
                      (N13)? data_i[403] : 
                      (N8)? data_i[531] : 
                      (N10)? data_i[659] : 
                      (N12)? data_i[787] : 
                      (N14)? data_i[915] : 1'b0;
  assign data_o[18] = (N7)? data_i[18] : 
                      (N9)? data_i[146] : 
                      (N11)? data_i[274] : 
                      (N13)? data_i[402] : 
                      (N8)? data_i[530] : 
                      (N10)? data_i[658] : 
                      (N12)? data_i[786] : 
                      (N14)? data_i[914] : 1'b0;
  assign data_o[17] = (N7)? data_i[17] : 
                      (N9)? data_i[145] : 
                      (N11)? data_i[273] : 
                      (N13)? data_i[401] : 
                      (N8)? data_i[529] : 
                      (N10)? data_i[657] : 
                      (N12)? data_i[785] : 
                      (N14)? data_i[913] : 1'b0;
  assign data_o[16] = (N7)? data_i[16] : 
                      (N9)? data_i[144] : 
                      (N11)? data_i[272] : 
                      (N13)? data_i[400] : 
                      (N8)? data_i[528] : 
                      (N10)? data_i[656] : 
                      (N12)? data_i[784] : 
                      (N14)? data_i[912] : 1'b0;
  assign data_o[15] = (N7)? data_i[15] : 
                      (N9)? data_i[143] : 
                      (N11)? data_i[271] : 
                      (N13)? data_i[399] : 
                      (N8)? data_i[527] : 
                      (N10)? data_i[655] : 
                      (N12)? data_i[783] : 
                      (N14)? data_i[911] : 1'b0;
  assign data_o[14] = (N7)? data_i[14] : 
                      (N9)? data_i[142] : 
                      (N11)? data_i[270] : 
                      (N13)? data_i[398] : 
                      (N8)? data_i[526] : 
                      (N10)? data_i[654] : 
                      (N12)? data_i[782] : 
                      (N14)? data_i[910] : 1'b0;
  assign data_o[13] = (N7)? data_i[13] : 
                      (N9)? data_i[141] : 
                      (N11)? data_i[269] : 
                      (N13)? data_i[397] : 
                      (N8)? data_i[525] : 
                      (N10)? data_i[653] : 
                      (N12)? data_i[781] : 
                      (N14)? data_i[909] : 1'b0;
  assign data_o[12] = (N7)? data_i[12] : 
                      (N9)? data_i[140] : 
                      (N11)? data_i[268] : 
                      (N13)? data_i[396] : 
                      (N8)? data_i[524] : 
                      (N10)? data_i[652] : 
                      (N12)? data_i[780] : 
                      (N14)? data_i[908] : 1'b0;
  assign data_o[11] = (N7)? data_i[11] : 
                      (N9)? data_i[139] : 
                      (N11)? data_i[267] : 
                      (N13)? data_i[395] : 
                      (N8)? data_i[523] : 
                      (N10)? data_i[651] : 
                      (N12)? data_i[779] : 
                      (N14)? data_i[907] : 1'b0;
  assign data_o[10] = (N7)? data_i[10] : 
                      (N9)? data_i[138] : 
                      (N11)? data_i[266] : 
                      (N13)? data_i[394] : 
                      (N8)? data_i[522] : 
                      (N10)? data_i[650] : 
                      (N12)? data_i[778] : 
                      (N14)? data_i[906] : 1'b0;
  assign data_o[9] = (N7)? data_i[9] : 
                     (N9)? data_i[137] : 
                     (N11)? data_i[265] : 
                     (N13)? data_i[393] : 
                     (N8)? data_i[521] : 
                     (N10)? data_i[649] : 
                     (N12)? data_i[777] : 
                     (N14)? data_i[905] : 1'b0;
  assign data_o[8] = (N7)? data_i[8] : 
                     (N9)? data_i[136] : 
                     (N11)? data_i[264] : 
                     (N13)? data_i[392] : 
                     (N8)? data_i[520] : 
                     (N10)? data_i[648] : 
                     (N12)? data_i[776] : 
                     (N14)? data_i[904] : 1'b0;
  assign data_o[7] = (N7)? data_i[7] : 
                     (N9)? data_i[135] : 
                     (N11)? data_i[263] : 
                     (N13)? data_i[391] : 
                     (N8)? data_i[519] : 
                     (N10)? data_i[647] : 
                     (N12)? data_i[775] : 
                     (N14)? data_i[903] : 1'b0;
  assign data_o[6] = (N7)? data_i[6] : 
                     (N9)? data_i[134] : 
                     (N11)? data_i[262] : 
                     (N13)? data_i[390] : 
                     (N8)? data_i[518] : 
                     (N10)? data_i[646] : 
                     (N12)? data_i[774] : 
                     (N14)? data_i[902] : 1'b0;
  assign data_o[5] = (N7)? data_i[5] : 
                     (N9)? data_i[133] : 
                     (N11)? data_i[261] : 
                     (N13)? data_i[389] : 
                     (N8)? data_i[517] : 
                     (N10)? data_i[645] : 
                     (N12)? data_i[773] : 
                     (N14)? data_i[901] : 1'b0;
  assign data_o[4] = (N7)? data_i[4] : 
                     (N9)? data_i[132] : 
                     (N11)? data_i[260] : 
                     (N13)? data_i[388] : 
                     (N8)? data_i[516] : 
                     (N10)? data_i[644] : 
                     (N12)? data_i[772] : 
                     (N14)? data_i[900] : 1'b0;
  assign data_o[3] = (N7)? data_i[3] : 
                     (N9)? data_i[131] : 
                     (N11)? data_i[259] : 
                     (N13)? data_i[387] : 
                     (N8)? data_i[515] : 
                     (N10)? data_i[643] : 
                     (N12)? data_i[771] : 
                     (N14)? data_i[899] : 1'b0;
  assign data_o[2] = (N7)? data_i[2] : 
                     (N9)? data_i[130] : 
                     (N11)? data_i[258] : 
                     (N13)? data_i[386] : 
                     (N8)? data_i[514] : 
                     (N10)? data_i[642] : 
                     (N12)? data_i[770] : 
                     (N14)? data_i[898] : 1'b0;
  assign data_o[1] = (N7)? data_i[1] : 
                     (N9)? data_i[129] : 
                     (N11)? data_i[257] : 
                     (N13)? data_i[385] : 
                     (N8)? data_i[513] : 
                     (N10)? data_i[641] : 
                     (N12)? data_i[769] : 
                     (N14)? data_i[897] : 1'b0;
  assign data_o[0] = (N7)? data_i[0] : 
                     (N9)? data_i[128] : 
                     (N11)? data_i[256] : 
                     (N13)? data_i[384] : 
                     (N8)? data_i[512] : 
                     (N10)? data_i[640] : 
                     (N12)? data_i[768] : 
                     (N14)? data_i[896] : 1'b0;
  assign data_o[255] = (N22)? data_i[127] : 
                       (N24)? data_i[255] : 
                       (N26)? data_i[383] : 
                       (N28)? data_i[511] : 
                       (N23)? data_i[639] : 
                       (N25)? data_i[767] : 
                       (N27)? data_i[895] : 
                       (N29)? data_i[1023] : 1'b0;
  assign data_o[254] = (N22)? data_i[126] : 
                       (N24)? data_i[254] : 
                       (N26)? data_i[382] : 
                       (N28)? data_i[510] : 
                       (N23)? data_i[638] : 
                       (N25)? data_i[766] : 
                       (N27)? data_i[894] : 
                       (N29)? data_i[1022] : 1'b0;
  assign data_o[253] = (N22)? data_i[125] : 
                       (N24)? data_i[253] : 
                       (N26)? data_i[381] : 
                       (N28)? data_i[509] : 
                       (N23)? data_i[637] : 
                       (N25)? data_i[765] : 
                       (N27)? data_i[893] : 
                       (N29)? data_i[1021] : 1'b0;
  assign data_o[252] = (N22)? data_i[124] : 
                       (N24)? data_i[252] : 
                       (N26)? data_i[380] : 
                       (N28)? data_i[508] : 
                       (N23)? data_i[636] : 
                       (N25)? data_i[764] : 
                       (N27)? data_i[892] : 
                       (N29)? data_i[1020] : 1'b0;
  assign data_o[251] = (N22)? data_i[123] : 
                       (N24)? data_i[251] : 
                       (N26)? data_i[379] : 
                       (N28)? data_i[507] : 
                       (N23)? data_i[635] : 
                       (N25)? data_i[763] : 
                       (N27)? data_i[891] : 
                       (N29)? data_i[1019] : 1'b0;
  assign data_o[250] = (N22)? data_i[122] : 
                       (N24)? data_i[250] : 
                       (N26)? data_i[378] : 
                       (N28)? data_i[506] : 
                       (N23)? data_i[634] : 
                       (N25)? data_i[762] : 
                       (N27)? data_i[890] : 
                       (N29)? data_i[1018] : 1'b0;
  assign data_o[249] = (N22)? data_i[121] : 
                       (N24)? data_i[249] : 
                       (N26)? data_i[377] : 
                       (N28)? data_i[505] : 
                       (N23)? data_i[633] : 
                       (N25)? data_i[761] : 
                       (N27)? data_i[889] : 
                       (N29)? data_i[1017] : 1'b0;
  assign data_o[248] = (N22)? data_i[120] : 
                       (N24)? data_i[248] : 
                       (N26)? data_i[376] : 
                       (N28)? data_i[504] : 
                       (N23)? data_i[632] : 
                       (N25)? data_i[760] : 
                       (N27)? data_i[888] : 
                       (N29)? data_i[1016] : 1'b0;
  assign data_o[247] = (N22)? data_i[119] : 
                       (N24)? data_i[247] : 
                       (N26)? data_i[375] : 
                       (N28)? data_i[503] : 
                       (N23)? data_i[631] : 
                       (N25)? data_i[759] : 
                       (N27)? data_i[887] : 
                       (N29)? data_i[1015] : 1'b0;
  assign data_o[246] = (N22)? data_i[118] : 
                       (N24)? data_i[246] : 
                       (N26)? data_i[374] : 
                       (N28)? data_i[502] : 
                       (N23)? data_i[630] : 
                       (N25)? data_i[758] : 
                       (N27)? data_i[886] : 
                       (N29)? data_i[1014] : 1'b0;
  assign data_o[245] = (N22)? data_i[117] : 
                       (N24)? data_i[245] : 
                       (N26)? data_i[373] : 
                       (N28)? data_i[501] : 
                       (N23)? data_i[629] : 
                       (N25)? data_i[757] : 
                       (N27)? data_i[885] : 
                       (N29)? data_i[1013] : 1'b0;
  assign data_o[244] = (N22)? data_i[116] : 
                       (N24)? data_i[244] : 
                       (N26)? data_i[372] : 
                       (N28)? data_i[500] : 
                       (N23)? data_i[628] : 
                       (N25)? data_i[756] : 
                       (N27)? data_i[884] : 
                       (N29)? data_i[1012] : 1'b0;
  assign data_o[243] = (N22)? data_i[115] : 
                       (N24)? data_i[243] : 
                       (N26)? data_i[371] : 
                       (N28)? data_i[499] : 
                       (N23)? data_i[627] : 
                       (N25)? data_i[755] : 
                       (N27)? data_i[883] : 
                       (N29)? data_i[1011] : 1'b0;
  assign data_o[242] = (N22)? data_i[114] : 
                       (N24)? data_i[242] : 
                       (N26)? data_i[370] : 
                       (N28)? data_i[498] : 
                       (N23)? data_i[626] : 
                       (N25)? data_i[754] : 
                       (N27)? data_i[882] : 
                       (N29)? data_i[1010] : 1'b0;
  assign data_o[241] = (N22)? data_i[113] : 
                       (N24)? data_i[241] : 
                       (N26)? data_i[369] : 
                       (N28)? data_i[497] : 
                       (N23)? data_i[625] : 
                       (N25)? data_i[753] : 
                       (N27)? data_i[881] : 
                       (N29)? data_i[1009] : 1'b0;
  assign data_o[240] = (N22)? data_i[112] : 
                       (N24)? data_i[240] : 
                       (N26)? data_i[368] : 
                       (N28)? data_i[496] : 
                       (N23)? data_i[624] : 
                       (N25)? data_i[752] : 
                       (N27)? data_i[880] : 
                       (N29)? data_i[1008] : 1'b0;
  assign data_o[239] = (N22)? data_i[111] : 
                       (N24)? data_i[239] : 
                       (N26)? data_i[367] : 
                       (N28)? data_i[495] : 
                       (N23)? data_i[623] : 
                       (N25)? data_i[751] : 
                       (N27)? data_i[879] : 
                       (N29)? data_i[1007] : 1'b0;
  assign data_o[238] = (N22)? data_i[110] : 
                       (N24)? data_i[238] : 
                       (N26)? data_i[366] : 
                       (N28)? data_i[494] : 
                       (N23)? data_i[622] : 
                       (N25)? data_i[750] : 
                       (N27)? data_i[878] : 
                       (N29)? data_i[1006] : 1'b0;
  assign data_o[237] = (N22)? data_i[109] : 
                       (N24)? data_i[237] : 
                       (N26)? data_i[365] : 
                       (N28)? data_i[493] : 
                       (N23)? data_i[621] : 
                       (N25)? data_i[749] : 
                       (N27)? data_i[877] : 
                       (N29)? data_i[1005] : 1'b0;
  assign data_o[236] = (N22)? data_i[108] : 
                       (N24)? data_i[236] : 
                       (N26)? data_i[364] : 
                       (N28)? data_i[492] : 
                       (N23)? data_i[620] : 
                       (N25)? data_i[748] : 
                       (N27)? data_i[876] : 
                       (N29)? data_i[1004] : 1'b0;
  assign data_o[235] = (N22)? data_i[107] : 
                       (N24)? data_i[235] : 
                       (N26)? data_i[363] : 
                       (N28)? data_i[491] : 
                       (N23)? data_i[619] : 
                       (N25)? data_i[747] : 
                       (N27)? data_i[875] : 
                       (N29)? data_i[1003] : 1'b0;
  assign data_o[234] = (N22)? data_i[106] : 
                       (N24)? data_i[234] : 
                       (N26)? data_i[362] : 
                       (N28)? data_i[490] : 
                       (N23)? data_i[618] : 
                       (N25)? data_i[746] : 
                       (N27)? data_i[874] : 
                       (N29)? data_i[1002] : 1'b0;
  assign data_o[233] = (N22)? data_i[105] : 
                       (N24)? data_i[233] : 
                       (N26)? data_i[361] : 
                       (N28)? data_i[489] : 
                       (N23)? data_i[617] : 
                       (N25)? data_i[745] : 
                       (N27)? data_i[873] : 
                       (N29)? data_i[1001] : 1'b0;
  assign data_o[232] = (N22)? data_i[104] : 
                       (N24)? data_i[232] : 
                       (N26)? data_i[360] : 
                       (N28)? data_i[488] : 
                       (N23)? data_i[616] : 
                       (N25)? data_i[744] : 
                       (N27)? data_i[872] : 
                       (N29)? data_i[1000] : 1'b0;
  assign data_o[231] = (N22)? data_i[103] : 
                       (N24)? data_i[231] : 
                       (N26)? data_i[359] : 
                       (N28)? data_i[487] : 
                       (N23)? data_i[615] : 
                       (N25)? data_i[743] : 
                       (N27)? data_i[871] : 
                       (N29)? data_i[999] : 1'b0;
  assign data_o[230] = (N22)? data_i[102] : 
                       (N24)? data_i[230] : 
                       (N26)? data_i[358] : 
                       (N28)? data_i[486] : 
                       (N23)? data_i[614] : 
                       (N25)? data_i[742] : 
                       (N27)? data_i[870] : 
                       (N29)? data_i[998] : 1'b0;
  assign data_o[229] = (N22)? data_i[101] : 
                       (N24)? data_i[229] : 
                       (N26)? data_i[357] : 
                       (N28)? data_i[485] : 
                       (N23)? data_i[613] : 
                       (N25)? data_i[741] : 
                       (N27)? data_i[869] : 
                       (N29)? data_i[997] : 1'b0;
  assign data_o[228] = (N22)? data_i[100] : 
                       (N24)? data_i[228] : 
                       (N26)? data_i[356] : 
                       (N28)? data_i[484] : 
                       (N23)? data_i[612] : 
                       (N25)? data_i[740] : 
                       (N27)? data_i[868] : 
                       (N29)? data_i[996] : 1'b0;
  assign data_o[227] = (N22)? data_i[99] : 
                       (N24)? data_i[227] : 
                       (N26)? data_i[355] : 
                       (N28)? data_i[483] : 
                       (N23)? data_i[611] : 
                       (N25)? data_i[739] : 
                       (N27)? data_i[867] : 
                       (N29)? data_i[995] : 1'b0;
  assign data_o[226] = (N22)? data_i[98] : 
                       (N24)? data_i[226] : 
                       (N26)? data_i[354] : 
                       (N28)? data_i[482] : 
                       (N23)? data_i[610] : 
                       (N25)? data_i[738] : 
                       (N27)? data_i[866] : 
                       (N29)? data_i[994] : 1'b0;
  assign data_o[225] = (N22)? data_i[97] : 
                       (N24)? data_i[225] : 
                       (N26)? data_i[353] : 
                       (N28)? data_i[481] : 
                       (N23)? data_i[609] : 
                       (N25)? data_i[737] : 
                       (N27)? data_i[865] : 
                       (N29)? data_i[993] : 1'b0;
  assign data_o[224] = (N22)? data_i[96] : 
                       (N24)? data_i[224] : 
                       (N26)? data_i[352] : 
                       (N28)? data_i[480] : 
                       (N23)? data_i[608] : 
                       (N25)? data_i[736] : 
                       (N27)? data_i[864] : 
                       (N29)? data_i[992] : 1'b0;
  assign data_o[223] = (N22)? data_i[95] : 
                       (N24)? data_i[223] : 
                       (N26)? data_i[351] : 
                       (N28)? data_i[479] : 
                       (N23)? data_i[607] : 
                       (N25)? data_i[735] : 
                       (N27)? data_i[863] : 
                       (N29)? data_i[991] : 1'b0;
  assign data_o[222] = (N22)? data_i[94] : 
                       (N24)? data_i[222] : 
                       (N26)? data_i[350] : 
                       (N28)? data_i[478] : 
                       (N23)? data_i[606] : 
                       (N25)? data_i[734] : 
                       (N27)? data_i[862] : 
                       (N29)? data_i[990] : 1'b0;
  assign data_o[221] = (N22)? data_i[93] : 
                       (N24)? data_i[221] : 
                       (N26)? data_i[349] : 
                       (N28)? data_i[477] : 
                       (N23)? data_i[605] : 
                       (N25)? data_i[733] : 
                       (N27)? data_i[861] : 
                       (N29)? data_i[989] : 1'b0;
  assign data_o[220] = (N22)? data_i[92] : 
                       (N24)? data_i[220] : 
                       (N26)? data_i[348] : 
                       (N28)? data_i[476] : 
                       (N23)? data_i[604] : 
                       (N25)? data_i[732] : 
                       (N27)? data_i[860] : 
                       (N29)? data_i[988] : 1'b0;
  assign data_o[219] = (N22)? data_i[91] : 
                       (N24)? data_i[219] : 
                       (N26)? data_i[347] : 
                       (N28)? data_i[475] : 
                       (N23)? data_i[603] : 
                       (N25)? data_i[731] : 
                       (N27)? data_i[859] : 
                       (N29)? data_i[987] : 1'b0;
  assign data_o[218] = (N22)? data_i[90] : 
                       (N24)? data_i[218] : 
                       (N26)? data_i[346] : 
                       (N28)? data_i[474] : 
                       (N23)? data_i[602] : 
                       (N25)? data_i[730] : 
                       (N27)? data_i[858] : 
                       (N29)? data_i[986] : 1'b0;
  assign data_o[217] = (N22)? data_i[89] : 
                       (N24)? data_i[217] : 
                       (N26)? data_i[345] : 
                       (N28)? data_i[473] : 
                       (N23)? data_i[601] : 
                       (N25)? data_i[729] : 
                       (N27)? data_i[857] : 
                       (N29)? data_i[985] : 1'b0;
  assign data_o[216] = (N22)? data_i[88] : 
                       (N24)? data_i[216] : 
                       (N26)? data_i[344] : 
                       (N28)? data_i[472] : 
                       (N23)? data_i[600] : 
                       (N25)? data_i[728] : 
                       (N27)? data_i[856] : 
                       (N29)? data_i[984] : 1'b0;
  assign data_o[215] = (N22)? data_i[87] : 
                       (N24)? data_i[215] : 
                       (N26)? data_i[343] : 
                       (N28)? data_i[471] : 
                       (N23)? data_i[599] : 
                       (N25)? data_i[727] : 
                       (N27)? data_i[855] : 
                       (N29)? data_i[983] : 1'b0;
  assign data_o[214] = (N22)? data_i[86] : 
                       (N24)? data_i[214] : 
                       (N26)? data_i[342] : 
                       (N28)? data_i[470] : 
                       (N23)? data_i[598] : 
                       (N25)? data_i[726] : 
                       (N27)? data_i[854] : 
                       (N29)? data_i[982] : 1'b0;
  assign data_o[213] = (N22)? data_i[85] : 
                       (N24)? data_i[213] : 
                       (N26)? data_i[341] : 
                       (N28)? data_i[469] : 
                       (N23)? data_i[597] : 
                       (N25)? data_i[725] : 
                       (N27)? data_i[853] : 
                       (N29)? data_i[981] : 1'b0;
  assign data_o[212] = (N22)? data_i[84] : 
                       (N24)? data_i[212] : 
                       (N26)? data_i[340] : 
                       (N28)? data_i[468] : 
                       (N23)? data_i[596] : 
                       (N25)? data_i[724] : 
                       (N27)? data_i[852] : 
                       (N29)? data_i[980] : 1'b0;
  assign data_o[211] = (N22)? data_i[83] : 
                       (N24)? data_i[211] : 
                       (N26)? data_i[339] : 
                       (N28)? data_i[467] : 
                       (N23)? data_i[595] : 
                       (N25)? data_i[723] : 
                       (N27)? data_i[851] : 
                       (N29)? data_i[979] : 1'b0;
  assign data_o[210] = (N22)? data_i[82] : 
                       (N24)? data_i[210] : 
                       (N26)? data_i[338] : 
                       (N28)? data_i[466] : 
                       (N23)? data_i[594] : 
                       (N25)? data_i[722] : 
                       (N27)? data_i[850] : 
                       (N29)? data_i[978] : 1'b0;
  assign data_o[209] = (N22)? data_i[81] : 
                       (N24)? data_i[209] : 
                       (N26)? data_i[337] : 
                       (N28)? data_i[465] : 
                       (N23)? data_i[593] : 
                       (N25)? data_i[721] : 
                       (N27)? data_i[849] : 
                       (N29)? data_i[977] : 1'b0;
  assign data_o[208] = (N22)? data_i[80] : 
                       (N24)? data_i[208] : 
                       (N26)? data_i[336] : 
                       (N28)? data_i[464] : 
                       (N23)? data_i[592] : 
                       (N25)? data_i[720] : 
                       (N27)? data_i[848] : 
                       (N29)? data_i[976] : 1'b0;
  assign data_o[207] = (N22)? data_i[79] : 
                       (N24)? data_i[207] : 
                       (N26)? data_i[335] : 
                       (N28)? data_i[463] : 
                       (N23)? data_i[591] : 
                       (N25)? data_i[719] : 
                       (N27)? data_i[847] : 
                       (N29)? data_i[975] : 1'b0;
  assign data_o[206] = (N22)? data_i[78] : 
                       (N24)? data_i[206] : 
                       (N26)? data_i[334] : 
                       (N28)? data_i[462] : 
                       (N23)? data_i[590] : 
                       (N25)? data_i[718] : 
                       (N27)? data_i[846] : 
                       (N29)? data_i[974] : 1'b0;
  assign data_o[205] = (N22)? data_i[77] : 
                       (N24)? data_i[205] : 
                       (N26)? data_i[333] : 
                       (N28)? data_i[461] : 
                       (N23)? data_i[589] : 
                       (N25)? data_i[717] : 
                       (N27)? data_i[845] : 
                       (N29)? data_i[973] : 1'b0;
  assign data_o[204] = (N22)? data_i[76] : 
                       (N24)? data_i[204] : 
                       (N26)? data_i[332] : 
                       (N28)? data_i[460] : 
                       (N23)? data_i[588] : 
                       (N25)? data_i[716] : 
                       (N27)? data_i[844] : 
                       (N29)? data_i[972] : 1'b0;
  assign data_o[203] = (N22)? data_i[75] : 
                       (N24)? data_i[203] : 
                       (N26)? data_i[331] : 
                       (N28)? data_i[459] : 
                       (N23)? data_i[587] : 
                       (N25)? data_i[715] : 
                       (N27)? data_i[843] : 
                       (N29)? data_i[971] : 1'b0;
  assign data_o[202] = (N22)? data_i[74] : 
                       (N24)? data_i[202] : 
                       (N26)? data_i[330] : 
                       (N28)? data_i[458] : 
                       (N23)? data_i[586] : 
                       (N25)? data_i[714] : 
                       (N27)? data_i[842] : 
                       (N29)? data_i[970] : 1'b0;
  assign data_o[201] = (N22)? data_i[73] : 
                       (N24)? data_i[201] : 
                       (N26)? data_i[329] : 
                       (N28)? data_i[457] : 
                       (N23)? data_i[585] : 
                       (N25)? data_i[713] : 
                       (N27)? data_i[841] : 
                       (N29)? data_i[969] : 1'b0;
  assign data_o[200] = (N22)? data_i[72] : 
                       (N24)? data_i[200] : 
                       (N26)? data_i[328] : 
                       (N28)? data_i[456] : 
                       (N23)? data_i[584] : 
                       (N25)? data_i[712] : 
                       (N27)? data_i[840] : 
                       (N29)? data_i[968] : 1'b0;
  assign data_o[199] = (N22)? data_i[71] : 
                       (N24)? data_i[199] : 
                       (N26)? data_i[327] : 
                       (N28)? data_i[455] : 
                       (N23)? data_i[583] : 
                       (N25)? data_i[711] : 
                       (N27)? data_i[839] : 
                       (N29)? data_i[967] : 1'b0;
  assign data_o[198] = (N22)? data_i[70] : 
                       (N24)? data_i[198] : 
                       (N26)? data_i[326] : 
                       (N28)? data_i[454] : 
                       (N23)? data_i[582] : 
                       (N25)? data_i[710] : 
                       (N27)? data_i[838] : 
                       (N29)? data_i[966] : 1'b0;
  assign data_o[197] = (N22)? data_i[69] : 
                       (N24)? data_i[197] : 
                       (N26)? data_i[325] : 
                       (N28)? data_i[453] : 
                       (N23)? data_i[581] : 
                       (N25)? data_i[709] : 
                       (N27)? data_i[837] : 
                       (N29)? data_i[965] : 1'b0;
  assign data_o[196] = (N22)? data_i[68] : 
                       (N24)? data_i[196] : 
                       (N26)? data_i[324] : 
                       (N28)? data_i[452] : 
                       (N23)? data_i[580] : 
                       (N25)? data_i[708] : 
                       (N27)? data_i[836] : 
                       (N29)? data_i[964] : 1'b0;
  assign data_o[195] = (N22)? data_i[67] : 
                       (N24)? data_i[195] : 
                       (N26)? data_i[323] : 
                       (N28)? data_i[451] : 
                       (N23)? data_i[579] : 
                       (N25)? data_i[707] : 
                       (N27)? data_i[835] : 
                       (N29)? data_i[963] : 1'b0;
  assign data_o[194] = (N22)? data_i[66] : 
                       (N24)? data_i[194] : 
                       (N26)? data_i[322] : 
                       (N28)? data_i[450] : 
                       (N23)? data_i[578] : 
                       (N25)? data_i[706] : 
                       (N27)? data_i[834] : 
                       (N29)? data_i[962] : 1'b0;
  assign data_o[193] = (N22)? data_i[65] : 
                       (N24)? data_i[193] : 
                       (N26)? data_i[321] : 
                       (N28)? data_i[449] : 
                       (N23)? data_i[577] : 
                       (N25)? data_i[705] : 
                       (N27)? data_i[833] : 
                       (N29)? data_i[961] : 1'b0;
  assign data_o[192] = (N22)? data_i[64] : 
                       (N24)? data_i[192] : 
                       (N26)? data_i[320] : 
                       (N28)? data_i[448] : 
                       (N23)? data_i[576] : 
                       (N25)? data_i[704] : 
                       (N27)? data_i[832] : 
                       (N29)? data_i[960] : 1'b0;
  assign data_o[191] = (N22)? data_i[63] : 
                       (N24)? data_i[191] : 
                       (N26)? data_i[319] : 
                       (N28)? data_i[447] : 
                       (N23)? data_i[575] : 
                       (N25)? data_i[703] : 
                       (N27)? data_i[831] : 
                       (N29)? data_i[959] : 1'b0;
  assign data_o[190] = (N22)? data_i[62] : 
                       (N24)? data_i[190] : 
                       (N26)? data_i[318] : 
                       (N28)? data_i[446] : 
                       (N23)? data_i[574] : 
                       (N25)? data_i[702] : 
                       (N27)? data_i[830] : 
                       (N29)? data_i[958] : 1'b0;
  assign data_o[189] = (N22)? data_i[61] : 
                       (N24)? data_i[189] : 
                       (N26)? data_i[317] : 
                       (N28)? data_i[445] : 
                       (N23)? data_i[573] : 
                       (N25)? data_i[701] : 
                       (N27)? data_i[829] : 
                       (N29)? data_i[957] : 1'b0;
  assign data_o[188] = (N22)? data_i[60] : 
                       (N24)? data_i[188] : 
                       (N26)? data_i[316] : 
                       (N28)? data_i[444] : 
                       (N23)? data_i[572] : 
                       (N25)? data_i[700] : 
                       (N27)? data_i[828] : 
                       (N29)? data_i[956] : 1'b0;
  assign data_o[187] = (N22)? data_i[59] : 
                       (N24)? data_i[187] : 
                       (N26)? data_i[315] : 
                       (N28)? data_i[443] : 
                       (N23)? data_i[571] : 
                       (N25)? data_i[699] : 
                       (N27)? data_i[827] : 
                       (N29)? data_i[955] : 1'b0;
  assign data_o[186] = (N22)? data_i[58] : 
                       (N24)? data_i[186] : 
                       (N26)? data_i[314] : 
                       (N28)? data_i[442] : 
                       (N23)? data_i[570] : 
                       (N25)? data_i[698] : 
                       (N27)? data_i[826] : 
                       (N29)? data_i[954] : 1'b0;
  assign data_o[185] = (N22)? data_i[57] : 
                       (N24)? data_i[185] : 
                       (N26)? data_i[313] : 
                       (N28)? data_i[441] : 
                       (N23)? data_i[569] : 
                       (N25)? data_i[697] : 
                       (N27)? data_i[825] : 
                       (N29)? data_i[953] : 1'b0;
  assign data_o[184] = (N22)? data_i[56] : 
                       (N24)? data_i[184] : 
                       (N26)? data_i[312] : 
                       (N28)? data_i[440] : 
                       (N23)? data_i[568] : 
                       (N25)? data_i[696] : 
                       (N27)? data_i[824] : 
                       (N29)? data_i[952] : 1'b0;
  assign data_o[183] = (N22)? data_i[55] : 
                       (N24)? data_i[183] : 
                       (N26)? data_i[311] : 
                       (N28)? data_i[439] : 
                       (N23)? data_i[567] : 
                       (N25)? data_i[695] : 
                       (N27)? data_i[823] : 
                       (N29)? data_i[951] : 1'b0;
  assign data_o[182] = (N22)? data_i[54] : 
                       (N24)? data_i[182] : 
                       (N26)? data_i[310] : 
                       (N28)? data_i[438] : 
                       (N23)? data_i[566] : 
                       (N25)? data_i[694] : 
                       (N27)? data_i[822] : 
                       (N29)? data_i[950] : 1'b0;
  assign data_o[181] = (N22)? data_i[53] : 
                       (N24)? data_i[181] : 
                       (N26)? data_i[309] : 
                       (N28)? data_i[437] : 
                       (N23)? data_i[565] : 
                       (N25)? data_i[693] : 
                       (N27)? data_i[821] : 
                       (N29)? data_i[949] : 1'b0;
  assign data_o[180] = (N22)? data_i[52] : 
                       (N24)? data_i[180] : 
                       (N26)? data_i[308] : 
                       (N28)? data_i[436] : 
                       (N23)? data_i[564] : 
                       (N25)? data_i[692] : 
                       (N27)? data_i[820] : 
                       (N29)? data_i[948] : 1'b0;
  assign data_o[179] = (N22)? data_i[51] : 
                       (N24)? data_i[179] : 
                       (N26)? data_i[307] : 
                       (N28)? data_i[435] : 
                       (N23)? data_i[563] : 
                       (N25)? data_i[691] : 
                       (N27)? data_i[819] : 
                       (N29)? data_i[947] : 1'b0;
  assign data_o[178] = (N22)? data_i[50] : 
                       (N24)? data_i[178] : 
                       (N26)? data_i[306] : 
                       (N28)? data_i[434] : 
                       (N23)? data_i[562] : 
                       (N25)? data_i[690] : 
                       (N27)? data_i[818] : 
                       (N29)? data_i[946] : 1'b0;
  assign data_o[177] = (N22)? data_i[49] : 
                       (N24)? data_i[177] : 
                       (N26)? data_i[305] : 
                       (N28)? data_i[433] : 
                       (N23)? data_i[561] : 
                       (N25)? data_i[689] : 
                       (N27)? data_i[817] : 
                       (N29)? data_i[945] : 1'b0;
  assign data_o[176] = (N22)? data_i[48] : 
                       (N24)? data_i[176] : 
                       (N26)? data_i[304] : 
                       (N28)? data_i[432] : 
                       (N23)? data_i[560] : 
                       (N25)? data_i[688] : 
                       (N27)? data_i[816] : 
                       (N29)? data_i[944] : 1'b0;
  assign data_o[175] = (N22)? data_i[47] : 
                       (N24)? data_i[175] : 
                       (N26)? data_i[303] : 
                       (N28)? data_i[431] : 
                       (N23)? data_i[559] : 
                       (N25)? data_i[687] : 
                       (N27)? data_i[815] : 
                       (N29)? data_i[943] : 1'b0;
  assign data_o[174] = (N22)? data_i[46] : 
                       (N24)? data_i[174] : 
                       (N26)? data_i[302] : 
                       (N28)? data_i[430] : 
                       (N23)? data_i[558] : 
                       (N25)? data_i[686] : 
                       (N27)? data_i[814] : 
                       (N29)? data_i[942] : 1'b0;
  assign data_o[173] = (N22)? data_i[45] : 
                       (N24)? data_i[173] : 
                       (N26)? data_i[301] : 
                       (N28)? data_i[429] : 
                       (N23)? data_i[557] : 
                       (N25)? data_i[685] : 
                       (N27)? data_i[813] : 
                       (N29)? data_i[941] : 1'b0;
  assign data_o[172] = (N22)? data_i[44] : 
                       (N24)? data_i[172] : 
                       (N26)? data_i[300] : 
                       (N28)? data_i[428] : 
                       (N23)? data_i[556] : 
                       (N25)? data_i[684] : 
                       (N27)? data_i[812] : 
                       (N29)? data_i[940] : 1'b0;
  assign data_o[171] = (N22)? data_i[43] : 
                       (N24)? data_i[171] : 
                       (N26)? data_i[299] : 
                       (N28)? data_i[427] : 
                       (N23)? data_i[555] : 
                       (N25)? data_i[683] : 
                       (N27)? data_i[811] : 
                       (N29)? data_i[939] : 1'b0;
  assign data_o[170] = (N22)? data_i[42] : 
                       (N24)? data_i[170] : 
                       (N26)? data_i[298] : 
                       (N28)? data_i[426] : 
                       (N23)? data_i[554] : 
                       (N25)? data_i[682] : 
                       (N27)? data_i[810] : 
                       (N29)? data_i[938] : 1'b0;
  assign data_o[169] = (N22)? data_i[41] : 
                       (N24)? data_i[169] : 
                       (N26)? data_i[297] : 
                       (N28)? data_i[425] : 
                       (N23)? data_i[553] : 
                       (N25)? data_i[681] : 
                       (N27)? data_i[809] : 
                       (N29)? data_i[937] : 1'b0;
  assign data_o[168] = (N22)? data_i[40] : 
                       (N24)? data_i[168] : 
                       (N26)? data_i[296] : 
                       (N28)? data_i[424] : 
                       (N23)? data_i[552] : 
                       (N25)? data_i[680] : 
                       (N27)? data_i[808] : 
                       (N29)? data_i[936] : 1'b0;
  assign data_o[167] = (N22)? data_i[39] : 
                       (N24)? data_i[167] : 
                       (N26)? data_i[295] : 
                       (N28)? data_i[423] : 
                       (N23)? data_i[551] : 
                       (N25)? data_i[679] : 
                       (N27)? data_i[807] : 
                       (N29)? data_i[935] : 1'b0;
  assign data_o[166] = (N22)? data_i[38] : 
                       (N24)? data_i[166] : 
                       (N26)? data_i[294] : 
                       (N28)? data_i[422] : 
                       (N23)? data_i[550] : 
                       (N25)? data_i[678] : 
                       (N27)? data_i[806] : 
                       (N29)? data_i[934] : 1'b0;
  assign data_o[165] = (N22)? data_i[37] : 
                       (N24)? data_i[165] : 
                       (N26)? data_i[293] : 
                       (N28)? data_i[421] : 
                       (N23)? data_i[549] : 
                       (N25)? data_i[677] : 
                       (N27)? data_i[805] : 
                       (N29)? data_i[933] : 1'b0;
  assign data_o[164] = (N22)? data_i[36] : 
                       (N24)? data_i[164] : 
                       (N26)? data_i[292] : 
                       (N28)? data_i[420] : 
                       (N23)? data_i[548] : 
                       (N25)? data_i[676] : 
                       (N27)? data_i[804] : 
                       (N29)? data_i[932] : 1'b0;
  assign data_o[163] = (N22)? data_i[35] : 
                       (N24)? data_i[163] : 
                       (N26)? data_i[291] : 
                       (N28)? data_i[419] : 
                       (N23)? data_i[547] : 
                       (N25)? data_i[675] : 
                       (N27)? data_i[803] : 
                       (N29)? data_i[931] : 1'b0;
  assign data_o[162] = (N22)? data_i[34] : 
                       (N24)? data_i[162] : 
                       (N26)? data_i[290] : 
                       (N28)? data_i[418] : 
                       (N23)? data_i[546] : 
                       (N25)? data_i[674] : 
                       (N27)? data_i[802] : 
                       (N29)? data_i[930] : 1'b0;
  assign data_o[161] = (N22)? data_i[33] : 
                       (N24)? data_i[161] : 
                       (N26)? data_i[289] : 
                       (N28)? data_i[417] : 
                       (N23)? data_i[545] : 
                       (N25)? data_i[673] : 
                       (N27)? data_i[801] : 
                       (N29)? data_i[929] : 1'b0;
  assign data_o[160] = (N22)? data_i[32] : 
                       (N24)? data_i[160] : 
                       (N26)? data_i[288] : 
                       (N28)? data_i[416] : 
                       (N23)? data_i[544] : 
                       (N25)? data_i[672] : 
                       (N27)? data_i[800] : 
                       (N29)? data_i[928] : 1'b0;
  assign data_o[159] = (N22)? data_i[31] : 
                       (N24)? data_i[159] : 
                       (N26)? data_i[287] : 
                       (N28)? data_i[415] : 
                       (N23)? data_i[543] : 
                       (N25)? data_i[671] : 
                       (N27)? data_i[799] : 
                       (N29)? data_i[927] : 1'b0;
  assign data_o[158] = (N22)? data_i[30] : 
                       (N24)? data_i[158] : 
                       (N26)? data_i[286] : 
                       (N28)? data_i[414] : 
                       (N23)? data_i[542] : 
                       (N25)? data_i[670] : 
                       (N27)? data_i[798] : 
                       (N29)? data_i[926] : 1'b0;
  assign data_o[157] = (N22)? data_i[29] : 
                       (N24)? data_i[157] : 
                       (N26)? data_i[285] : 
                       (N28)? data_i[413] : 
                       (N23)? data_i[541] : 
                       (N25)? data_i[669] : 
                       (N27)? data_i[797] : 
                       (N29)? data_i[925] : 1'b0;
  assign data_o[156] = (N22)? data_i[28] : 
                       (N24)? data_i[156] : 
                       (N26)? data_i[284] : 
                       (N28)? data_i[412] : 
                       (N23)? data_i[540] : 
                       (N25)? data_i[668] : 
                       (N27)? data_i[796] : 
                       (N29)? data_i[924] : 1'b0;
  assign data_o[155] = (N22)? data_i[27] : 
                       (N24)? data_i[155] : 
                       (N26)? data_i[283] : 
                       (N28)? data_i[411] : 
                       (N23)? data_i[539] : 
                       (N25)? data_i[667] : 
                       (N27)? data_i[795] : 
                       (N29)? data_i[923] : 1'b0;
  assign data_o[154] = (N22)? data_i[26] : 
                       (N24)? data_i[154] : 
                       (N26)? data_i[282] : 
                       (N28)? data_i[410] : 
                       (N23)? data_i[538] : 
                       (N25)? data_i[666] : 
                       (N27)? data_i[794] : 
                       (N29)? data_i[922] : 1'b0;
  assign data_o[153] = (N22)? data_i[25] : 
                       (N24)? data_i[153] : 
                       (N26)? data_i[281] : 
                       (N28)? data_i[409] : 
                       (N23)? data_i[537] : 
                       (N25)? data_i[665] : 
                       (N27)? data_i[793] : 
                       (N29)? data_i[921] : 1'b0;
  assign data_o[152] = (N22)? data_i[24] : 
                       (N24)? data_i[152] : 
                       (N26)? data_i[280] : 
                       (N28)? data_i[408] : 
                       (N23)? data_i[536] : 
                       (N25)? data_i[664] : 
                       (N27)? data_i[792] : 
                       (N29)? data_i[920] : 1'b0;
  assign data_o[151] = (N22)? data_i[23] : 
                       (N24)? data_i[151] : 
                       (N26)? data_i[279] : 
                       (N28)? data_i[407] : 
                       (N23)? data_i[535] : 
                       (N25)? data_i[663] : 
                       (N27)? data_i[791] : 
                       (N29)? data_i[919] : 1'b0;
  assign data_o[150] = (N22)? data_i[22] : 
                       (N24)? data_i[150] : 
                       (N26)? data_i[278] : 
                       (N28)? data_i[406] : 
                       (N23)? data_i[534] : 
                       (N25)? data_i[662] : 
                       (N27)? data_i[790] : 
                       (N29)? data_i[918] : 1'b0;
  assign data_o[149] = (N22)? data_i[21] : 
                       (N24)? data_i[149] : 
                       (N26)? data_i[277] : 
                       (N28)? data_i[405] : 
                       (N23)? data_i[533] : 
                       (N25)? data_i[661] : 
                       (N27)? data_i[789] : 
                       (N29)? data_i[917] : 1'b0;
  assign data_o[148] = (N22)? data_i[20] : 
                       (N24)? data_i[148] : 
                       (N26)? data_i[276] : 
                       (N28)? data_i[404] : 
                       (N23)? data_i[532] : 
                       (N25)? data_i[660] : 
                       (N27)? data_i[788] : 
                       (N29)? data_i[916] : 1'b0;
  assign data_o[147] = (N22)? data_i[19] : 
                       (N24)? data_i[147] : 
                       (N26)? data_i[275] : 
                       (N28)? data_i[403] : 
                       (N23)? data_i[531] : 
                       (N25)? data_i[659] : 
                       (N27)? data_i[787] : 
                       (N29)? data_i[915] : 1'b0;
  assign data_o[146] = (N22)? data_i[18] : 
                       (N24)? data_i[146] : 
                       (N26)? data_i[274] : 
                       (N28)? data_i[402] : 
                       (N23)? data_i[530] : 
                       (N25)? data_i[658] : 
                       (N27)? data_i[786] : 
                       (N29)? data_i[914] : 1'b0;
  assign data_o[145] = (N22)? data_i[17] : 
                       (N24)? data_i[145] : 
                       (N26)? data_i[273] : 
                       (N28)? data_i[401] : 
                       (N23)? data_i[529] : 
                       (N25)? data_i[657] : 
                       (N27)? data_i[785] : 
                       (N29)? data_i[913] : 1'b0;
  assign data_o[144] = (N22)? data_i[16] : 
                       (N24)? data_i[144] : 
                       (N26)? data_i[272] : 
                       (N28)? data_i[400] : 
                       (N23)? data_i[528] : 
                       (N25)? data_i[656] : 
                       (N27)? data_i[784] : 
                       (N29)? data_i[912] : 1'b0;
  assign data_o[143] = (N22)? data_i[15] : 
                       (N24)? data_i[143] : 
                       (N26)? data_i[271] : 
                       (N28)? data_i[399] : 
                       (N23)? data_i[527] : 
                       (N25)? data_i[655] : 
                       (N27)? data_i[783] : 
                       (N29)? data_i[911] : 1'b0;
  assign data_o[142] = (N22)? data_i[14] : 
                       (N24)? data_i[142] : 
                       (N26)? data_i[270] : 
                       (N28)? data_i[398] : 
                       (N23)? data_i[526] : 
                       (N25)? data_i[654] : 
                       (N27)? data_i[782] : 
                       (N29)? data_i[910] : 1'b0;
  assign data_o[141] = (N22)? data_i[13] : 
                       (N24)? data_i[141] : 
                       (N26)? data_i[269] : 
                       (N28)? data_i[397] : 
                       (N23)? data_i[525] : 
                       (N25)? data_i[653] : 
                       (N27)? data_i[781] : 
                       (N29)? data_i[909] : 1'b0;
  assign data_o[140] = (N22)? data_i[12] : 
                       (N24)? data_i[140] : 
                       (N26)? data_i[268] : 
                       (N28)? data_i[396] : 
                       (N23)? data_i[524] : 
                       (N25)? data_i[652] : 
                       (N27)? data_i[780] : 
                       (N29)? data_i[908] : 1'b0;
  assign data_o[139] = (N22)? data_i[11] : 
                       (N24)? data_i[139] : 
                       (N26)? data_i[267] : 
                       (N28)? data_i[395] : 
                       (N23)? data_i[523] : 
                       (N25)? data_i[651] : 
                       (N27)? data_i[779] : 
                       (N29)? data_i[907] : 1'b0;
  assign data_o[138] = (N22)? data_i[10] : 
                       (N24)? data_i[138] : 
                       (N26)? data_i[266] : 
                       (N28)? data_i[394] : 
                       (N23)? data_i[522] : 
                       (N25)? data_i[650] : 
                       (N27)? data_i[778] : 
                       (N29)? data_i[906] : 1'b0;
  assign data_o[137] = (N22)? data_i[9] : 
                       (N24)? data_i[137] : 
                       (N26)? data_i[265] : 
                       (N28)? data_i[393] : 
                       (N23)? data_i[521] : 
                       (N25)? data_i[649] : 
                       (N27)? data_i[777] : 
                       (N29)? data_i[905] : 1'b0;
  assign data_o[136] = (N22)? data_i[8] : 
                       (N24)? data_i[136] : 
                       (N26)? data_i[264] : 
                       (N28)? data_i[392] : 
                       (N23)? data_i[520] : 
                       (N25)? data_i[648] : 
                       (N27)? data_i[776] : 
                       (N29)? data_i[904] : 1'b0;
  assign data_o[135] = (N22)? data_i[7] : 
                       (N24)? data_i[135] : 
                       (N26)? data_i[263] : 
                       (N28)? data_i[391] : 
                       (N23)? data_i[519] : 
                       (N25)? data_i[647] : 
                       (N27)? data_i[775] : 
                       (N29)? data_i[903] : 1'b0;
  assign data_o[134] = (N22)? data_i[6] : 
                       (N24)? data_i[134] : 
                       (N26)? data_i[262] : 
                       (N28)? data_i[390] : 
                       (N23)? data_i[518] : 
                       (N25)? data_i[646] : 
                       (N27)? data_i[774] : 
                       (N29)? data_i[902] : 1'b0;
  assign data_o[133] = (N22)? data_i[5] : 
                       (N24)? data_i[133] : 
                       (N26)? data_i[261] : 
                       (N28)? data_i[389] : 
                       (N23)? data_i[517] : 
                       (N25)? data_i[645] : 
                       (N27)? data_i[773] : 
                       (N29)? data_i[901] : 1'b0;
  assign data_o[132] = (N22)? data_i[4] : 
                       (N24)? data_i[132] : 
                       (N26)? data_i[260] : 
                       (N28)? data_i[388] : 
                       (N23)? data_i[516] : 
                       (N25)? data_i[644] : 
                       (N27)? data_i[772] : 
                       (N29)? data_i[900] : 1'b0;
  assign data_o[131] = (N22)? data_i[3] : 
                       (N24)? data_i[131] : 
                       (N26)? data_i[259] : 
                       (N28)? data_i[387] : 
                       (N23)? data_i[515] : 
                       (N25)? data_i[643] : 
                       (N27)? data_i[771] : 
                       (N29)? data_i[899] : 1'b0;
  assign data_o[130] = (N22)? data_i[2] : 
                       (N24)? data_i[130] : 
                       (N26)? data_i[258] : 
                       (N28)? data_i[386] : 
                       (N23)? data_i[514] : 
                       (N25)? data_i[642] : 
                       (N27)? data_i[770] : 
                       (N29)? data_i[898] : 1'b0;
  assign data_o[129] = (N22)? data_i[1] : 
                       (N24)? data_i[129] : 
                       (N26)? data_i[257] : 
                       (N28)? data_i[385] : 
                       (N23)? data_i[513] : 
                       (N25)? data_i[641] : 
                       (N27)? data_i[769] : 
                       (N29)? data_i[897] : 1'b0;
  assign data_o[128] = (N22)? data_i[0] : 
                       (N24)? data_i[128] : 
                       (N26)? data_i[256] : 
                       (N28)? data_i[384] : 
                       (N23)? data_i[512] : 
                       (N25)? data_i[640] : 
                       (N27)? data_i[768] : 
                       (N29)? data_i[896] : 1'b0;
  assign data_o[383] = (N37)? data_i[127] : 
                       (N39)? data_i[255] : 
                       (N41)? data_i[383] : 
                       (N43)? data_i[511] : 
                       (N38)? data_i[639] : 
                       (N40)? data_i[767] : 
                       (N42)? data_i[895] : 
                       (N44)? data_i[1023] : 1'b0;
  assign data_o[382] = (N37)? data_i[126] : 
                       (N39)? data_i[254] : 
                       (N41)? data_i[382] : 
                       (N43)? data_i[510] : 
                       (N38)? data_i[638] : 
                       (N40)? data_i[766] : 
                       (N42)? data_i[894] : 
                       (N44)? data_i[1022] : 1'b0;
  assign data_o[381] = (N37)? data_i[125] : 
                       (N39)? data_i[253] : 
                       (N41)? data_i[381] : 
                       (N43)? data_i[509] : 
                       (N38)? data_i[637] : 
                       (N40)? data_i[765] : 
                       (N42)? data_i[893] : 
                       (N44)? data_i[1021] : 1'b0;
  assign data_o[380] = (N37)? data_i[124] : 
                       (N39)? data_i[252] : 
                       (N41)? data_i[380] : 
                       (N43)? data_i[508] : 
                       (N38)? data_i[636] : 
                       (N40)? data_i[764] : 
                       (N42)? data_i[892] : 
                       (N44)? data_i[1020] : 1'b0;
  assign data_o[379] = (N37)? data_i[123] : 
                       (N39)? data_i[251] : 
                       (N41)? data_i[379] : 
                       (N43)? data_i[507] : 
                       (N38)? data_i[635] : 
                       (N40)? data_i[763] : 
                       (N42)? data_i[891] : 
                       (N44)? data_i[1019] : 1'b0;
  assign data_o[378] = (N37)? data_i[122] : 
                       (N39)? data_i[250] : 
                       (N41)? data_i[378] : 
                       (N43)? data_i[506] : 
                       (N38)? data_i[634] : 
                       (N40)? data_i[762] : 
                       (N42)? data_i[890] : 
                       (N44)? data_i[1018] : 1'b0;
  assign data_o[377] = (N37)? data_i[121] : 
                       (N39)? data_i[249] : 
                       (N41)? data_i[377] : 
                       (N43)? data_i[505] : 
                       (N38)? data_i[633] : 
                       (N40)? data_i[761] : 
                       (N42)? data_i[889] : 
                       (N44)? data_i[1017] : 1'b0;
  assign data_o[376] = (N37)? data_i[120] : 
                       (N39)? data_i[248] : 
                       (N41)? data_i[376] : 
                       (N43)? data_i[504] : 
                       (N38)? data_i[632] : 
                       (N40)? data_i[760] : 
                       (N42)? data_i[888] : 
                       (N44)? data_i[1016] : 1'b0;
  assign data_o[375] = (N37)? data_i[119] : 
                       (N39)? data_i[247] : 
                       (N41)? data_i[375] : 
                       (N43)? data_i[503] : 
                       (N38)? data_i[631] : 
                       (N40)? data_i[759] : 
                       (N42)? data_i[887] : 
                       (N44)? data_i[1015] : 1'b0;
  assign data_o[374] = (N37)? data_i[118] : 
                       (N39)? data_i[246] : 
                       (N41)? data_i[374] : 
                       (N43)? data_i[502] : 
                       (N38)? data_i[630] : 
                       (N40)? data_i[758] : 
                       (N42)? data_i[886] : 
                       (N44)? data_i[1014] : 1'b0;
  assign data_o[373] = (N37)? data_i[117] : 
                       (N39)? data_i[245] : 
                       (N41)? data_i[373] : 
                       (N43)? data_i[501] : 
                       (N38)? data_i[629] : 
                       (N40)? data_i[757] : 
                       (N42)? data_i[885] : 
                       (N44)? data_i[1013] : 1'b0;
  assign data_o[372] = (N37)? data_i[116] : 
                       (N39)? data_i[244] : 
                       (N41)? data_i[372] : 
                       (N43)? data_i[500] : 
                       (N38)? data_i[628] : 
                       (N40)? data_i[756] : 
                       (N42)? data_i[884] : 
                       (N44)? data_i[1012] : 1'b0;
  assign data_o[371] = (N37)? data_i[115] : 
                       (N39)? data_i[243] : 
                       (N41)? data_i[371] : 
                       (N43)? data_i[499] : 
                       (N38)? data_i[627] : 
                       (N40)? data_i[755] : 
                       (N42)? data_i[883] : 
                       (N44)? data_i[1011] : 1'b0;
  assign data_o[370] = (N37)? data_i[114] : 
                       (N39)? data_i[242] : 
                       (N41)? data_i[370] : 
                       (N43)? data_i[498] : 
                       (N38)? data_i[626] : 
                       (N40)? data_i[754] : 
                       (N42)? data_i[882] : 
                       (N44)? data_i[1010] : 1'b0;
  assign data_o[369] = (N37)? data_i[113] : 
                       (N39)? data_i[241] : 
                       (N41)? data_i[369] : 
                       (N43)? data_i[497] : 
                       (N38)? data_i[625] : 
                       (N40)? data_i[753] : 
                       (N42)? data_i[881] : 
                       (N44)? data_i[1009] : 1'b0;
  assign data_o[368] = (N37)? data_i[112] : 
                       (N39)? data_i[240] : 
                       (N41)? data_i[368] : 
                       (N43)? data_i[496] : 
                       (N38)? data_i[624] : 
                       (N40)? data_i[752] : 
                       (N42)? data_i[880] : 
                       (N44)? data_i[1008] : 1'b0;
  assign data_o[367] = (N37)? data_i[111] : 
                       (N39)? data_i[239] : 
                       (N41)? data_i[367] : 
                       (N43)? data_i[495] : 
                       (N38)? data_i[623] : 
                       (N40)? data_i[751] : 
                       (N42)? data_i[879] : 
                       (N44)? data_i[1007] : 1'b0;
  assign data_o[366] = (N37)? data_i[110] : 
                       (N39)? data_i[238] : 
                       (N41)? data_i[366] : 
                       (N43)? data_i[494] : 
                       (N38)? data_i[622] : 
                       (N40)? data_i[750] : 
                       (N42)? data_i[878] : 
                       (N44)? data_i[1006] : 1'b0;
  assign data_o[365] = (N37)? data_i[109] : 
                       (N39)? data_i[237] : 
                       (N41)? data_i[365] : 
                       (N43)? data_i[493] : 
                       (N38)? data_i[621] : 
                       (N40)? data_i[749] : 
                       (N42)? data_i[877] : 
                       (N44)? data_i[1005] : 1'b0;
  assign data_o[364] = (N37)? data_i[108] : 
                       (N39)? data_i[236] : 
                       (N41)? data_i[364] : 
                       (N43)? data_i[492] : 
                       (N38)? data_i[620] : 
                       (N40)? data_i[748] : 
                       (N42)? data_i[876] : 
                       (N44)? data_i[1004] : 1'b0;
  assign data_o[363] = (N37)? data_i[107] : 
                       (N39)? data_i[235] : 
                       (N41)? data_i[363] : 
                       (N43)? data_i[491] : 
                       (N38)? data_i[619] : 
                       (N40)? data_i[747] : 
                       (N42)? data_i[875] : 
                       (N44)? data_i[1003] : 1'b0;
  assign data_o[362] = (N37)? data_i[106] : 
                       (N39)? data_i[234] : 
                       (N41)? data_i[362] : 
                       (N43)? data_i[490] : 
                       (N38)? data_i[618] : 
                       (N40)? data_i[746] : 
                       (N42)? data_i[874] : 
                       (N44)? data_i[1002] : 1'b0;
  assign data_o[361] = (N37)? data_i[105] : 
                       (N39)? data_i[233] : 
                       (N41)? data_i[361] : 
                       (N43)? data_i[489] : 
                       (N38)? data_i[617] : 
                       (N40)? data_i[745] : 
                       (N42)? data_i[873] : 
                       (N44)? data_i[1001] : 1'b0;
  assign data_o[360] = (N37)? data_i[104] : 
                       (N39)? data_i[232] : 
                       (N41)? data_i[360] : 
                       (N43)? data_i[488] : 
                       (N38)? data_i[616] : 
                       (N40)? data_i[744] : 
                       (N42)? data_i[872] : 
                       (N44)? data_i[1000] : 1'b0;
  assign data_o[359] = (N37)? data_i[103] : 
                       (N39)? data_i[231] : 
                       (N41)? data_i[359] : 
                       (N43)? data_i[487] : 
                       (N38)? data_i[615] : 
                       (N40)? data_i[743] : 
                       (N42)? data_i[871] : 
                       (N44)? data_i[999] : 1'b0;
  assign data_o[358] = (N37)? data_i[102] : 
                       (N39)? data_i[230] : 
                       (N41)? data_i[358] : 
                       (N43)? data_i[486] : 
                       (N38)? data_i[614] : 
                       (N40)? data_i[742] : 
                       (N42)? data_i[870] : 
                       (N44)? data_i[998] : 1'b0;
  assign data_o[357] = (N37)? data_i[101] : 
                       (N39)? data_i[229] : 
                       (N41)? data_i[357] : 
                       (N43)? data_i[485] : 
                       (N38)? data_i[613] : 
                       (N40)? data_i[741] : 
                       (N42)? data_i[869] : 
                       (N44)? data_i[997] : 1'b0;
  assign data_o[356] = (N37)? data_i[100] : 
                       (N39)? data_i[228] : 
                       (N41)? data_i[356] : 
                       (N43)? data_i[484] : 
                       (N38)? data_i[612] : 
                       (N40)? data_i[740] : 
                       (N42)? data_i[868] : 
                       (N44)? data_i[996] : 1'b0;
  assign data_o[355] = (N37)? data_i[99] : 
                       (N39)? data_i[227] : 
                       (N41)? data_i[355] : 
                       (N43)? data_i[483] : 
                       (N38)? data_i[611] : 
                       (N40)? data_i[739] : 
                       (N42)? data_i[867] : 
                       (N44)? data_i[995] : 1'b0;
  assign data_o[354] = (N37)? data_i[98] : 
                       (N39)? data_i[226] : 
                       (N41)? data_i[354] : 
                       (N43)? data_i[482] : 
                       (N38)? data_i[610] : 
                       (N40)? data_i[738] : 
                       (N42)? data_i[866] : 
                       (N44)? data_i[994] : 1'b0;
  assign data_o[353] = (N37)? data_i[97] : 
                       (N39)? data_i[225] : 
                       (N41)? data_i[353] : 
                       (N43)? data_i[481] : 
                       (N38)? data_i[609] : 
                       (N40)? data_i[737] : 
                       (N42)? data_i[865] : 
                       (N44)? data_i[993] : 1'b0;
  assign data_o[352] = (N37)? data_i[96] : 
                       (N39)? data_i[224] : 
                       (N41)? data_i[352] : 
                       (N43)? data_i[480] : 
                       (N38)? data_i[608] : 
                       (N40)? data_i[736] : 
                       (N42)? data_i[864] : 
                       (N44)? data_i[992] : 1'b0;
  assign data_o[351] = (N37)? data_i[95] : 
                       (N39)? data_i[223] : 
                       (N41)? data_i[351] : 
                       (N43)? data_i[479] : 
                       (N38)? data_i[607] : 
                       (N40)? data_i[735] : 
                       (N42)? data_i[863] : 
                       (N44)? data_i[991] : 1'b0;
  assign data_o[350] = (N37)? data_i[94] : 
                       (N39)? data_i[222] : 
                       (N41)? data_i[350] : 
                       (N43)? data_i[478] : 
                       (N38)? data_i[606] : 
                       (N40)? data_i[734] : 
                       (N42)? data_i[862] : 
                       (N44)? data_i[990] : 1'b0;
  assign data_o[349] = (N37)? data_i[93] : 
                       (N39)? data_i[221] : 
                       (N41)? data_i[349] : 
                       (N43)? data_i[477] : 
                       (N38)? data_i[605] : 
                       (N40)? data_i[733] : 
                       (N42)? data_i[861] : 
                       (N44)? data_i[989] : 1'b0;
  assign data_o[348] = (N37)? data_i[92] : 
                       (N39)? data_i[220] : 
                       (N41)? data_i[348] : 
                       (N43)? data_i[476] : 
                       (N38)? data_i[604] : 
                       (N40)? data_i[732] : 
                       (N42)? data_i[860] : 
                       (N44)? data_i[988] : 1'b0;
  assign data_o[347] = (N37)? data_i[91] : 
                       (N39)? data_i[219] : 
                       (N41)? data_i[347] : 
                       (N43)? data_i[475] : 
                       (N38)? data_i[603] : 
                       (N40)? data_i[731] : 
                       (N42)? data_i[859] : 
                       (N44)? data_i[987] : 1'b0;
  assign data_o[346] = (N37)? data_i[90] : 
                       (N39)? data_i[218] : 
                       (N41)? data_i[346] : 
                       (N43)? data_i[474] : 
                       (N38)? data_i[602] : 
                       (N40)? data_i[730] : 
                       (N42)? data_i[858] : 
                       (N44)? data_i[986] : 1'b0;
  assign data_o[345] = (N37)? data_i[89] : 
                       (N39)? data_i[217] : 
                       (N41)? data_i[345] : 
                       (N43)? data_i[473] : 
                       (N38)? data_i[601] : 
                       (N40)? data_i[729] : 
                       (N42)? data_i[857] : 
                       (N44)? data_i[985] : 1'b0;
  assign data_o[344] = (N37)? data_i[88] : 
                       (N39)? data_i[216] : 
                       (N41)? data_i[344] : 
                       (N43)? data_i[472] : 
                       (N38)? data_i[600] : 
                       (N40)? data_i[728] : 
                       (N42)? data_i[856] : 
                       (N44)? data_i[984] : 1'b0;
  assign data_o[343] = (N37)? data_i[87] : 
                       (N39)? data_i[215] : 
                       (N41)? data_i[343] : 
                       (N43)? data_i[471] : 
                       (N38)? data_i[599] : 
                       (N40)? data_i[727] : 
                       (N42)? data_i[855] : 
                       (N44)? data_i[983] : 1'b0;
  assign data_o[342] = (N37)? data_i[86] : 
                       (N39)? data_i[214] : 
                       (N41)? data_i[342] : 
                       (N43)? data_i[470] : 
                       (N38)? data_i[598] : 
                       (N40)? data_i[726] : 
                       (N42)? data_i[854] : 
                       (N44)? data_i[982] : 1'b0;
  assign data_o[341] = (N37)? data_i[85] : 
                       (N39)? data_i[213] : 
                       (N41)? data_i[341] : 
                       (N43)? data_i[469] : 
                       (N38)? data_i[597] : 
                       (N40)? data_i[725] : 
                       (N42)? data_i[853] : 
                       (N44)? data_i[981] : 1'b0;
  assign data_o[340] = (N37)? data_i[84] : 
                       (N39)? data_i[212] : 
                       (N41)? data_i[340] : 
                       (N43)? data_i[468] : 
                       (N38)? data_i[596] : 
                       (N40)? data_i[724] : 
                       (N42)? data_i[852] : 
                       (N44)? data_i[980] : 1'b0;
  assign data_o[339] = (N37)? data_i[83] : 
                       (N39)? data_i[211] : 
                       (N41)? data_i[339] : 
                       (N43)? data_i[467] : 
                       (N38)? data_i[595] : 
                       (N40)? data_i[723] : 
                       (N42)? data_i[851] : 
                       (N44)? data_i[979] : 1'b0;
  assign data_o[338] = (N37)? data_i[82] : 
                       (N39)? data_i[210] : 
                       (N41)? data_i[338] : 
                       (N43)? data_i[466] : 
                       (N38)? data_i[594] : 
                       (N40)? data_i[722] : 
                       (N42)? data_i[850] : 
                       (N44)? data_i[978] : 1'b0;
  assign data_o[337] = (N37)? data_i[81] : 
                       (N39)? data_i[209] : 
                       (N41)? data_i[337] : 
                       (N43)? data_i[465] : 
                       (N38)? data_i[593] : 
                       (N40)? data_i[721] : 
                       (N42)? data_i[849] : 
                       (N44)? data_i[977] : 1'b0;
  assign data_o[336] = (N37)? data_i[80] : 
                       (N39)? data_i[208] : 
                       (N41)? data_i[336] : 
                       (N43)? data_i[464] : 
                       (N38)? data_i[592] : 
                       (N40)? data_i[720] : 
                       (N42)? data_i[848] : 
                       (N44)? data_i[976] : 1'b0;
  assign data_o[335] = (N37)? data_i[79] : 
                       (N39)? data_i[207] : 
                       (N41)? data_i[335] : 
                       (N43)? data_i[463] : 
                       (N38)? data_i[591] : 
                       (N40)? data_i[719] : 
                       (N42)? data_i[847] : 
                       (N44)? data_i[975] : 1'b0;
  assign data_o[334] = (N37)? data_i[78] : 
                       (N39)? data_i[206] : 
                       (N41)? data_i[334] : 
                       (N43)? data_i[462] : 
                       (N38)? data_i[590] : 
                       (N40)? data_i[718] : 
                       (N42)? data_i[846] : 
                       (N44)? data_i[974] : 1'b0;
  assign data_o[333] = (N37)? data_i[77] : 
                       (N39)? data_i[205] : 
                       (N41)? data_i[333] : 
                       (N43)? data_i[461] : 
                       (N38)? data_i[589] : 
                       (N40)? data_i[717] : 
                       (N42)? data_i[845] : 
                       (N44)? data_i[973] : 1'b0;
  assign data_o[332] = (N37)? data_i[76] : 
                       (N39)? data_i[204] : 
                       (N41)? data_i[332] : 
                       (N43)? data_i[460] : 
                       (N38)? data_i[588] : 
                       (N40)? data_i[716] : 
                       (N42)? data_i[844] : 
                       (N44)? data_i[972] : 1'b0;
  assign data_o[331] = (N37)? data_i[75] : 
                       (N39)? data_i[203] : 
                       (N41)? data_i[331] : 
                       (N43)? data_i[459] : 
                       (N38)? data_i[587] : 
                       (N40)? data_i[715] : 
                       (N42)? data_i[843] : 
                       (N44)? data_i[971] : 1'b0;
  assign data_o[330] = (N37)? data_i[74] : 
                       (N39)? data_i[202] : 
                       (N41)? data_i[330] : 
                       (N43)? data_i[458] : 
                       (N38)? data_i[586] : 
                       (N40)? data_i[714] : 
                       (N42)? data_i[842] : 
                       (N44)? data_i[970] : 1'b0;
  assign data_o[329] = (N37)? data_i[73] : 
                       (N39)? data_i[201] : 
                       (N41)? data_i[329] : 
                       (N43)? data_i[457] : 
                       (N38)? data_i[585] : 
                       (N40)? data_i[713] : 
                       (N42)? data_i[841] : 
                       (N44)? data_i[969] : 1'b0;
  assign data_o[328] = (N37)? data_i[72] : 
                       (N39)? data_i[200] : 
                       (N41)? data_i[328] : 
                       (N43)? data_i[456] : 
                       (N38)? data_i[584] : 
                       (N40)? data_i[712] : 
                       (N42)? data_i[840] : 
                       (N44)? data_i[968] : 1'b0;
  assign data_o[327] = (N37)? data_i[71] : 
                       (N39)? data_i[199] : 
                       (N41)? data_i[327] : 
                       (N43)? data_i[455] : 
                       (N38)? data_i[583] : 
                       (N40)? data_i[711] : 
                       (N42)? data_i[839] : 
                       (N44)? data_i[967] : 1'b0;
  assign data_o[326] = (N37)? data_i[70] : 
                       (N39)? data_i[198] : 
                       (N41)? data_i[326] : 
                       (N43)? data_i[454] : 
                       (N38)? data_i[582] : 
                       (N40)? data_i[710] : 
                       (N42)? data_i[838] : 
                       (N44)? data_i[966] : 1'b0;
  assign data_o[325] = (N37)? data_i[69] : 
                       (N39)? data_i[197] : 
                       (N41)? data_i[325] : 
                       (N43)? data_i[453] : 
                       (N38)? data_i[581] : 
                       (N40)? data_i[709] : 
                       (N42)? data_i[837] : 
                       (N44)? data_i[965] : 1'b0;
  assign data_o[324] = (N37)? data_i[68] : 
                       (N39)? data_i[196] : 
                       (N41)? data_i[324] : 
                       (N43)? data_i[452] : 
                       (N38)? data_i[580] : 
                       (N40)? data_i[708] : 
                       (N42)? data_i[836] : 
                       (N44)? data_i[964] : 1'b0;
  assign data_o[323] = (N37)? data_i[67] : 
                       (N39)? data_i[195] : 
                       (N41)? data_i[323] : 
                       (N43)? data_i[451] : 
                       (N38)? data_i[579] : 
                       (N40)? data_i[707] : 
                       (N42)? data_i[835] : 
                       (N44)? data_i[963] : 1'b0;
  assign data_o[322] = (N37)? data_i[66] : 
                       (N39)? data_i[194] : 
                       (N41)? data_i[322] : 
                       (N43)? data_i[450] : 
                       (N38)? data_i[578] : 
                       (N40)? data_i[706] : 
                       (N42)? data_i[834] : 
                       (N44)? data_i[962] : 1'b0;
  assign data_o[321] = (N37)? data_i[65] : 
                       (N39)? data_i[193] : 
                       (N41)? data_i[321] : 
                       (N43)? data_i[449] : 
                       (N38)? data_i[577] : 
                       (N40)? data_i[705] : 
                       (N42)? data_i[833] : 
                       (N44)? data_i[961] : 1'b0;
  assign data_o[320] = (N37)? data_i[64] : 
                       (N39)? data_i[192] : 
                       (N41)? data_i[320] : 
                       (N43)? data_i[448] : 
                       (N38)? data_i[576] : 
                       (N40)? data_i[704] : 
                       (N42)? data_i[832] : 
                       (N44)? data_i[960] : 1'b0;
  assign data_o[319] = (N37)? data_i[63] : 
                       (N39)? data_i[191] : 
                       (N41)? data_i[319] : 
                       (N43)? data_i[447] : 
                       (N38)? data_i[575] : 
                       (N40)? data_i[703] : 
                       (N42)? data_i[831] : 
                       (N44)? data_i[959] : 1'b0;
  assign data_o[318] = (N37)? data_i[62] : 
                       (N39)? data_i[190] : 
                       (N41)? data_i[318] : 
                       (N43)? data_i[446] : 
                       (N38)? data_i[574] : 
                       (N40)? data_i[702] : 
                       (N42)? data_i[830] : 
                       (N44)? data_i[958] : 1'b0;
  assign data_o[317] = (N37)? data_i[61] : 
                       (N39)? data_i[189] : 
                       (N41)? data_i[317] : 
                       (N43)? data_i[445] : 
                       (N38)? data_i[573] : 
                       (N40)? data_i[701] : 
                       (N42)? data_i[829] : 
                       (N44)? data_i[957] : 1'b0;
  assign data_o[316] = (N37)? data_i[60] : 
                       (N39)? data_i[188] : 
                       (N41)? data_i[316] : 
                       (N43)? data_i[444] : 
                       (N38)? data_i[572] : 
                       (N40)? data_i[700] : 
                       (N42)? data_i[828] : 
                       (N44)? data_i[956] : 1'b0;
  assign data_o[315] = (N37)? data_i[59] : 
                       (N39)? data_i[187] : 
                       (N41)? data_i[315] : 
                       (N43)? data_i[443] : 
                       (N38)? data_i[571] : 
                       (N40)? data_i[699] : 
                       (N42)? data_i[827] : 
                       (N44)? data_i[955] : 1'b0;
  assign data_o[314] = (N37)? data_i[58] : 
                       (N39)? data_i[186] : 
                       (N41)? data_i[314] : 
                       (N43)? data_i[442] : 
                       (N38)? data_i[570] : 
                       (N40)? data_i[698] : 
                       (N42)? data_i[826] : 
                       (N44)? data_i[954] : 1'b0;
  assign data_o[313] = (N37)? data_i[57] : 
                       (N39)? data_i[185] : 
                       (N41)? data_i[313] : 
                       (N43)? data_i[441] : 
                       (N38)? data_i[569] : 
                       (N40)? data_i[697] : 
                       (N42)? data_i[825] : 
                       (N44)? data_i[953] : 1'b0;
  assign data_o[312] = (N37)? data_i[56] : 
                       (N39)? data_i[184] : 
                       (N41)? data_i[312] : 
                       (N43)? data_i[440] : 
                       (N38)? data_i[568] : 
                       (N40)? data_i[696] : 
                       (N42)? data_i[824] : 
                       (N44)? data_i[952] : 1'b0;
  assign data_o[311] = (N37)? data_i[55] : 
                       (N39)? data_i[183] : 
                       (N41)? data_i[311] : 
                       (N43)? data_i[439] : 
                       (N38)? data_i[567] : 
                       (N40)? data_i[695] : 
                       (N42)? data_i[823] : 
                       (N44)? data_i[951] : 1'b0;
  assign data_o[310] = (N37)? data_i[54] : 
                       (N39)? data_i[182] : 
                       (N41)? data_i[310] : 
                       (N43)? data_i[438] : 
                       (N38)? data_i[566] : 
                       (N40)? data_i[694] : 
                       (N42)? data_i[822] : 
                       (N44)? data_i[950] : 1'b0;
  assign data_o[309] = (N37)? data_i[53] : 
                       (N39)? data_i[181] : 
                       (N41)? data_i[309] : 
                       (N43)? data_i[437] : 
                       (N38)? data_i[565] : 
                       (N40)? data_i[693] : 
                       (N42)? data_i[821] : 
                       (N44)? data_i[949] : 1'b0;
  assign data_o[308] = (N37)? data_i[52] : 
                       (N39)? data_i[180] : 
                       (N41)? data_i[308] : 
                       (N43)? data_i[436] : 
                       (N38)? data_i[564] : 
                       (N40)? data_i[692] : 
                       (N42)? data_i[820] : 
                       (N44)? data_i[948] : 1'b0;
  assign data_o[307] = (N37)? data_i[51] : 
                       (N39)? data_i[179] : 
                       (N41)? data_i[307] : 
                       (N43)? data_i[435] : 
                       (N38)? data_i[563] : 
                       (N40)? data_i[691] : 
                       (N42)? data_i[819] : 
                       (N44)? data_i[947] : 1'b0;
  assign data_o[306] = (N37)? data_i[50] : 
                       (N39)? data_i[178] : 
                       (N41)? data_i[306] : 
                       (N43)? data_i[434] : 
                       (N38)? data_i[562] : 
                       (N40)? data_i[690] : 
                       (N42)? data_i[818] : 
                       (N44)? data_i[946] : 1'b0;
  assign data_o[305] = (N37)? data_i[49] : 
                       (N39)? data_i[177] : 
                       (N41)? data_i[305] : 
                       (N43)? data_i[433] : 
                       (N38)? data_i[561] : 
                       (N40)? data_i[689] : 
                       (N42)? data_i[817] : 
                       (N44)? data_i[945] : 1'b0;
  assign data_o[304] = (N37)? data_i[48] : 
                       (N39)? data_i[176] : 
                       (N41)? data_i[304] : 
                       (N43)? data_i[432] : 
                       (N38)? data_i[560] : 
                       (N40)? data_i[688] : 
                       (N42)? data_i[816] : 
                       (N44)? data_i[944] : 1'b0;
  assign data_o[303] = (N37)? data_i[47] : 
                       (N39)? data_i[175] : 
                       (N41)? data_i[303] : 
                       (N43)? data_i[431] : 
                       (N38)? data_i[559] : 
                       (N40)? data_i[687] : 
                       (N42)? data_i[815] : 
                       (N44)? data_i[943] : 1'b0;
  assign data_o[302] = (N37)? data_i[46] : 
                       (N39)? data_i[174] : 
                       (N41)? data_i[302] : 
                       (N43)? data_i[430] : 
                       (N38)? data_i[558] : 
                       (N40)? data_i[686] : 
                       (N42)? data_i[814] : 
                       (N44)? data_i[942] : 1'b0;
  assign data_o[301] = (N37)? data_i[45] : 
                       (N39)? data_i[173] : 
                       (N41)? data_i[301] : 
                       (N43)? data_i[429] : 
                       (N38)? data_i[557] : 
                       (N40)? data_i[685] : 
                       (N42)? data_i[813] : 
                       (N44)? data_i[941] : 1'b0;
  assign data_o[300] = (N37)? data_i[44] : 
                       (N39)? data_i[172] : 
                       (N41)? data_i[300] : 
                       (N43)? data_i[428] : 
                       (N38)? data_i[556] : 
                       (N40)? data_i[684] : 
                       (N42)? data_i[812] : 
                       (N44)? data_i[940] : 1'b0;
  assign data_o[299] = (N37)? data_i[43] : 
                       (N39)? data_i[171] : 
                       (N41)? data_i[299] : 
                       (N43)? data_i[427] : 
                       (N38)? data_i[555] : 
                       (N40)? data_i[683] : 
                       (N42)? data_i[811] : 
                       (N44)? data_i[939] : 1'b0;
  assign data_o[298] = (N37)? data_i[42] : 
                       (N39)? data_i[170] : 
                       (N41)? data_i[298] : 
                       (N43)? data_i[426] : 
                       (N38)? data_i[554] : 
                       (N40)? data_i[682] : 
                       (N42)? data_i[810] : 
                       (N44)? data_i[938] : 1'b0;
  assign data_o[297] = (N37)? data_i[41] : 
                       (N39)? data_i[169] : 
                       (N41)? data_i[297] : 
                       (N43)? data_i[425] : 
                       (N38)? data_i[553] : 
                       (N40)? data_i[681] : 
                       (N42)? data_i[809] : 
                       (N44)? data_i[937] : 1'b0;
  assign data_o[296] = (N37)? data_i[40] : 
                       (N39)? data_i[168] : 
                       (N41)? data_i[296] : 
                       (N43)? data_i[424] : 
                       (N38)? data_i[552] : 
                       (N40)? data_i[680] : 
                       (N42)? data_i[808] : 
                       (N44)? data_i[936] : 1'b0;
  assign data_o[295] = (N37)? data_i[39] : 
                       (N39)? data_i[167] : 
                       (N41)? data_i[295] : 
                       (N43)? data_i[423] : 
                       (N38)? data_i[551] : 
                       (N40)? data_i[679] : 
                       (N42)? data_i[807] : 
                       (N44)? data_i[935] : 1'b0;
  assign data_o[294] = (N37)? data_i[38] : 
                       (N39)? data_i[166] : 
                       (N41)? data_i[294] : 
                       (N43)? data_i[422] : 
                       (N38)? data_i[550] : 
                       (N40)? data_i[678] : 
                       (N42)? data_i[806] : 
                       (N44)? data_i[934] : 1'b0;
  assign data_o[293] = (N37)? data_i[37] : 
                       (N39)? data_i[165] : 
                       (N41)? data_i[293] : 
                       (N43)? data_i[421] : 
                       (N38)? data_i[549] : 
                       (N40)? data_i[677] : 
                       (N42)? data_i[805] : 
                       (N44)? data_i[933] : 1'b0;
  assign data_o[292] = (N37)? data_i[36] : 
                       (N39)? data_i[164] : 
                       (N41)? data_i[292] : 
                       (N43)? data_i[420] : 
                       (N38)? data_i[548] : 
                       (N40)? data_i[676] : 
                       (N42)? data_i[804] : 
                       (N44)? data_i[932] : 1'b0;
  assign data_o[291] = (N37)? data_i[35] : 
                       (N39)? data_i[163] : 
                       (N41)? data_i[291] : 
                       (N43)? data_i[419] : 
                       (N38)? data_i[547] : 
                       (N40)? data_i[675] : 
                       (N42)? data_i[803] : 
                       (N44)? data_i[931] : 1'b0;
  assign data_o[290] = (N37)? data_i[34] : 
                       (N39)? data_i[162] : 
                       (N41)? data_i[290] : 
                       (N43)? data_i[418] : 
                       (N38)? data_i[546] : 
                       (N40)? data_i[674] : 
                       (N42)? data_i[802] : 
                       (N44)? data_i[930] : 1'b0;
  assign data_o[289] = (N37)? data_i[33] : 
                       (N39)? data_i[161] : 
                       (N41)? data_i[289] : 
                       (N43)? data_i[417] : 
                       (N38)? data_i[545] : 
                       (N40)? data_i[673] : 
                       (N42)? data_i[801] : 
                       (N44)? data_i[929] : 1'b0;
  assign data_o[288] = (N37)? data_i[32] : 
                       (N39)? data_i[160] : 
                       (N41)? data_i[288] : 
                       (N43)? data_i[416] : 
                       (N38)? data_i[544] : 
                       (N40)? data_i[672] : 
                       (N42)? data_i[800] : 
                       (N44)? data_i[928] : 1'b0;
  assign data_o[287] = (N37)? data_i[31] : 
                       (N39)? data_i[159] : 
                       (N41)? data_i[287] : 
                       (N43)? data_i[415] : 
                       (N38)? data_i[543] : 
                       (N40)? data_i[671] : 
                       (N42)? data_i[799] : 
                       (N44)? data_i[927] : 1'b0;
  assign data_o[286] = (N37)? data_i[30] : 
                       (N39)? data_i[158] : 
                       (N41)? data_i[286] : 
                       (N43)? data_i[414] : 
                       (N38)? data_i[542] : 
                       (N40)? data_i[670] : 
                       (N42)? data_i[798] : 
                       (N44)? data_i[926] : 1'b0;
  assign data_o[285] = (N37)? data_i[29] : 
                       (N39)? data_i[157] : 
                       (N41)? data_i[285] : 
                       (N43)? data_i[413] : 
                       (N38)? data_i[541] : 
                       (N40)? data_i[669] : 
                       (N42)? data_i[797] : 
                       (N44)? data_i[925] : 1'b0;
  assign data_o[284] = (N37)? data_i[28] : 
                       (N39)? data_i[156] : 
                       (N41)? data_i[284] : 
                       (N43)? data_i[412] : 
                       (N38)? data_i[540] : 
                       (N40)? data_i[668] : 
                       (N42)? data_i[796] : 
                       (N44)? data_i[924] : 1'b0;
  assign data_o[283] = (N37)? data_i[27] : 
                       (N39)? data_i[155] : 
                       (N41)? data_i[283] : 
                       (N43)? data_i[411] : 
                       (N38)? data_i[539] : 
                       (N40)? data_i[667] : 
                       (N42)? data_i[795] : 
                       (N44)? data_i[923] : 1'b0;
  assign data_o[282] = (N37)? data_i[26] : 
                       (N39)? data_i[154] : 
                       (N41)? data_i[282] : 
                       (N43)? data_i[410] : 
                       (N38)? data_i[538] : 
                       (N40)? data_i[666] : 
                       (N42)? data_i[794] : 
                       (N44)? data_i[922] : 1'b0;
  assign data_o[281] = (N37)? data_i[25] : 
                       (N39)? data_i[153] : 
                       (N41)? data_i[281] : 
                       (N43)? data_i[409] : 
                       (N38)? data_i[537] : 
                       (N40)? data_i[665] : 
                       (N42)? data_i[793] : 
                       (N44)? data_i[921] : 1'b0;
  assign data_o[280] = (N37)? data_i[24] : 
                       (N39)? data_i[152] : 
                       (N41)? data_i[280] : 
                       (N43)? data_i[408] : 
                       (N38)? data_i[536] : 
                       (N40)? data_i[664] : 
                       (N42)? data_i[792] : 
                       (N44)? data_i[920] : 1'b0;
  assign data_o[279] = (N37)? data_i[23] : 
                       (N39)? data_i[151] : 
                       (N41)? data_i[279] : 
                       (N43)? data_i[407] : 
                       (N38)? data_i[535] : 
                       (N40)? data_i[663] : 
                       (N42)? data_i[791] : 
                       (N44)? data_i[919] : 1'b0;
  assign data_o[278] = (N37)? data_i[22] : 
                       (N39)? data_i[150] : 
                       (N41)? data_i[278] : 
                       (N43)? data_i[406] : 
                       (N38)? data_i[534] : 
                       (N40)? data_i[662] : 
                       (N42)? data_i[790] : 
                       (N44)? data_i[918] : 1'b0;
  assign data_o[277] = (N37)? data_i[21] : 
                       (N39)? data_i[149] : 
                       (N41)? data_i[277] : 
                       (N43)? data_i[405] : 
                       (N38)? data_i[533] : 
                       (N40)? data_i[661] : 
                       (N42)? data_i[789] : 
                       (N44)? data_i[917] : 1'b0;
  assign data_o[276] = (N37)? data_i[20] : 
                       (N39)? data_i[148] : 
                       (N41)? data_i[276] : 
                       (N43)? data_i[404] : 
                       (N38)? data_i[532] : 
                       (N40)? data_i[660] : 
                       (N42)? data_i[788] : 
                       (N44)? data_i[916] : 1'b0;
  assign data_o[275] = (N37)? data_i[19] : 
                       (N39)? data_i[147] : 
                       (N41)? data_i[275] : 
                       (N43)? data_i[403] : 
                       (N38)? data_i[531] : 
                       (N40)? data_i[659] : 
                       (N42)? data_i[787] : 
                       (N44)? data_i[915] : 1'b0;
  assign data_o[274] = (N37)? data_i[18] : 
                       (N39)? data_i[146] : 
                       (N41)? data_i[274] : 
                       (N43)? data_i[402] : 
                       (N38)? data_i[530] : 
                       (N40)? data_i[658] : 
                       (N42)? data_i[786] : 
                       (N44)? data_i[914] : 1'b0;
  assign data_o[273] = (N37)? data_i[17] : 
                       (N39)? data_i[145] : 
                       (N41)? data_i[273] : 
                       (N43)? data_i[401] : 
                       (N38)? data_i[529] : 
                       (N40)? data_i[657] : 
                       (N42)? data_i[785] : 
                       (N44)? data_i[913] : 1'b0;
  assign data_o[272] = (N37)? data_i[16] : 
                       (N39)? data_i[144] : 
                       (N41)? data_i[272] : 
                       (N43)? data_i[400] : 
                       (N38)? data_i[528] : 
                       (N40)? data_i[656] : 
                       (N42)? data_i[784] : 
                       (N44)? data_i[912] : 1'b0;
  assign data_o[271] = (N37)? data_i[15] : 
                       (N39)? data_i[143] : 
                       (N41)? data_i[271] : 
                       (N43)? data_i[399] : 
                       (N38)? data_i[527] : 
                       (N40)? data_i[655] : 
                       (N42)? data_i[783] : 
                       (N44)? data_i[911] : 1'b0;
  assign data_o[270] = (N37)? data_i[14] : 
                       (N39)? data_i[142] : 
                       (N41)? data_i[270] : 
                       (N43)? data_i[398] : 
                       (N38)? data_i[526] : 
                       (N40)? data_i[654] : 
                       (N42)? data_i[782] : 
                       (N44)? data_i[910] : 1'b0;
  assign data_o[269] = (N37)? data_i[13] : 
                       (N39)? data_i[141] : 
                       (N41)? data_i[269] : 
                       (N43)? data_i[397] : 
                       (N38)? data_i[525] : 
                       (N40)? data_i[653] : 
                       (N42)? data_i[781] : 
                       (N44)? data_i[909] : 1'b0;
  assign data_o[268] = (N37)? data_i[12] : 
                       (N39)? data_i[140] : 
                       (N41)? data_i[268] : 
                       (N43)? data_i[396] : 
                       (N38)? data_i[524] : 
                       (N40)? data_i[652] : 
                       (N42)? data_i[780] : 
                       (N44)? data_i[908] : 1'b0;
  assign data_o[267] = (N37)? data_i[11] : 
                       (N39)? data_i[139] : 
                       (N41)? data_i[267] : 
                       (N43)? data_i[395] : 
                       (N38)? data_i[523] : 
                       (N40)? data_i[651] : 
                       (N42)? data_i[779] : 
                       (N44)? data_i[907] : 1'b0;
  assign data_o[266] = (N37)? data_i[10] : 
                       (N39)? data_i[138] : 
                       (N41)? data_i[266] : 
                       (N43)? data_i[394] : 
                       (N38)? data_i[522] : 
                       (N40)? data_i[650] : 
                       (N42)? data_i[778] : 
                       (N44)? data_i[906] : 1'b0;
  assign data_o[265] = (N37)? data_i[9] : 
                       (N39)? data_i[137] : 
                       (N41)? data_i[265] : 
                       (N43)? data_i[393] : 
                       (N38)? data_i[521] : 
                       (N40)? data_i[649] : 
                       (N42)? data_i[777] : 
                       (N44)? data_i[905] : 1'b0;
  assign data_o[264] = (N37)? data_i[8] : 
                       (N39)? data_i[136] : 
                       (N41)? data_i[264] : 
                       (N43)? data_i[392] : 
                       (N38)? data_i[520] : 
                       (N40)? data_i[648] : 
                       (N42)? data_i[776] : 
                       (N44)? data_i[904] : 1'b0;
  assign data_o[263] = (N37)? data_i[7] : 
                       (N39)? data_i[135] : 
                       (N41)? data_i[263] : 
                       (N43)? data_i[391] : 
                       (N38)? data_i[519] : 
                       (N40)? data_i[647] : 
                       (N42)? data_i[775] : 
                       (N44)? data_i[903] : 1'b0;
  assign data_o[262] = (N37)? data_i[6] : 
                       (N39)? data_i[134] : 
                       (N41)? data_i[262] : 
                       (N43)? data_i[390] : 
                       (N38)? data_i[518] : 
                       (N40)? data_i[646] : 
                       (N42)? data_i[774] : 
                       (N44)? data_i[902] : 1'b0;
  assign data_o[261] = (N37)? data_i[5] : 
                       (N39)? data_i[133] : 
                       (N41)? data_i[261] : 
                       (N43)? data_i[389] : 
                       (N38)? data_i[517] : 
                       (N40)? data_i[645] : 
                       (N42)? data_i[773] : 
                       (N44)? data_i[901] : 1'b0;
  assign data_o[260] = (N37)? data_i[4] : 
                       (N39)? data_i[132] : 
                       (N41)? data_i[260] : 
                       (N43)? data_i[388] : 
                       (N38)? data_i[516] : 
                       (N40)? data_i[644] : 
                       (N42)? data_i[772] : 
                       (N44)? data_i[900] : 1'b0;
  assign data_o[259] = (N37)? data_i[3] : 
                       (N39)? data_i[131] : 
                       (N41)? data_i[259] : 
                       (N43)? data_i[387] : 
                       (N38)? data_i[515] : 
                       (N40)? data_i[643] : 
                       (N42)? data_i[771] : 
                       (N44)? data_i[899] : 1'b0;
  assign data_o[258] = (N37)? data_i[2] : 
                       (N39)? data_i[130] : 
                       (N41)? data_i[258] : 
                       (N43)? data_i[386] : 
                       (N38)? data_i[514] : 
                       (N40)? data_i[642] : 
                       (N42)? data_i[770] : 
                       (N44)? data_i[898] : 1'b0;
  assign data_o[257] = (N37)? data_i[1] : 
                       (N39)? data_i[129] : 
                       (N41)? data_i[257] : 
                       (N43)? data_i[385] : 
                       (N38)? data_i[513] : 
                       (N40)? data_i[641] : 
                       (N42)? data_i[769] : 
                       (N44)? data_i[897] : 1'b0;
  assign data_o[256] = (N37)? data_i[0] : 
                       (N39)? data_i[128] : 
                       (N41)? data_i[256] : 
                       (N43)? data_i[384] : 
                       (N38)? data_i[512] : 
                       (N40)? data_i[640] : 
                       (N42)? data_i[768] : 
                       (N44)? data_i[896] : 1'b0;
  assign data_o[511] = (N52)? data_i[127] : 
                       (N54)? data_i[255] : 
                       (N56)? data_i[383] : 
                       (N58)? data_i[511] : 
                       (N53)? data_i[639] : 
                       (N55)? data_i[767] : 
                       (N57)? data_i[895] : 
                       (N59)? data_i[1023] : 1'b0;
  assign data_o[510] = (N52)? data_i[126] : 
                       (N54)? data_i[254] : 
                       (N56)? data_i[382] : 
                       (N58)? data_i[510] : 
                       (N53)? data_i[638] : 
                       (N55)? data_i[766] : 
                       (N57)? data_i[894] : 
                       (N59)? data_i[1022] : 1'b0;
  assign data_o[509] = (N52)? data_i[125] : 
                       (N54)? data_i[253] : 
                       (N56)? data_i[381] : 
                       (N58)? data_i[509] : 
                       (N53)? data_i[637] : 
                       (N55)? data_i[765] : 
                       (N57)? data_i[893] : 
                       (N59)? data_i[1021] : 1'b0;
  assign data_o[508] = (N52)? data_i[124] : 
                       (N54)? data_i[252] : 
                       (N56)? data_i[380] : 
                       (N58)? data_i[508] : 
                       (N53)? data_i[636] : 
                       (N55)? data_i[764] : 
                       (N57)? data_i[892] : 
                       (N59)? data_i[1020] : 1'b0;
  assign data_o[507] = (N52)? data_i[123] : 
                       (N54)? data_i[251] : 
                       (N56)? data_i[379] : 
                       (N58)? data_i[507] : 
                       (N53)? data_i[635] : 
                       (N55)? data_i[763] : 
                       (N57)? data_i[891] : 
                       (N59)? data_i[1019] : 1'b0;
  assign data_o[506] = (N52)? data_i[122] : 
                       (N54)? data_i[250] : 
                       (N56)? data_i[378] : 
                       (N58)? data_i[506] : 
                       (N53)? data_i[634] : 
                       (N55)? data_i[762] : 
                       (N57)? data_i[890] : 
                       (N59)? data_i[1018] : 1'b0;
  assign data_o[505] = (N52)? data_i[121] : 
                       (N54)? data_i[249] : 
                       (N56)? data_i[377] : 
                       (N58)? data_i[505] : 
                       (N53)? data_i[633] : 
                       (N55)? data_i[761] : 
                       (N57)? data_i[889] : 
                       (N59)? data_i[1017] : 1'b0;
  assign data_o[504] = (N52)? data_i[120] : 
                       (N54)? data_i[248] : 
                       (N56)? data_i[376] : 
                       (N58)? data_i[504] : 
                       (N53)? data_i[632] : 
                       (N55)? data_i[760] : 
                       (N57)? data_i[888] : 
                       (N59)? data_i[1016] : 1'b0;
  assign data_o[503] = (N52)? data_i[119] : 
                       (N54)? data_i[247] : 
                       (N56)? data_i[375] : 
                       (N58)? data_i[503] : 
                       (N53)? data_i[631] : 
                       (N55)? data_i[759] : 
                       (N57)? data_i[887] : 
                       (N59)? data_i[1015] : 1'b0;
  assign data_o[502] = (N52)? data_i[118] : 
                       (N54)? data_i[246] : 
                       (N56)? data_i[374] : 
                       (N58)? data_i[502] : 
                       (N53)? data_i[630] : 
                       (N55)? data_i[758] : 
                       (N57)? data_i[886] : 
                       (N59)? data_i[1014] : 1'b0;
  assign data_o[501] = (N52)? data_i[117] : 
                       (N54)? data_i[245] : 
                       (N56)? data_i[373] : 
                       (N58)? data_i[501] : 
                       (N53)? data_i[629] : 
                       (N55)? data_i[757] : 
                       (N57)? data_i[885] : 
                       (N59)? data_i[1013] : 1'b0;
  assign data_o[500] = (N52)? data_i[116] : 
                       (N54)? data_i[244] : 
                       (N56)? data_i[372] : 
                       (N58)? data_i[500] : 
                       (N53)? data_i[628] : 
                       (N55)? data_i[756] : 
                       (N57)? data_i[884] : 
                       (N59)? data_i[1012] : 1'b0;
  assign data_o[499] = (N52)? data_i[115] : 
                       (N54)? data_i[243] : 
                       (N56)? data_i[371] : 
                       (N58)? data_i[499] : 
                       (N53)? data_i[627] : 
                       (N55)? data_i[755] : 
                       (N57)? data_i[883] : 
                       (N59)? data_i[1011] : 1'b0;
  assign data_o[498] = (N52)? data_i[114] : 
                       (N54)? data_i[242] : 
                       (N56)? data_i[370] : 
                       (N58)? data_i[498] : 
                       (N53)? data_i[626] : 
                       (N55)? data_i[754] : 
                       (N57)? data_i[882] : 
                       (N59)? data_i[1010] : 1'b0;
  assign data_o[497] = (N52)? data_i[113] : 
                       (N54)? data_i[241] : 
                       (N56)? data_i[369] : 
                       (N58)? data_i[497] : 
                       (N53)? data_i[625] : 
                       (N55)? data_i[753] : 
                       (N57)? data_i[881] : 
                       (N59)? data_i[1009] : 1'b0;
  assign data_o[496] = (N52)? data_i[112] : 
                       (N54)? data_i[240] : 
                       (N56)? data_i[368] : 
                       (N58)? data_i[496] : 
                       (N53)? data_i[624] : 
                       (N55)? data_i[752] : 
                       (N57)? data_i[880] : 
                       (N59)? data_i[1008] : 1'b0;
  assign data_o[495] = (N52)? data_i[111] : 
                       (N54)? data_i[239] : 
                       (N56)? data_i[367] : 
                       (N58)? data_i[495] : 
                       (N53)? data_i[623] : 
                       (N55)? data_i[751] : 
                       (N57)? data_i[879] : 
                       (N59)? data_i[1007] : 1'b0;
  assign data_o[494] = (N52)? data_i[110] : 
                       (N54)? data_i[238] : 
                       (N56)? data_i[366] : 
                       (N58)? data_i[494] : 
                       (N53)? data_i[622] : 
                       (N55)? data_i[750] : 
                       (N57)? data_i[878] : 
                       (N59)? data_i[1006] : 1'b0;
  assign data_o[493] = (N52)? data_i[109] : 
                       (N54)? data_i[237] : 
                       (N56)? data_i[365] : 
                       (N58)? data_i[493] : 
                       (N53)? data_i[621] : 
                       (N55)? data_i[749] : 
                       (N57)? data_i[877] : 
                       (N59)? data_i[1005] : 1'b0;
  assign data_o[492] = (N52)? data_i[108] : 
                       (N54)? data_i[236] : 
                       (N56)? data_i[364] : 
                       (N58)? data_i[492] : 
                       (N53)? data_i[620] : 
                       (N55)? data_i[748] : 
                       (N57)? data_i[876] : 
                       (N59)? data_i[1004] : 1'b0;
  assign data_o[491] = (N52)? data_i[107] : 
                       (N54)? data_i[235] : 
                       (N56)? data_i[363] : 
                       (N58)? data_i[491] : 
                       (N53)? data_i[619] : 
                       (N55)? data_i[747] : 
                       (N57)? data_i[875] : 
                       (N59)? data_i[1003] : 1'b0;
  assign data_o[490] = (N52)? data_i[106] : 
                       (N54)? data_i[234] : 
                       (N56)? data_i[362] : 
                       (N58)? data_i[490] : 
                       (N53)? data_i[618] : 
                       (N55)? data_i[746] : 
                       (N57)? data_i[874] : 
                       (N59)? data_i[1002] : 1'b0;
  assign data_o[489] = (N52)? data_i[105] : 
                       (N54)? data_i[233] : 
                       (N56)? data_i[361] : 
                       (N58)? data_i[489] : 
                       (N53)? data_i[617] : 
                       (N55)? data_i[745] : 
                       (N57)? data_i[873] : 
                       (N59)? data_i[1001] : 1'b0;
  assign data_o[488] = (N52)? data_i[104] : 
                       (N54)? data_i[232] : 
                       (N56)? data_i[360] : 
                       (N58)? data_i[488] : 
                       (N53)? data_i[616] : 
                       (N55)? data_i[744] : 
                       (N57)? data_i[872] : 
                       (N59)? data_i[1000] : 1'b0;
  assign data_o[487] = (N52)? data_i[103] : 
                       (N54)? data_i[231] : 
                       (N56)? data_i[359] : 
                       (N58)? data_i[487] : 
                       (N53)? data_i[615] : 
                       (N55)? data_i[743] : 
                       (N57)? data_i[871] : 
                       (N59)? data_i[999] : 1'b0;
  assign data_o[486] = (N52)? data_i[102] : 
                       (N54)? data_i[230] : 
                       (N56)? data_i[358] : 
                       (N58)? data_i[486] : 
                       (N53)? data_i[614] : 
                       (N55)? data_i[742] : 
                       (N57)? data_i[870] : 
                       (N59)? data_i[998] : 1'b0;
  assign data_o[485] = (N52)? data_i[101] : 
                       (N54)? data_i[229] : 
                       (N56)? data_i[357] : 
                       (N58)? data_i[485] : 
                       (N53)? data_i[613] : 
                       (N55)? data_i[741] : 
                       (N57)? data_i[869] : 
                       (N59)? data_i[997] : 1'b0;
  assign data_o[484] = (N52)? data_i[100] : 
                       (N54)? data_i[228] : 
                       (N56)? data_i[356] : 
                       (N58)? data_i[484] : 
                       (N53)? data_i[612] : 
                       (N55)? data_i[740] : 
                       (N57)? data_i[868] : 
                       (N59)? data_i[996] : 1'b0;
  assign data_o[483] = (N52)? data_i[99] : 
                       (N54)? data_i[227] : 
                       (N56)? data_i[355] : 
                       (N58)? data_i[483] : 
                       (N53)? data_i[611] : 
                       (N55)? data_i[739] : 
                       (N57)? data_i[867] : 
                       (N59)? data_i[995] : 1'b0;
  assign data_o[482] = (N52)? data_i[98] : 
                       (N54)? data_i[226] : 
                       (N56)? data_i[354] : 
                       (N58)? data_i[482] : 
                       (N53)? data_i[610] : 
                       (N55)? data_i[738] : 
                       (N57)? data_i[866] : 
                       (N59)? data_i[994] : 1'b0;
  assign data_o[481] = (N52)? data_i[97] : 
                       (N54)? data_i[225] : 
                       (N56)? data_i[353] : 
                       (N58)? data_i[481] : 
                       (N53)? data_i[609] : 
                       (N55)? data_i[737] : 
                       (N57)? data_i[865] : 
                       (N59)? data_i[993] : 1'b0;
  assign data_o[480] = (N52)? data_i[96] : 
                       (N54)? data_i[224] : 
                       (N56)? data_i[352] : 
                       (N58)? data_i[480] : 
                       (N53)? data_i[608] : 
                       (N55)? data_i[736] : 
                       (N57)? data_i[864] : 
                       (N59)? data_i[992] : 1'b0;
  assign data_o[479] = (N52)? data_i[95] : 
                       (N54)? data_i[223] : 
                       (N56)? data_i[351] : 
                       (N58)? data_i[479] : 
                       (N53)? data_i[607] : 
                       (N55)? data_i[735] : 
                       (N57)? data_i[863] : 
                       (N59)? data_i[991] : 1'b0;
  assign data_o[478] = (N52)? data_i[94] : 
                       (N54)? data_i[222] : 
                       (N56)? data_i[350] : 
                       (N58)? data_i[478] : 
                       (N53)? data_i[606] : 
                       (N55)? data_i[734] : 
                       (N57)? data_i[862] : 
                       (N59)? data_i[990] : 1'b0;
  assign data_o[477] = (N52)? data_i[93] : 
                       (N54)? data_i[221] : 
                       (N56)? data_i[349] : 
                       (N58)? data_i[477] : 
                       (N53)? data_i[605] : 
                       (N55)? data_i[733] : 
                       (N57)? data_i[861] : 
                       (N59)? data_i[989] : 1'b0;
  assign data_o[476] = (N52)? data_i[92] : 
                       (N54)? data_i[220] : 
                       (N56)? data_i[348] : 
                       (N58)? data_i[476] : 
                       (N53)? data_i[604] : 
                       (N55)? data_i[732] : 
                       (N57)? data_i[860] : 
                       (N59)? data_i[988] : 1'b0;
  assign data_o[475] = (N52)? data_i[91] : 
                       (N54)? data_i[219] : 
                       (N56)? data_i[347] : 
                       (N58)? data_i[475] : 
                       (N53)? data_i[603] : 
                       (N55)? data_i[731] : 
                       (N57)? data_i[859] : 
                       (N59)? data_i[987] : 1'b0;
  assign data_o[474] = (N52)? data_i[90] : 
                       (N54)? data_i[218] : 
                       (N56)? data_i[346] : 
                       (N58)? data_i[474] : 
                       (N53)? data_i[602] : 
                       (N55)? data_i[730] : 
                       (N57)? data_i[858] : 
                       (N59)? data_i[986] : 1'b0;
  assign data_o[473] = (N52)? data_i[89] : 
                       (N54)? data_i[217] : 
                       (N56)? data_i[345] : 
                       (N58)? data_i[473] : 
                       (N53)? data_i[601] : 
                       (N55)? data_i[729] : 
                       (N57)? data_i[857] : 
                       (N59)? data_i[985] : 1'b0;
  assign data_o[472] = (N52)? data_i[88] : 
                       (N54)? data_i[216] : 
                       (N56)? data_i[344] : 
                       (N58)? data_i[472] : 
                       (N53)? data_i[600] : 
                       (N55)? data_i[728] : 
                       (N57)? data_i[856] : 
                       (N59)? data_i[984] : 1'b0;
  assign data_o[471] = (N52)? data_i[87] : 
                       (N54)? data_i[215] : 
                       (N56)? data_i[343] : 
                       (N58)? data_i[471] : 
                       (N53)? data_i[599] : 
                       (N55)? data_i[727] : 
                       (N57)? data_i[855] : 
                       (N59)? data_i[983] : 1'b0;
  assign data_o[470] = (N52)? data_i[86] : 
                       (N54)? data_i[214] : 
                       (N56)? data_i[342] : 
                       (N58)? data_i[470] : 
                       (N53)? data_i[598] : 
                       (N55)? data_i[726] : 
                       (N57)? data_i[854] : 
                       (N59)? data_i[982] : 1'b0;
  assign data_o[469] = (N52)? data_i[85] : 
                       (N54)? data_i[213] : 
                       (N56)? data_i[341] : 
                       (N58)? data_i[469] : 
                       (N53)? data_i[597] : 
                       (N55)? data_i[725] : 
                       (N57)? data_i[853] : 
                       (N59)? data_i[981] : 1'b0;
  assign data_o[468] = (N52)? data_i[84] : 
                       (N54)? data_i[212] : 
                       (N56)? data_i[340] : 
                       (N58)? data_i[468] : 
                       (N53)? data_i[596] : 
                       (N55)? data_i[724] : 
                       (N57)? data_i[852] : 
                       (N59)? data_i[980] : 1'b0;
  assign data_o[467] = (N52)? data_i[83] : 
                       (N54)? data_i[211] : 
                       (N56)? data_i[339] : 
                       (N58)? data_i[467] : 
                       (N53)? data_i[595] : 
                       (N55)? data_i[723] : 
                       (N57)? data_i[851] : 
                       (N59)? data_i[979] : 1'b0;
  assign data_o[466] = (N52)? data_i[82] : 
                       (N54)? data_i[210] : 
                       (N56)? data_i[338] : 
                       (N58)? data_i[466] : 
                       (N53)? data_i[594] : 
                       (N55)? data_i[722] : 
                       (N57)? data_i[850] : 
                       (N59)? data_i[978] : 1'b0;
  assign data_o[465] = (N52)? data_i[81] : 
                       (N54)? data_i[209] : 
                       (N56)? data_i[337] : 
                       (N58)? data_i[465] : 
                       (N53)? data_i[593] : 
                       (N55)? data_i[721] : 
                       (N57)? data_i[849] : 
                       (N59)? data_i[977] : 1'b0;
  assign data_o[464] = (N52)? data_i[80] : 
                       (N54)? data_i[208] : 
                       (N56)? data_i[336] : 
                       (N58)? data_i[464] : 
                       (N53)? data_i[592] : 
                       (N55)? data_i[720] : 
                       (N57)? data_i[848] : 
                       (N59)? data_i[976] : 1'b0;
  assign data_o[463] = (N52)? data_i[79] : 
                       (N54)? data_i[207] : 
                       (N56)? data_i[335] : 
                       (N58)? data_i[463] : 
                       (N53)? data_i[591] : 
                       (N55)? data_i[719] : 
                       (N57)? data_i[847] : 
                       (N59)? data_i[975] : 1'b0;
  assign data_o[462] = (N52)? data_i[78] : 
                       (N54)? data_i[206] : 
                       (N56)? data_i[334] : 
                       (N58)? data_i[462] : 
                       (N53)? data_i[590] : 
                       (N55)? data_i[718] : 
                       (N57)? data_i[846] : 
                       (N59)? data_i[974] : 1'b0;
  assign data_o[461] = (N52)? data_i[77] : 
                       (N54)? data_i[205] : 
                       (N56)? data_i[333] : 
                       (N58)? data_i[461] : 
                       (N53)? data_i[589] : 
                       (N55)? data_i[717] : 
                       (N57)? data_i[845] : 
                       (N59)? data_i[973] : 1'b0;
  assign data_o[460] = (N52)? data_i[76] : 
                       (N54)? data_i[204] : 
                       (N56)? data_i[332] : 
                       (N58)? data_i[460] : 
                       (N53)? data_i[588] : 
                       (N55)? data_i[716] : 
                       (N57)? data_i[844] : 
                       (N59)? data_i[972] : 1'b0;
  assign data_o[459] = (N52)? data_i[75] : 
                       (N54)? data_i[203] : 
                       (N56)? data_i[331] : 
                       (N58)? data_i[459] : 
                       (N53)? data_i[587] : 
                       (N55)? data_i[715] : 
                       (N57)? data_i[843] : 
                       (N59)? data_i[971] : 1'b0;
  assign data_o[458] = (N52)? data_i[74] : 
                       (N54)? data_i[202] : 
                       (N56)? data_i[330] : 
                       (N58)? data_i[458] : 
                       (N53)? data_i[586] : 
                       (N55)? data_i[714] : 
                       (N57)? data_i[842] : 
                       (N59)? data_i[970] : 1'b0;
  assign data_o[457] = (N52)? data_i[73] : 
                       (N54)? data_i[201] : 
                       (N56)? data_i[329] : 
                       (N58)? data_i[457] : 
                       (N53)? data_i[585] : 
                       (N55)? data_i[713] : 
                       (N57)? data_i[841] : 
                       (N59)? data_i[969] : 1'b0;
  assign data_o[456] = (N52)? data_i[72] : 
                       (N54)? data_i[200] : 
                       (N56)? data_i[328] : 
                       (N58)? data_i[456] : 
                       (N53)? data_i[584] : 
                       (N55)? data_i[712] : 
                       (N57)? data_i[840] : 
                       (N59)? data_i[968] : 1'b0;
  assign data_o[455] = (N52)? data_i[71] : 
                       (N54)? data_i[199] : 
                       (N56)? data_i[327] : 
                       (N58)? data_i[455] : 
                       (N53)? data_i[583] : 
                       (N55)? data_i[711] : 
                       (N57)? data_i[839] : 
                       (N59)? data_i[967] : 1'b0;
  assign data_o[454] = (N52)? data_i[70] : 
                       (N54)? data_i[198] : 
                       (N56)? data_i[326] : 
                       (N58)? data_i[454] : 
                       (N53)? data_i[582] : 
                       (N55)? data_i[710] : 
                       (N57)? data_i[838] : 
                       (N59)? data_i[966] : 1'b0;
  assign data_o[453] = (N52)? data_i[69] : 
                       (N54)? data_i[197] : 
                       (N56)? data_i[325] : 
                       (N58)? data_i[453] : 
                       (N53)? data_i[581] : 
                       (N55)? data_i[709] : 
                       (N57)? data_i[837] : 
                       (N59)? data_i[965] : 1'b0;
  assign data_o[452] = (N52)? data_i[68] : 
                       (N54)? data_i[196] : 
                       (N56)? data_i[324] : 
                       (N58)? data_i[452] : 
                       (N53)? data_i[580] : 
                       (N55)? data_i[708] : 
                       (N57)? data_i[836] : 
                       (N59)? data_i[964] : 1'b0;
  assign data_o[451] = (N52)? data_i[67] : 
                       (N54)? data_i[195] : 
                       (N56)? data_i[323] : 
                       (N58)? data_i[451] : 
                       (N53)? data_i[579] : 
                       (N55)? data_i[707] : 
                       (N57)? data_i[835] : 
                       (N59)? data_i[963] : 1'b0;
  assign data_o[450] = (N52)? data_i[66] : 
                       (N54)? data_i[194] : 
                       (N56)? data_i[322] : 
                       (N58)? data_i[450] : 
                       (N53)? data_i[578] : 
                       (N55)? data_i[706] : 
                       (N57)? data_i[834] : 
                       (N59)? data_i[962] : 1'b0;
  assign data_o[449] = (N52)? data_i[65] : 
                       (N54)? data_i[193] : 
                       (N56)? data_i[321] : 
                       (N58)? data_i[449] : 
                       (N53)? data_i[577] : 
                       (N55)? data_i[705] : 
                       (N57)? data_i[833] : 
                       (N59)? data_i[961] : 1'b0;
  assign data_o[448] = (N52)? data_i[64] : 
                       (N54)? data_i[192] : 
                       (N56)? data_i[320] : 
                       (N58)? data_i[448] : 
                       (N53)? data_i[576] : 
                       (N55)? data_i[704] : 
                       (N57)? data_i[832] : 
                       (N59)? data_i[960] : 1'b0;
  assign data_o[447] = (N52)? data_i[63] : 
                       (N54)? data_i[191] : 
                       (N56)? data_i[319] : 
                       (N58)? data_i[447] : 
                       (N53)? data_i[575] : 
                       (N55)? data_i[703] : 
                       (N57)? data_i[831] : 
                       (N59)? data_i[959] : 1'b0;
  assign data_o[446] = (N52)? data_i[62] : 
                       (N54)? data_i[190] : 
                       (N56)? data_i[318] : 
                       (N58)? data_i[446] : 
                       (N53)? data_i[574] : 
                       (N55)? data_i[702] : 
                       (N57)? data_i[830] : 
                       (N59)? data_i[958] : 1'b0;
  assign data_o[445] = (N52)? data_i[61] : 
                       (N54)? data_i[189] : 
                       (N56)? data_i[317] : 
                       (N58)? data_i[445] : 
                       (N53)? data_i[573] : 
                       (N55)? data_i[701] : 
                       (N57)? data_i[829] : 
                       (N59)? data_i[957] : 1'b0;
  assign data_o[444] = (N52)? data_i[60] : 
                       (N54)? data_i[188] : 
                       (N56)? data_i[316] : 
                       (N58)? data_i[444] : 
                       (N53)? data_i[572] : 
                       (N55)? data_i[700] : 
                       (N57)? data_i[828] : 
                       (N59)? data_i[956] : 1'b0;
  assign data_o[443] = (N52)? data_i[59] : 
                       (N54)? data_i[187] : 
                       (N56)? data_i[315] : 
                       (N58)? data_i[443] : 
                       (N53)? data_i[571] : 
                       (N55)? data_i[699] : 
                       (N57)? data_i[827] : 
                       (N59)? data_i[955] : 1'b0;
  assign data_o[442] = (N52)? data_i[58] : 
                       (N54)? data_i[186] : 
                       (N56)? data_i[314] : 
                       (N58)? data_i[442] : 
                       (N53)? data_i[570] : 
                       (N55)? data_i[698] : 
                       (N57)? data_i[826] : 
                       (N59)? data_i[954] : 1'b0;
  assign data_o[441] = (N52)? data_i[57] : 
                       (N54)? data_i[185] : 
                       (N56)? data_i[313] : 
                       (N58)? data_i[441] : 
                       (N53)? data_i[569] : 
                       (N55)? data_i[697] : 
                       (N57)? data_i[825] : 
                       (N59)? data_i[953] : 1'b0;
  assign data_o[440] = (N52)? data_i[56] : 
                       (N54)? data_i[184] : 
                       (N56)? data_i[312] : 
                       (N58)? data_i[440] : 
                       (N53)? data_i[568] : 
                       (N55)? data_i[696] : 
                       (N57)? data_i[824] : 
                       (N59)? data_i[952] : 1'b0;
  assign data_o[439] = (N52)? data_i[55] : 
                       (N54)? data_i[183] : 
                       (N56)? data_i[311] : 
                       (N58)? data_i[439] : 
                       (N53)? data_i[567] : 
                       (N55)? data_i[695] : 
                       (N57)? data_i[823] : 
                       (N59)? data_i[951] : 1'b0;
  assign data_o[438] = (N52)? data_i[54] : 
                       (N54)? data_i[182] : 
                       (N56)? data_i[310] : 
                       (N58)? data_i[438] : 
                       (N53)? data_i[566] : 
                       (N55)? data_i[694] : 
                       (N57)? data_i[822] : 
                       (N59)? data_i[950] : 1'b0;
  assign data_o[437] = (N52)? data_i[53] : 
                       (N54)? data_i[181] : 
                       (N56)? data_i[309] : 
                       (N58)? data_i[437] : 
                       (N53)? data_i[565] : 
                       (N55)? data_i[693] : 
                       (N57)? data_i[821] : 
                       (N59)? data_i[949] : 1'b0;
  assign data_o[436] = (N52)? data_i[52] : 
                       (N54)? data_i[180] : 
                       (N56)? data_i[308] : 
                       (N58)? data_i[436] : 
                       (N53)? data_i[564] : 
                       (N55)? data_i[692] : 
                       (N57)? data_i[820] : 
                       (N59)? data_i[948] : 1'b0;
  assign data_o[435] = (N52)? data_i[51] : 
                       (N54)? data_i[179] : 
                       (N56)? data_i[307] : 
                       (N58)? data_i[435] : 
                       (N53)? data_i[563] : 
                       (N55)? data_i[691] : 
                       (N57)? data_i[819] : 
                       (N59)? data_i[947] : 1'b0;
  assign data_o[434] = (N52)? data_i[50] : 
                       (N54)? data_i[178] : 
                       (N56)? data_i[306] : 
                       (N58)? data_i[434] : 
                       (N53)? data_i[562] : 
                       (N55)? data_i[690] : 
                       (N57)? data_i[818] : 
                       (N59)? data_i[946] : 1'b0;
  assign data_o[433] = (N52)? data_i[49] : 
                       (N54)? data_i[177] : 
                       (N56)? data_i[305] : 
                       (N58)? data_i[433] : 
                       (N53)? data_i[561] : 
                       (N55)? data_i[689] : 
                       (N57)? data_i[817] : 
                       (N59)? data_i[945] : 1'b0;
  assign data_o[432] = (N52)? data_i[48] : 
                       (N54)? data_i[176] : 
                       (N56)? data_i[304] : 
                       (N58)? data_i[432] : 
                       (N53)? data_i[560] : 
                       (N55)? data_i[688] : 
                       (N57)? data_i[816] : 
                       (N59)? data_i[944] : 1'b0;
  assign data_o[431] = (N52)? data_i[47] : 
                       (N54)? data_i[175] : 
                       (N56)? data_i[303] : 
                       (N58)? data_i[431] : 
                       (N53)? data_i[559] : 
                       (N55)? data_i[687] : 
                       (N57)? data_i[815] : 
                       (N59)? data_i[943] : 1'b0;
  assign data_o[430] = (N52)? data_i[46] : 
                       (N54)? data_i[174] : 
                       (N56)? data_i[302] : 
                       (N58)? data_i[430] : 
                       (N53)? data_i[558] : 
                       (N55)? data_i[686] : 
                       (N57)? data_i[814] : 
                       (N59)? data_i[942] : 1'b0;
  assign data_o[429] = (N52)? data_i[45] : 
                       (N54)? data_i[173] : 
                       (N56)? data_i[301] : 
                       (N58)? data_i[429] : 
                       (N53)? data_i[557] : 
                       (N55)? data_i[685] : 
                       (N57)? data_i[813] : 
                       (N59)? data_i[941] : 1'b0;
  assign data_o[428] = (N52)? data_i[44] : 
                       (N54)? data_i[172] : 
                       (N56)? data_i[300] : 
                       (N58)? data_i[428] : 
                       (N53)? data_i[556] : 
                       (N55)? data_i[684] : 
                       (N57)? data_i[812] : 
                       (N59)? data_i[940] : 1'b0;
  assign data_o[427] = (N52)? data_i[43] : 
                       (N54)? data_i[171] : 
                       (N56)? data_i[299] : 
                       (N58)? data_i[427] : 
                       (N53)? data_i[555] : 
                       (N55)? data_i[683] : 
                       (N57)? data_i[811] : 
                       (N59)? data_i[939] : 1'b0;
  assign data_o[426] = (N52)? data_i[42] : 
                       (N54)? data_i[170] : 
                       (N56)? data_i[298] : 
                       (N58)? data_i[426] : 
                       (N53)? data_i[554] : 
                       (N55)? data_i[682] : 
                       (N57)? data_i[810] : 
                       (N59)? data_i[938] : 1'b0;
  assign data_o[425] = (N52)? data_i[41] : 
                       (N54)? data_i[169] : 
                       (N56)? data_i[297] : 
                       (N58)? data_i[425] : 
                       (N53)? data_i[553] : 
                       (N55)? data_i[681] : 
                       (N57)? data_i[809] : 
                       (N59)? data_i[937] : 1'b0;
  assign data_o[424] = (N52)? data_i[40] : 
                       (N54)? data_i[168] : 
                       (N56)? data_i[296] : 
                       (N58)? data_i[424] : 
                       (N53)? data_i[552] : 
                       (N55)? data_i[680] : 
                       (N57)? data_i[808] : 
                       (N59)? data_i[936] : 1'b0;
  assign data_o[423] = (N52)? data_i[39] : 
                       (N54)? data_i[167] : 
                       (N56)? data_i[295] : 
                       (N58)? data_i[423] : 
                       (N53)? data_i[551] : 
                       (N55)? data_i[679] : 
                       (N57)? data_i[807] : 
                       (N59)? data_i[935] : 1'b0;
  assign data_o[422] = (N52)? data_i[38] : 
                       (N54)? data_i[166] : 
                       (N56)? data_i[294] : 
                       (N58)? data_i[422] : 
                       (N53)? data_i[550] : 
                       (N55)? data_i[678] : 
                       (N57)? data_i[806] : 
                       (N59)? data_i[934] : 1'b0;
  assign data_o[421] = (N52)? data_i[37] : 
                       (N54)? data_i[165] : 
                       (N56)? data_i[293] : 
                       (N58)? data_i[421] : 
                       (N53)? data_i[549] : 
                       (N55)? data_i[677] : 
                       (N57)? data_i[805] : 
                       (N59)? data_i[933] : 1'b0;
  assign data_o[420] = (N52)? data_i[36] : 
                       (N54)? data_i[164] : 
                       (N56)? data_i[292] : 
                       (N58)? data_i[420] : 
                       (N53)? data_i[548] : 
                       (N55)? data_i[676] : 
                       (N57)? data_i[804] : 
                       (N59)? data_i[932] : 1'b0;
  assign data_o[419] = (N52)? data_i[35] : 
                       (N54)? data_i[163] : 
                       (N56)? data_i[291] : 
                       (N58)? data_i[419] : 
                       (N53)? data_i[547] : 
                       (N55)? data_i[675] : 
                       (N57)? data_i[803] : 
                       (N59)? data_i[931] : 1'b0;
  assign data_o[418] = (N52)? data_i[34] : 
                       (N54)? data_i[162] : 
                       (N56)? data_i[290] : 
                       (N58)? data_i[418] : 
                       (N53)? data_i[546] : 
                       (N55)? data_i[674] : 
                       (N57)? data_i[802] : 
                       (N59)? data_i[930] : 1'b0;
  assign data_o[417] = (N52)? data_i[33] : 
                       (N54)? data_i[161] : 
                       (N56)? data_i[289] : 
                       (N58)? data_i[417] : 
                       (N53)? data_i[545] : 
                       (N55)? data_i[673] : 
                       (N57)? data_i[801] : 
                       (N59)? data_i[929] : 1'b0;
  assign data_o[416] = (N52)? data_i[32] : 
                       (N54)? data_i[160] : 
                       (N56)? data_i[288] : 
                       (N58)? data_i[416] : 
                       (N53)? data_i[544] : 
                       (N55)? data_i[672] : 
                       (N57)? data_i[800] : 
                       (N59)? data_i[928] : 1'b0;
  assign data_o[415] = (N52)? data_i[31] : 
                       (N54)? data_i[159] : 
                       (N56)? data_i[287] : 
                       (N58)? data_i[415] : 
                       (N53)? data_i[543] : 
                       (N55)? data_i[671] : 
                       (N57)? data_i[799] : 
                       (N59)? data_i[927] : 1'b0;
  assign data_o[414] = (N52)? data_i[30] : 
                       (N54)? data_i[158] : 
                       (N56)? data_i[286] : 
                       (N58)? data_i[414] : 
                       (N53)? data_i[542] : 
                       (N55)? data_i[670] : 
                       (N57)? data_i[798] : 
                       (N59)? data_i[926] : 1'b0;
  assign data_o[413] = (N52)? data_i[29] : 
                       (N54)? data_i[157] : 
                       (N56)? data_i[285] : 
                       (N58)? data_i[413] : 
                       (N53)? data_i[541] : 
                       (N55)? data_i[669] : 
                       (N57)? data_i[797] : 
                       (N59)? data_i[925] : 1'b0;
  assign data_o[412] = (N52)? data_i[28] : 
                       (N54)? data_i[156] : 
                       (N56)? data_i[284] : 
                       (N58)? data_i[412] : 
                       (N53)? data_i[540] : 
                       (N55)? data_i[668] : 
                       (N57)? data_i[796] : 
                       (N59)? data_i[924] : 1'b0;
  assign data_o[411] = (N52)? data_i[27] : 
                       (N54)? data_i[155] : 
                       (N56)? data_i[283] : 
                       (N58)? data_i[411] : 
                       (N53)? data_i[539] : 
                       (N55)? data_i[667] : 
                       (N57)? data_i[795] : 
                       (N59)? data_i[923] : 1'b0;
  assign data_o[410] = (N52)? data_i[26] : 
                       (N54)? data_i[154] : 
                       (N56)? data_i[282] : 
                       (N58)? data_i[410] : 
                       (N53)? data_i[538] : 
                       (N55)? data_i[666] : 
                       (N57)? data_i[794] : 
                       (N59)? data_i[922] : 1'b0;
  assign data_o[409] = (N52)? data_i[25] : 
                       (N54)? data_i[153] : 
                       (N56)? data_i[281] : 
                       (N58)? data_i[409] : 
                       (N53)? data_i[537] : 
                       (N55)? data_i[665] : 
                       (N57)? data_i[793] : 
                       (N59)? data_i[921] : 1'b0;
  assign data_o[408] = (N52)? data_i[24] : 
                       (N54)? data_i[152] : 
                       (N56)? data_i[280] : 
                       (N58)? data_i[408] : 
                       (N53)? data_i[536] : 
                       (N55)? data_i[664] : 
                       (N57)? data_i[792] : 
                       (N59)? data_i[920] : 1'b0;
  assign data_o[407] = (N52)? data_i[23] : 
                       (N54)? data_i[151] : 
                       (N56)? data_i[279] : 
                       (N58)? data_i[407] : 
                       (N53)? data_i[535] : 
                       (N55)? data_i[663] : 
                       (N57)? data_i[791] : 
                       (N59)? data_i[919] : 1'b0;
  assign data_o[406] = (N52)? data_i[22] : 
                       (N54)? data_i[150] : 
                       (N56)? data_i[278] : 
                       (N58)? data_i[406] : 
                       (N53)? data_i[534] : 
                       (N55)? data_i[662] : 
                       (N57)? data_i[790] : 
                       (N59)? data_i[918] : 1'b0;
  assign data_o[405] = (N52)? data_i[21] : 
                       (N54)? data_i[149] : 
                       (N56)? data_i[277] : 
                       (N58)? data_i[405] : 
                       (N53)? data_i[533] : 
                       (N55)? data_i[661] : 
                       (N57)? data_i[789] : 
                       (N59)? data_i[917] : 1'b0;
  assign data_o[404] = (N52)? data_i[20] : 
                       (N54)? data_i[148] : 
                       (N56)? data_i[276] : 
                       (N58)? data_i[404] : 
                       (N53)? data_i[532] : 
                       (N55)? data_i[660] : 
                       (N57)? data_i[788] : 
                       (N59)? data_i[916] : 1'b0;
  assign data_o[403] = (N52)? data_i[19] : 
                       (N54)? data_i[147] : 
                       (N56)? data_i[275] : 
                       (N58)? data_i[403] : 
                       (N53)? data_i[531] : 
                       (N55)? data_i[659] : 
                       (N57)? data_i[787] : 
                       (N59)? data_i[915] : 1'b0;
  assign data_o[402] = (N52)? data_i[18] : 
                       (N54)? data_i[146] : 
                       (N56)? data_i[274] : 
                       (N58)? data_i[402] : 
                       (N53)? data_i[530] : 
                       (N55)? data_i[658] : 
                       (N57)? data_i[786] : 
                       (N59)? data_i[914] : 1'b0;
  assign data_o[401] = (N52)? data_i[17] : 
                       (N54)? data_i[145] : 
                       (N56)? data_i[273] : 
                       (N58)? data_i[401] : 
                       (N53)? data_i[529] : 
                       (N55)? data_i[657] : 
                       (N57)? data_i[785] : 
                       (N59)? data_i[913] : 1'b0;
  assign data_o[400] = (N52)? data_i[16] : 
                       (N54)? data_i[144] : 
                       (N56)? data_i[272] : 
                       (N58)? data_i[400] : 
                       (N53)? data_i[528] : 
                       (N55)? data_i[656] : 
                       (N57)? data_i[784] : 
                       (N59)? data_i[912] : 1'b0;
  assign data_o[399] = (N52)? data_i[15] : 
                       (N54)? data_i[143] : 
                       (N56)? data_i[271] : 
                       (N58)? data_i[399] : 
                       (N53)? data_i[527] : 
                       (N55)? data_i[655] : 
                       (N57)? data_i[783] : 
                       (N59)? data_i[911] : 1'b0;
  assign data_o[398] = (N52)? data_i[14] : 
                       (N54)? data_i[142] : 
                       (N56)? data_i[270] : 
                       (N58)? data_i[398] : 
                       (N53)? data_i[526] : 
                       (N55)? data_i[654] : 
                       (N57)? data_i[782] : 
                       (N59)? data_i[910] : 1'b0;
  assign data_o[397] = (N52)? data_i[13] : 
                       (N54)? data_i[141] : 
                       (N56)? data_i[269] : 
                       (N58)? data_i[397] : 
                       (N53)? data_i[525] : 
                       (N55)? data_i[653] : 
                       (N57)? data_i[781] : 
                       (N59)? data_i[909] : 1'b0;
  assign data_o[396] = (N52)? data_i[12] : 
                       (N54)? data_i[140] : 
                       (N56)? data_i[268] : 
                       (N58)? data_i[396] : 
                       (N53)? data_i[524] : 
                       (N55)? data_i[652] : 
                       (N57)? data_i[780] : 
                       (N59)? data_i[908] : 1'b0;
  assign data_o[395] = (N52)? data_i[11] : 
                       (N54)? data_i[139] : 
                       (N56)? data_i[267] : 
                       (N58)? data_i[395] : 
                       (N53)? data_i[523] : 
                       (N55)? data_i[651] : 
                       (N57)? data_i[779] : 
                       (N59)? data_i[907] : 1'b0;
  assign data_o[394] = (N52)? data_i[10] : 
                       (N54)? data_i[138] : 
                       (N56)? data_i[266] : 
                       (N58)? data_i[394] : 
                       (N53)? data_i[522] : 
                       (N55)? data_i[650] : 
                       (N57)? data_i[778] : 
                       (N59)? data_i[906] : 1'b0;
  assign data_o[393] = (N52)? data_i[9] : 
                       (N54)? data_i[137] : 
                       (N56)? data_i[265] : 
                       (N58)? data_i[393] : 
                       (N53)? data_i[521] : 
                       (N55)? data_i[649] : 
                       (N57)? data_i[777] : 
                       (N59)? data_i[905] : 1'b0;
  assign data_o[392] = (N52)? data_i[8] : 
                       (N54)? data_i[136] : 
                       (N56)? data_i[264] : 
                       (N58)? data_i[392] : 
                       (N53)? data_i[520] : 
                       (N55)? data_i[648] : 
                       (N57)? data_i[776] : 
                       (N59)? data_i[904] : 1'b0;
  assign data_o[391] = (N52)? data_i[7] : 
                       (N54)? data_i[135] : 
                       (N56)? data_i[263] : 
                       (N58)? data_i[391] : 
                       (N53)? data_i[519] : 
                       (N55)? data_i[647] : 
                       (N57)? data_i[775] : 
                       (N59)? data_i[903] : 1'b0;
  assign data_o[390] = (N52)? data_i[6] : 
                       (N54)? data_i[134] : 
                       (N56)? data_i[262] : 
                       (N58)? data_i[390] : 
                       (N53)? data_i[518] : 
                       (N55)? data_i[646] : 
                       (N57)? data_i[774] : 
                       (N59)? data_i[902] : 1'b0;
  assign data_o[389] = (N52)? data_i[5] : 
                       (N54)? data_i[133] : 
                       (N56)? data_i[261] : 
                       (N58)? data_i[389] : 
                       (N53)? data_i[517] : 
                       (N55)? data_i[645] : 
                       (N57)? data_i[773] : 
                       (N59)? data_i[901] : 1'b0;
  assign data_o[388] = (N52)? data_i[4] : 
                       (N54)? data_i[132] : 
                       (N56)? data_i[260] : 
                       (N58)? data_i[388] : 
                       (N53)? data_i[516] : 
                       (N55)? data_i[644] : 
                       (N57)? data_i[772] : 
                       (N59)? data_i[900] : 1'b0;
  assign data_o[387] = (N52)? data_i[3] : 
                       (N54)? data_i[131] : 
                       (N56)? data_i[259] : 
                       (N58)? data_i[387] : 
                       (N53)? data_i[515] : 
                       (N55)? data_i[643] : 
                       (N57)? data_i[771] : 
                       (N59)? data_i[899] : 1'b0;
  assign data_o[386] = (N52)? data_i[2] : 
                       (N54)? data_i[130] : 
                       (N56)? data_i[258] : 
                       (N58)? data_i[386] : 
                       (N53)? data_i[514] : 
                       (N55)? data_i[642] : 
                       (N57)? data_i[770] : 
                       (N59)? data_i[898] : 1'b0;
  assign data_o[385] = (N52)? data_i[1] : 
                       (N54)? data_i[129] : 
                       (N56)? data_i[257] : 
                       (N58)? data_i[385] : 
                       (N53)? data_i[513] : 
                       (N55)? data_i[641] : 
                       (N57)? data_i[769] : 
                       (N59)? data_i[897] : 1'b0;
  assign data_o[384] = (N52)? data_i[0] : 
                       (N54)? data_i[128] : 
                       (N56)? data_i[256] : 
                       (N58)? data_i[384] : 
                       (N53)? data_i[512] : 
                       (N55)? data_i[640] : 
                       (N57)? data_i[768] : 
                       (N59)? data_i[896] : 1'b0;
  assign data_o[639] = (N67)? data_i[127] : 
                       (N69)? data_i[255] : 
                       (N71)? data_i[383] : 
                       (N73)? data_i[511] : 
                       (N68)? data_i[639] : 
                       (N70)? data_i[767] : 
                       (N72)? data_i[895] : 
                       (N74)? data_i[1023] : 1'b0;
  assign data_o[638] = (N67)? data_i[126] : 
                       (N69)? data_i[254] : 
                       (N71)? data_i[382] : 
                       (N73)? data_i[510] : 
                       (N68)? data_i[638] : 
                       (N70)? data_i[766] : 
                       (N72)? data_i[894] : 
                       (N74)? data_i[1022] : 1'b0;
  assign data_o[637] = (N67)? data_i[125] : 
                       (N69)? data_i[253] : 
                       (N71)? data_i[381] : 
                       (N73)? data_i[509] : 
                       (N68)? data_i[637] : 
                       (N70)? data_i[765] : 
                       (N72)? data_i[893] : 
                       (N74)? data_i[1021] : 1'b0;
  assign data_o[636] = (N67)? data_i[124] : 
                       (N69)? data_i[252] : 
                       (N71)? data_i[380] : 
                       (N73)? data_i[508] : 
                       (N68)? data_i[636] : 
                       (N70)? data_i[764] : 
                       (N72)? data_i[892] : 
                       (N74)? data_i[1020] : 1'b0;
  assign data_o[635] = (N67)? data_i[123] : 
                       (N69)? data_i[251] : 
                       (N71)? data_i[379] : 
                       (N73)? data_i[507] : 
                       (N68)? data_i[635] : 
                       (N70)? data_i[763] : 
                       (N72)? data_i[891] : 
                       (N74)? data_i[1019] : 1'b0;
  assign data_o[634] = (N67)? data_i[122] : 
                       (N69)? data_i[250] : 
                       (N71)? data_i[378] : 
                       (N73)? data_i[506] : 
                       (N68)? data_i[634] : 
                       (N70)? data_i[762] : 
                       (N72)? data_i[890] : 
                       (N74)? data_i[1018] : 1'b0;
  assign data_o[633] = (N67)? data_i[121] : 
                       (N69)? data_i[249] : 
                       (N71)? data_i[377] : 
                       (N73)? data_i[505] : 
                       (N68)? data_i[633] : 
                       (N70)? data_i[761] : 
                       (N72)? data_i[889] : 
                       (N74)? data_i[1017] : 1'b0;
  assign data_o[632] = (N67)? data_i[120] : 
                       (N69)? data_i[248] : 
                       (N71)? data_i[376] : 
                       (N73)? data_i[504] : 
                       (N68)? data_i[632] : 
                       (N70)? data_i[760] : 
                       (N72)? data_i[888] : 
                       (N74)? data_i[1016] : 1'b0;
  assign data_o[631] = (N67)? data_i[119] : 
                       (N69)? data_i[247] : 
                       (N71)? data_i[375] : 
                       (N73)? data_i[503] : 
                       (N68)? data_i[631] : 
                       (N70)? data_i[759] : 
                       (N72)? data_i[887] : 
                       (N74)? data_i[1015] : 1'b0;
  assign data_o[630] = (N67)? data_i[118] : 
                       (N69)? data_i[246] : 
                       (N71)? data_i[374] : 
                       (N73)? data_i[502] : 
                       (N68)? data_i[630] : 
                       (N70)? data_i[758] : 
                       (N72)? data_i[886] : 
                       (N74)? data_i[1014] : 1'b0;
  assign data_o[629] = (N67)? data_i[117] : 
                       (N69)? data_i[245] : 
                       (N71)? data_i[373] : 
                       (N73)? data_i[501] : 
                       (N68)? data_i[629] : 
                       (N70)? data_i[757] : 
                       (N72)? data_i[885] : 
                       (N74)? data_i[1013] : 1'b0;
  assign data_o[628] = (N67)? data_i[116] : 
                       (N69)? data_i[244] : 
                       (N71)? data_i[372] : 
                       (N73)? data_i[500] : 
                       (N68)? data_i[628] : 
                       (N70)? data_i[756] : 
                       (N72)? data_i[884] : 
                       (N74)? data_i[1012] : 1'b0;
  assign data_o[627] = (N67)? data_i[115] : 
                       (N69)? data_i[243] : 
                       (N71)? data_i[371] : 
                       (N73)? data_i[499] : 
                       (N68)? data_i[627] : 
                       (N70)? data_i[755] : 
                       (N72)? data_i[883] : 
                       (N74)? data_i[1011] : 1'b0;
  assign data_o[626] = (N67)? data_i[114] : 
                       (N69)? data_i[242] : 
                       (N71)? data_i[370] : 
                       (N73)? data_i[498] : 
                       (N68)? data_i[626] : 
                       (N70)? data_i[754] : 
                       (N72)? data_i[882] : 
                       (N74)? data_i[1010] : 1'b0;
  assign data_o[625] = (N67)? data_i[113] : 
                       (N69)? data_i[241] : 
                       (N71)? data_i[369] : 
                       (N73)? data_i[497] : 
                       (N68)? data_i[625] : 
                       (N70)? data_i[753] : 
                       (N72)? data_i[881] : 
                       (N74)? data_i[1009] : 1'b0;
  assign data_o[624] = (N67)? data_i[112] : 
                       (N69)? data_i[240] : 
                       (N71)? data_i[368] : 
                       (N73)? data_i[496] : 
                       (N68)? data_i[624] : 
                       (N70)? data_i[752] : 
                       (N72)? data_i[880] : 
                       (N74)? data_i[1008] : 1'b0;
  assign data_o[623] = (N67)? data_i[111] : 
                       (N69)? data_i[239] : 
                       (N71)? data_i[367] : 
                       (N73)? data_i[495] : 
                       (N68)? data_i[623] : 
                       (N70)? data_i[751] : 
                       (N72)? data_i[879] : 
                       (N74)? data_i[1007] : 1'b0;
  assign data_o[622] = (N67)? data_i[110] : 
                       (N69)? data_i[238] : 
                       (N71)? data_i[366] : 
                       (N73)? data_i[494] : 
                       (N68)? data_i[622] : 
                       (N70)? data_i[750] : 
                       (N72)? data_i[878] : 
                       (N74)? data_i[1006] : 1'b0;
  assign data_o[621] = (N67)? data_i[109] : 
                       (N69)? data_i[237] : 
                       (N71)? data_i[365] : 
                       (N73)? data_i[493] : 
                       (N68)? data_i[621] : 
                       (N70)? data_i[749] : 
                       (N72)? data_i[877] : 
                       (N74)? data_i[1005] : 1'b0;
  assign data_o[620] = (N67)? data_i[108] : 
                       (N69)? data_i[236] : 
                       (N71)? data_i[364] : 
                       (N73)? data_i[492] : 
                       (N68)? data_i[620] : 
                       (N70)? data_i[748] : 
                       (N72)? data_i[876] : 
                       (N74)? data_i[1004] : 1'b0;
  assign data_o[619] = (N67)? data_i[107] : 
                       (N69)? data_i[235] : 
                       (N71)? data_i[363] : 
                       (N73)? data_i[491] : 
                       (N68)? data_i[619] : 
                       (N70)? data_i[747] : 
                       (N72)? data_i[875] : 
                       (N74)? data_i[1003] : 1'b0;
  assign data_o[618] = (N67)? data_i[106] : 
                       (N69)? data_i[234] : 
                       (N71)? data_i[362] : 
                       (N73)? data_i[490] : 
                       (N68)? data_i[618] : 
                       (N70)? data_i[746] : 
                       (N72)? data_i[874] : 
                       (N74)? data_i[1002] : 1'b0;
  assign data_o[617] = (N67)? data_i[105] : 
                       (N69)? data_i[233] : 
                       (N71)? data_i[361] : 
                       (N73)? data_i[489] : 
                       (N68)? data_i[617] : 
                       (N70)? data_i[745] : 
                       (N72)? data_i[873] : 
                       (N74)? data_i[1001] : 1'b0;
  assign data_o[616] = (N67)? data_i[104] : 
                       (N69)? data_i[232] : 
                       (N71)? data_i[360] : 
                       (N73)? data_i[488] : 
                       (N68)? data_i[616] : 
                       (N70)? data_i[744] : 
                       (N72)? data_i[872] : 
                       (N74)? data_i[1000] : 1'b0;
  assign data_o[615] = (N67)? data_i[103] : 
                       (N69)? data_i[231] : 
                       (N71)? data_i[359] : 
                       (N73)? data_i[487] : 
                       (N68)? data_i[615] : 
                       (N70)? data_i[743] : 
                       (N72)? data_i[871] : 
                       (N74)? data_i[999] : 1'b0;
  assign data_o[614] = (N67)? data_i[102] : 
                       (N69)? data_i[230] : 
                       (N71)? data_i[358] : 
                       (N73)? data_i[486] : 
                       (N68)? data_i[614] : 
                       (N70)? data_i[742] : 
                       (N72)? data_i[870] : 
                       (N74)? data_i[998] : 1'b0;
  assign data_o[613] = (N67)? data_i[101] : 
                       (N69)? data_i[229] : 
                       (N71)? data_i[357] : 
                       (N73)? data_i[485] : 
                       (N68)? data_i[613] : 
                       (N70)? data_i[741] : 
                       (N72)? data_i[869] : 
                       (N74)? data_i[997] : 1'b0;
  assign data_o[612] = (N67)? data_i[100] : 
                       (N69)? data_i[228] : 
                       (N71)? data_i[356] : 
                       (N73)? data_i[484] : 
                       (N68)? data_i[612] : 
                       (N70)? data_i[740] : 
                       (N72)? data_i[868] : 
                       (N74)? data_i[996] : 1'b0;
  assign data_o[611] = (N67)? data_i[99] : 
                       (N69)? data_i[227] : 
                       (N71)? data_i[355] : 
                       (N73)? data_i[483] : 
                       (N68)? data_i[611] : 
                       (N70)? data_i[739] : 
                       (N72)? data_i[867] : 
                       (N74)? data_i[995] : 1'b0;
  assign data_o[610] = (N67)? data_i[98] : 
                       (N69)? data_i[226] : 
                       (N71)? data_i[354] : 
                       (N73)? data_i[482] : 
                       (N68)? data_i[610] : 
                       (N70)? data_i[738] : 
                       (N72)? data_i[866] : 
                       (N74)? data_i[994] : 1'b0;
  assign data_o[609] = (N67)? data_i[97] : 
                       (N69)? data_i[225] : 
                       (N71)? data_i[353] : 
                       (N73)? data_i[481] : 
                       (N68)? data_i[609] : 
                       (N70)? data_i[737] : 
                       (N72)? data_i[865] : 
                       (N74)? data_i[993] : 1'b0;
  assign data_o[608] = (N67)? data_i[96] : 
                       (N69)? data_i[224] : 
                       (N71)? data_i[352] : 
                       (N73)? data_i[480] : 
                       (N68)? data_i[608] : 
                       (N70)? data_i[736] : 
                       (N72)? data_i[864] : 
                       (N74)? data_i[992] : 1'b0;
  assign data_o[607] = (N67)? data_i[95] : 
                       (N69)? data_i[223] : 
                       (N71)? data_i[351] : 
                       (N73)? data_i[479] : 
                       (N68)? data_i[607] : 
                       (N70)? data_i[735] : 
                       (N72)? data_i[863] : 
                       (N74)? data_i[991] : 1'b0;
  assign data_o[606] = (N67)? data_i[94] : 
                       (N69)? data_i[222] : 
                       (N71)? data_i[350] : 
                       (N73)? data_i[478] : 
                       (N68)? data_i[606] : 
                       (N70)? data_i[734] : 
                       (N72)? data_i[862] : 
                       (N74)? data_i[990] : 1'b0;
  assign data_o[605] = (N67)? data_i[93] : 
                       (N69)? data_i[221] : 
                       (N71)? data_i[349] : 
                       (N73)? data_i[477] : 
                       (N68)? data_i[605] : 
                       (N70)? data_i[733] : 
                       (N72)? data_i[861] : 
                       (N74)? data_i[989] : 1'b0;
  assign data_o[604] = (N67)? data_i[92] : 
                       (N69)? data_i[220] : 
                       (N71)? data_i[348] : 
                       (N73)? data_i[476] : 
                       (N68)? data_i[604] : 
                       (N70)? data_i[732] : 
                       (N72)? data_i[860] : 
                       (N74)? data_i[988] : 1'b0;
  assign data_o[603] = (N67)? data_i[91] : 
                       (N69)? data_i[219] : 
                       (N71)? data_i[347] : 
                       (N73)? data_i[475] : 
                       (N68)? data_i[603] : 
                       (N70)? data_i[731] : 
                       (N72)? data_i[859] : 
                       (N74)? data_i[987] : 1'b0;
  assign data_o[602] = (N67)? data_i[90] : 
                       (N69)? data_i[218] : 
                       (N71)? data_i[346] : 
                       (N73)? data_i[474] : 
                       (N68)? data_i[602] : 
                       (N70)? data_i[730] : 
                       (N72)? data_i[858] : 
                       (N74)? data_i[986] : 1'b0;
  assign data_o[601] = (N67)? data_i[89] : 
                       (N69)? data_i[217] : 
                       (N71)? data_i[345] : 
                       (N73)? data_i[473] : 
                       (N68)? data_i[601] : 
                       (N70)? data_i[729] : 
                       (N72)? data_i[857] : 
                       (N74)? data_i[985] : 1'b0;
  assign data_o[600] = (N67)? data_i[88] : 
                       (N69)? data_i[216] : 
                       (N71)? data_i[344] : 
                       (N73)? data_i[472] : 
                       (N68)? data_i[600] : 
                       (N70)? data_i[728] : 
                       (N72)? data_i[856] : 
                       (N74)? data_i[984] : 1'b0;
  assign data_o[599] = (N67)? data_i[87] : 
                       (N69)? data_i[215] : 
                       (N71)? data_i[343] : 
                       (N73)? data_i[471] : 
                       (N68)? data_i[599] : 
                       (N70)? data_i[727] : 
                       (N72)? data_i[855] : 
                       (N74)? data_i[983] : 1'b0;
  assign data_o[598] = (N67)? data_i[86] : 
                       (N69)? data_i[214] : 
                       (N71)? data_i[342] : 
                       (N73)? data_i[470] : 
                       (N68)? data_i[598] : 
                       (N70)? data_i[726] : 
                       (N72)? data_i[854] : 
                       (N74)? data_i[982] : 1'b0;
  assign data_o[597] = (N67)? data_i[85] : 
                       (N69)? data_i[213] : 
                       (N71)? data_i[341] : 
                       (N73)? data_i[469] : 
                       (N68)? data_i[597] : 
                       (N70)? data_i[725] : 
                       (N72)? data_i[853] : 
                       (N74)? data_i[981] : 1'b0;
  assign data_o[596] = (N67)? data_i[84] : 
                       (N69)? data_i[212] : 
                       (N71)? data_i[340] : 
                       (N73)? data_i[468] : 
                       (N68)? data_i[596] : 
                       (N70)? data_i[724] : 
                       (N72)? data_i[852] : 
                       (N74)? data_i[980] : 1'b0;
  assign data_o[595] = (N67)? data_i[83] : 
                       (N69)? data_i[211] : 
                       (N71)? data_i[339] : 
                       (N73)? data_i[467] : 
                       (N68)? data_i[595] : 
                       (N70)? data_i[723] : 
                       (N72)? data_i[851] : 
                       (N74)? data_i[979] : 1'b0;
  assign data_o[594] = (N67)? data_i[82] : 
                       (N69)? data_i[210] : 
                       (N71)? data_i[338] : 
                       (N73)? data_i[466] : 
                       (N68)? data_i[594] : 
                       (N70)? data_i[722] : 
                       (N72)? data_i[850] : 
                       (N74)? data_i[978] : 1'b0;
  assign data_o[593] = (N67)? data_i[81] : 
                       (N69)? data_i[209] : 
                       (N71)? data_i[337] : 
                       (N73)? data_i[465] : 
                       (N68)? data_i[593] : 
                       (N70)? data_i[721] : 
                       (N72)? data_i[849] : 
                       (N74)? data_i[977] : 1'b0;
  assign data_o[592] = (N67)? data_i[80] : 
                       (N69)? data_i[208] : 
                       (N71)? data_i[336] : 
                       (N73)? data_i[464] : 
                       (N68)? data_i[592] : 
                       (N70)? data_i[720] : 
                       (N72)? data_i[848] : 
                       (N74)? data_i[976] : 1'b0;
  assign data_o[591] = (N67)? data_i[79] : 
                       (N69)? data_i[207] : 
                       (N71)? data_i[335] : 
                       (N73)? data_i[463] : 
                       (N68)? data_i[591] : 
                       (N70)? data_i[719] : 
                       (N72)? data_i[847] : 
                       (N74)? data_i[975] : 1'b0;
  assign data_o[590] = (N67)? data_i[78] : 
                       (N69)? data_i[206] : 
                       (N71)? data_i[334] : 
                       (N73)? data_i[462] : 
                       (N68)? data_i[590] : 
                       (N70)? data_i[718] : 
                       (N72)? data_i[846] : 
                       (N74)? data_i[974] : 1'b0;
  assign data_o[589] = (N67)? data_i[77] : 
                       (N69)? data_i[205] : 
                       (N71)? data_i[333] : 
                       (N73)? data_i[461] : 
                       (N68)? data_i[589] : 
                       (N70)? data_i[717] : 
                       (N72)? data_i[845] : 
                       (N74)? data_i[973] : 1'b0;
  assign data_o[588] = (N67)? data_i[76] : 
                       (N69)? data_i[204] : 
                       (N71)? data_i[332] : 
                       (N73)? data_i[460] : 
                       (N68)? data_i[588] : 
                       (N70)? data_i[716] : 
                       (N72)? data_i[844] : 
                       (N74)? data_i[972] : 1'b0;
  assign data_o[587] = (N67)? data_i[75] : 
                       (N69)? data_i[203] : 
                       (N71)? data_i[331] : 
                       (N73)? data_i[459] : 
                       (N68)? data_i[587] : 
                       (N70)? data_i[715] : 
                       (N72)? data_i[843] : 
                       (N74)? data_i[971] : 1'b0;
  assign data_o[586] = (N67)? data_i[74] : 
                       (N69)? data_i[202] : 
                       (N71)? data_i[330] : 
                       (N73)? data_i[458] : 
                       (N68)? data_i[586] : 
                       (N70)? data_i[714] : 
                       (N72)? data_i[842] : 
                       (N74)? data_i[970] : 1'b0;
  assign data_o[585] = (N67)? data_i[73] : 
                       (N69)? data_i[201] : 
                       (N71)? data_i[329] : 
                       (N73)? data_i[457] : 
                       (N68)? data_i[585] : 
                       (N70)? data_i[713] : 
                       (N72)? data_i[841] : 
                       (N74)? data_i[969] : 1'b0;
  assign data_o[584] = (N67)? data_i[72] : 
                       (N69)? data_i[200] : 
                       (N71)? data_i[328] : 
                       (N73)? data_i[456] : 
                       (N68)? data_i[584] : 
                       (N70)? data_i[712] : 
                       (N72)? data_i[840] : 
                       (N74)? data_i[968] : 1'b0;
  assign data_o[583] = (N67)? data_i[71] : 
                       (N69)? data_i[199] : 
                       (N71)? data_i[327] : 
                       (N73)? data_i[455] : 
                       (N68)? data_i[583] : 
                       (N70)? data_i[711] : 
                       (N72)? data_i[839] : 
                       (N74)? data_i[967] : 1'b0;
  assign data_o[582] = (N67)? data_i[70] : 
                       (N69)? data_i[198] : 
                       (N71)? data_i[326] : 
                       (N73)? data_i[454] : 
                       (N68)? data_i[582] : 
                       (N70)? data_i[710] : 
                       (N72)? data_i[838] : 
                       (N74)? data_i[966] : 1'b0;
  assign data_o[581] = (N67)? data_i[69] : 
                       (N69)? data_i[197] : 
                       (N71)? data_i[325] : 
                       (N73)? data_i[453] : 
                       (N68)? data_i[581] : 
                       (N70)? data_i[709] : 
                       (N72)? data_i[837] : 
                       (N74)? data_i[965] : 1'b0;
  assign data_o[580] = (N67)? data_i[68] : 
                       (N69)? data_i[196] : 
                       (N71)? data_i[324] : 
                       (N73)? data_i[452] : 
                       (N68)? data_i[580] : 
                       (N70)? data_i[708] : 
                       (N72)? data_i[836] : 
                       (N74)? data_i[964] : 1'b0;
  assign data_o[579] = (N67)? data_i[67] : 
                       (N69)? data_i[195] : 
                       (N71)? data_i[323] : 
                       (N73)? data_i[451] : 
                       (N68)? data_i[579] : 
                       (N70)? data_i[707] : 
                       (N72)? data_i[835] : 
                       (N74)? data_i[963] : 1'b0;
  assign data_o[578] = (N67)? data_i[66] : 
                       (N69)? data_i[194] : 
                       (N71)? data_i[322] : 
                       (N73)? data_i[450] : 
                       (N68)? data_i[578] : 
                       (N70)? data_i[706] : 
                       (N72)? data_i[834] : 
                       (N74)? data_i[962] : 1'b0;
  assign data_o[577] = (N67)? data_i[65] : 
                       (N69)? data_i[193] : 
                       (N71)? data_i[321] : 
                       (N73)? data_i[449] : 
                       (N68)? data_i[577] : 
                       (N70)? data_i[705] : 
                       (N72)? data_i[833] : 
                       (N74)? data_i[961] : 1'b0;
  assign data_o[576] = (N67)? data_i[64] : 
                       (N69)? data_i[192] : 
                       (N71)? data_i[320] : 
                       (N73)? data_i[448] : 
                       (N68)? data_i[576] : 
                       (N70)? data_i[704] : 
                       (N72)? data_i[832] : 
                       (N74)? data_i[960] : 1'b0;
  assign data_o[575] = (N67)? data_i[63] : 
                       (N69)? data_i[191] : 
                       (N71)? data_i[319] : 
                       (N73)? data_i[447] : 
                       (N68)? data_i[575] : 
                       (N70)? data_i[703] : 
                       (N72)? data_i[831] : 
                       (N74)? data_i[959] : 1'b0;
  assign data_o[574] = (N67)? data_i[62] : 
                       (N69)? data_i[190] : 
                       (N71)? data_i[318] : 
                       (N73)? data_i[446] : 
                       (N68)? data_i[574] : 
                       (N70)? data_i[702] : 
                       (N72)? data_i[830] : 
                       (N74)? data_i[958] : 1'b0;
  assign data_o[573] = (N67)? data_i[61] : 
                       (N69)? data_i[189] : 
                       (N71)? data_i[317] : 
                       (N73)? data_i[445] : 
                       (N68)? data_i[573] : 
                       (N70)? data_i[701] : 
                       (N72)? data_i[829] : 
                       (N74)? data_i[957] : 1'b0;
  assign data_o[572] = (N67)? data_i[60] : 
                       (N69)? data_i[188] : 
                       (N71)? data_i[316] : 
                       (N73)? data_i[444] : 
                       (N68)? data_i[572] : 
                       (N70)? data_i[700] : 
                       (N72)? data_i[828] : 
                       (N74)? data_i[956] : 1'b0;
  assign data_o[571] = (N67)? data_i[59] : 
                       (N69)? data_i[187] : 
                       (N71)? data_i[315] : 
                       (N73)? data_i[443] : 
                       (N68)? data_i[571] : 
                       (N70)? data_i[699] : 
                       (N72)? data_i[827] : 
                       (N74)? data_i[955] : 1'b0;
  assign data_o[570] = (N67)? data_i[58] : 
                       (N69)? data_i[186] : 
                       (N71)? data_i[314] : 
                       (N73)? data_i[442] : 
                       (N68)? data_i[570] : 
                       (N70)? data_i[698] : 
                       (N72)? data_i[826] : 
                       (N74)? data_i[954] : 1'b0;
  assign data_o[569] = (N67)? data_i[57] : 
                       (N69)? data_i[185] : 
                       (N71)? data_i[313] : 
                       (N73)? data_i[441] : 
                       (N68)? data_i[569] : 
                       (N70)? data_i[697] : 
                       (N72)? data_i[825] : 
                       (N74)? data_i[953] : 1'b0;
  assign data_o[568] = (N67)? data_i[56] : 
                       (N69)? data_i[184] : 
                       (N71)? data_i[312] : 
                       (N73)? data_i[440] : 
                       (N68)? data_i[568] : 
                       (N70)? data_i[696] : 
                       (N72)? data_i[824] : 
                       (N74)? data_i[952] : 1'b0;
  assign data_o[567] = (N67)? data_i[55] : 
                       (N69)? data_i[183] : 
                       (N71)? data_i[311] : 
                       (N73)? data_i[439] : 
                       (N68)? data_i[567] : 
                       (N70)? data_i[695] : 
                       (N72)? data_i[823] : 
                       (N74)? data_i[951] : 1'b0;
  assign data_o[566] = (N67)? data_i[54] : 
                       (N69)? data_i[182] : 
                       (N71)? data_i[310] : 
                       (N73)? data_i[438] : 
                       (N68)? data_i[566] : 
                       (N70)? data_i[694] : 
                       (N72)? data_i[822] : 
                       (N74)? data_i[950] : 1'b0;
  assign data_o[565] = (N67)? data_i[53] : 
                       (N69)? data_i[181] : 
                       (N71)? data_i[309] : 
                       (N73)? data_i[437] : 
                       (N68)? data_i[565] : 
                       (N70)? data_i[693] : 
                       (N72)? data_i[821] : 
                       (N74)? data_i[949] : 1'b0;
  assign data_o[564] = (N67)? data_i[52] : 
                       (N69)? data_i[180] : 
                       (N71)? data_i[308] : 
                       (N73)? data_i[436] : 
                       (N68)? data_i[564] : 
                       (N70)? data_i[692] : 
                       (N72)? data_i[820] : 
                       (N74)? data_i[948] : 1'b0;
  assign data_o[563] = (N67)? data_i[51] : 
                       (N69)? data_i[179] : 
                       (N71)? data_i[307] : 
                       (N73)? data_i[435] : 
                       (N68)? data_i[563] : 
                       (N70)? data_i[691] : 
                       (N72)? data_i[819] : 
                       (N74)? data_i[947] : 1'b0;
  assign data_o[562] = (N67)? data_i[50] : 
                       (N69)? data_i[178] : 
                       (N71)? data_i[306] : 
                       (N73)? data_i[434] : 
                       (N68)? data_i[562] : 
                       (N70)? data_i[690] : 
                       (N72)? data_i[818] : 
                       (N74)? data_i[946] : 1'b0;
  assign data_o[561] = (N67)? data_i[49] : 
                       (N69)? data_i[177] : 
                       (N71)? data_i[305] : 
                       (N73)? data_i[433] : 
                       (N68)? data_i[561] : 
                       (N70)? data_i[689] : 
                       (N72)? data_i[817] : 
                       (N74)? data_i[945] : 1'b0;
  assign data_o[560] = (N67)? data_i[48] : 
                       (N69)? data_i[176] : 
                       (N71)? data_i[304] : 
                       (N73)? data_i[432] : 
                       (N68)? data_i[560] : 
                       (N70)? data_i[688] : 
                       (N72)? data_i[816] : 
                       (N74)? data_i[944] : 1'b0;
  assign data_o[559] = (N67)? data_i[47] : 
                       (N69)? data_i[175] : 
                       (N71)? data_i[303] : 
                       (N73)? data_i[431] : 
                       (N68)? data_i[559] : 
                       (N70)? data_i[687] : 
                       (N72)? data_i[815] : 
                       (N74)? data_i[943] : 1'b0;
  assign data_o[558] = (N67)? data_i[46] : 
                       (N69)? data_i[174] : 
                       (N71)? data_i[302] : 
                       (N73)? data_i[430] : 
                       (N68)? data_i[558] : 
                       (N70)? data_i[686] : 
                       (N72)? data_i[814] : 
                       (N74)? data_i[942] : 1'b0;
  assign data_o[557] = (N67)? data_i[45] : 
                       (N69)? data_i[173] : 
                       (N71)? data_i[301] : 
                       (N73)? data_i[429] : 
                       (N68)? data_i[557] : 
                       (N70)? data_i[685] : 
                       (N72)? data_i[813] : 
                       (N74)? data_i[941] : 1'b0;
  assign data_o[556] = (N67)? data_i[44] : 
                       (N69)? data_i[172] : 
                       (N71)? data_i[300] : 
                       (N73)? data_i[428] : 
                       (N68)? data_i[556] : 
                       (N70)? data_i[684] : 
                       (N72)? data_i[812] : 
                       (N74)? data_i[940] : 1'b0;
  assign data_o[555] = (N67)? data_i[43] : 
                       (N69)? data_i[171] : 
                       (N71)? data_i[299] : 
                       (N73)? data_i[427] : 
                       (N68)? data_i[555] : 
                       (N70)? data_i[683] : 
                       (N72)? data_i[811] : 
                       (N74)? data_i[939] : 1'b0;
  assign data_o[554] = (N67)? data_i[42] : 
                       (N69)? data_i[170] : 
                       (N71)? data_i[298] : 
                       (N73)? data_i[426] : 
                       (N68)? data_i[554] : 
                       (N70)? data_i[682] : 
                       (N72)? data_i[810] : 
                       (N74)? data_i[938] : 1'b0;
  assign data_o[553] = (N67)? data_i[41] : 
                       (N69)? data_i[169] : 
                       (N71)? data_i[297] : 
                       (N73)? data_i[425] : 
                       (N68)? data_i[553] : 
                       (N70)? data_i[681] : 
                       (N72)? data_i[809] : 
                       (N74)? data_i[937] : 1'b0;
  assign data_o[552] = (N67)? data_i[40] : 
                       (N69)? data_i[168] : 
                       (N71)? data_i[296] : 
                       (N73)? data_i[424] : 
                       (N68)? data_i[552] : 
                       (N70)? data_i[680] : 
                       (N72)? data_i[808] : 
                       (N74)? data_i[936] : 1'b0;
  assign data_o[551] = (N67)? data_i[39] : 
                       (N69)? data_i[167] : 
                       (N71)? data_i[295] : 
                       (N73)? data_i[423] : 
                       (N68)? data_i[551] : 
                       (N70)? data_i[679] : 
                       (N72)? data_i[807] : 
                       (N74)? data_i[935] : 1'b0;
  assign data_o[550] = (N67)? data_i[38] : 
                       (N69)? data_i[166] : 
                       (N71)? data_i[294] : 
                       (N73)? data_i[422] : 
                       (N68)? data_i[550] : 
                       (N70)? data_i[678] : 
                       (N72)? data_i[806] : 
                       (N74)? data_i[934] : 1'b0;
  assign data_o[549] = (N67)? data_i[37] : 
                       (N69)? data_i[165] : 
                       (N71)? data_i[293] : 
                       (N73)? data_i[421] : 
                       (N68)? data_i[549] : 
                       (N70)? data_i[677] : 
                       (N72)? data_i[805] : 
                       (N74)? data_i[933] : 1'b0;
  assign data_o[548] = (N67)? data_i[36] : 
                       (N69)? data_i[164] : 
                       (N71)? data_i[292] : 
                       (N73)? data_i[420] : 
                       (N68)? data_i[548] : 
                       (N70)? data_i[676] : 
                       (N72)? data_i[804] : 
                       (N74)? data_i[932] : 1'b0;
  assign data_o[547] = (N67)? data_i[35] : 
                       (N69)? data_i[163] : 
                       (N71)? data_i[291] : 
                       (N73)? data_i[419] : 
                       (N68)? data_i[547] : 
                       (N70)? data_i[675] : 
                       (N72)? data_i[803] : 
                       (N74)? data_i[931] : 1'b0;
  assign data_o[546] = (N67)? data_i[34] : 
                       (N69)? data_i[162] : 
                       (N71)? data_i[290] : 
                       (N73)? data_i[418] : 
                       (N68)? data_i[546] : 
                       (N70)? data_i[674] : 
                       (N72)? data_i[802] : 
                       (N74)? data_i[930] : 1'b0;
  assign data_o[545] = (N67)? data_i[33] : 
                       (N69)? data_i[161] : 
                       (N71)? data_i[289] : 
                       (N73)? data_i[417] : 
                       (N68)? data_i[545] : 
                       (N70)? data_i[673] : 
                       (N72)? data_i[801] : 
                       (N74)? data_i[929] : 1'b0;
  assign data_o[544] = (N67)? data_i[32] : 
                       (N69)? data_i[160] : 
                       (N71)? data_i[288] : 
                       (N73)? data_i[416] : 
                       (N68)? data_i[544] : 
                       (N70)? data_i[672] : 
                       (N72)? data_i[800] : 
                       (N74)? data_i[928] : 1'b0;
  assign data_o[543] = (N67)? data_i[31] : 
                       (N69)? data_i[159] : 
                       (N71)? data_i[287] : 
                       (N73)? data_i[415] : 
                       (N68)? data_i[543] : 
                       (N70)? data_i[671] : 
                       (N72)? data_i[799] : 
                       (N74)? data_i[927] : 1'b0;
  assign data_o[542] = (N67)? data_i[30] : 
                       (N69)? data_i[158] : 
                       (N71)? data_i[286] : 
                       (N73)? data_i[414] : 
                       (N68)? data_i[542] : 
                       (N70)? data_i[670] : 
                       (N72)? data_i[798] : 
                       (N74)? data_i[926] : 1'b0;
  assign data_o[541] = (N67)? data_i[29] : 
                       (N69)? data_i[157] : 
                       (N71)? data_i[285] : 
                       (N73)? data_i[413] : 
                       (N68)? data_i[541] : 
                       (N70)? data_i[669] : 
                       (N72)? data_i[797] : 
                       (N74)? data_i[925] : 1'b0;
  assign data_o[540] = (N67)? data_i[28] : 
                       (N69)? data_i[156] : 
                       (N71)? data_i[284] : 
                       (N73)? data_i[412] : 
                       (N68)? data_i[540] : 
                       (N70)? data_i[668] : 
                       (N72)? data_i[796] : 
                       (N74)? data_i[924] : 1'b0;
  assign data_o[539] = (N67)? data_i[27] : 
                       (N69)? data_i[155] : 
                       (N71)? data_i[283] : 
                       (N73)? data_i[411] : 
                       (N68)? data_i[539] : 
                       (N70)? data_i[667] : 
                       (N72)? data_i[795] : 
                       (N74)? data_i[923] : 1'b0;
  assign data_o[538] = (N67)? data_i[26] : 
                       (N69)? data_i[154] : 
                       (N71)? data_i[282] : 
                       (N73)? data_i[410] : 
                       (N68)? data_i[538] : 
                       (N70)? data_i[666] : 
                       (N72)? data_i[794] : 
                       (N74)? data_i[922] : 1'b0;
  assign data_o[537] = (N67)? data_i[25] : 
                       (N69)? data_i[153] : 
                       (N71)? data_i[281] : 
                       (N73)? data_i[409] : 
                       (N68)? data_i[537] : 
                       (N70)? data_i[665] : 
                       (N72)? data_i[793] : 
                       (N74)? data_i[921] : 1'b0;
  assign data_o[536] = (N67)? data_i[24] : 
                       (N69)? data_i[152] : 
                       (N71)? data_i[280] : 
                       (N73)? data_i[408] : 
                       (N68)? data_i[536] : 
                       (N70)? data_i[664] : 
                       (N72)? data_i[792] : 
                       (N74)? data_i[920] : 1'b0;
  assign data_o[535] = (N67)? data_i[23] : 
                       (N69)? data_i[151] : 
                       (N71)? data_i[279] : 
                       (N73)? data_i[407] : 
                       (N68)? data_i[535] : 
                       (N70)? data_i[663] : 
                       (N72)? data_i[791] : 
                       (N74)? data_i[919] : 1'b0;
  assign data_o[534] = (N67)? data_i[22] : 
                       (N69)? data_i[150] : 
                       (N71)? data_i[278] : 
                       (N73)? data_i[406] : 
                       (N68)? data_i[534] : 
                       (N70)? data_i[662] : 
                       (N72)? data_i[790] : 
                       (N74)? data_i[918] : 1'b0;
  assign data_o[533] = (N67)? data_i[21] : 
                       (N69)? data_i[149] : 
                       (N71)? data_i[277] : 
                       (N73)? data_i[405] : 
                       (N68)? data_i[533] : 
                       (N70)? data_i[661] : 
                       (N72)? data_i[789] : 
                       (N74)? data_i[917] : 1'b0;
  assign data_o[532] = (N67)? data_i[20] : 
                       (N69)? data_i[148] : 
                       (N71)? data_i[276] : 
                       (N73)? data_i[404] : 
                       (N68)? data_i[532] : 
                       (N70)? data_i[660] : 
                       (N72)? data_i[788] : 
                       (N74)? data_i[916] : 1'b0;
  assign data_o[531] = (N67)? data_i[19] : 
                       (N69)? data_i[147] : 
                       (N71)? data_i[275] : 
                       (N73)? data_i[403] : 
                       (N68)? data_i[531] : 
                       (N70)? data_i[659] : 
                       (N72)? data_i[787] : 
                       (N74)? data_i[915] : 1'b0;
  assign data_o[530] = (N67)? data_i[18] : 
                       (N69)? data_i[146] : 
                       (N71)? data_i[274] : 
                       (N73)? data_i[402] : 
                       (N68)? data_i[530] : 
                       (N70)? data_i[658] : 
                       (N72)? data_i[786] : 
                       (N74)? data_i[914] : 1'b0;
  assign data_o[529] = (N67)? data_i[17] : 
                       (N69)? data_i[145] : 
                       (N71)? data_i[273] : 
                       (N73)? data_i[401] : 
                       (N68)? data_i[529] : 
                       (N70)? data_i[657] : 
                       (N72)? data_i[785] : 
                       (N74)? data_i[913] : 1'b0;
  assign data_o[528] = (N67)? data_i[16] : 
                       (N69)? data_i[144] : 
                       (N71)? data_i[272] : 
                       (N73)? data_i[400] : 
                       (N68)? data_i[528] : 
                       (N70)? data_i[656] : 
                       (N72)? data_i[784] : 
                       (N74)? data_i[912] : 1'b0;
  assign data_o[527] = (N67)? data_i[15] : 
                       (N69)? data_i[143] : 
                       (N71)? data_i[271] : 
                       (N73)? data_i[399] : 
                       (N68)? data_i[527] : 
                       (N70)? data_i[655] : 
                       (N72)? data_i[783] : 
                       (N74)? data_i[911] : 1'b0;
  assign data_o[526] = (N67)? data_i[14] : 
                       (N69)? data_i[142] : 
                       (N71)? data_i[270] : 
                       (N73)? data_i[398] : 
                       (N68)? data_i[526] : 
                       (N70)? data_i[654] : 
                       (N72)? data_i[782] : 
                       (N74)? data_i[910] : 1'b0;
  assign data_o[525] = (N67)? data_i[13] : 
                       (N69)? data_i[141] : 
                       (N71)? data_i[269] : 
                       (N73)? data_i[397] : 
                       (N68)? data_i[525] : 
                       (N70)? data_i[653] : 
                       (N72)? data_i[781] : 
                       (N74)? data_i[909] : 1'b0;
  assign data_o[524] = (N67)? data_i[12] : 
                       (N69)? data_i[140] : 
                       (N71)? data_i[268] : 
                       (N73)? data_i[396] : 
                       (N68)? data_i[524] : 
                       (N70)? data_i[652] : 
                       (N72)? data_i[780] : 
                       (N74)? data_i[908] : 1'b0;
  assign data_o[523] = (N67)? data_i[11] : 
                       (N69)? data_i[139] : 
                       (N71)? data_i[267] : 
                       (N73)? data_i[395] : 
                       (N68)? data_i[523] : 
                       (N70)? data_i[651] : 
                       (N72)? data_i[779] : 
                       (N74)? data_i[907] : 1'b0;
  assign data_o[522] = (N67)? data_i[10] : 
                       (N69)? data_i[138] : 
                       (N71)? data_i[266] : 
                       (N73)? data_i[394] : 
                       (N68)? data_i[522] : 
                       (N70)? data_i[650] : 
                       (N72)? data_i[778] : 
                       (N74)? data_i[906] : 1'b0;
  assign data_o[521] = (N67)? data_i[9] : 
                       (N69)? data_i[137] : 
                       (N71)? data_i[265] : 
                       (N73)? data_i[393] : 
                       (N68)? data_i[521] : 
                       (N70)? data_i[649] : 
                       (N72)? data_i[777] : 
                       (N74)? data_i[905] : 1'b0;
  assign data_o[520] = (N67)? data_i[8] : 
                       (N69)? data_i[136] : 
                       (N71)? data_i[264] : 
                       (N73)? data_i[392] : 
                       (N68)? data_i[520] : 
                       (N70)? data_i[648] : 
                       (N72)? data_i[776] : 
                       (N74)? data_i[904] : 1'b0;
  assign data_o[519] = (N67)? data_i[7] : 
                       (N69)? data_i[135] : 
                       (N71)? data_i[263] : 
                       (N73)? data_i[391] : 
                       (N68)? data_i[519] : 
                       (N70)? data_i[647] : 
                       (N72)? data_i[775] : 
                       (N74)? data_i[903] : 1'b0;
  assign data_o[518] = (N67)? data_i[6] : 
                       (N69)? data_i[134] : 
                       (N71)? data_i[262] : 
                       (N73)? data_i[390] : 
                       (N68)? data_i[518] : 
                       (N70)? data_i[646] : 
                       (N72)? data_i[774] : 
                       (N74)? data_i[902] : 1'b0;
  assign data_o[517] = (N67)? data_i[5] : 
                       (N69)? data_i[133] : 
                       (N71)? data_i[261] : 
                       (N73)? data_i[389] : 
                       (N68)? data_i[517] : 
                       (N70)? data_i[645] : 
                       (N72)? data_i[773] : 
                       (N74)? data_i[901] : 1'b0;
  assign data_o[516] = (N67)? data_i[4] : 
                       (N69)? data_i[132] : 
                       (N71)? data_i[260] : 
                       (N73)? data_i[388] : 
                       (N68)? data_i[516] : 
                       (N70)? data_i[644] : 
                       (N72)? data_i[772] : 
                       (N74)? data_i[900] : 1'b0;
  assign data_o[515] = (N67)? data_i[3] : 
                       (N69)? data_i[131] : 
                       (N71)? data_i[259] : 
                       (N73)? data_i[387] : 
                       (N68)? data_i[515] : 
                       (N70)? data_i[643] : 
                       (N72)? data_i[771] : 
                       (N74)? data_i[899] : 1'b0;
  assign data_o[514] = (N67)? data_i[2] : 
                       (N69)? data_i[130] : 
                       (N71)? data_i[258] : 
                       (N73)? data_i[386] : 
                       (N68)? data_i[514] : 
                       (N70)? data_i[642] : 
                       (N72)? data_i[770] : 
                       (N74)? data_i[898] : 1'b0;
  assign data_o[513] = (N67)? data_i[1] : 
                       (N69)? data_i[129] : 
                       (N71)? data_i[257] : 
                       (N73)? data_i[385] : 
                       (N68)? data_i[513] : 
                       (N70)? data_i[641] : 
                       (N72)? data_i[769] : 
                       (N74)? data_i[897] : 1'b0;
  assign data_o[512] = (N67)? data_i[0] : 
                       (N69)? data_i[128] : 
                       (N71)? data_i[256] : 
                       (N73)? data_i[384] : 
                       (N68)? data_i[512] : 
                       (N70)? data_i[640] : 
                       (N72)? data_i[768] : 
                       (N74)? data_i[896] : 1'b0;
  assign data_o[767] = (N82)? data_i[127] : 
                       (N84)? data_i[255] : 
                       (N86)? data_i[383] : 
                       (N88)? data_i[511] : 
                       (N83)? data_i[639] : 
                       (N85)? data_i[767] : 
                       (N87)? data_i[895] : 
                       (N89)? data_i[1023] : 1'b0;
  assign data_o[766] = (N82)? data_i[126] : 
                       (N84)? data_i[254] : 
                       (N86)? data_i[382] : 
                       (N88)? data_i[510] : 
                       (N83)? data_i[638] : 
                       (N85)? data_i[766] : 
                       (N87)? data_i[894] : 
                       (N89)? data_i[1022] : 1'b0;
  assign data_o[765] = (N82)? data_i[125] : 
                       (N84)? data_i[253] : 
                       (N86)? data_i[381] : 
                       (N88)? data_i[509] : 
                       (N83)? data_i[637] : 
                       (N85)? data_i[765] : 
                       (N87)? data_i[893] : 
                       (N89)? data_i[1021] : 1'b0;
  assign data_o[764] = (N82)? data_i[124] : 
                       (N84)? data_i[252] : 
                       (N86)? data_i[380] : 
                       (N88)? data_i[508] : 
                       (N83)? data_i[636] : 
                       (N85)? data_i[764] : 
                       (N87)? data_i[892] : 
                       (N89)? data_i[1020] : 1'b0;
  assign data_o[763] = (N82)? data_i[123] : 
                       (N84)? data_i[251] : 
                       (N86)? data_i[379] : 
                       (N88)? data_i[507] : 
                       (N83)? data_i[635] : 
                       (N85)? data_i[763] : 
                       (N87)? data_i[891] : 
                       (N89)? data_i[1019] : 1'b0;
  assign data_o[762] = (N82)? data_i[122] : 
                       (N84)? data_i[250] : 
                       (N86)? data_i[378] : 
                       (N88)? data_i[506] : 
                       (N83)? data_i[634] : 
                       (N85)? data_i[762] : 
                       (N87)? data_i[890] : 
                       (N89)? data_i[1018] : 1'b0;
  assign data_o[761] = (N82)? data_i[121] : 
                       (N84)? data_i[249] : 
                       (N86)? data_i[377] : 
                       (N88)? data_i[505] : 
                       (N83)? data_i[633] : 
                       (N85)? data_i[761] : 
                       (N87)? data_i[889] : 
                       (N89)? data_i[1017] : 1'b0;
  assign data_o[760] = (N82)? data_i[120] : 
                       (N84)? data_i[248] : 
                       (N86)? data_i[376] : 
                       (N88)? data_i[504] : 
                       (N83)? data_i[632] : 
                       (N85)? data_i[760] : 
                       (N87)? data_i[888] : 
                       (N89)? data_i[1016] : 1'b0;
  assign data_o[759] = (N82)? data_i[119] : 
                       (N84)? data_i[247] : 
                       (N86)? data_i[375] : 
                       (N88)? data_i[503] : 
                       (N83)? data_i[631] : 
                       (N85)? data_i[759] : 
                       (N87)? data_i[887] : 
                       (N89)? data_i[1015] : 1'b0;
  assign data_o[758] = (N82)? data_i[118] : 
                       (N84)? data_i[246] : 
                       (N86)? data_i[374] : 
                       (N88)? data_i[502] : 
                       (N83)? data_i[630] : 
                       (N85)? data_i[758] : 
                       (N87)? data_i[886] : 
                       (N89)? data_i[1014] : 1'b0;
  assign data_o[757] = (N82)? data_i[117] : 
                       (N84)? data_i[245] : 
                       (N86)? data_i[373] : 
                       (N88)? data_i[501] : 
                       (N83)? data_i[629] : 
                       (N85)? data_i[757] : 
                       (N87)? data_i[885] : 
                       (N89)? data_i[1013] : 1'b0;
  assign data_o[756] = (N82)? data_i[116] : 
                       (N84)? data_i[244] : 
                       (N86)? data_i[372] : 
                       (N88)? data_i[500] : 
                       (N83)? data_i[628] : 
                       (N85)? data_i[756] : 
                       (N87)? data_i[884] : 
                       (N89)? data_i[1012] : 1'b0;
  assign data_o[755] = (N82)? data_i[115] : 
                       (N84)? data_i[243] : 
                       (N86)? data_i[371] : 
                       (N88)? data_i[499] : 
                       (N83)? data_i[627] : 
                       (N85)? data_i[755] : 
                       (N87)? data_i[883] : 
                       (N89)? data_i[1011] : 1'b0;
  assign data_o[754] = (N82)? data_i[114] : 
                       (N84)? data_i[242] : 
                       (N86)? data_i[370] : 
                       (N88)? data_i[498] : 
                       (N83)? data_i[626] : 
                       (N85)? data_i[754] : 
                       (N87)? data_i[882] : 
                       (N89)? data_i[1010] : 1'b0;
  assign data_o[753] = (N82)? data_i[113] : 
                       (N84)? data_i[241] : 
                       (N86)? data_i[369] : 
                       (N88)? data_i[497] : 
                       (N83)? data_i[625] : 
                       (N85)? data_i[753] : 
                       (N87)? data_i[881] : 
                       (N89)? data_i[1009] : 1'b0;
  assign data_o[752] = (N82)? data_i[112] : 
                       (N84)? data_i[240] : 
                       (N86)? data_i[368] : 
                       (N88)? data_i[496] : 
                       (N83)? data_i[624] : 
                       (N85)? data_i[752] : 
                       (N87)? data_i[880] : 
                       (N89)? data_i[1008] : 1'b0;
  assign data_o[751] = (N82)? data_i[111] : 
                       (N84)? data_i[239] : 
                       (N86)? data_i[367] : 
                       (N88)? data_i[495] : 
                       (N83)? data_i[623] : 
                       (N85)? data_i[751] : 
                       (N87)? data_i[879] : 
                       (N89)? data_i[1007] : 1'b0;
  assign data_o[750] = (N82)? data_i[110] : 
                       (N84)? data_i[238] : 
                       (N86)? data_i[366] : 
                       (N88)? data_i[494] : 
                       (N83)? data_i[622] : 
                       (N85)? data_i[750] : 
                       (N87)? data_i[878] : 
                       (N89)? data_i[1006] : 1'b0;
  assign data_o[749] = (N82)? data_i[109] : 
                       (N84)? data_i[237] : 
                       (N86)? data_i[365] : 
                       (N88)? data_i[493] : 
                       (N83)? data_i[621] : 
                       (N85)? data_i[749] : 
                       (N87)? data_i[877] : 
                       (N89)? data_i[1005] : 1'b0;
  assign data_o[748] = (N82)? data_i[108] : 
                       (N84)? data_i[236] : 
                       (N86)? data_i[364] : 
                       (N88)? data_i[492] : 
                       (N83)? data_i[620] : 
                       (N85)? data_i[748] : 
                       (N87)? data_i[876] : 
                       (N89)? data_i[1004] : 1'b0;
  assign data_o[747] = (N82)? data_i[107] : 
                       (N84)? data_i[235] : 
                       (N86)? data_i[363] : 
                       (N88)? data_i[491] : 
                       (N83)? data_i[619] : 
                       (N85)? data_i[747] : 
                       (N87)? data_i[875] : 
                       (N89)? data_i[1003] : 1'b0;
  assign data_o[746] = (N82)? data_i[106] : 
                       (N84)? data_i[234] : 
                       (N86)? data_i[362] : 
                       (N88)? data_i[490] : 
                       (N83)? data_i[618] : 
                       (N85)? data_i[746] : 
                       (N87)? data_i[874] : 
                       (N89)? data_i[1002] : 1'b0;
  assign data_o[745] = (N82)? data_i[105] : 
                       (N84)? data_i[233] : 
                       (N86)? data_i[361] : 
                       (N88)? data_i[489] : 
                       (N83)? data_i[617] : 
                       (N85)? data_i[745] : 
                       (N87)? data_i[873] : 
                       (N89)? data_i[1001] : 1'b0;
  assign data_o[744] = (N82)? data_i[104] : 
                       (N84)? data_i[232] : 
                       (N86)? data_i[360] : 
                       (N88)? data_i[488] : 
                       (N83)? data_i[616] : 
                       (N85)? data_i[744] : 
                       (N87)? data_i[872] : 
                       (N89)? data_i[1000] : 1'b0;
  assign data_o[743] = (N82)? data_i[103] : 
                       (N84)? data_i[231] : 
                       (N86)? data_i[359] : 
                       (N88)? data_i[487] : 
                       (N83)? data_i[615] : 
                       (N85)? data_i[743] : 
                       (N87)? data_i[871] : 
                       (N89)? data_i[999] : 1'b0;
  assign data_o[742] = (N82)? data_i[102] : 
                       (N84)? data_i[230] : 
                       (N86)? data_i[358] : 
                       (N88)? data_i[486] : 
                       (N83)? data_i[614] : 
                       (N85)? data_i[742] : 
                       (N87)? data_i[870] : 
                       (N89)? data_i[998] : 1'b0;
  assign data_o[741] = (N82)? data_i[101] : 
                       (N84)? data_i[229] : 
                       (N86)? data_i[357] : 
                       (N88)? data_i[485] : 
                       (N83)? data_i[613] : 
                       (N85)? data_i[741] : 
                       (N87)? data_i[869] : 
                       (N89)? data_i[997] : 1'b0;
  assign data_o[740] = (N82)? data_i[100] : 
                       (N84)? data_i[228] : 
                       (N86)? data_i[356] : 
                       (N88)? data_i[484] : 
                       (N83)? data_i[612] : 
                       (N85)? data_i[740] : 
                       (N87)? data_i[868] : 
                       (N89)? data_i[996] : 1'b0;
  assign data_o[739] = (N82)? data_i[99] : 
                       (N84)? data_i[227] : 
                       (N86)? data_i[355] : 
                       (N88)? data_i[483] : 
                       (N83)? data_i[611] : 
                       (N85)? data_i[739] : 
                       (N87)? data_i[867] : 
                       (N89)? data_i[995] : 1'b0;
  assign data_o[738] = (N82)? data_i[98] : 
                       (N84)? data_i[226] : 
                       (N86)? data_i[354] : 
                       (N88)? data_i[482] : 
                       (N83)? data_i[610] : 
                       (N85)? data_i[738] : 
                       (N87)? data_i[866] : 
                       (N89)? data_i[994] : 1'b0;
  assign data_o[737] = (N82)? data_i[97] : 
                       (N84)? data_i[225] : 
                       (N86)? data_i[353] : 
                       (N88)? data_i[481] : 
                       (N83)? data_i[609] : 
                       (N85)? data_i[737] : 
                       (N87)? data_i[865] : 
                       (N89)? data_i[993] : 1'b0;
  assign data_o[736] = (N82)? data_i[96] : 
                       (N84)? data_i[224] : 
                       (N86)? data_i[352] : 
                       (N88)? data_i[480] : 
                       (N83)? data_i[608] : 
                       (N85)? data_i[736] : 
                       (N87)? data_i[864] : 
                       (N89)? data_i[992] : 1'b0;
  assign data_o[735] = (N82)? data_i[95] : 
                       (N84)? data_i[223] : 
                       (N86)? data_i[351] : 
                       (N88)? data_i[479] : 
                       (N83)? data_i[607] : 
                       (N85)? data_i[735] : 
                       (N87)? data_i[863] : 
                       (N89)? data_i[991] : 1'b0;
  assign data_o[734] = (N82)? data_i[94] : 
                       (N84)? data_i[222] : 
                       (N86)? data_i[350] : 
                       (N88)? data_i[478] : 
                       (N83)? data_i[606] : 
                       (N85)? data_i[734] : 
                       (N87)? data_i[862] : 
                       (N89)? data_i[990] : 1'b0;
  assign data_o[733] = (N82)? data_i[93] : 
                       (N84)? data_i[221] : 
                       (N86)? data_i[349] : 
                       (N88)? data_i[477] : 
                       (N83)? data_i[605] : 
                       (N85)? data_i[733] : 
                       (N87)? data_i[861] : 
                       (N89)? data_i[989] : 1'b0;
  assign data_o[732] = (N82)? data_i[92] : 
                       (N84)? data_i[220] : 
                       (N86)? data_i[348] : 
                       (N88)? data_i[476] : 
                       (N83)? data_i[604] : 
                       (N85)? data_i[732] : 
                       (N87)? data_i[860] : 
                       (N89)? data_i[988] : 1'b0;
  assign data_o[731] = (N82)? data_i[91] : 
                       (N84)? data_i[219] : 
                       (N86)? data_i[347] : 
                       (N88)? data_i[475] : 
                       (N83)? data_i[603] : 
                       (N85)? data_i[731] : 
                       (N87)? data_i[859] : 
                       (N89)? data_i[987] : 1'b0;
  assign data_o[730] = (N82)? data_i[90] : 
                       (N84)? data_i[218] : 
                       (N86)? data_i[346] : 
                       (N88)? data_i[474] : 
                       (N83)? data_i[602] : 
                       (N85)? data_i[730] : 
                       (N87)? data_i[858] : 
                       (N89)? data_i[986] : 1'b0;
  assign data_o[729] = (N82)? data_i[89] : 
                       (N84)? data_i[217] : 
                       (N86)? data_i[345] : 
                       (N88)? data_i[473] : 
                       (N83)? data_i[601] : 
                       (N85)? data_i[729] : 
                       (N87)? data_i[857] : 
                       (N89)? data_i[985] : 1'b0;
  assign data_o[728] = (N82)? data_i[88] : 
                       (N84)? data_i[216] : 
                       (N86)? data_i[344] : 
                       (N88)? data_i[472] : 
                       (N83)? data_i[600] : 
                       (N85)? data_i[728] : 
                       (N87)? data_i[856] : 
                       (N89)? data_i[984] : 1'b0;
  assign data_o[727] = (N82)? data_i[87] : 
                       (N84)? data_i[215] : 
                       (N86)? data_i[343] : 
                       (N88)? data_i[471] : 
                       (N83)? data_i[599] : 
                       (N85)? data_i[727] : 
                       (N87)? data_i[855] : 
                       (N89)? data_i[983] : 1'b0;
  assign data_o[726] = (N82)? data_i[86] : 
                       (N84)? data_i[214] : 
                       (N86)? data_i[342] : 
                       (N88)? data_i[470] : 
                       (N83)? data_i[598] : 
                       (N85)? data_i[726] : 
                       (N87)? data_i[854] : 
                       (N89)? data_i[982] : 1'b0;
  assign data_o[725] = (N82)? data_i[85] : 
                       (N84)? data_i[213] : 
                       (N86)? data_i[341] : 
                       (N88)? data_i[469] : 
                       (N83)? data_i[597] : 
                       (N85)? data_i[725] : 
                       (N87)? data_i[853] : 
                       (N89)? data_i[981] : 1'b0;
  assign data_o[724] = (N82)? data_i[84] : 
                       (N84)? data_i[212] : 
                       (N86)? data_i[340] : 
                       (N88)? data_i[468] : 
                       (N83)? data_i[596] : 
                       (N85)? data_i[724] : 
                       (N87)? data_i[852] : 
                       (N89)? data_i[980] : 1'b0;
  assign data_o[723] = (N82)? data_i[83] : 
                       (N84)? data_i[211] : 
                       (N86)? data_i[339] : 
                       (N88)? data_i[467] : 
                       (N83)? data_i[595] : 
                       (N85)? data_i[723] : 
                       (N87)? data_i[851] : 
                       (N89)? data_i[979] : 1'b0;
  assign data_o[722] = (N82)? data_i[82] : 
                       (N84)? data_i[210] : 
                       (N86)? data_i[338] : 
                       (N88)? data_i[466] : 
                       (N83)? data_i[594] : 
                       (N85)? data_i[722] : 
                       (N87)? data_i[850] : 
                       (N89)? data_i[978] : 1'b0;
  assign data_o[721] = (N82)? data_i[81] : 
                       (N84)? data_i[209] : 
                       (N86)? data_i[337] : 
                       (N88)? data_i[465] : 
                       (N83)? data_i[593] : 
                       (N85)? data_i[721] : 
                       (N87)? data_i[849] : 
                       (N89)? data_i[977] : 1'b0;
  assign data_o[720] = (N82)? data_i[80] : 
                       (N84)? data_i[208] : 
                       (N86)? data_i[336] : 
                       (N88)? data_i[464] : 
                       (N83)? data_i[592] : 
                       (N85)? data_i[720] : 
                       (N87)? data_i[848] : 
                       (N89)? data_i[976] : 1'b0;
  assign data_o[719] = (N82)? data_i[79] : 
                       (N84)? data_i[207] : 
                       (N86)? data_i[335] : 
                       (N88)? data_i[463] : 
                       (N83)? data_i[591] : 
                       (N85)? data_i[719] : 
                       (N87)? data_i[847] : 
                       (N89)? data_i[975] : 1'b0;
  assign data_o[718] = (N82)? data_i[78] : 
                       (N84)? data_i[206] : 
                       (N86)? data_i[334] : 
                       (N88)? data_i[462] : 
                       (N83)? data_i[590] : 
                       (N85)? data_i[718] : 
                       (N87)? data_i[846] : 
                       (N89)? data_i[974] : 1'b0;
  assign data_o[717] = (N82)? data_i[77] : 
                       (N84)? data_i[205] : 
                       (N86)? data_i[333] : 
                       (N88)? data_i[461] : 
                       (N83)? data_i[589] : 
                       (N85)? data_i[717] : 
                       (N87)? data_i[845] : 
                       (N89)? data_i[973] : 1'b0;
  assign data_o[716] = (N82)? data_i[76] : 
                       (N84)? data_i[204] : 
                       (N86)? data_i[332] : 
                       (N88)? data_i[460] : 
                       (N83)? data_i[588] : 
                       (N85)? data_i[716] : 
                       (N87)? data_i[844] : 
                       (N89)? data_i[972] : 1'b0;
  assign data_o[715] = (N82)? data_i[75] : 
                       (N84)? data_i[203] : 
                       (N86)? data_i[331] : 
                       (N88)? data_i[459] : 
                       (N83)? data_i[587] : 
                       (N85)? data_i[715] : 
                       (N87)? data_i[843] : 
                       (N89)? data_i[971] : 1'b0;
  assign data_o[714] = (N82)? data_i[74] : 
                       (N84)? data_i[202] : 
                       (N86)? data_i[330] : 
                       (N88)? data_i[458] : 
                       (N83)? data_i[586] : 
                       (N85)? data_i[714] : 
                       (N87)? data_i[842] : 
                       (N89)? data_i[970] : 1'b0;
  assign data_o[713] = (N82)? data_i[73] : 
                       (N84)? data_i[201] : 
                       (N86)? data_i[329] : 
                       (N88)? data_i[457] : 
                       (N83)? data_i[585] : 
                       (N85)? data_i[713] : 
                       (N87)? data_i[841] : 
                       (N89)? data_i[969] : 1'b0;
  assign data_o[712] = (N82)? data_i[72] : 
                       (N84)? data_i[200] : 
                       (N86)? data_i[328] : 
                       (N88)? data_i[456] : 
                       (N83)? data_i[584] : 
                       (N85)? data_i[712] : 
                       (N87)? data_i[840] : 
                       (N89)? data_i[968] : 1'b0;
  assign data_o[711] = (N82)? data_i[71] : 
                       (N84)? data_i[199] : 
                       (N86)? data_i[327] : 
                       (N88)? data_i[455] : 
                       (N83)? data_i[583] : 
                       (N85)? data_i[711] : 
                       (N87)? data_i[839] : 
                       (N89)? data_i[967] : 1'b0;
  assign data_o[710] = (N82)? data_i[70] : 
                       (N84)? data_i[198] : 
                       (N86)? data_i[326] : 
                       (N88)? data_i[454] : 
                       (N83)? data_i[582] : 
                       (N85)? data_i[710] : 
                       (N87)? data_i[838] : 
                       (N89)? data_i[966] : 1'b0;
  assign data_o[709] = (N82)? data_i[69] : 
                       (N84)? data_i[197] : 
                       (N86)? data_i[325] : 
                       (N88)? data_i[453] : 
                       (N83)? data_i[581] : 
                       (N85)? data_i[709] : 
                       (N87)? data_i[837] : 
                       (N89)? data_i[965] : 1'b0;
  assign data_o[708] = (N82)? data_i[68] : 
                       (N84)? data_i[196] : 
                       (N86)? data_i[324] : 
                       (N88)? data_i[452] : 
                       (N83)? data_i[580] : 
                       (N85)? data_i[708] : 
                       (N87)? data_i[836] : 
                       (N89)? data_i[964] : 1'b0;
  assign data_o[707] = (N82)? data_i[67] : 
                       (N84)? data_i[195] : 
                       (N86)? data_i[323] : 
                       (N88)? data_i[451] : 
                       (N83)? data_i[579] : 
                       (N85)? data_i[707] : 
                       (N87)? data_i[835] : 
                       (N89)? data_i[963] : 1'b0;
  assign data_o[706] = (N82)? data_i[66] : 
                       (N84)? data_i[194] : 
                       (N86)? data_i[322] : 
                       (N88)? data_i[450] : 
                       (N83)? data_i[578] : 
                       (N85)? data_i[706] : 
                       (N87)? data_i[834] : 
                       (N89)? data_i[962] : 1'b0;
  assign data_o[705] = (N82)? data_i[65] : 
                       (N84)? data_i[193] : 
                       (N86)? data_i[321] : 
                       (N88)? data_i[449] : 
                       (N83)? data_i[577] : 
                       (N85)? data_i[705] : 
                       (N87)? data_i[833] : 
                       (N89)? data_i[961] : 1'b0;
  assign data_o[704] = (N82)? data_i[64] : 
                       (N84)? data_i[192] : 
                       (N86)? data_i[320] : 
                       (N88)? data_i[448] : 
                       (N83)? data_i[576] : 
                       (N85)? data_i[704] : 
                       (N87)? data_i[832] : 
                       (N89)? data_i[960] : 1'b0;
  assign data_o[703] = (N82)? data_i[63] : 
                       (N84)? data_i[191] : 
                       (N86)? data_i[319] : 
                       (N88)? data_i[447] : 
                       (N83)? data_i[575] : 
                       (N85)? data_i[703] : 
                       (N87)? data_i[831] : 
                       (N89)? data_i[959] : 1'b0;
  assign data_o[702] = (N82)? data_i[62] : 
                       (N84)? data_i[190] : 
                       (N86)? data_i[318] : 
                       (N88)? data_i[446] : 
                       (N83)? data_i[574] : 
                       (N85)? data_i[702] : 
                       (N87)? data_i[830] : 
                       (N89)? data_i[958] : 1'b0;
  assign data_o[701] = (N82)? data_i[61] : 
                       (N84)? data_i[189] : 
                       (N86)? data_i[317] : 
                       (N88)? data_i[445] : 
                       (N83)? data_i[573] : 
                       (N85)? data_i[701] : 
                       (N87)? data_i[829] : 
                       (N89)? data_i[957] : 1'b0;
  assign data_o[700] = (N82)? data_i[60] : 
                       (N84)? data_i[188] : 
                       (N86)? data_i[316] : 
                       (N88)? data_i[444] : 
                       (N83)? data_i[572] : 
                       (N85)? data_i[700] : 
                       (N87)? data_i[828] : 
                       (N89)? data_i[956] : 1'b0;
  assign data_o[699] = (N82)? data_i[59] : 
                       (N84)? data_i[187] : 
                       (N86)? data_i[315] : 
                       (N88)? data_i[443] : 
                       (N83)? data_i[571] : 
                       (N85)? data_i[699] : 
                       (N87)? data_i[827] : 
                       (N89)? data_i[955] : 1'b0;
  assign data_o[698] = (N82)? data_i[58] : 
                       (N84)? data_i[186] : 
                       (N86)? data_i[314] : 
                       (N88)? data_i[442] : 
                       (N83)? data_i[570] : 
                       (N85)? data_i[698] : 
                       (N87)? data_i[826] : 
                       (N89)? data_i[954] : 1'b0;
  assign data_o[697] = (N82)? data_i[57] : 
                       (N84)? data_i[185] : 
                       (N86)? data_i[313] : 
                       (N88)? data_i[441] : 
                       (N83)? data_i[569] : 
                       (N85)? data_i[697] : 
                       (N87)? data_i[825] : 
                       (N89)? data_i[953] : 1'b0;
  assign data_o[696] = (N82)? data_i[56] : 
                       (N84)? data_i[184] : 
                       (N86)? data_i[312] : 
                       (N88)? data_i[440] : 
                       (N83)? data_i[568] : 
                       (N85)? data_i[696] : 
                       (N87)? data_i[824] : 
                       (N89)? data_i[952] : 1'b0;
  assign data_o[695] = (N82)? data_i[55] : 
                       (N84)? data_i[183] : 
                       (N86)? data_i[311] : 
                       (N88)? data_i[439] : 
                       (N83)? data_i[567] : 
                       (N85)? data_i[695] : 
                       (N87)? data_i[823] : 
                       (N89)? data_i[951] : 1'b0;
  assign data_o[694] = (N82)? data_i[54] : 
                       (N84)? data_i[182] : 
                       (N86)? data_i[310] : 
                       (N88)? data_i[438] : 
                       (N83)? data_i[566] : 
                       (N85)? data_i[694] : 
                       (N87)? data_i[822] : 
                       (N89)? data_i[950] : 1'b0;
  assign data_o[693] = (N82)? data_i[53] : 
                       (N84)? data_i[181] : 
                       (N86)? data_i[309] : 
                       (N88)? data_i[437] : 
                       (N83)? data_i[565] : 
                       (N85)? data_i[693] : 
                       (N87)? data_i[821] : 
                       (N89)? data_i[949] : 1'b0;
  assign data_o[692] = (N82)? data_i[52] : 
                       (N84)? data_i[180] : 
                       (N86)? data_i[308] : 
                       (N88)? data_i[436] : 
                       (N83)? data_i[564] : 
                       (N85)? data_i[692] : 
                       (N87)? data_i[820] : 
                       (N89)? data_i[948] : 1'b0;
  assign data_o[691] = (N82)? data_i[51] : 
                       (N84)? data_i[179] : 
                       (N86)? data_i[307] : 
                       (N88)? data_i[435] : 
                       (N83)? data_i[563] : 
                       (N85)? data_i[691] : 
                       (N87)? data_i[819] : 
                       (N89)? data_i[947] : 1'b0;
  assign data_o[690] = (N82)? data_i[50] : 
                       (N84)? data_i[178] : 
                       (N86)? data_i[306] : 
                       (N88)? data_i[434] : 
                       (N83)? data_i[562] : 
                       (N85)? data_i[690] : 
                       (N87)? data_i[818] : 
                       (N89)? data_i[946] : 1'b0;
  assign data_o[689] = (N82)? data_i[49] : 
                       (N84)? data_i[177] : 
                       (N86)? data_i[305] : 
                       (N88)? data_i[433] : 
                       (N83)? data_i[561] : 
                       (N85)? data_i[689] : 
                       (N87)? data_i[817] : 
                       (N89)? data_i[945] : 1'b0;
  assign data_o[688] = (N82)? data_i[48] : 
                       (N84)? data_i[176] : 
                       (N86)? data_i[304] : 
                       (N88)? data_i[432] : 
                       (N83)? data_i[560] : 
                       (N85)? data_i[688] : 
                       (N87)? data_i[816] : 
                       (N89)? data_i[944] : 1'b0;
  assign data_o[687] = (N82)? data_i[47] : 
                       (N84)? data_i[175] : 
                       (N86)? data_i[303] : 
                       (N88)? data_i[431] : 
                       (N83)? data_i[559] : 
                       (N85)? data_i[687] : 
                       (N87)? data_i[815] : 
                       (N89)? data_i[943] : 1'b0;
  assign data_o[686] = (N82)? data_i[46] : 
                       (N84)? data_i[174] : 
                       (N86)? data_i[302] : 
                       (N88)? data_i[430] : 
                       (N83)? data_i[558] : 
                       (N85)? data_i[686] : 
                       (N87)? data_i[814] : 
                       (N89)? data_i[942] : 1'b0;
  assign data_o[685] = (N82)? data_i[45] : 
                       (N84)? data_i[173] : 
                       (N86)? data_i[301] : 
                       (N88)? data_i[429] : 
                       (N83)? data_i[557] : 
                       (N85)? data_i[685] : 
                       (N87)? data_i[813] : 
                       (N89)? data_i[941] : 1'b0;
  assign data_o[684] = (N82)? data_i[44] : 
                       (N84)? data_i[172] : 
                       (N86)? data_i[300] : 
                       (N88)? data_i[428] : 
                       (N83)? data_i[556] : 
                       (N85)? data_i[684] : 
                       (N87)? data_i[812] : 
                       (N89)? data_i[940] : 1'b0;
  assign data_o[683] = (N82)? data_i[43] : 
                       (N84)? data_i[171] : 
                       (N86)? data_i[299] : 
                       (N88)? data_i[427] : 
                       (N83)? data_i[555] : 
                       (N85)? data_i[683] : 
                       (N87)? data_i[811] : 
                       (N89)? data_i[939] : 1'b0;
  assign data_o[682] = (N82)? data_i[42] : 
                       (N84)? data_i[170] : 
                       (N86)? data_i[298] : 
                       (N88)? data_i[426] : 
                       (N83)? data_i[554] : 
                       (N85)? data_i[682] : 
                       (N87)? data_i[810] : 
                       (N89)? data_i[938] : 1'b0;
  assign data_o[681] = (N82)? data_i[41] : 
                       (N84)? data_i[169] : 
                       (N86)? data_i[297] : 
                       (N88)? data_i[425] : 
                       (N83)? data_i[553] : 
                       (N85)? data_i[681] : 
                       (N87)? data_i[809] : 
                       (N89)? data_i[937] : 1'b0;
  assign data_o[680] = (N82)? data_i[40] : 
                       (N84)? data_i[168] : 
                       (N86)? data_i[296] : 
                       (N88)? data_i[424] : 
                       (N83)? data_i[552] : 
                       (N85)? data_i[680] : 
                       (N87)? data_i[808] : 
                       (N89)? data_i[936] : 1'b0;
  assign data_o[679] = (N82)? data_i[39] : 
                       (N84)? data_i[167] : 
                       (N86)? data_i[295] : 
                       (N88)? data_i[423] : 
                       (N83)? data_i[551] : 
                       (N85)? data_i[679] : 
                       (N87)? data_i[807] : 
                       (N89)? data_i[935] : 1'b0;
  assign data_o[678] = (N82)? data_i[38] : 
                       (N84)? data_i[166] : 
                       (N86)? data_i[294] : 
                       (N88)? data_i[422] : 
                       (N83)? data_i[550] : 
                       (N85)? data_i[678] : 
                       (N87)? data_i[806] : 
                       (N89)? data_i[934] : 1'b0;
  assign data_o[677] = (N82)? data_i[37] : 
                       (N84)? data_i[165] : 
                       (N86)? data_i[293] : 
                       (N88)? data_i[421] : 
                       (N83)? data_i[549] : 
                       (N85)? data_i[677] : 
                       (N87)? data_i[805] : 
                       (N89)? data_i[933] : 1'b0;
  assign data_o[676] = (N82)? data_i[36] : 
                       (N84)? data_i[164] : 
                       (N86)? data_i[292] : 
                       (N88)? data_i[420] : 
                       (N83)? data_i[548] : 
                       (N85)? data_i[676] : 
                       (N87)? data_i[804] : 
                       (N89)? data_i[932] : 1'b0;
  assign data_o[675] = (N82)? data_i[35] : 
                       (N84)? data_i[163] : 
                       (N86)? data_i[291] : 
                       (N88)? data_i[419] : 
                       (N83)? data_i[547] : 
                       (N85)? data_i[675] : 
                       (N87)? data_i[803] : 
                       (N89)? data_i[931] : 1'b0;
  assign data_o[674] = (N82)? data_i[34] : 
                       (N84)? data_i[162] : 
                       (N86)? data_i[290] : 
                       (N88)? data_i[418] : 
                       (N83)? data_i[546] : 
                       (N85)? data_i[674] : 
                       (N87)? data_i[802] : 
                       (N89)? data_i[930] : 1'b0;
  assign data_o[673] = (N82)? data_i[33] : 
                       (N84)? data_i[161] : 
                       (N86)? data_i[289] : 
                       (N88)? data_i[417] : 
                       (N83)? data_i[545] : 
                       (N85)? data_i[673] : 
                       (N87)? data_i[801] : 
                       (N89)? data_i[929] : 1'b0;
  assign data_o[672] = (N82)? data_i[32] : 
                       (N84)? data_i[160] : 
                       (N86)? data_i[288] : 
                       (N88)? data_i[416] : 
                       (N83)? data_i[544] : 
                       (N85)? data_i[672] : 
                       (N87)? data_i[800] : 
                       (N89)? data_i[928] : 1'b0;
  assign data_o[671] = (N82)? data_i[31] : 
                       (N84)? data_i[159] : 
                       (N86)? data_i[287] : 
                       (N88)? data_i[415] : 
                       (N83)? data_i[543] : 
                       (N85)? data_i[671] : 
                       (N87)? data_i[799] : 
                       (N89)? data_i[927] : 1'b0;
  assign data_o[670] = (N82)? data_i[30] : 
                       (N84)? data_i[158] : 
                       (N86)? data_i[286] : 
                       (N88)? data_i[414] : 
                       (N83)? data_i[542] : 
                       (N85)? data_i[670] : 
                       (N87)? data_i[798] : 
                       (N89)? data_i[926] : 1'b0;
  assign data_o[669] = (N82)? data_i[29] : 
                       (N84)? data_i[157] : 
                       (N86)? data_i[285] : 
                       (N88)? data_i[413] : 
                       (N83)? data_i[541] : 
                       (N85)? data_i[669] : 
                       (N87)? data_i[797] : 
                       (N89)? data_i[925] : 1'b0;
  assign data_o[668] = (N82)? data_i[28] : 
                       (N84)? data_i[156] : 
                       (N86)? data_i[284] : 
                       (N88)? data_i[412] : 
                       (N83)? data_i[540] : 
                       (N85)? data_i[668] : 
                       (N87)? data_i[796] : 
                       (N89)? data_i[924] : 1'b0;
  assign data_o[667] = (N82)? data_i[27] : 
                       (N84)? data_i[155] : 
                       (N86)? data_i[283] : 
                       (N88)? data_i[411] : 
                       (N83)? data_i[539] : 
                       (N85)? data_i[667] : 
                       (N87)? data_i[795] : 
                       (N89)? data_i[923] : 1'b0;
  assign data_o[666] = (N82)? data_i[26] : 
                       (N84)? data_i[154] : 
                       (N86)? data_i[282] : 
                       (N88)? data_i[410] : 
                       (N83)? data_i[538] : 
                       (N85)? data_i[666] : 
                       (N87)? data_i[794] : 
                       (N89)? data_i[922] : 1'b0;
  assign data_o[665] = (N82)? data_i[25] : 
                       (N84)? data_i[153] : 
                       (N86)? data_i[281] : 
                       (N88)? data_i[409] : 
                       (N83)? data_i[537] : 
                       (N85)? data_i[665] : 
                       (N87)? data_i[793] : 
                       (N89)? data_i[921] : 1'b0;
  assign data_o[664] = (N82)? data_i[24] : 
                       (N84)? data_i[152] : 
                       (N86)? data_i[280] : 
                       (N88)? data_i[408] : 
                       (N83)? data_i[536] : 
                       (N85)? data_i[664] : 
                       (N87)? data_i[792] : 
                       (N89)? data_i[920] : 1'b0;
  assign data_o[663] = (N82)? data_i[23] : 
                       (N84)? data_i[151] : 
                       (N86)? data_i[279] : 
                       (N88)? data_i[407] : 
                       (N83)? data_i[535] : 
                       (N85)? data_i[663] : 
                       (N87)? data_i[791] : 
                       (N89)? data_i[919] : 1'b0;
  assign data_o[662] = (N82)? data_i[22] : 
                       (N84)? data_i[150] : 
                       (N86)? data_i[278] : 
                       (N88)? data_i[406] : 
                       (N83)? data_i[534] : 
                       (N85)? data_i[662] : 
                       (N87)? data_i[790] : 
                       (N89)? data_i[918] : 1'b0;
  assign data_o[661] = (N82)? data_i[21] : 
                       (N84)? data_i[149] : 
                       (N86)? data_i[277] : 
                       (N88)? data_i[405] : 
                       (N83)? data_i[533] : 
                       (N85)? data_i[661] : 
                       (N87)? data_i[789] : 
                       (N89)? data_i[917] : 1'b0;
  assign data_o[660] = (N82)? data_i[20] : 
                       (N84)? data_i[148] : 
                       (N86)? data_i[276] : 
                       (N88)? data_i[404] : 
                       (N83)? data_i[532] : 
                       (N85)? data_i[660] : 
                       (N87)? data_i[788] : 
                       (N89)? data_i[916] : 1'b0;
  assign data_o[659] = (N82)? data_i[19] : 
                       (N84)? data_i[147] : 
                       (N86)? data_i[275] : 
                       (N88)? data_i[403] : 
                       (N83)? data_i[531] : 
                       (N85)? data_i[659] : 
                       (N87)? data_i[787] : 
                       (N89)? data_i[915] : 1'b0;
  assign data_o[658] = (N82)? data_i[18] : 
                       (N84)? data_i[146] : 
                       (N86)? data_i[274] : 
                       (N88)? data_i[402] : 
                       (N83)? data_i[530] : 
                       (N85)? data_i[658] : 
                       (N87)? data_i[786] : 
                       (N89)? data_i[914] : 1'b0;
  assign data_o[657] = (N82)? data_i[17] : 
                       (N84)? data_i[145] : 
                       (N86)? data_i[273] : 
                       (N88)? data_i[401] : 
                       (N83)? data_i[529] : 
                       (N85)? data_i[657] : 
                       (N87)? data_i[785] : 
                       (N89)? data_i[913] : 1'b0;
  assign data_o[656] = (N82)? data_i[16] : 
                       (N84)? data_i[144] : 
                       (N86)? data_i[272] : 
                       (N88)? data_i[400] : 
                       (N83)? data_i[528] : 
                       (N85)? data_i[656] : 
                       (N87)? data_i[784] : 
                       (N89)? data_i[912] : 1'b0;
  assign data_o[655] = (N82)? data_i[15] : 
                       (N84)? data_i[143] : 
                       (N86)? data_i[271] : 
                       (N88)? data_i[399] : 
                       (N83)? data_i[527] : 
                       (N85)? data_i[655] : 
                       (N87)? data_i[783] : 
                       (N89)? data_i[911] : 1'b0;
  assign data_o[654] = (N82)? data_i[14] : 
                       (N84)? data_i[142] : 
                       (N86)? data_i[270] : 
                       (N88)? data_i[398] : 
                       (N83)? data_i[526] : 
                       (N85)? data_i[654] : 
                       (N87)? data_i[782] : 
                       (N89)? data_i[910] : 1'b0;
  assign data_o[653] = (N82)? data_i[13] : 
                       (N84)? data_i[141] : 
                       (N86)? data_i[269] : 
                       (N88)? data_i[397] : 
                       (N83)? data_i[525] : 
                       (N85)? data_i[653] : 
                       (N87)? data_i[781] : 
                       (N89)? data_i[909] : 1'b0;
  assign data_o[652] = (N82)? data_i[12] : 
                       (N84)? data_i[140] : 
                       (N86)? data_i[268] : 
                       (N88)? data_i[396] : 
                       (N83)? data_i[524] : 
                       (N85)? data_i[652] : 
                       (N87)? data_i[780] : 
                       (N89)? data_i[908] : 1'b0;
  assign data_o[651] = (N82)? data_i[11] : 
                       (N84)? data_i[139] : 
                       (N86)? data_i[267] : 
                       (N88)? data_i[395] : 
                       (N83)? data_i[523] : 
                       (N85)? data_i[651] : 
                       (N87)? data_i[779] : 
                       (N89)? data_i[907] : 1'b0;
  assign data_o[650] = (N82)? data_i[10] : 
                       (N84)? data_i[138] : 
                       (N86)? data_i[266] : 
                       (N88)? data_i[394] : 
                       (N83)? data_i[522] : 
                       (N85)? data_i[650] : 
                       (N87)? data_i[778] : 
                       (N89)? data_i[906] : 1'b0;
  assign data_o[649] = (N82)? data_i[9] : 
                       (N84)? data_i[137] : 
                       (N86)? data_i[265] : 
                       (N88)? data_i[393] : 
                       (N83)? data_i[521] : 
                       (N85)? data_i[649] : 
                       (N87)? data_i[777] : 
                       (N89)? data_i[905] : 1'b0;
  assign data_o[648] = (N82)? data_i[8] : 
                       (N84)? data_i[136] : 
                       (N86)? data_i[264] : 
                       (N88)? data_i[392] : 
                       (N83)? data_i[520] : 
                       (N85)? data_i[648] : 
                       (N87)? data_i[776] : 
                       (N89)? data_i[904] : 1'b0;
  assign data_o[647] = (N82)? data_i[7] : 
                       (N84)? data_i[135] : 
                       (N86)? data_i[263] : 
                       (N88)? data_i[391] : 
                       (N83)? data_i[519] : 
                       (N85)? data_i[647] : 
                       (N87)? data_i[775] : 
                       (N89)? data_i[903] : 1'b0;
  assign data_o[646] = (N82)? data_i[6] : 
                       (N84)? data_i[134] : 
                       (N86)? data_i[262] : 
                       (N88)? data_i[390] : 
                       (N83)? data_i[518] : 
                       (N85)? data_i[646] : 
                       (N87)? data_i[774] : 
                       (N89)? data_i[902] : 1'b0;
  assign data_o[645] = (N82)? data_i[5] : 
                       (N84)? data_i[133] : 
                       (N86)? data_i[261] : 
                       (N88)? data_i[389] : 
                       (N83)? data_i[517] : 
                       (N85)? data_i[645] : 
                       (N87)? data_i[773] : 
                       (N89)? data_i[901] : 1'b0;
  assign data_o[644] = (N82)? data_i[4] : 
                       (N84)? data_i[132] : 
                       (N86)? data_i[260] : 
                       (N88)? data_i[388] : 
                       (N83)? data_i[516] : 
                       (N85)? data_i[644] : 
                       (N87)? data_i[772] : 
                       (N89)? data_i[900] : 1'b0;
  assign data_o[643] = (N82)? data_i[3] : 
                       (N84)? data_i[131] : 
                       (N86)? data_i[259] : 
                       (N88)? data_i[387] : 
                       (N83)? data_i[515] : 
                       (N85)? data_i[643] : 
                       (N87)? data_i[771] : 
                       (N89)? data_i[899] : 1'b0;
  assign data_o[642] = (N82)? data_i[2] : 
                       (N84)? data_i[130] : 
                       (N86)? data_i[258] : 
                       (N88)? data_i[386] : 
                       (N83)? data_i[514] : 
                       (N85)? data_i[642] : 
                       (N87)? data_i[770] : 
                       (N89)? data_i[898] : 1'b0;
  assign data_o[641] = (N82)? data_i[1] : 
                       (N84)? data_i[129] : 
                       (N86)? data_i[257] : 
                       (N88)? data_i[385] : 
                       (N83)? data_i[513] : 
                       (N85)? data_i[641] : 
                       (N87)? data_i[769] : 
                       (N89)? data_i[897] : 1'b0;
  assign data_o[640] = (N82)? data_i[0] : 
                       (N84)? data_i[128] : 
                       (N86)? data_i[256] : 
                       (N88)? data_i[384] : 
                       (N83)? data_i[512] : 
                       (N85)? data_i[640] : 
                       (N87)? data_i[768] : 
                       (N89)? data_i[896] : 1'b0;
  assign data_o[895] = (N97)? data_i[127] : 
                       (N99)? data_i[255] : 
                       (N101)? data_i[383] : 
                       (N103)? data_i[511] : 
                       (N98)? data_i[639] : 
                       (N100)? data_i[767] : 
                       (N102)? data_i[895] : 
                       (N104)? data_i[1023] : 1'b0;
  assign data_o[894] = (N97)? data_i[126] : 
                       (N99)? data_i[254] : 
                       (N101)? data_i[382] : 
                       (N103)? data_i[510] : 
                       (N98)? data_i[638] : 
                       (N100)? data_i[766] : 
                       (N102)? data_i[894] : 
                       (N104)? data_i[1022] : 1'b0;
  assign data_o[893] = (N97)? data_i[125] : 
                       (N99)? data_i[253] : 
                       (N101)? data_i[381] : 
                       (N103)? data_i[509] : 
                       (N98)? data_i[637] : 
                       (N100)? data_i[765] : 
                       (N102)? data_i[893] : 
                       (N104)? data_i[1021] : 1'b0;
  assign data_o[892] = (N97)? data_i[124] : 
                       (N99)? data_i[252] : 
                       (N101)? data_i[380] : 
                       (N103)? data_i[508] : 
                       (N98)? data_i[636] : 
                       (N100)? data_i[764] : 
                       (N102)? data_i[892] : 
                       (N104)? data_i[1020] : 1'b0;
  assign data_o[891] = (N97)? data_i[123] : 
                       (N99)? data_i[251] : 
                       (N101)? data_i[379] : 
                       (N103)? data_i[507] : 
                       (N98)? data_i[635] : 
                       (N100)? data_i[763] : 
                       (N102)? data_i[891] : 
                       (N104)? data_i[1019] : 1'b0;
  assign data_o[890] = (N97)? data_i[122] : 
                       (N99)? data_i[250] : 
                       (N101)? data_i[378] : 
                       (N103)? data_i[506] : 
                       (N98)? data_i[634] : 
                       (N100)? data_i[762] : 
                       (N102)? data_i[890] : 
                       (N104)? data_i[1018] : 1'b0;
  assign data_o[889] = (N97)? data_i[121] : 
                       (N99)? data_i[249] : 
                       (N101)? data_i[377] : 
                       (N103)? data_i[505] : 
                       (N98)? data_i[633] : 
                       (N100)? data_i[761] : 
                       (N102)? data_i[889] : 
                       (N104)? data_i[1017] : 1'b0;
  assign data_o[888] = (N97)? data_i[120] : 
                       (N99)? data_i[248] : 
                       (N101)? data_i[376] : 
                       (N103)? data_i[504] : 
                       (N98)? data_i[632] : 
                       (N100)? data_i[760] : 
                       (N102)? data_i[888] : 
                       (N104)? data_i[1016] : 1'b0;
  assign data_o[887] = (N97)? data_i[119] : 
                       (N99)? data_i[247] : 
                       (N101)? data_i[375] : 
                       (N103)? data_i[503] : 
                       (N98)? data_i[631] : 
                       (N100)? data_i[759] : 
                       (N102)? data_i[887] : 
                       (N104)? data_i[1015] : 1'b0;
  assign data_o[886] = (N97)? data_i[118] : 
                       (N99)? data_i[246] : 
                       (N101)? data_i[374] : 
                       (N103)? data_i[502] : 
                       (N98)? data_i[630] : 
                       (N100)? data_i[758] : 
                       (N102)? data_i[886] : 
                       (N104)? data_i[1014] : 1'b0;
  assign data_o[885] = (N97)? data_i[117] : 
                       (N99)? data_i[245] : 
                       (N101)? data_i[373] : 
                       (N103)? data_i[501] : 
                       (N98)? data_i[629] : 
                       (N100)? data_i[757] : 
                       (N102)? data_i[885] : 
                       (N104)? data_i[1013] : 1'b0;
  assign data_o[884] = (N97)? data_i[116] : 
                       (N99)? data_i[244] : 
                       (N101)? data_i[372] : 
                       (N103)? data_i[500] : 
                       (N98)? data_i[628] : 
                       (N100)? data_i[756] : 
                       (N102)? data_i[884] : 
                       (N104)? data_i[1012] : 1'b0;
  assign data_o[883] = (N97)? data_i[115] : 
                       (N99)? data_i[243] : 
                       (N101)? data_i[371] : 
                       (N103)? data_i[499] : 
                       (N98)? data_i[627] : 
                       (N100)? data_i[755] : 
                       (N102)? data_i[883] : 
                       (N104)? data_i[1011] : 1'b0;
  assign data_o[882] = (N97)? data_i[114] : 
                       (N99)? data_i[242] : 
                       (N101)? data_i[370] : 
                       (N103)? data_i[498] : 
                       (N98)? data_i[626] : 
                       (N100)? data_i[754] : 
                       (N102)? data_i[882] : 
                       (N104)? data_i[1010] : 1'b0;
  assign data_o[881] = (N97)? data_i[113] : 
                       (N99)? data_i[241] : 
                       (N101)? data_i[369] : 
                       (N103)? data_i[497] : 
                       (N98)? data_i[625] : 
                       (N100)? data_i[753] : 
                       (N102)? data_i[881] : 
                       (N104)? data_i[1009] : 1'b0;
  assign data_o[880] = (N97)? data_i[112] : 
                       (N99)? data_i[240] : 
                       (N101)? data_i[368] : 
                       (N103)? data_i[496] : 
                       (N98)? data_i[624] : 
                       (N100)? data_i[752] : 
                       (N102)? data_i[880] : 
                       (N104)? data_i[1008] : 1'b0;
  assign data_o[879] = (N97)? data_i[111] : 
                       (N99)? data_i[239] : 
                       (N101)? data_i[367] : 
                       (N103)? data_i[495] : 
                       (N98)? data_i[623] : 
                       (N100)? data_i[751] : 
                       (N102)? data_i[879] : 
                       (N104)? data_i[1007] : 1'b0;
  assign data_o[878] = (N97)? data_i[110] : 
                       (N99)? data_i[238] : 
                       (N101)? data_i[366] : 
                       (N103)? data_i[494] : 
                       (N98)? data_i[622] : 
                       (N100)? data_i[750] : 
                       (N102)? data_i[878] : 
                       (N104)? data_i[1006] : 1'b0;
  assign data_o[877] = (N97)? data_i[109] : 
                       (N99)? data_i[237] : 
                       (N101)? data_i[365] : 
                       (N103)? data_i[493] : 
                       (N98)? data_i[621] : 
                       (N100)? data_i[749] : 
                       (N102)? data_i[877] : 
                       (N104)? data_i[1005] : 1'b0;
  assign data_o[876] = (N97)? data_i[108] : 
                       (N99)? data_i[236] : 
                       (N101)? data_i[364] : 
                       (N103)? data_i[492] : 
                       (N98)? data_i[620] : 
                       (N100)? data_i[748] : 
                       (N102)? data_i[876] : 
                       (N104)? data_i[1004] : 1'b0;
  assign data_o[875] = (N97)? data_i[107] : 
                       (N99)? data_i[235] : 
                       (N101)? data_i[363] : 
                       (N103)? data_i[491] : 
                       (N98)? data_i[619] : 
                       (N100)? data_i[747] : 
                       (N102)? data_i[875] : 
                       (N104)? data_i[1003] : 1'b0;
  assign data_o[874] = (N97)? data_i[106] : 
                       (N99)? data_i[234] : 
                       (N101)? data_i[362] : 
                       (N103)? data_i[490] : 
                       (N98)? data_i[618] : 
                       (N100)? data_i[746] : 
                       (N102)? data_i[874] : 
                       (N104)? data_i[1002] : 1'b0;
  assign data_o[873] = (N97)? data_i[105] : 
                       (N99)? data_i[233] : 
                       (N101)? data_i[361] : 
                       (N103)? data_i[489] : 
                       (N98)? data_i[617] : 
                       (N100)? data_i[745] : 
                       (N102)? data_i[873] : 
                       (N104)? data_i[1001] : 1'b0;
  assign data_o[872] = (N97)? data_i[104] : 
                       (N99)? data_i[232] : 
                       (N101)? data_i[360] : 
                       (N103)? data_i[488] : 
                       (N98)? data_i[616] : 
                       (N100)? data_i[744] : 
                       (N102)? data_i[872] : 
                       (N104)? data_i[1000] : 1'b0;
  assign data_o[871] = (N97)? data_i[103] : 
                       (N99)? data_i[231] : 
                       (N101)? data_i[359] : 
                       (N103)? data_i[487] : 
                       (N98)? data_i[615] : 
                       (N100)? data_i[743] : 
                       (N102)? data_i[871] : 
                       (N104)? data_i[999] : 1'b0;
  assign data_o[870] = (N97)? data_i[102] : 
                       (N99)? data_i[230] : 
                       (N101)? data_i[358] : 
                       (N103)? data_i[486] : 
                       (N98)? data_i[614] : 
                       (N100)? data_i[742] : 
                       (N102)? data_i[870] : 
                       (N104)? data_i[998] : 1'b0;
  assign data_o[869] = (N97)? data_i[101] : 
                       (N99)? data_i[229] : 
                       (N101)? data_i[357] : 
                       (N103)? data_i[485] : 
                       (N98)? data_i[613] : 
                       (N100)? data_i[741] : 
                       (N102)? data_i[869] : 
                       (N104)? data_i[997] : 1'b0;
  assign data_o[868] = (N97)? data_i[100] : 
                       (N99)? data_i[228] : 
                       (N101)? data_i[356] : 
                       (N103)? data_i[484] : 
                       (N98)? data_i[612] : 
                       (N100)? data_i[740] : 
                       (N102)? data_i[868] : 
                       (N104)? data_i[996] : 1'b0;
  assign data_o[867] = (N97)? data_i[99] : 
                       (N99)? data_i[227] : 
                       (N101)? data_i[355] : 
                       (N103)? data_i[483] : 
                       (N98)? data_i[611] : 
                       (N100)? data_i[739] : 
                       (N102)? data_i[867] : 
                       (N104)? data_i[995] : 1'b0;
  assign data_o[866] = (N97)? data_i[98] : 
                       (N99)? data_i[226] : 
                       (N101)? data_i[354] : 
                       (N103)? data_i[482] : 
                       (N98)? data_i[610] : 
                       (N100)? data_i[738] : 
                       (N102)? data_i[866] : 
                       (N104)? data_i[994] : 1'b0;
  assign data_o[865] = (N97)? data_i[97] : 
                       (N99)? data_i[225] : 
                       (N101)? data_i[353] : 
                       (N103)? data_i[481] : 
                       (N98)? data_i[609] : 
                       (N100)? data_i[737] : 
                       (N102)? data_i[865] : 
                       (N104)? data_i[993] : 1'b0;
  assign data_o[864] = (N97)? data_i[96] : 
                       (N99)? data_i[224] : 
                       (N101)? data_i[352] : 
                       (N103)? data_i[480] : 
                       (N98)? data_i[608] : 
                       (N100)? data_i[736] : 
                       (N102)? data_i[864] : 
                       (N104)? data_i[992] : 1'b0;
  assign data_o[863] = (N97)? data_i[95] : 
                       (N99)? data_i[223] : 
                       (N101)? data_i[351] : 
                       (N103)? data_i[479] : 
                       (N98)? data_i[607] : 
                       (N100)? data_i[735] : 
                       (N102)? data_i[863] : 
                       (N104)? data_i[991] : 1'b0;
  assign data_o[862] = (N97)? data_i[94] : 
                       (N99)? data_i[222] : 
                       (N101)? data_i[350] : 
                       (N103)? data_i[478] : 
                       (N98)? data_i[606] : 
                       (N100)? data_i[734] : 
                       (N102)? data_i[862] : 
                       (N104)? data_i[990] : 1'b0;
  assign data_o[861] = (N97)? data_i[93] : 
                       (N99)? data_i[221] : 
                       (N101)? data_i[349] : 
                       (N103)? data_i[477] : 
                       (N98)? data_i[605] : 
                       (N100)? data_i[733] : 
                       (N102)? data_i[861] : 
                       (N104)? data_i[989] : 1'b0;
  assign data_o[860] = (N97)? data_i[92] : 
                       (N99)? data_i[220] : 
                       (N101)? data_i[348] : 
                       (N103)? data_i[476] : 
                       (N98)? data_i[604] : 
                       (N100)? data_i[732] : 
                       (N102)? data_i[860] : 
                       (N104)? data_i[988] : 1'b0;
  assign data_o[859] = (N97)? data_i[91] : 
                       (N99)? data_i[219] : 
                       (N101)? data_i[347] : 
                       (N103)? data_i[475] : 
                       (N98)? data_i[603] : 
                       (N100)? data_i[731] : 
                       (N102)? data_i[859] : 
                       (N104)? data_i[987] : 1'b0;
  assign data_o[858] = (N97)? data_i[90] : 
                       (N99)? data_i[218] : 
                       (N101)? data_i[346] : 
                       (N103)? data_i[474] : 
                       (N98)? data_i[602] : 
                       (N100)? data_i[730] : 
                       (N102)? data_i[858] : 
                       (N104)? data_i[986] : 1'b0;
  assign data_o[857] = (N97)? data_i[89] : 
                       (N99)? data_i[217] : 
                       (N101)? data_i[345] : 
                       (N103)? data_i[473] : 
                       (N98)? data_i[601] : 
                       (N100)? data_i[729] : 
                       (N102)? data_i[857] : 
                       (N104)? data_i[985] : 1'b0;
  assign data_o[856] = (N97)? data_i[88] : 
                       (N99)? data_i[216] : 
                       (N101)? data_i[344] : 
                       (N103)? data_i[472] : 
                       (N98)? data_i[600] : 
                       (N100)? data_i[728] : 
                       (N102)? data_i[856] : 
                       (N104)? data_i[984] : 1'b0;
  assign data_o[855] = (N97)? data_i[87] : 
                       (N99)? data_i[215] : 
                       (N101)? data_i[343] : 
                       (N103)? data_i[471] : 
                       (N98)? data_i[599] : 
                       (N100)? data_i[727] : 
                       (N102)? data_i[855] : 
                       (N104)? data_i[983] : 1'b0;
  assign data_o[854] = (N97)? data_i[86] : 
                       (N99)? data_i[214] : 
                       (N101)? data_i[342] : 
                       (N103)? data_i[470] : 
                       (N98)? data_i[598] : 
                       (N100)? data_i[726] : 
                       (N102)? data_i[854] : 
                       (N104)? data_i[982] : 1'b0;
  assign data_o[853] = (N97)? data_i[85] : 
                       (N99)? data_i[213] : 
                       (N101)? data_i[341] : 
                       (N103)? data_i[469] : 
                       (N98)? data_i[597] : 
                       (N100)? data_i[725] : 
                       (N102)? data_i[853] : 
                       (N104)? data_i[981] : 1'b0;
  assign data_o[852] = (N97)? data_i[84] : 
                       (N99)? data_i[212] : 
                       (N101)? data_i[340] : 
                       (N103)? data_i[468] : 
                       (N98)? data_i[596] : 
                       (N100)? data_i[724] : 
                       (N102)? data_i[852] : 
                       (N104)? data_i[980] : 1'b0;
  assign data_o[851] = (N97)? data_i[83] : 
                       (N99)? data_i[211] : 
                       (N101)? data_i[339] : 
                       (N103)? data_i[467] : 
                       (N98)? data_i[595] : 
                       (N100)? data_i[723] : 
                       (N102)? data_i[851] : 
                       (N104)? data_i[979] : 1'b0;
  assign data_o[850] = (N97)? data_i[82] : 
                       (N99)? data_i[210] : 
                       (N101)? data_i[338] : 
                       (N103)? data_i[466] : 
                       (N98)? data_i[594] : 
                       (N100)? data_i[722] : 
                       (N102)? data_i[850] : 
                       (N104)? data_i[978] : 1'b0;
  assign data_o[849] = (N97)? data_i[81] : 
                       (N99)? data_i[209] : 
                       (N101)? data_i[337] : 
                       (N103)? data_i[465] : 
                       (N98)? data_i[593] : 
                       (N100)? data_i[721] : 
                       (N102)? data_i[849] : 
                       (N104)? data_i[977] : 1'b0;
  assign data_o[848] = (N97)? data_i[80] : 
                       (N99)? data_i[208] : 
                       (N101)? data_i[336] : 
                       (N103)? data_i[464] : 
                       (N98)? data_i[592] : 
                       (N100)? data_i[720] : 
                       (N102)? data_i[848] : 
                       (N104)? data_i[976] : 1'b0;
  assign data_o[847] = (N97)? data_i[79] : 
                       (N99)? data_i[207] : 
                       (N101)? data_i[335] : 
                       (N103)? data_i[463] : 
                       (N98)? data_i[591] : 
                       (N100)? data_i[719] : 
                       (N102)? data_i[847] : 
                       (N104)? data_i[975] : 1'b0;
  assign data_o[846] = (N97)? data_i[78] : 
                       (N99)? data_i[206] : 
                       (N101)? data_i[334] : 
                       (N103)? data_i[462] : 
                       (N98)? data_i[590] : 
                       (N100)? data_i[718] : 
                       (N102)? data_i[846] : 
                       (N104)? data_i[974] : 1'b0;
  assign data_o[845] = (N97)? data_i[77] : 
                       (N99)? data_i[205] : 
                       (N101)? data_i[333] : 
                       (N103)? data_i[461] : 
                       (N98)? data_i[589] : 
                       (N100)? data_i[717] : 
                       (N102)? data_i[845] : 
                       (N104)? data_i[973] : 1'b0;
  assign data_o[844] = (N97)? data_i[76] : 
                       (N99)? data_i[204] : 
                       (N101)? data_i[332] : 
                       (N103)? data_i[460] : 
                       (N98)? data_i[588] : 
                       (N100)? data_i[716] : 
                       (N102)? data_i[844] : 
                       (N104)? data_i[972] : 1'b0;
  assign data_o[843] = (N97)? data_i[75] : 
                       (N99)? data_i[203] : 
                       (N101)? data_i[331] : 
                       (N103)? data_i[459] : 
                       (N98)? data_i[587] : 
                       (N100)? data_i[715] : 
                       (N102)? data_i[843] : 
                       (N104)? data_i[971] : 1'b0;
  assign data_o[842] = (N97)? data_i[74] : 
                       (N99)? data_i[202] : 
                       (N101)? data_i[330] : 
                       (N103)? data_i[458] : 
                       (N98)? data_i[586] : 
                       (N100)? data_i[714] : 
                       (N102)? data_i[842] : 
                       (N104)? data_i[970] : 1'b0;
  assign data_o[841] = (N97)? data_i[73] : 
                       (N99)? data_i[201] : 
                       (N101)? data_i[329] : 
                       (N103)? data_i[457] : 
                       (N98)? data_i[585] : 
                       (N100)? data_i[713] : 
                       (N102)? data_i[841] : 
                       (N104)? data_i[969] : 1'b0;
  assign data_o[840] = (N97)? data_i[72] : 
                       (N99)? data_i[200] : 
                       (N101)? data_i[328] : 
                       (N103)? data_i[456] : 
                       (N98)? data_i[584] : 
                       (N100)? data_i[712] : 
                       (N102)? data_i[840] : 
                       (N104)? data_i[968] : 1'b0;
  assign data_o[839] = (N97)? data_i[71] : 
                       (N99)? data_i[199] : 
                       (N101)? data_i[327] : 
                       (N103)? data_i[455] : 
                       (N98)? data_i[583] : 
                       (N100)? data_i[711] : 
                       (N102)? data_i[839] : 
                       (N104)? data_i[967] : 1'b0;
  assign data_o[838] = (N97)? data_i[70] : 
                       (N99)? data_i[198] : 
                       (N101)? data_i[326] : 
                       (N103)? data_i[454] : 
                       (N98)? data_i[582] : 
                       (N100)? data_i[710] : 
                       (N102)? data_i[838] : 
                       (N104)? data_i[966] : 1'b0;
  assign data_o[837] = (N97)? data_i[69] : 
                       (N99)? data_i[197] : 
                       (N101)? data_i[325] : 
                       (N103)? data_i[453] : 
                       (N98)? data_i[581] : 
                       (N100)? data_i[709] : 
                       (N102)? data_i[837] : 
                       (N104)? data_i[965] : 1'b0;
  assign data_o[836] = (N97)? data_i[68] : 
                       (N99)? data_i[196] : 
                       (N101)? data_i[324] : 
                       (N103)? data_i[452] : 
                       (N98)? data_i[580] : 
                       (N100)? data_i[708] : 
                       (N102)? data_i[836] : 
                       (N104)? data_i[964] : 1'b0;
  assign data_o[835] = (N97)? data_i[67] : 
                       (N99)? data_i[195] : 
                       (N101)? data_i[323] : 
                       (N103)? data_i[451] : 
                       (N98)? data_i[579] : 
                       (N100)? data_i[707] : 
                       (N102)? data_i[835] : 
                       (N104)? data_i[963] : 1'b0;
  assign data_o[834] = (N97)? data_i[66] : 
                       (N99)? data_i[194] : 
                       (N101)? data_i[322] : 
                       (N103)? data_i[450] : 
                       (N98)? data_i[578] : 
                       (N100)? data_i[706] : 
                       (N102)? data_i[834] : 
                       (N104)? data_i[962] : 1'b0;
  assign data_o[833] = (N97)? data_i[65] : 
                       (N99)? data_i[193] : 
                       (N101)? data_i[321] : 
                       (N103)? data_i[449] : 
                       (N98)? data_i[577] : 
                       (N100)? data_i[705] : 
                       (N102)? data_i[833] : 
                       (N104)? data_i[961] : 1'b0;
  assign data_o[832] = (N97)? data_i[64] : 
                       (N99)? data_i[192] : 
                       (N101)? data_i[320] : 
                       (N103)? data_i[448] : 
                       (N98)? data_i[576] : 
                       (N100)? data_i[704] : 
                       (N102)? data_i[832] : 
                       (N104)? data_i[960] : 1'b0;
  assign data_o[831] = (N97)? data_i[63] : 
                       (N99)? data_i[191] : 
                       (N101)? data_i[319] : 
                       (N103)? data_i[447] : 
                       (N98)? data_i[575] : 
                       (N100)? data_i[703] : 
                       (N102)? data_i[831] : 
                       (N104)? data_i[959] : 1'b0;
  assign data_o[830] = (N97)? data_i[62] : 
                       (N99)? data_i[190] : 
                       (N101)? data_i[318] : 
                       (N103)? data_i[446] : 
                       (N98)? data_i[574] : 
                       (N100)? data_i[702] : 
                       (N102)? data_i[830] : 
                       (N104)? data_i[958] : 1'b0;
  assign data_o[829] = (N97)? data_i[61] : 
                       (N99)? data_i[189] : 
                       (N101)? data_i[317] : 
                       (N103)? data_i[445] : 
                       (N98)? data_i[573] : 
                       (N100)? data_i[701] : 
                       (N102)? data_i[829] : 
                       (N104)? data_i[957] : 1'b0;
  assign data_o[828] = (N97)? data_i[60] : 
                       (N99)? data_i[188] : 
                       (N101)? data_i[316] : 
                       (N103)? data_i[444] : 
                       (N98)? data_i[572] : 
                       (N100)? data_i[700] : 
                       (N102)? data_i[828] : 
                       (N104)? data_i[956] : 1'b0;
  assign data_o[827] = (N97)? data_i[59] : 
                       (N99)? data_i[187] : 
                       (N101)? data_i[315] : 
                       (N103)? data_i[443] : 
                       (N98)? data_i[571] : 
                       (N100)? data_i[699] : 
                       (N102)? data_i[827] : 
                       (N104)? data_i[955] : 1'b0;
  assign data_o[826] = (N97)? data_i[58] : 
                       (N99)? data_i[186] : 
                       (N101)? data_i[314] : 
                       (N103)? data_i[442] : 
                       (N98)? data_i[570] : 
                       (N100)? data_i[698] : 
                       (N102)? data_i[826] : 
                       (N104)? data_i[954] : 1'b0;
  assign data_o[825] = (N97)? data_i[57] : 
                       (N99)? data_i[185] : 
                       (N101)? data_i[313] : 
                       (N103)? data_i[441] : 
                       (N98)? data_i[569] : 
                       (N100)? data_i[697] : 
                       (N102)? data_i[825] : 
                       (N104)? data_i[953] : 1'b0;
  assign data_o[824] = (N97)? data_i[56] : 
                       (N99)? data_i[184] : 
                       (N101)? data_i[312] : 
                       (N103)? data_i[440] : 
                       (N98)? data_i[568] : 
                       (N100)? data_i[696] : 
                       (N102)? data_i[824] : 
                       (N104)? data_i[952] : 1'b0;
  assign data_o[823] = (N97)? data_i[55] : 
                       (N99)? data_i[183] : 
                       (N101)? data_i[311] : 
                       (N103)? data_i[439] : 
                       (N98)? data_i[567] : 
                       (N100)? data_i[695] : 
                       (N102)? data_i[823] : 
                       (N104)? data_i[951] : 1'b0;
  assign data_o[822] = (N97)? data_i[54] : 
                       (N99)? data_i[182] : 
                       (N101)? data_i[310] : 
                       (N103)? data_i[438] : 
                       (N98)? data_i[566] : 
                       (N100)? data_i[694] : 
                       (N102)? data_i[822] : 
                       (N104)? data_i[950] : 1'b0;
  assign data_o[821] = (N97)? data_i[53] : 
                       (N99)? data_i[181] : 
                       (N101)? data_i[309] : 
                       (N103)? data_i[437] : 
                       (N98)? data_i[565] : 
                       (N100)? data_i[693] : 
                       (N102)? data_i[821] : 
                       (N104)? data_i[949] : 1'b0;
  assign data_o[820] = (N97)? data_i[52] : 
                       (N99)? data_i[180] : 
                       (N101)? data_i[308] : 
                       (N103)? data_i[436] : 
                       (N98)? data_i[564] : 
                       (N100)? data_i[692] : 
                       (N102)? data_i[820] : 
                       (N104)? data_i[948] : 1'b0;
  assign data_o[819] = (N97)? data_i[51] : 
                       (N99)? data_i[179] : 
                       (N101)? data_i[307] : 
                       (N103)? data_i[435] : 
                       (N98)? data_i[563] : 
                       (N100)? data_i[691] : 
                       (N102)? data_i[819] : 
                       (N104)? data_i[947] : 1'b0;
  assign data_o[818] = (N97)? data_i[50] : 
                       (N99)? data_i[178] : 
                       (N101)? data_i[306] : 
                       (N103)? data_i[434] : 
                       (N98)? data_i[562] : 
                       (N100)? data_i[690] : 
                       (N102)? data_i[818] : 
                       (N104)? data_i[946] : 1'b0;
  assign data_o[817] = (N97)? data_i[49] : 
                       (N99)? data_i[177] : 
                       (N101)? data_i[305] : 
                       (N103)? data_i[433] : 
                       (N98)? data_i[561] : 
                       (N100)? data_i[689] : 
                       (N102)? data_i[817] : 
                       (N104)? data_i[945] : 1'b0;
  assign data_o[816] = (N97)? data_i[48] : 
                       (N99)? data_i[176] : 
                       (N101)? data_i[304] : 
                       (N103)? data_i[432] : 
                       (N98)? data_i[560] : 
                       (N100)? data_i[688] : 
                       (N102)? data_i[816] : 
                       (N104)? data_i[944] : 1'b0;
  assign data_o[815] = (N97)? data_i[47] : 
                       (N99)? data_i[175] : 
                       (N101)? data_i[303] : 
                       (N103)? data_i[431] : 
                       (N98)? data_i[559] : 
                       (N100)? data_i[687] : 
                       (N102)? data_i[815] : 
                       (N104)? data_i[943] : 1'b0;
  assign data_o[814] = (N97)? data_i[46] : 
                       (N99)? data_i[174] : 
                       (N101)? data_i[302] : 
                       (N103)? data_i[430] : 
                       (N98)? data_i[558] : 
                       (N100)? data_i[686] : 
                       (N102)? data_i[814] : 
                       (N104)? data_i[942] : 1'b0;
  assign data_o[813] = (N97)? data_i[45] : 
                       (N99)? data_i[173] : 
                       (N101)? data_i[301] : 
                       (N103)? data_i[429] : 
                       (N98)? data_i[557] : 
                       (N100)? data_i[685] : 
                       (N102)? data_i[813] : 
                       (N104)? data_i[941] : 1'b0;
  assign data_o[812] = (N97)? data_i[44] : 
                       (N99)? data_i[172] : 
                       (N101)? data_i[300] : 
                       (N103)? data_i[428] : 
                       (N98)? data_i[556] : 
                       (N100)? data_i[684] : 
                       (N102)? data_i[812] : 
                       (N104)? data_i[940] : 1'b0;
  assign data_o[811] = (N97)? data_i[43] : 
                       (N99)? data_i[171] : 
                       (N101)? data_i[299] : 
                       (N103)? data_i[427] : 
                       (N98)? data_i[555] : 
                       (N100)? data_i[683] : 
                       (N102)? data_i[811] : 
                       (N104)? data_i[939] : 1'b0;
  assign data_o[810] = (N97)? data_i[42] : 
                       (N99)? data_i[170] : 
                       (N101)? data_i[298] : 
                       (N103)? data_i[426] : 
                       (N98)? data_i[554] : 
                       (N100)? data_i[682] : 
                       (N102)? data_i[810] : 
                       (N104)? data_i[938] : 1'b0;
  assign data_o[809] = (N97)? data_i[41] : 
                       (N99)? data_i[169] : 
                       (N101)? data_i[297] : 
                       (N103)? data_i[425] : 
                       (N98)? data_i[553] : 
                       (N100)? data_i[681] : 
                       (N102)? data_i[809] : 
                       (N104)? data_i[937] : 1'b0;
  assign data_o[808] = (N97)? data_i[40] : 
                       (N99)? data_i[168] : 
                       (N101)? data_i[296] : 
                       (N103)? data_i[424] : 
                       (N98)? data_i[552] : 
                       (N100)? data_i[680] : 
                       (N102)? data_i[808] : 
                       (N104)? data_i[936] : 1'b0;
  assign data_o[807] = (N97)? data_i[39] : 
                       (N99)? data_i[167] : 
                       (N101)? data_i[295] : 
                       (N103)? data_i[423] : 
                       (N98)? data_i[551] : 
                       (N100)? data_i[679] : 
                       (N102)? data_i[807] : 
                       (N104)? data_i[935] : 1'b0;
  assign data_o[806] = (N97)? data_i[38] : 
                       (N99)? data_i[166] : 
                       (N101)? data_i[294] : 
                       (N103)? data_i[422] : 
                       (N98)? data_i[550] : 
                       (N100)? data_i[678] : 
                       (N102)? data_i[806] : 
                       (N104)? data_i[934] : 1'b0;
  assign data_o[805] = (N97)? data_i[37] : 
                       (N99)? data_i[165] : 
                       (N101)? data_i[293] : 
                       (N103)? data_i[421] : 
                       (N98)? data_i[549] : 
                       (N100)? data_i[677] : 
                       (N102)? data_i[805] : 
                       (N104)? data_i[933] : 1'b0;
  assign data_o[804] = (N97)? data_i[36] : 
                       (N99)? data_i[164] : 
                       (N101)? data_i[292] : 
                       (N103)? data_i[420] : 
                       (N98)? data_i[548] : 
                       (N100)? data_i[676] : 
                       (N102)? data_i[804] : 
                       (N104)? data_i[932] : 1'b0;
  assign data_o[803] = (N97)? data_i[35] : 
                       (N99)? data_i[163] : 
                       (N101)? data_i[291] : 
                       (N103)? data_i[419] : 
                       (N98)? data_i[547] : 
                       (N100)? data_i[675] : 
                       (N102)? data_i[803] : 
                       (N104)? data_i[931] : 1'b0;
  assign data_o[802] = (N97)? data_i[34] : 
                       (N99)? data_i[162] : 
                       (N101)? data_i[290] : 
                       (N103)? data_i[418] : 
                       (N98)? data_i[546] : 
                       (N100)? data_i[674] : 
                       (N102)? data_i[802] : 
                       (N104)? data_i[930] : 1'b0;
  assign data_o[801] = (N97)? data_i[33] : 
                       (N99)? data_i[161] : 
                       (N101)? data_i[289] : 
                       (N103)? data_i[417] : 
                       (N98)? data_i[545] : 
                       (N100)? data_i[673] : 
                       (N102)? data_i[801] : 
                       (N104)? data_i[929] : 1'b0;
  assign data_o[800] = (N97)? data_i[32] : 
                       (N99)? data_i[160] : 
                       (N101)? data_i[288] : 
                       (N103)? data_i[416] : 
                       (N98)? data_i[544] : 
                       (N100)? data_i[672] : 
                       (N102)? data_i[800] : 
                       (N104)? data_i[928] : 1'b0;
  assign data_o[799] = (N97)? data_i[31] : 
                       (N99)? data_i[159] : 
                       (N101)? data_i[287] : 
                       (N103)? data_i[415] : 
                       (N98)? data_i[543] : 
                       (N100)? data_i[671] : 
                       (N102)? data_i[799] : 
                       (N104)? data_i[927] : 1'b0;
  assign data_o[798] = (N97)? data_i[30] : 
                       (N99)? data_i[158] : 
                       (N101)? data_i[286] : 
                       (N103)? data_i[414] : 
                       (N98)? data_i[542] : 
                       (N100)? data_i[670] : 
                       (N102)? data_i[798] : 
                       (N104)? data_i[926] : 1'b0;
  assign data_o[797] = (N97)? data_i[29] : 
                       (N99)? data_i[157] : 
                       (N101)? data_i[285] : 
                       (N103)? data_i[413] : 
                       (N98)? data_i[541] : 
                       (N100)? data_i[669] : 
                       (N102)? data_i[797] : 
                       (N104)? data_i[925] : 1'b0;
  assign data_o[796] = (N97)? data_i[28] : 
                       (N99)? data_i[156] : 
                       (N101)? data_i[284] : 
                       (N103)? data_i[412] : 
                       (N98)? data_i[540] : 
                       (N100)? data_i[668] : 
                       (N102)? data_i[796] : 
                       (N104)? data_i[924] : 1'b0;
  assign data_o[795] = (N97)? data_i[27] : 
                       (N99)? data_i[155] : 
                       (N101)? data_i[283] : 
                       (N103)? data_i[411] : 
                       (N98)? data_i[539] : 
                       (N100)? data_i[667] : 
                       (N102)? data_i[795] : 
                       (N104)? data_i[923] : 1'b0;
  assign data_o[794] = (N97)? data_i[26] : 
                       (N99)? data_i[154] : 
                       (N101)? data_i[282] : 
                       (N103)? data_i[410] : 
                       (N98)? data_i[538] : 
                       (N100)? data_i[666] : 
                       (N102)? data_i[794] : 
                       (N104)? data_i[922] : 1'b0;
  assign data_o[793] = (N97)? data_i[25] : 
                       (N99)? data_i[153] : 
                       (N101)? data_i[281] : 
                       (N103)? data_i[409] : 
                       (N98)? data_i[537] : 
                       (N100)? data_i[665] : 
                       (N102)? data_i[793] : 
                       (N104)? data_i[921] : 1'b0;
  assign data_o[792] = (N97)? data_i[24] : 
                       (N99)? data_i[152] : 
                       (N101)? data_i[280] : 
                       (N103)? data_i[408] : 
                       (N98)? data_i[536] : 
                       (N100)? data_i[664] : 
                       (N102)? data_i[792] : 
                       (N104)? data_i[920] : 1'b0;
  assign data_o[791] = (N97)? data_i[23] : 
                       (N99)? data_i[151] : 
                       (N101)? data_i[279] : 
                       (N103)? data_i[407] : 
                       (N98)? data_i[535] : 
                       (N100)? data_i[663] : 
                       (N102)? data_i[791] : 
                       (N104)? data_i[919] : 1'b0;
  assign data_o[790] = (N97)? data_i[22] : 
                       (N99)? data_i[150] : 
                       (N101)? data_i[278] : 
                       (N103)? data_i[406] : 
                       (N98)? data_i[534] : 
                       (N100)? data_i[662] : 
                       (N102)? data_i[790] : 
                       (N104)? data_i[918] : 1'b0;
  assign data_o[789] = (N97)? data_i[21] : 
                       (N99)? data_i[149] : 
                       (N101)? data_i[277] : 
                       (N103)? data_i[405] : 
                       (N98)? data_i[533] : 
                       (N100)? data_i[661] : 
                       (N102)? data_i[789] : 
                       (N104)? data_i[917] : 1'b0;
  assign data_o[788] = (N97)? data_i[20] : 
                       (N99)? data_i[148] : 
                       (N101)? data_i[276] : 
                       (N103)? data_i[404] : 
                       (N98)? data_i[532] : 
                       (N100)? data_i[660] : 
                       (N102)? data_i[788] : 
                       (N104)? data_i[916] : 1'b0;
  assign data_o[787] = (N97)? data_i[19] : 
                       (N99)? data_i[147] : 
                       (N101)? data_i[275] : 
                       (N103)? data_i[403] : 
                       (N98)? data_i[531] : 
                       (N100)? data_i[659] : 
                       (N102)? data_i[787] : 
                       (N104)? data_i[915] : 1'b0;
  assign data_o[786] = (N97)? data_i[18] : 
                       (N99)? data_i[146] : 
                       (N101)? data_i[274] : 
                       (N103)? data_i[402] : 
                       (N98)? data_i[530] : 
                       (N100)? data_i[658] : 
                       (N102)? data_i[786] : 
                       (N104)? data_i[914] : 1'b0;
  assign data_o[785] = (N97)? data_i[17] : 
                       (N99)? data_i[145] : 
                       (N101)? data_i[273] : 
                       (N103)? data_i[401] : 
                       (N98)? data_i[529] : 
                       (N100)? data_i[657] : 
                       (N102)? data_i[785] : 
                       (N104)? data_i[913] : 1'b0;
  assign data_o[784] = (N97)? data_i[16] : 
                       (N99)? data_i[144] : 
                       (N101)? data_i[272] : 
                       (N103)? data_i[400] : 
                       (N98)? data_i[528] : 
                       (N100)? data_i[656] : 
                       (N102)? data_i[784] : 
                       (N104)? data_i[912] : 1'b0;
  assign data_o[783] = (N97)? data_i[15] : 
                       (N99)? data_i[143] : 
                       (N101)? data_i[271] : 
                       (N103)? data_i[399] : 
                       (N98)? data_i[527] : 
                       (N100)? data_i[655] : 
                       (N102)? data_i[783] : 
                       (N104)? data_i[911] : 1'b0;
  assign data_o[782] = (N97)? data_i[14] : 
                       (N99)? data_i[142] : 
                       (N101)? data_i[270] : 
                       (N103)? data_i[398] : 
                       (N98)? data_i[526] : 
                       (N100)? data_i[654] : 
                       (N102)? data_i[782] : 
                       (N104)? data_i[910] : 1'b0;
  assign data_o[781] = (N97)? data_i[13] : 
                       (N99)? data_i[141] : 
                       (N101)? data_i[269] : 
                       (N103)? data_i[397] : 
                       (N98)? data_i[525] : 
                       (N100)? data_i[653] : 
                       (N102)? data_i[781] : 
                       (N104)? data_i[909] : 1'b0;
  assign data_o[780] = (N97)? data_i[12] : 
                       (N99)? data_i[140] : 
                       (N101)? data_i[268] : 
                       (N103)? data_i[396] : 
                       (N98)? data_i[524] : 
                       (N100)? data_i[652] : 
                       (N102)? data_i[780] : 
                       (N104)? data_i[908] : 1'b0;
  assign data_o[779] = (N97)? data_i[11] : 
                       (N99)? data_i[139] : 
                       (N101)? data_i[267] : 
                       (N103)? data_i[395] : 
                       (N98)? data_i[523] : 
                       (N100)? data_i[651] : 
                       (N102)? data_i[779] : 
                       (N104)? data_i[907] : 1'b0;
  assign data_o[778] = (N97)? data_i[10] : 
                       (N99)? data_i[138] : 
                       (N101)? data_i[266] : 
                       (N103)? data_i[394] : 
                       (N98)? data_i[522] : 
                       (N100)? data_i[650] : 
                       (N102)? data_i[778] : 
                       (N104)? data_i[906] : 1'b0;
  assign data_o[777] = (N97)? data_i[9] : 
                       (N99)? data_i[137] : 
                       (N101)? data_i[265] : 
                       (N103)? data_i[393] : 
                       (N98)? data_i[521] : 
                       (N100)? data_i[649] : 
                       (N102)? data_i[777] : 
                       (N104)? data_i[905] : 1'b0;
  assign data_o[776] = (N97)? data_i[8] : 
                       (N99)? data_i[136] : 
                       (N101)? data_i[264] : 
                       (N103)? data_i[392] : 
                       (N98)? data_i[520] : 
                       (N100)? data_i[648] : 
                       (N102)? data_i[776] : 
                       (N104)? data_i[904] : 1'b0;
  assign data_o[775] = (N97)? data_i[7] : 
                       (N99)? data_i[135] : 
                       (N101)? data_i[263] : 
                       (N103)? data_i[391] : 
                       (N98)? data_i[519] : 
                       (N100)? data_i[647] : 
                       (N102)? data_i[775] : 
                       (N104)? data_i[903] : 1'b0;
  assign data_o[774] = (N97)? data_i[6] : 
                       (N99)? data_i[134] : 
                       (N101)? data_i[262] : 
                       (N103)? data_i[390] : 
                       (N98)? data_i[518] : 
                       (N100)? data_i[646] : 
                       (N102)? data_i[774] : 
                       (N104)? data_i[902] : 1'b0;
  assign data_o[773] = (N97)? data_i[5] : 
                       (N99)? data_i[133] : 
                       (N101)? data_i[261] : 
                       (N103)? data_i[389] : 
                       (N98)? data_i[517] : 
                       (N100)? data_i[645] : 
                       (N102)? data_i[773] : 
                       (N104)? data_i[901] : 1'b0;
  assign data_o[772] = (N97)? data_i[4] : 
                       (N99)? data_i[132] : 
                       (N101)? data_i[260] : 
                       (N103)? data_i[388] : 
                       (N98)? data_i[516] : 
                       (N100)? data_i[644] : 
                       (N102)? data_i[772] : 
                       (N104)? data_i[900] : 1'b0;
  assign data_o[771] = (N97)? data_i[3] : 
                       (N99)? data_i[131] : 
                       (N101)? data_i[259] : 
                       (N103)? data_i[387] : 
                       (N98)? data_i[515] : 
                       (N100)? data_i[643] : 
                       (N102)? data_i[771] : 
                       (N104)? data_i[899] : 1'b0;
  assign data_o[770] = (N97)? data_i[2] : 
                       (N99)? data_i[130] : 
                       (N101)? data_i[258] : 
                       (N103)? data_i[386] : 
                       (N98)? data_i[514] : 
                       (N100)? data_i[642] : 
                       (N102)? data_i[770] : 
                       (N104)? data_i[898] : 1'b0;
  assign data_o[769] = (N97)? data_i[1] : 
                       (N99)? data_i[129] : 
                       (N101)? data_i[257] : 
                       (N103)? data_i[385] : 
                       (N98)? data_i[513] : 
                       (N100)? data_i[641] : 
                       (N102)? data_i[769] : 
                       (N104)? data_i[897] : 1'b0;
  assign data_o[768] = (N97)? data_i[0] : 
                       (N99)? data_i[128] : 
                       (N101)? data_i[256] : 
                       (N103)? data_i[384] : 
                       (N98)? data_i[512] : 
                       (N100)? data_i[640] : 
                       (N102)? data_i[768] : 
                       (N104)? data_i[896] : 1'b0;
  assign data_o[1023] = (N112)? data_i[127] : 
                        (N114)? data_i[255] : 
                        (N116)? data_i[383] : 
                        (N118)? data_i[511] : 
                        (N113)? data_i[639] : 
                        (N115)? data_i[767] : 
                        (N117)? data_i[895] : 
                        (N119)? data_i[1023] : 1'b0;
  assign data_o[1022] = (N112)? data_i[126] : 
                        (N114)? data_i[254] : 
                        (N116)? data_i[382] : 
                        (N118)? data_i[510] : 
                        (N113)? data_i[638] : 
                        (N115)? data_i[766] : 
                        (N117)? data_i[894] : 
                        (N119)? data_i[1022] : 1'b0;
  assign data_o[1021] = (N112)? data_i[125] : 
                        (N114)? data_i[253] : 
                        (N116)? data_i[381] : 
                        (N118)? data_i[509] : 
                        (N113)? data_i[637] : 
                        (N115)? data_i[765] : 
                        (N117)? data_i[893] : 
                        (N119)? data_i[1021] : 1'b0;
  assign data_o[1020] = (N112)? data_i[124] : 
                        (N114)? data_i[252] : 
                        (N116)? data_i[380] : 
                        (N118)? data_i[508] : 
                        (N113)? data_i[636] : 
                        (N115)? data_i[764] : 
                        (N117)? data_i[892] : 
                        (N119)? data_i[1020] : 1'b0;
  assign data_o[1019] = (N112)? data_i[123] : 
                        (N114)? data_i[251] : 
                        (N116)? data_i[379] : 
                        (N118)? data_i[507] : 
                        (N113)? data_i[635] : 
                        (N115)? data_i[763] : 
                        (N117)? data_i[891] : 
                        (N119)? data_i[1019] : 1'b0;
  assign data_o[1018] = (N112)? data_i[122] : 
                        (N114)? data_i[250] : 
                        (N116)? data_i[378] : 
                        (N118)? data_i[506] : 
                        (N113)? data_i[634] : 
                        (N115)? data_i[762] : 
                        (N117)? data_i[890] : 
                        (N119)? data_i[1018] : 1'b0;
  assign data_o[1017] = (N112)? data_i[121] : 
                        (N114)? data_i[249] : 
                        (N116)? data_i[377] : 
                        (N118)? data_i[505] : 
                        (N113)? data_i[633] : 
                        (N115)? data_i[761] : 
                        (N117)? data_i[889] : 
                        (N119)? data_i[1017] : 1'b0;
  assign data_o[1016] = (N112)? data_i[120] : 
                        (N114)? data_i[248] : 
                        (N116)? data_i[376] : 
                        (N118)? data_i[504] : 
                        (N113)? data_i[632] : 
                        (N115)? data_i[760] : 
                        (N117)? data_i[888] : 
                        (N119)? data_i[1016] : 1'b0;
  assign data_o[1015] = (N112)? data_i[119] : 
                        (N114)? data_i[247] : 
                        (N116)? data_i[375] : 
                        (N118)? data_i[503] : 
                        (N113)? data_i[631] : 
                        (N115)? data_i[759] : 
                        (N117)? data_i[887] : 
                        (N119)? data_i[1015] : 1'b0;
  assign data_o[1014] = (N112)? data_i[118] : 
                        (N114)? data_i[246] : 
                        (N116)? data_i[374] : 
                        (N118)? data_i[502] : 
                        (N113)? data_i[630] : 
                        (N115)? data_i[758] : 
                        (N117)? data_i[886] : 
                        (N119)? data_i[1014] : 1'b0;
  assign data_o[1013] = (N112)? data_i[117] : 
                        (N114)? data_i[245] : 
                        (N116)? data_i[373] : 
                        (N118)? data_i[501] : 
                        (N113)? data_i[629] : 
                        (N115)? data_i[757] : 
                        (N117)? data_i[885] : 
                        (N119)? data_i[1013] : 1'b0;
  assign data_o[1012] = (N112)? data_i[116] : 
                        (N114)? data_i[244] : 
                        (N116)? data_i[372] : 
                        (N118)? data_i[500] : 
                        (N113)? data_i[628] : 
                        (N115)? data_i[756] : 
                        (N117)? data_i[884] : 
                        (N119)? data_i[1012] : 1'b0;
  assign data_o[1011] = (N112)? data_i[115] : 
                        (N114)? data_i[243] : 
                        (N116)? data_i[371] : 
                        (N118)? data_i[499] : 
                        (N113)? data_i[627] : 
                        (N115)? data_i[755] : 
                        (N117)? data_i[883] : 
                        (N119)? data_i[1011] : 1'b0;
  assign data_o[1010] = (N112)? data_i[114] : 
                        (N114)? data_i[242] : 
                        (N116)? data_i[370] : 
                        (N118)? data_i[498] : 
                        (N113)? data_i[626] : 
                        (N115)? data_i[754] : 
                        (N117)? data_i[882] : 
                        (N119)? data_i[1010] : 1'b0;
  assign data_o[1009] = (N112)? data_i[113] : 
                        (N114)? data_i[241] : 
                        (N116)? data_i[369] : 
                        (N118)? data_i[497] : 
                        (N113)? data_i[625] : 
                        (N115)? data_i[753] : 
                        (N117)? data_i[881] : 
                        (N119)? data_i[1009] : 1'b0;
  assign data_o[1008] = (N112)? data_i[112] : 
                        (N114)? data_i[240] : 
                        (N116)? data_i[368] : 
                        (N118)? data_i[496] : 
                        (N113)? data_i[624] : 
                        (N115)? data_i[752] : 
                        (N117)? data_i[880] : 
                        (N119)? data_i[1008] : 1'b0;
  assign data_o[1007] = (N112)? data_i[111] : 
                        (N114)? data_i[239] : 
                        (N116)? data_i[367] : 
                        (N118)? data_i[495] : 
                        (N113)? data_i[623] : 
                        (N115)? data_i[751] : 
                        (N117)? data_i[879] : 
                        (N119)? data_i[1007] : 1'b0;
  assign data_o[1006] = (N112)? data_i[110] : 
                        (N114)? data_i[238] : 
                        (N116)? data_i[366] : 
                        (N118)? data_i[494] : 
                        (N113)? data_i[622] : 
                        (N115)? data_i[750] : 
                        (N117)? data_i[878] : 
                        (N119)? data_i[1006] : 1'b0;
  assign data_o[1005] = (N112)? data_i[109] : 
                        (N114)? data_i[237] : 
                        (N116)? data_i[365] : 
                        (N118)? data_i[493] : 
                        (N113)? data_i[621] : 
                        (N115)? data_i[749] : 
                        (N117)? data_i[877] : 
                        (N119)? data_i[1005] : 1'b0;
  assign data_o[1004] = (N112)? data_i[108] : 
                        (N114)? data_i[236] : 
                        (N116)? data_i[364] : 
                        (N118)? data_i[492] : 
                        (N113)? data_i[620] : 
                        (N115)? data_i[748] : 
                        (N117)? data_i[876] : 
                        (N119)? data_i[1004] : 1'b0;
  assign data_o[1003] = (N112)? data_i[107] : 
                        (N114)? data_i[235] : 
                        (N116)? data_i[363] : 
                        (N118)? data_i[491] : 
                        (N113)? data_i[619] : 
                        (N115)? data_i[747] : 
                        (N117)? data_i[875] : 
                        (N119)? data_i[1003] : 1'b0;
  assign data_o[1002] = (N112)? data_i[106] : 
                        (N114)? data_i[234] : 
                        (N116)? data_i[362] : 
                        (N118)? data_i[490] : 
                        (N113)? data_i[618] : 
                        (N115)? data_i[746] : 
                        (N117)? data_i[874] : 
                        (N119)? data_i[1002] : 1'b0;
  assign data_o[1001] = (N112)? data_i[105] : 
                        (N114)? data_i[233] : 
                        (N116)? data_i[361] : 
                        (N118)? data_i[489] : 
                        (N113)? data_i[617] : 
                        (N115)? data_i[745] : 
                        (N117)? data_i[873] : 
                        (N119)? data_i[1001] : 1'b0;
  assign data_o[1000] = (N112)? data_i[104] : 
                        (N114)? data_i[232] : 
                        (N116)? data_i[360] : 
                        (N118)? data_i[488] : 
                        (N113)? data_i[616] : 
                        (N115)? data_i[744] : 
                        (N117)? data_i[872] : 
                        (N119)? data_i[1000] : 1'b0;
  assign data_o[999] = (N112)? data_i[103] : 
                       (N114)? data_i[231] : 
                       (N116)? data_i[359] : 
                       (N118)? data_i[487] : 
                       (N113)? data_i[615] : 
                       (N115)? data_i[743] : 
                       (N117)? data_i[871] : 
                       (N119)? data_i[999] : 1'b0;
  assign data_o[998] = (N112)? data_i[102] : 
                       (N114)? data_i[230] : 
                       (N116)? data_i[358] : 
                       (N118)? data_i[486] : 
                       (N113)? data_i[614] : 
                       (N115)? data_i[742] : 
                       (N117)? data_i[870] : 
                       (N119)? data_i[998] : 1'b0;
  assign data_o[997] = (N112)? data_i[101] : 
                       (N114)? data_i[229] : 
                       (N116)? data_i[357] : 
                       (N118)? data_i[485] : 
                       (N113)? data_i[613] : 
                       (N115)? data_i[741] : 
                       (N117)? data_i[869] : 
                       (N119)? data_i[997] : 1'b0;
  assign data_o[996] = (N112)? data_i[100] : 
                       (N114)? data_i[228] : 
                       (N116)? data_i[356] : 
                       (N118)? data_i[484] : 
                       (N113)? data_i[612] : 
                       (N115)? data_i[740] : 
                       (N117)? data_i[868] : 
                       (N119)? data_i[996] : 1'b0;
  assign data_o[995] = (N112)? data_i[99] : 
                       (N114)? data_i[227] : 
                       (N116)? data_i[355] : 
                       (N118)? data_i[483] : 
                       (N113)? data_i[611] : 
                       (N115)? data_i[739] : 
                       (N117)? data_i[867] : 
                       (N119)? data_i[995] : 1'b0;
  assign data_o[994] = (N112)? data_i[98] : 
                       (N114)? data_i[226] : 
                       (N116)? data_i[354] : 
                       (N118)? data_i[482] : 
                       (N113)? data_i[610] : 
                       (N115)? data_i[738] : 
                       (N117)? data_i[866] : 
                       (N119)? data_i[994] : 1'b0;
  assign data_o[993] = (N112)? data_i[97] : 
                       (N114)? data_i[225] : 
                       (N116)? data_i[353] : 
                       (N118)? data_i[481] : 
                       (N113)? data_i[609] : 
                       (N115)? data_i[737] : 
                       (N117)? data_i[865] : 
                       (N119)? data_i[993] : 1'b0;
  assign data_o[992] = (N112)? data_i[96] : 
                       (N114)? data_i[224] : 
                       (N116)? data_i[352] : 
                       (N118)? data_i[480] : 
                       (N113)? data_i[608] : 
                       (N115)? data_i[736] : 
                       (N117)? data_i[864] : 
                       (N119)? data_i[992] : 1'b0;
  assign data_o[991] = (N112)? data_i[95] : 
                       (N114)? data_i[223] : 
                       (N116)? data_i[351] : 
                       (N118)? data_i[479] : 
                       (N113)? data_i[607] : 
                       (N115)? data_i[735] : 
                       (N117)? data_i[863] : 
                       (N119)? data_i[991] : 1'b0;
  assign data_o[990] = (N112)? data_i[94] : 
                       (N114)? data_i[222] : 
                       (N116)? data_i[350] : 
                       (N118)? data_i[478] : 
                       (N113)? data_i[606] : 
                       (N115)? data_i[734] : 
                       (N117)? data_i[862] : 
                       (N119)? data_i[990] : 1'b0;
  assign data_o[989] = (N112)? data_i[93] : 
                       (N114)? data_i[221] : 
                       (N116)? data_i[349] : 
                       (N118)? data_i[477] : 
                       (N113)? data_i[605] : 
                       (N115)? data_i[733] : 
                       (N117)? data_i[861] : 
                       (N119)? data_i[989] : 1'b0;
  assign data_o[988] = (N112)? data_i[92] : 
                       (N114)? data_i[220] : 
                       (N116)? data_i[348] : 
                       (N118)? data_i[476] : 
                       (N113)? data_i[604] : 
                       (N115)? data_i[732] : 
                       (N117)? data_i[860] : 
                       (N119)? data_i[988] : 1'b0;
  assign data_o[987] = (N112)? data_i[91] : 
                       (N114)? data_i[219] : 
                       (N116)? data_i[347] : 
                       (N118)? data_i[475] : 
                       (N113)? data_i[603] : 
                       (N115)? data_i[731] : 
                       (N117)? data_i[859] : 
                       (N119)? data_i[987] : 1'b0;
  assign data_o[986] = (N112)? data_i[90] : 
                       (N114)? data_i[218] : 
                       (N116)? data_i[346] : 
                       (N118)? data_i[474] : 
                       (N113)? data_i[602] : 
                       (N115)? data_i[730] : 
                       (N117)? data_i[858] : 
                       (N119)? data_i[986] : 1'b0;
  assign data_o[985] = (N112)? data_i[89] : 
                       (N114)? data_i[217] : 
                       (N116)? data_i[345] : 
                       (N118)? data_i[473] : 
                       (N113)? data_i[601] : 
                       (N115)? data_i[729] : 
                       (N117)? data_i[857] : 
                       (N119)? data_i[985] : 1'b0;
  assign data_o[984] = (N112)? data_i[88] : 
                       (N114)? data_i[216] : 
                       (N116)? data_i[344] : 
                       (N118)? data_i[472] : 
                       (N113)? data_i[600] : 
                       (N115)? data_i[728] : 
                       (N117)? data_i[856] : 
                       (N119)? data_i[984] : 1'b0;
  assign data_o[983] = (N112)? data_i[87] : 
                       (N114)? data_i[215] : 
                       (N116)? data_i[343] : 
                       (N118)? data_i[471] : 
                       (N113)? data_i[599] : 
                       (N115)? data_i[727] : 
                       (N117)? data_i[855] : 
                       (N119)? data_i[983] : 1'b0;
  assign data_o[982] = (N112)? data_i[86] : 
                       (N114)? data_i[214] : 
                       (N116)? data_i[342] : 
                       (N118)? data_i[470] : 
                       (N113)? data_i[598] : 
                       (N115)? data_i[726] : 
                       (N117)? data_i[854] : 
                       (N119)? data_i[982] : 1'b0;
  assign data_o[981] = (N112)? data_i[85] : 
                       (N114)? data_i[213] : 
                       (N116)? data_i[341] : 
                       (N118)? data_i[469] : 
                       (N113)? data_i[597] : 
                       (N115)? data_i[725] : 
                       (N117)? data_i[853] : 
                       (N119)? data_i[981] : 1'b0;
  assign data_o[980] = (N112)? data_i[84] : 
                       (N114)? data_i[212] : 
                       (N116)? data_i[340] : 
                       (N118)? data_i[468] : 
                       (N113)? data_i[596] : 
                       (N115)? data_i[724] : 
                       (N117)? data_i[852] : 
                       (N119)? data_i[980] : 1'b0;
  assign data_o[979] = (N112)? data_i[83] : 
                       (N114)? data_i[211] : 
                       (N116)? data_i[339] : 
                       (N118)? data_i[467] : 
                       (N113)? data_i[595] : 
                       (N115)? data_i[723] : 
                       (N117)? data_i[851] : 
                       (N119)? data_i[979] : 1'b0;
  assign data_o[978] = (N112)? data_i[82] : 
                       (N114)? data_i[210] : 
                       (N116)? data_i[338] : 
                       (N118)? data_i[466] : 
                       (N113)? data_i[594] : 
                       (N115)? data_i[722] : 
                       (N117)? data_i[850] : 
                       (N119)? data_i[978] : 1'b0;
  assign data_o[977] = (N112)? data_i[81] : 
                       (N114)? data_i[209] : 
                       (N116)? data_i[337] : 
                       (N118)? data_i[465] : 
                       (N113)? data_i[593] : 
                       (N115)? data_i[721] : 
                       (N117)? data_i[849] : 
                       (N119)? data_i[977] : 1'b0;
  assign data_o[976] = (N112)? data_i[80] : 
                       (N114)? data_i[208] : 
                       (N116)? data_i[336] : 
                       (N118)? data_i[464] : 
                       (N113)? data_i[592] : 
                       (N115)? data_i[720] : 
                       (N117)? data_i[848] : 
                       (N119)? data_i[976] : 1'b0;
  assign data_o[975] = (N112)? data_i[79] : 
                       (N114)? data_i[207] : 
                       (N116)? data_i[335] : 
                       (N118)? data_i[463] : 
                       (N113)? data_i[591] : 
                       (N115)? data_i[719] : 
                       (N117)? data_i[847] : 
                       (N119)? data_i[975] : 1'b0;
  assign data_o[974] = (N112)? data_i[78] : 
                       (N114)? data_i[206] : 
                       (N116)? data_i[334] : 
                       (N118)? data_i[462] : 
                       (N113)? data_i[590] : 
                       (N115)? data_i[718] : 
                       (N117)? data_i[846] : 
                       (N119)? data_i[974] : 1'b0;
  assign data_o[973] = (N112)? data_i[77] : 
                       (N114)? data_i[205] : 
                       (N116)? data_i[333] : 
                       (N118)? data_i[461] : 
                       (N113)? data_i[589] : 
                       (N115)? data_i[717] : 
                       (N117)? data_i[845] : 
                       (N119)? data_i[973] : 1'b0;
  assign data_o[972] = (N112)? data_i[76] : 
                       (N114)? data_i[204] : 
                       (N116)? data_i[332] : 
                       (N118)? data_i[460] : 
                       (N113)? data_i[588] : 
                       (N115)? data_i[716] : 
                       (N117)? data_i[844] : 
                       (N119)? data_i[972] : 1'b0;
  assign data_o[971] = (N112)? data_i[75] : 
                       (N114)? data_i[203] : 
                       (N116)? data_i[331] : 
                       (N118)? data_i[459] : 
                       (N113)? data_i[587] : 
                       (N115)? data_i[715] : 
                       (N117)? data_i[843] : 
                       (N119)? data_i[971] : 1'b0;
  assign data_o[970] = (N112)? data_i[74] : 
                       (N114)? data_i[202] : 
                       (N116)? data_i[330] : 
                       (N118)? data_i[458] : 
                       (N113)? data_i[586] : 
                       (N115)? data_i[714] : 
                       (N117)? data_i[842] : 
                       (N119)? data_i[970] : 1'b0;
  assign data_o[969] = (N112)? data_i[73] : 
                       (N114)? data_i[201] : 
                       (N116)? data_i[329] : 
                       (N118)? data_i[457] : 
                       (N113)? data_i[585] : 
                       (N115)? data_i[713] : 
                       (N117)? data_i[841] : 
                       (N119)? data_i[969] : 1'b0;
  assign data_o[968] = (N112)? data_i[72] : 
                       (N114)? data_i[200] : 
                       (N116)? data_i[328] : 
                       (N118)? data_i[456] : 
                       (N113)? data_i[584] : 
                       (N115)? data_i[712] : 
                       (N117)? data_i[840] : 
                       (N119)? data_i[968] : 1'b0;
  assign data_o[967] = (N112)? data_i[71] : 
                       (N114)? data_i[199] : 
                       (N116)? data_i[327] : 
                       (N118)? data_i[455] : 
                       (N113)? data_i[583] : 
                       (N115)? data_i[711] : 
                       (N117)? data_i[839] : 
                       (N119)? data_i[967] : 1'b0;
  assign data_o[966] = (N112)? data_i[70] : 
                       (N114)? data_i[198] : 
                       (N116)? data_i[326] : 
                       (N118)? data_i[454] : 
                       (N113)? data_i[582] : 
                       (N115)? data_i[710] : 
                       (N117)? data_i[838] : 
                       (N119)? data_i[966] : 1'b0;
  assign data_o[965] = (N112)? data_i[69] : 
                       (N114)? data_i[197] : 
                       (N116)? data_i[325] : 
                       (N118)? data_i[453] : 
                       (N113)? data_i[581] : 
                       (N115)? data_i[709] : 
                       (N117)? data_i[837] : 
                       (N119)? data_i[965] : 1'b0;
  assign data_o[964] = (N112)? data_i[68] : 
                       (N114)? data_i[196] : 
                       (N116)? data_i[324] : 
                       (N118)? data_i[452] : 
                       (N113)? data_i[580] : 
                       (N115)? data_i[708] : 
                       (N117)? data_i[836] : 
                       (N119)? data_i[964] : 1'b0;
  assign data_o[963] = (N112)? data_i[67] : 
                       (N114)? data_i[195] : 
                       (N116)? data_i[323] : 
                       (N118)? data_i[451] : 
                       (N113)? data_i[579] : 
                       (N115)? data_i[707] : 
                       (N117)? data_i[835] : 
                       (N119)? data_i[963] : 1'b0;
  assign data_o[962] = (N112)? data_i[66] : 
                       (N114)? data_i[194] : 
                       (N116)? data_i[322] : 
                       (N118)? data_i[450] : 
                       (N113)? data_i[578] : 
                       (N115)? data_i[706] : 
                       (N117)? data_i[834] : 
                       (N119)? data_i[962] : 1'b0;
  assign data_o[961] = (N112)? data_i[65] : 
                       (N114)? data_i[193] : 
                       (N116)? data_i[321] : 
                       (N118)? data_i[449] : 
                       (N113)? data_i[577] : 
                       (N115)? data_i[705] : 
                       (N117)? data_i[833] : 
                       (N119)? data_i[961] : 1'b0;
  assign data_o[960] = (N112)? data_i[64] : 
                       (N114)? data_i[192] : 
                       (N116)? data_i[320] : 
                       (N118)? data_i[448] : 
                       (N113)? data_i[576] : 
                       (N115)? data_i[704] : 
                       (N117)? data_i[832] : 
                       (N119)? data_i[960] : 1'b0;
  assign data_o[959] = (N112)? data_i[63] : 
                       (N114)? data_i[191] : 
                       (N116)? data_i[319] : 
                       (N118)? data_i[447] : 
                       (N113)? data_i[575] : 
                       (N115)? data_i[703] : 
                       (N117)? data_i[831] : 
                       (N119)? data_i[959] : 1'b0;
  assign data_o[958] = (N112)? data_i[62] : 
                       (N114)? data_i[190] : 
                       (N116)? data_i[318] : 
                       (N118)? data_i[446] : 
                       (N113)? data_i[574] : 
                       (N115)? data_i[702] : 
                       (N117)? data_i[830] : 
                       (N119)? data_i[958] : 1'b0;
  assign data_o[957] = (N112)? data_i[61] : 
                       (N114)? data_i[189] : 
                       (N116)? data_i[317] : 
                       (N118)? data_i[445] : 
                       (N113)? data_i[573] : 
                       (N115)? data_i[701] : 
                       (N117)? data_i[829] : 
                       (N119)? data_i[957] : 1'b0;
  assign data_o[956] = (N112)? data_i[60] : 
                       (N114)? data_i[188] : 
                       (N116)? data_i[316] : 
                       (N118)? data_i[444] : 
                       (N113)? data_i[572] : 
                       (N115)? data_i[700] : 
                       (N117)? data_i[828] : 
                       (N119)? data_i[956] : 1'b0;
  assign data_o[955] = (N112)? data_i[59] : 
                       (N114)? data_i[187] : 
                       (N116)? data_i[315] : 
                       (N118)? data_i[443] : 
                       (N113)? data_i[571] : 
                       (N115)? data_i[699] : 
                       (N117)? data_i[827] : 
                       (N119)? data_i[955] : 1'b0;
  assign data_o[954] = (N112)? data_i[58] : 
                       (N114)? data_i[186] : 
                       (N116)? data_i[314] : 
                       (N118)? data_i[442] : 
                       (N113)? data_i[570] : 
                       (N115)? data_i[698] : 
                       (N117)? data_i[826] : 
                       (N119)? data_i[954] : 1'b0;
  assign data_o[953] = (N112)? data_i[57] : 
                       (N114)? data_i[185] : 
                       (N116)? data_i[313] : 
                       (N118)? data_i[441] : 
                       (N113)? data_i[569] : 
                       (N115)? data_i[697] : 
                       (N117)? data_i[825] : 
                       (N119)? data_i[953] : 1'b0;
  assign data_o[952] = (N112)? data_i[56] : 
                       (N114)? data_i[184] : 
                       (N116)? data_i[312] : 
                       (N118)? data_i[440] : 
                       (N113)? data_i[568] : 
                       (N115)? data_i[696] : 
                       (N117)? data_i[824] : 
                       (N119)? data_i[952] : 1'b0;
  assign data_o[951] = (N112)? data_i[55] : 
                       (N114)? data_i[183] : 
                       (N116)? data_i[311] : 
                       (N118)? data_i[439] : 
                       (N113)? data_i[567] : 
                       (N115)? data_i[695] : 
                       (N117)? data_i[823] : 
                       (N119)? data_i[951] : 1'b0;
  assign data_o[950] = (N112)? data_i[54] : 
                       (N114)? data_i[182] : 
                       (N116)? data_i[310] : 
                       (N118)? data_i[438] : 
                       (N113)? data_i[566] : 
                       (N115)? data_i[694] : 
                       (N117)? data_i[822] : 
                       (N119)? data_i[950] : 1'b0;
  assign data_o[949] = (N112)? data_i[53] : 
                       (N114)? data_i[181] : 
                       (N116)? data_i[309] : 
                       (N118)? data_i[437] : 
                       (N113)? data_i[565] : 
                       (N115)? data_i[693] : 
                       (N117)? data_i[821] : 
                       (N119)? data_i[949] : 1'b0;
  assign data_o[948] = (N112)? data_i[52] : 
                       (N114)? data_i[180] : 
                       (N116)? data_i[308] : 
                       (N118)? data_i[436] : 
                       (N113)? data_i[564] : 
                       (N115)? data_i[692] : 
                       (N117)? data_i[820] : 
                       (N119)? data_i[948] : 1'b0;
  assign data_o[947] = (N112)? data_i[51] : 
                       (N114)? data_i[179] : 
                       (N116)? data_i[307] : 
                       (N118)? data_i[435] : 
                       (N113)? data_i[563] : 
                       (N115)? data_i[691] : 
                       (N117)? data_i[819] : 
                       (N119)? data_i[947] : 1'b0;
  assign data_o[946] = (N112)? data_i[50] : 
                       (N114)? data_i[178] : 
                       (N116)? data_i[306] : 
                       (N118)? data_i[434] : 
                       (N113)? data_i[562] : 
                       (N115)? data_i[690] : 
                       (N117)? data_i[818] : 
                       (N119)? data_i[946] : 1'b0;
  assign data_o[945] = (N112)? data_i[49] : 
                       (N114)? data_i[177] : 
                       (N116)? data_i[305] : 
                       (N118)? data_i[433] : 
                       (N113)? data_i[561] : 
                       (N115)? data_i[689] : 
                       (N117)? data_i[817] : 
                       (N119)? data_i[945] : 1'b0;
  assign data_o[944] = (N112)? data_i[48] : 
                       (N114)? data_i[176] : 
                       (N116)? data_i[304] : 
                       (N118)? data_i[432] : 
                       (N113)? data_i[560] : 
                       (N115)? data_i[688] : 
                       (N117)? data_i[816] : 
                       (N119)? data_i[944] : 1'b0;
  assign data_o[943] = (N112)? data_i[47] : 
                       (N114)? data_i[175] : 
                       (N116)? data_i[303] : 
                       (N118)? data_i[431] : 
                       (N113)? data_i[559] : 
                       (N115)? data_i[687] : 
                       (N117)? data_i[815] : 
                       (N119)? data_i[943] : 1'b0;
  assign data_o[942] = (N112)? data_i[46] : 
                       (N114)? data_i[174] : 
                       (N116)? data_i[302] : 
                       (N118)? data_i[430] : 
                       (N113)? data_i[558] : 
                       (N115)? data_i[686] : 
                       (N117)? data_i[814] : 
                       (N119)? data_i[942] : 1'b0;
  assign data_o[941] = (N112)? data_i[45] : 
                       (N114)? data_i[173] : 
                       (N116)? data_i[301] : 
                       (N118)? data_i[429] : 
                       (N113)? data_i[557] : 
                       (N115)? data_i[685] : 
                       (N117)? data_i[813] : 
                       (N119)? data_i[941] : 1'b0;
  assign data_o[940] = (N112)? data_i[44] : 
                       (N114)? data_i[172] : 
                       (N116)? data_i[300] : 
                       (N118)? data_i[428] : 
                       (N113)? data_i[556] : 
                       (N115)? data_i[684] : 
                       (N117)? data_i[812] : 
                       (N119)? data_i[940] : 1'b0;
  assign data_o[939] = (N112)? data_i[43] : 
                       (N114)? data_i[171] : 
                       (N116)? data_i[299] : 
                       (N118)? data_i[427] : 
                       (N113)? data_i[555] : 
                       (N115)? data_i[683] : 
                       (N117)? data_i[811] : 
                       (N119)? data_i[939] : 1'b0;
  assign data_o[938] = (N112)? data_i[42] : 
                       (N114)? data_i[170] : 
                       (N116)? data_i[298] : 
                       (N118)? data_i[426] : 
                       (N113)? data_i[554] : 
                       (N115)? data_i[682] : 
                       (N117)? data_i[810] : 
                       (N119)? data_i[938] : 1'b0;
  assign data_o[937] = (N112)? data_i[41] : 
                       (N114)? data_i[169] : 
                       (N116)? data_i[297] : 
                       (N118)? data_i[425] : 
                       (N113)? data_i[553] : 
                       (N115)? data_i[681] : 
                       (N117)? data_i[809] : 
                       (N119)? data_i[937] : 1'b0;
  assign data_o[936] = (N112)? data_i[40] : 
                       (N114)? data_i[168] : 
                       (N116)? data_i[296] : 
                       (N118)? data_i[424] : 
                       (N113)? data_i[552] : 
                       (N115)? data_i[680] : 
                       (N117)? data_i[808] : 
                       (N119)? data_i[936] : 1'b0;
  assign data_o[935] = (N112)? data_i[39] : 
                       (N114)? data_i[167] : 
                       (N116)? data_i[295] : 
                       (N118)? data_i[423] : 
                       (N113)? data_i[551] : 
                       (N115)? data_i[679] : 
                       (N117)? data_i[807] : 
                       (N119)? data_i[935] : 1'b0;
  assign data_o[934] = (N112)? data_i[38] : 
                       (N114)? data_i[166] : 
                       (N116)? data_i[294] : 
                       (N118)? data_i[422] : 
                       (N113)? data_i[550] : 
                       (N115)? data_i[678] : 
                       (N117)? data_i[806] : 
                       (N119)? data_i[934] : 1'b0;
  assign data_o[933] = (N112)? data_i[37] : 
                       (N114)? data_i[165] : 
                       (N116)? data_i[293] : 
                       (N118)? data_i[421] : 
                       (N113)? data_i[549] : 
                       (N115)? data_i[677] : 
                       (N117)? data_i[805] : 
                       (N119)? data_i[933] : 1'b0;
  assign data_o[932] = (N112)? data_i[36] : 
                       (N114)? data_i[164] : 
                       (N116)? data_i[292] : 
                       (N118)? data_i[420] : 
                       (N113)? data_i[548] : 
                       (N115)? data_i[676] : 
                       (N117)? data_i[804] : 
                       (N119)? data_i[932] : 1'b0;
  assign data_o[931] = (N112)? data_i[35] : 
                       (N114)? data_i[163] : 
                       (N116)? data_i[291] : 
                       (N118)? data_i[419] : 
                       (N113)? data_i[547] : 
                       (N115)? data_i[675] : 
                       (N117)? data_i[803] : 
                       (N119)? data_i[931] : 1'b0;
  assign data_o[930] = (N112)? data_i[34] : 
                       (N114)? data_i[162] : 
                       (N116)? data_i[290] : 
                       (N118)? data_i[418] : 
                       (N113)? data_i[546] : 
                       (N115)? data_i[674] : 
                       (N117)? data_i[802] : 
                       (N119)? data_i[930] : 1'b0;
  assign data_o[929] = (N112)? data_i[33] : 
                       (N114)? data_i[161] : 
                       (N116)? data_i[289] : 
                       (N118)? data_i[417] : 
                       (N113)? data_i[545] : 
                       (N115)? data_i[673] : 
                       (N117)? data_i[801] : 
                       (N119)? data_i[929] : 1'b0;
  assign data_o[928] = (N112)? data_i[32] : 
                       (N114)? data_i[160] : 
                       (N116)? data_i[288] : 
                       (N118)? data_i[416] : 
                       (N113)? data_i[544] : 
                       (N115)? data_i[672] : 
                       (N117)? data_i[800] : 
                       (N119)? data_i[928] : 1'b0;
  assign data_o[927] = (N112)? data_i[31] : 
                       (N114)? data_i[159] : 
                       (N116)? data_i[287] : 
                       (N118)? data_i[415] : 
                       (N113)? data_i[543] : 
                       (N115)? data_i[671] : 
                       (N117)? data_i[799] : 
                       (N119)? data_i[927] : 1'b0;
  assign data_o[926] = (N112)? data_i[30] : 
                       (N114)? data_i[158] : 
                       (N116)? data_i[286] : 
                       (N118)? data_i[414] : 
                       (N113)? data_i[542] : 
                       (N115)? data_i[670] : 
                       (N117)? data_i[798] : 
                       (N119)? data_i[926] : 1'b0;
  assign data_o[925] = (N112)? data_i[29] : 
                       (N114)? data_i[157] : 
                       (N116)? data_i[285] : 
                       (N118)? data_i[413] : 
                       (N113)? data_i[541] : 
                       (N115)? data_i[669] : 
                       (N117)? data_i[797] : 
                       (N119)? data_i[925] : 1'b0;
  assign data_o[924] = (N112)? data_i[28] : 
                       (N114)? data_i[156] : 
                       (N116)? data_i[284] : 
                       (N118)? data_i[412] : 
                       (N113)? data_i[540] : 
                       (N115)? data_i[668] : 
                       (N117)? data_i[796] : 
                       (N119)? data_i[924] : 1'b0;
  assign data_o[923] = (N112)? data_i[27] : 
                       (N114)? data_i[155] : 
                       (N116)? data_i[283] : 
                       (N118)? data_i[411] : 
                       (N113)? data_i[539] : 
                       (N115)? data_i[667] : 
                       (N117)? data_i[795] : 
                       (N119)? data_i[923] : 1'b0;
  assign data_o[922] = (N112)? data_i[26] : 
                       (N114)? data_i[154] : 
                       (N116)? data_i[282] : 
                       (N118)? data_i[410] : 
                       (N113)? data_i[538] : 
                       (N115)? data_i[666] : 
                       (N117)? data_i[794] : 
                       (N119)? data_i[922] : 1'b0;
  assign data_o[921] = (N112)? data_i[25] : 
                       (N114)? data_i[153] : 
                       (N116)? data_i[281] : 
                       (N118)? data_i[409] : 
                       (N113)? data_i[537] : 
                       (N115)? data_i[665] : 
                       (N117)? data_i[793] : 
                       (N119)? data_i[921] : 1'b0;
  assign data_o[920] = (N112)? data_i[24] : 
                       (N114)? data_i[152] : 
                       (N116)? data_i[280] : 
                       (N118)? data_i[408] : 
                       (N113)? data_i[536] : 
                       (N115)? data_i[664] : 
                       (N117)? data_i[792] : 
                       (N119)? data_i[920] : 1'b0;
  assign data_o[919] = (N112)? data_i[23] : 
                       (N114)? data_i[151] : 
                       (N116)? data_i[279] : 
                       (N118)? data_i[407] : 
                       (N113)? data_i[535] : 
                       (N115)? data_i[663] : 
                       (N117)? data_i[791] : 
                       (N119)? data_i[919] : 1'b0;
  assign data_o[918] = (N112)? data_i[22] : 
                       (N114)? data_i[150] : 
                       (N116)? data_i[278] : 
                       (N118)? data_i[406] : 
                       (N113)? data_i[534] : 
                       (N115)? data_i[662] : 
                       (N117)? data_i[790] : 
                       (N119)? data_i[918] : 1'b0;
  assign data_o[917] = (N112)? data_i[21] : 
                       (N114)? data_i[149] : 
                       (N116)? data_i[277] : 
                       (N118)? data_i[405] : 
                       (N113)? data_i[533] : 
                       (N115)? data_i[661] : 
                       (N117)? data_i[789] : 
                       (N119)? data_i[917] : 1'b0;
  assign data_o[916] = (N112)? data_i[20] : 
                       (N114)? data_i[148] : 
                       (N116)? data_i[276] : 
                       (N118)? data_i[404] : 
                       (N113)? data_i[532] : 
                       (N115)? data_i[660] : 
                       (N117)? data_i[788] : 
                       (N119)? data_i[916] : 1'b0;
  assign data_o[915] = (N112)? data_i[19] : 
                       (N114)? data_i[147] : 
                       (N116)? data_i[275] : 
                       (N118)? data_i[403] : 
                       (N113)? data_i[531] : 
                       (N115)? data_i[659] : 
                       (N117)? data_i[787] : 
                       (N119)? data_i[915] : 1'b0;
  assign data_o[914] = (N112)? data_i[18] : 
                       (N114)? data_i[146] : 
                       (N116)? data_i[274] : 
                       (N118)? data_i[402] : 
                       (N113)? data_i[530] : 
                       (N115)? data_i[658] : 
                       (N117)? data_i[786] : 
                       (N119)? data_i[914] : 1'b0;
  assign data_o[913] = (N112)? data_i[17] : 
                       (N114)? data_i[145] : 
                       (N116)? data_i[273] : 
                       (N118)? data_i[401] : 
                       (N113)? data_i[529] : 
                       (N115)? data_i[657] : 
                       (N117)? data_i[785] : 
                       (N119)? data_i[913] : 1'b0;
  assign data_o[912] = (N112)? data_i[16] : 
                       (N114)? data_i[144] : 
                       (N116)? data_i[272] : 
                       (N118)? data_i[400] : 
                       (N113)? data_i[528] : 
                       (N115)? data_i[656] : 
                       (N117)? data_i[784] : 
                       (N119)? data_i[912] : 1'b0;
  assign data_o[911] = (N112)? data_i[15] : 
                       (N114)? data_i[143] : 
                       (N116)? data_i[271] : 
                       (N118)? data_i[399] : 
                       (N113)? data_i[527] : 
                       (N115)? data_i[655] : 
                       (N117)? data_i[783] : 
                       (N119)? data_i[911] : 1'b0;
  assign data_o[910] = (N112)? data_i[14] : 
                       (N114)? data_i[142] : 
                       (N116)? data_i[270] : 
                       (N118)? data_i[398] : 
                       (N113)? data_i[526] : 
                       (N115)? data_i[654] : 
                       (N117)? data_i[782] : 
                       (N119)? data_i[910] : 1'b0;
  assign data_o[909] = (N112)? data_i[13] : 
                       (N114)? data_i[141] : 
                       (N116)? data_i[269] : 
                       (N118)? data_i[397] : 
                       (N113)? data_i[525] : 
                       (N115)? data_i[653] : 
                       (N117)? data_i[781] : 
                       (N119)? data_i[909] : 1'b0;
  assign data_o[908] = (N112)? data_i[12] : 
                       (N114)? data_i[140] : 
                       (N116)? data_i[268] : 
                       (N118)? data_i[396] : 
                       (N113)? data_i[524] : 
                       (N115)? data_i[652] : 
                       (N117)? data_i[780] : 
                       (N119)? data_i[908] : 1'b0;
  assign data_o[907] = (N112)? data_i[11] : 
                       (N114)? data_i[139] : 
                       (N116)? data_i[267] : 
                       (N118)? data_i[395] : 
                       (N113)? data_i[523] : 
                       (N115)? data_i[651] : 
                       (N117)? data_i[779] : 
                       (N119)? data_i[907] : 1'b0;
  assign data_o[906] = (N112)? data_i[10] : 
                       (N114)? data_i[138] : 
                       (N116)? data_i[266] : 
                       (N118)? data_i[394] : 
                       (N113)? data_i[522] : 
                       (N115)? data_i[650] : 
                       (N117)? data_i[778] : 
                       (N119)? data_i[906] : 1'b0;
  assign data_o[905] = (N112)? data_i[9] : 
                       (N114)? data_i[137] : 
                       (N116)? data_i[265] : 
                       (N118)? data_i[393] : 
                       (N113)? data_i[521] : 
                       (N115)? data_i[649] : 
                       (N117)? data_i[777] : 
                       (N119)? data_i[905] : 1'b0;
  assign data_o[904] = (N112)? data_i[8] : 
                       (N114)? data_i[136] : 
                       (N116)? data_i[264] : 
                       (N118)? data_i[392] : 
                       (N113)? data_i[520] : 
                       (N115)? data_i[648] : 
                       (N117)? data_i[776] : 
                       (N119)? data_i[904] : 1'b0;
  assign data_o[903] = (N112)? data_i[7] : 
                       (N114)? data_i[135] : 
                       (N116)? data_i[263] : 
                       (N118)? data_i[391] : 
                       (N113)? data_i[519] : 
                       (N115)? data_i[647] : 
                       (N117)? data_i[775] : 
                       (N119)? data_i[903] : 1'b0;
  assign data_o[902] = (N112)? data_i[6] : 
                       (N114)? data_i[134] : 
                       (N116)? data_i[262] : 
                       (N118)? data_i[390] : 
                       (N113)? data_i[518] : 
                       (N115)? data_i[646] : 
                       (N117)? data_i[774] : 
                       (N119)? data_i[902] : 1'b0;
  assign data_o[901] = (N112)? data_i[5] : 
                       (N114)? data_i[133] : 
                       (N116)? data_i[261] : 
                       (N118)? data_i[389] : 
                       (N113)? data_i[517] : 
                       (N115)? data_i[645] : 
                       (N117)? data_i[773] : 
                       (N119)? data_i[901] : 1'b0;
  assign data_o[900] = (N112)? data_i[4] : 
                       (N114)? data_i[132] : 
                       (N116)? data_i[260] : 
                       (N118)? data_i[388] : 
                       (N113)? data_i[516] : 
                       (N115)? data_i[644] : 
                       (N117)? data_i[772] : 
                       (N119)? data_i[900] : 1'b0;
  assign data_o[899] = (N112)? data_i[3] : 
                       (N114)? data_i[131] : 
                       (N116)? data_i[259] : 
                       (N118)? data_i[387] : 
                       (N113)? data_i[515] : 
                       (N115)? data_i[643] : 
                       (N117)? data_i[771] : 
                       (N119)? data_i[899] : 1'b0;
  assign data_o[898] = (N112)? data_i[2] : 
                       (N114)? data_i[130] : 
                       (N116)? data_i[258] : 
                       (N118)? data_i[386] : 
                       (N113)? data_i[514] : 
                       (N115)? data_i[642] : 
                       (N117)? data_i[770] : 
                       (N119)? data_i[898] : 1'b0;
  assign data_o[897] = (N112)? data_i[1] : 
                       (N114)? data_i[129] : 
                       (N116)? data_i[257] : 
                       (N118)? data_i[385] : 
                       (N113)? data_i[513] : 
                       (N115)? data_i[641] : 
                       (N117)? data_i[769] : 
                       (N119)? data_i[897] : 1'b0;
  assign data_o[896] = (N112)? data_i[0] : 
                       (N114)? data_i[128] : 
                       (N116)? data_i[256] : 
                       (N118)? data_i[384] : 
                       (N113)? data_i[512] : 
                       (N115)? data_i[640] : 
                       (N117)? data_i[768] : 
                       (N119)? data_i[896] : 1'b0;
  assign N0 = ~select_i[0];
  assign N1 = ~select_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & select_i[1];
  assign N4 = select_i[0] & N1;
  assign N5 = select_i[0] & select_i[1];
  assign N6 = ~select_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & select_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & select_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & select_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & select_i[2];
  assign N15 = ~select_i[32];
  assign N16 = ~select_i[33];
  assign N17 = N15 & N16;
  assign N18 = N15 & select_i[33];
  assign N19 = select_i[32] & N16;
  assign N20 = select_i[32] & select_i[33];
  assign N21 = ~select_i[34];
  assign N22 = N17 & N21;
  assign N23 = N17 & select_i[34];
  assign N24 = N19 & N21;
  assign N25 = N19 & select_i[34];
  assign N26 = N18 & N21;
  assign N27 = N18 & select_i[34];
  assign N28 = N20 & N21;
  assign N29 = N20 & select_i[34];
  assign N30 = ~select_i[64];
  assign N31 = ~select_i[65];
  assign N32 = N30 & N31;
  assign N33 = N30 & select_i[65];
  assign N34 = select_i[64] & N31;
  assign N35 = select_i[64] & select_i[65];
  assign N36 = ~select_i[66];
  assign N37 = N32 & N36;
  assign N38 = N32 & select_i[66];
  assign N39 = N34 & N36;
  assign N40 = N34 & select_i[66];
  assign N41 = N33 & N36;
  assign N42 = N33 & select_i[66];
  assign N43 = N35 & N36;
  assign N44 = N35 & select_i[66];
  assign N45 = ~select_i[96];
  assign N46 = ~select_i[97];
  assign N47 = N45 & N46;
  assign N48 = N45 & select_i[97];
  assign N49 = select_i[96] & N46;
  assign N50 = select_i[96] & select_i[97];
  assign N51 = ~select_i[98];
  assign N52 = N47 & N51;
  assign N53 = N47 & select_i[98];
  assign N54 = N49 & N51;
  assign N55 = N49 & select_i[98];
  assign N56 = N48 & N51;
  assign N57 = N48 & select_i[98];
  assign N58 = N50 & N51;
  assign N59 = N50 & select_i[98];
  assign N60 = ~select_i[128];
  assign N61 = ~select_i[129];
  assign N62 = N60 & N61;
  assign N63 = N60 & select_i[129];
  assign N64 = select_i[128] & N61;
  assign N65 = select_i[128] & select_i[129];
  assign N66 = ~select_i[130];
  assign N67 = N62 & N66;
  assign N68 = N62 & select_i[130];
  assign N69 = N64 & N66;
  assign N70 = N64 & select_i[130];
  assign N71 = N63 & N66;
  assign N72 = N63 & select_i[130];
  assign N73 = N65 & N66;
  assign N74 = N65 & select_i[130];
  assign N75 = ~select_i[160];
  assign N76 = ~select_i[161];
  assign N77 = N75 & N76;
  assign N78 = N75 & select_i[161];
  assign N79 = select_i[160] & N76;
  assign N80 = select_i[160] & select_i[161];
  assign N81 = ~select_i[162];
  assign N82 = N77 & N81;
  assign N83 = N77 & select_i[162];
  assign N84 = N79 & N81;
  assign N85 = N79 & select_i[162];
  assign N86 = N78 & N81;
  assign N87 = N78 & select_i[162];
  assign N88 = N80 & N81;
  assign N89 = N80 & select_i[162];
  assign N90 = ~select_i[192];
  assign N91 = ~select_i[193];
  assign N92 = N90 & N91;
  assign N93 = N90 & select_i[193];
  assign N94 = select_i[192] & N91;
  assign N95 = select_i[192] & select_i[193];
  assign N96 = ~select_i[194];
  assign N97 = N92 & N96;
  assign N98 = N92 & select_i[194];
  assign N99 = N94 & N96;
  assign N100 = N94 & select_i[194];
  assign N101 = N93 & N96;
  assign N102 = N93 & select_i[194];
  assign N103 = N95 & N96;
  assign N104 = N95 & select_i[194];
  assign N105 = ~select_i[224];
  assign N106 = ~select_i[225];
  assign N107 = N105 & N106;
  assign N108 = N105 & select_i[225];
  assign N109 = select_i[224] & N106;
  assign N110 = select_i[224] & select_i[225];
  assign N111 = ~select_i[226];
  assign N112 = N107 & N111;
  assign N113 = N107 & select_i[226];
  assign N114 = N109 & N111;
  assign N115 = N109 & select_i[226];
  assign N116 = N108 & N111;
  assign N117 = N108 & select_i[226];
  assign N118 = N110 & N111;
  assign N119 = N110 & select_i[226];

endmodule

