

module top
(
  i,
  o
);

  input [16383:0] i;
  output [16383:0] o;

  bsg_array_reverse
  wrapper
  (
    .i(i),
    .o(o)
  );


endmodule



module bsg_array_reverse
(
  i,
  o
);

  input [16383:0] i;
  output [16383:0] o;
  wire [16383:0] o;
  assign o[16383] = i[127];
  assign o[16382] = i[126];
  assign o[16381] = i[125];
  assign o[16380] = i[124];
  assign o[16379] = i[123];
  assign o[16378] = i[122];
  assign o[16377] = i[121];
  assign o[16376] = i[120];
  assign o[16375] = i[119];
  assign o[16374] = i[118];
  assign o[16373] = i[117];
  assign o[16372] = i[116];
  assign o[16371] = i[115];
  assign o[16370] = i[114];
  assign o[16369] = i[113];
  assign o[16368] = i[112];
  assign o[16367] = i[111];
  assign o[16366] = i[110];
  assign o[16365] = i[109];
  assign o[16364] = i[108];
  assign o[16363] = i[107];
  assign o[16362] = i[106];
  assign o[16361] = i[105];
  assign o[16360] = i[104];
  assign o[16359] = i[103];
  assign o[16358] = i[102];
  assign o[16357] = i[101];
  assign o[16356] = i[100];
  assign o[16355] = i[99];
  assign o[16354] = i[98];
  assign o[16353] = i[97];
  assign o[16352] = i[96];
  assign o[16351] = i[95];
  assign o[16350] = i[94];
  assign o[16349] = i[93];
  assign o[16348] = i[92];
  assign o[16347] = i[91];
  assign o[16346] = i[90];
  assign o[16345] = i[89];
  assign o[16344] = i[88];
  assign o[16343] = i[87];
  assign o[16342] = i[86];
  assign o[16341] = i[85];
  assign o[16340] = i[84];
  assign o[16339] = i[83];
  assign o[16338] = i[82];
  assign o[16337] = i[81];
  assign o[16336] = i[80];
  assign o[16335] = i[79];
  assign o[16334] = i[78];
  assign o[16333] = i[77];
  assign o[16332] = i[76];
  assign o[16331] = i[75];
  assign o[16330] = i[74];
  assign o[16329] = i[73];
  assign o[16328] = i[72];
  assign o[16327] = i[71];
  assign o[16326] = i[70];
  assign o[16325] = i[69];
  assign o[16324] = i[68];
  assign o[16323] = i[67];
  assign o[16322] = i[66];
  assign o[16321] = i[65];
  assign o[16320] = i[64];
  assign o[16319] = i[63];
  assign o[16318] = i[62];
  assign o[16317] = i[61];
  assign o[16316] = i[60];
  assign o[16315] = i[59];
  assign o[16314] = i[58];
  assign o[16313] = i[57];
  assign o[16312] = i[56];
  assign o[16311] = i[55];
  assign o[16310] = i[54];
  assign o[16309] = i[53];
  assign o[16308] = i[52];
  assign o[16307] = i[51];
  assign o[16306] = i[50];
  assign o[16305] = i[49];
  assign o[16304] = i[48];
  assign o[16303] = i[47];
  assign o[16302] = i[46];
  assign o[16301] = i[45];
  assign o[16300] = i[44];
  assign o[16299] = i[43];
  assign o[16298] = i[42];
  assign o[16297] = i[41];
  assign o[16296] = i[40];
  assign o[16295] = i[39];
  assign o[16294] = i[38];
  assign o[16293] = i[37];
  assign o[16292] = i[36];
  assign o[16291] = i[35];
  assign o[16290] = i[34];
  assign o[16289] = i[33];
  assign o[16288] = i[32];
  assign o[16287] = i[31];
  assign o[16286] = i[30];
  assign o[16285] = i[29];
  assign o[16284] = i[28];
  assign o[16283] = i[27];
  assign o[16282] = i[26];
  assign o[16281] = i[25];
  assign o[16280] = i[24];
  assign o[16279] = i[23];
  assign o[16278] = i[22];
  assign o[16277] = i[21];
  assign o[16276] = i[20];
  assign o[16275] = i[19];
  assign o[16274] = i[18];
  assign o[16273] = i[17];
  assign o[16272] = i[16];
  assign o[16271] = i[15];
  assign o[16270] = i[14];
  assign o[16269] = i[13];
  assign o[16268] = i[12];
  assign o[16267] = i[11];
  assign o[16266] = i[10];
  assign o[16265] = i[9];
  assign o[16264] = i[8];
  assign o[16263] = i[7];
  assign o[16262] = i[6];
  assign o[16261] = i[5];
  assign o[16260] = i[4];
  assign o[16259] = i[3];
  assign o[16258] = i[2];
  assign o[16257] = i[1];
  assign o[16256] = i[0];
  assign o[16255] = i[255];
  assign o[16254] = i[254];
  assign o[16253] = i[253];
  assign o[16252] = i[252];
  assign o[16251] = i[251];
  assign o[16250] = i[250];
  assign o[16249] = i[249];
  assign o[16248] = i[248];
  assign o[16247] = i[247];
  assign o[16246] = i[246];
  assign o[16245] = i[245];
  assign o[16244] = i[244];
  assign o[16243] = i[243];
  assign o[16242] = i[242];
  assign o[16241] = i[241];
  assign o[16240] = i[240];
  assign o[16239] = i[239];
  assign o[16238] = i[238];
  assign o[16237] = i[237];
  assign o[16236] = i[236];
  assign o[16235] = i[235];
  assign o[16234] = i[234];
  assign o[16233] = i[233];
  assign o[16232] = i[232];
  assign o[16231] = i[231];
  assign o[16230] = i[230];
  assign o[16229] = i[229];
  assign o[16228] = i[228];
  assign o[16227] = i[227];
  assign o[16226] = i[226];
  assign o[16225] = i[225];
  assign o[16224] = i[224];
  assign o[16223] = i[223];
  assign o[16222] = i[222];
  assign o[16221] = i[221];
  assign o[16220] = i[220];
  assign o[16219] = i[219];
  assign o[16218] = i[218];
  assign o[16217] = i[217];
  assign o[16216] = i[216];
  assign o[16215] = i[215];
  assign o[16214] = i[214];
  assign o[16213] = i[213];
  assign o[16212] = i[212];
  assign o[16211] = i[211];
  assign o[16210] = i[210];
  assign o[16209] = i[209];
  assign o[16208] = i[208];
  assign o[16207] = i[207];
  assign o[16206] = i[206];
  assign o[16205] = i[205];
  assign o[16204] = i[204];
  assign o[16203] = i[203];
  assign o[16202] = i[202];
  assign o[16201] = i[201];
  assign o[16200] = i[200];
  assign o[16199] = i[199];
  assign o[16198] = i[198];
  assign o[16197] = i[197];
  assign o[16196] = i[196];
  assign o[16195] = i[195];
  assign o[16194] = i[194];
  assign o[16193] = i[193];
  assign o[16192] = i[192];
  assign o[16191] = i[191];
  assign o[16190] = i[190];
  assign o[16189] = i[189];
  assign o[16188] = i[188];
  assign o[16187] = i[187];
  assign o[16186] = i[186];
  assign o[16185] = i[185];
  assign o[16184] = i[184];
  assign o[16183] = i[183];
  assign o[16182] = i[182];
  assign o[16181] = i[181];
  assign o[16180] = i[180];
  assign o[16179] = i[179];
  assign o[16178] = i[178];
  assign o[16177] = i[177];
  assign o[16176] = i[176];
  assign o[16175] = i[175];
  assign o[16174] = i[174];
  assign o[16173] = i[173];
  assign o[16172] = i[172];
  assign o[16171] = i[171];
  assign o[16170] = i[170];
  assign o[16169] = i[169];
  assign o[16168] = i[168];
  assign o[16167] = i[167];
  assign o[16166] = i[166];
  assign o[16165] = i[165];
  assign o[16164] = i[164];
  assign o[16163] = i[163];
  assign o[16162] = i[162];
  assign o[16161] = i[161];
  assign o[16160] = i[160];
  assign o[16159] = i[159];
  assign o[16158] = i[158];
  assign o[16157] = i[157];
  assign o[16156] = i[156];
  assign o[16155] = i[155];
  assign o[16154] = i[154];
  assign o[16153] = i[153];
  assign o[16152] = i[152];
  assign o[16151] = i[151];
  assign o[16150] = i[150];
  assign o[16149] = i[149];
  assign o[16148] = i[148];
  assign o[16147] = i[147];
  assign o[16146] = i[146];
  assign o[16145] = i[145];
  assign o[16144] = i[144];
  assign o[16143] = i[143];
  assign o[16142] = i[142];
  assign o[16141] = i[141];
  assign o[16140] = i[140];
  assign o[16139] = i[139];
  assign o[16138] = i[138];
  assign o[16137] = i[137];
  assign o[16136] = i[136];
  assign o[16135] = i[135];
  assign o[16134] = i[134];
  assign o[16133] = i[133];
  assign o[16132] = i[132];
  assign o[16131] = i[131];
  assign o[16130] = i[130];
  assign o[16129] = i[129];
  assign o[16128] = i[128];
  assign o[16127] = i[383];
  assign o[16126] = i[382];
  assign o[16125] = i[381];
  assign o[16124] = i[380];
  assign o[16123] = i[379];
  assign o[16122] = i[378];
  assign o[16121] = i[377];
  assign o[16120] = i[376];
  assign o[16119] = i[375];
  assign o[16118] = i[374];
  assign o[16117] = i[373];
  assign o[16116] = i[372];
  assign o[16115] = i[371];
  assign o[16114] = i[370];
  assign o[16113] = i[369];
  assign o[16112] = i[368];
  assign o[16111] = i[367];
  assign o[16110] = i[366];
  assign o[16109] = i[365];
  assign o[16108] = i[364];
  assign o[16107] = i[363];
  assign o[16106] = i[362];
  assign o[16105] = i[361];
  assign o[16104] = i[360];
  assign o[16103] = i[359];
  assign o[16102] = i[358];
  assign o[16101] = i[357];
  assign o[16100] = i[356];
  assign o[16099] = i[355];
  assign o[16098] = i[354];
  assign o[16097] = i[353];
  assign o[16096] = i[352];
  assign o[16095] = i[351];
  assign o[16094] = i[350];
  assign o[16093] = i[349];
  assign o[16092] = i[348];
  assign o[16091] = i[347];
  assign o[16090] = i[346];
  assign o[16089] = i[345];
  assign o[16088] = i[344];
  assign o[16087] = i[343];
  assign o[16086] = i[342];
  assign o[16085] = i[341];
  assign o[16084] = i[340];
  assign o[16083] = i[339];
  assign o[16082] = i[338];
  assign o[16081] = i[337];
  assign o[16080] = i[336];
  assign o[16079] = i[335];
  assign o[16078] = i[334];
  assign o[16077] = i[333];
  assign o[16076] = i[332];
  assign o[16075] = i[331];
  assign o[16074] = i[330];
  assign o[16073] = i[329];
  assign o[16072] = i[328];
  assign o[16071] = i[327];
  assign o[16070] = i[326];
  assign o[16069] = i[325];
  assign o[16068] = i[324];
  assign o[16067] = i[323];
  assign o[16066] = i[322];
  assign o[16065] = i[321];
  assign o[16064] = i[320];
  assign o[16063] = i[319];
  assign o[16062] = i[318];
  assign o[16061] = i[317];
  assign o[16060] = i[316];
  assign o[16059] = i[315];
  assign o[16058] = i[314];
  assign o[16057] = i[313];
  assign o[16056] = i[312];
  assign o[16055] = i[311];
  assign o[16054] = i[310];
  assign o[16053] = i[309];
  assign o[16052] = i[308];
  assign o[16051] = i[307];
  assign o[16050] = i[306];
  assign o[16049] = i[305];
  assign o[16048] = i[304];
  assign o[16047] = i[303];
  assign o[16046] = i[302];
  assign o[16045] = i[301];
  assign o[16044] = i[300];
  assign o[16043] = i[299];
  assign o[16042] = i[298];
  assign o[16041] = i[297];
  assign o[16040] = i[296];
  assign o[16039] = i[295];
  assign o[16038] = i[294];
  assign o[16037] = i[293];
  assign o[16036] = i[292];
  assign o[16035] = i[291];
  assign o[16034] = i[290];
  assign o[16033] = i[289];
  assign o[16032] = i[288];
  assign o[16031] = i[287];
  assign o[16030] = i[286];
  assign o[16029] = i[285];
  assign o[16028] = i[284];
  assign o[16027] = i[283];
  assign o[16026] = i[282];
  assign o[16025] = i[281];
  assign o[16024] = i[280];
  assign o[16023] = i[279];
  assign o[16022] = i[278];
  assign o[16021] = i[277];
  assign o[16020] = i[276];
  assign o[16019] = i[275];
  assign o[16018] = i[274];
  assign o[16017] = i[273];
  assign o[16016] = i[272];
  assign o[16015] = i[271];
  assign o[16014] = i[270];
  assign o[16013] = i[269];
  assign o[16012] = i[268];
  assign o[16011] = i[267];
  assign o[16010] = i[266];
  assign o[16009] = i[265];
  assign o[16008] = i[264];
  assign o[16007] = i[263];
  assign o[16006] = i[262];
  assign o[16005] = i[261];
  assign o[16004] = i[260];
  assign o[16003] = i[259];
  assign o[16002] = i[258];
  assign o[16001] = i[257];
  assign o[16000] = i[256];
  assign o[15999] = i[511];
  assign o[15998] = i[510];
  assign o[15997] = i[509];
  assign o[15996] = i[508];
  assign o[15995] = i[507];
  assign o[15994] = i[506];
  assign o[15993] = i[505];
  assign o[15992] = i[504];
  assign o[15991] = i[503];
  assign o[15990] = i[502];
  assign o[15989] = i[501];
  assign o[15988] = i[500];
  assign o[15987] = i[499];
  assign o[15986] = i[498];
  assign o[15985] = i[497];
  assign o[15984] = i[496];
  assign o[15983] = i[495];
  assign o[15982] = i[494];
  assign o[15981] = i[493];
  assign o[15980] = i[492];
  assign o[15979] = i[491];
  assign o[15978] = i[490];
  assign o[15977] = i[489];
  assign o[15976] = i[488];
  assign o[15975] = i[487];
  assign o[15974] = i[486];
  assign o[15973] = i[485];
  assign o[15972] = i[484];
  assign o[15971] = i[483];
  assign o[15970] = i[482];
  assign o[15969] = i[481];
  assign o[15968] = i[480];
  assign o[15967] = i[479];
  assign o[15966] = i[478];
  assign o[15965] = i[477];
  assign o[15964] = i[476];
  assign o[15963] = i[475];
  assign o[15962] = i[474];
  assign o[15961] = i[473];
  assign o[15960] = i[472];
  assign o[15959] = i[471];
  assign o[15958] = i[470];
  assign o[15957] = i[469];
  assign o[15956] = i[468];
  assign o[15955] = i[467];
  assign o[15954] = i[466];
  assign o[15953] = i[465];
  assign o[15952] = i[464];
  assign o[15951] = i[463];
  assign o[15950] = i[462];
  assign o[15949] = i[461];
  assign o[15948] = i[460];
  assign o[15947] = i[459];
  assign o[15946] = i[458];
  assign o[15945] = i[457];
  assign o[15944] = i[456];
  assign o[15943] = i[455];
  assign o[15942] = i[454];
  assign o[15941] = i[453];
  assign o[15940] = i[452];
  assign o[15939] = i[451];
  assign o[15938] = i[450];
  assign o[15937] = i[449];
  assign o[15936] = i[448];
  assign o[15935] = i[447];
  assign o[15934] = i[446];
  assign o[15933] = i[445];
  assign o[15932] = i[444];
  assign o[15931] = i[443];
  assign o[15930] = i[442];
  assign o[15929] = i[441];
  assign o[15928] = i[440];
  assign o[15927] = i[439];
  assign o[15926] = i[438];
  assign o[15925] = i[437];
  assign o[15924] = i[436];
  assign o[15923] = i[435];
  assign o[15922] = i[434];
  assign o[15921] = i[433];
  assign o[15920] = i[432];
  assign o[15919] = i[431];
  assign o[15918] = i[430];
  assign o[15917] = i[429];
  assign o[15916] = i[428];
  assign o[15915] = i[427];
  assign o[15914] = i[426];
  assign o[15913] = i[425];
  assign o[15912] = i[424];
  assign o[15911] = i[423];
  assign o[15910] = i[422];
  assign o[15909] = i[421];
  assign o[15908] = i[420];
  assign o[15907] = i[419];
  assign o[15906] = i[418];
  assign o[15905] = i[417];
  assign o[15904] = i[416];
  assign o[15903] = i[415];
  assign o[15902] = i[414];
  assign o[15901] = i[413];
  assign o[15900] = i[412];
  assign o[15899] = i[411];
  assign o[15898] = i[410];
  assign o[15897] = i[409];
  assign o[15896] = i[408];
  assign o[15895] = i[407];
  assign o[15894] = i[406];
  assign o[15893] = i[405];
  assign o[15892] = i[404];
  assign o[15891] = i[403];
  assign o[15890] = i[402];
  assign o[15889] = i[401];
  assign o[15888] = i[400];
  assign o[15887] = i[399];
  assign o[15886] = i[398];
  assign o[15885] = i[397];
  assign o[15884] = i[396];
  assign o[15883] = i[395];
  assign o[15882] = i[394];
  assign o[15881] = i[393];
  assign o[15880] = i[392];
  assign o[15879] = i[391];
  assign o[15878] = i[390];
  assign o[15877] = i[389];
  assign o[15876] = i[388];
  assign o[15875] = i[387];
  assign o[15874] = i[386];
  assign o[15873] = i[385];
  assign o[15872] = i[384];
  assign o[15871] = i[639];
  assign o[15870] = i[638];
  assign o[15869] = i[637];
  assign o[15868] = i[636];
  assign o[15867] = i[635];
  assign o[15866] = i[634];
  assign o[15865] = i[633];
  assign o[15864] = i[632];
  assign o[15863] = i[631];
  assign o[15862] = i[630];
  assign o[15861] = i[629];
  assign o[15860] = i[628];
  assign o[15859] = i[627];
  assign o[15858] = i[626];
  assign o[15857] = i[625];
  assign o[15856] = i[624];
  assign o[15855] = i[623];
  assign o[15854] = i[622];
  assign o[15853] = i[621];
  assign o[15852] = i[620];
  assign o[15851] = i[619];
  assign o[15850] = i[618];
  assign o[15849] = i[617];
  assign o[15848] = i[616];
  assign o[15847] = i[615];
  assign o[15846] = i[614];
  assign o[15845] = i[613];
  assign o[15844] = i[612];
  assign o[15843] = i[611];
  assign o[15842] = i[610];
  assign o[15841] = i[609];
  assign o[15840] = i[608];
  assign o[15839] = i[607];
  assign o[15838] = i[606];
  assign o[15837] = i[605];
  assign o[15836] = i[604];
  assign o[15835] = i[603];
  assign o[15834] = i[602];
  assign o[15833] = i[601];
  assign o[15832] = i[600];
  assign o[15831] = i[599];
  assign o[15830] = i[598];
  assign o[15829] = i[597];
  assign o[15828] = i[596];
  assign o[15827] = i[595];
  assign o[15826] = i[594];
  assign o[15825] = i[593];
  assign o[15824] = i[592];
  assign o[15823] = i[591];
  assign o[15822] = i[590];
  assign o[15821] = i[589];
  assign o[15820] = i[588];
  assign o[15819] = i[587];
  assign o[15818] = i[586];
  assign o[15817] = i[585];
  assign o[15816] = i[584];
  assign o[15815] = i[583];
  assign o[15814] = i[582];
  assign o[15813] = i[581];
  assign o[15812] = i[580];
  assign o[15811] = i[579];
  assign o[15810] = i[578];
  assign o[15809] = i[577];
  assign o[15808] = i[576];
  assign o[15807] = i[575];
  assign o[15806] = i[574];
  assign o[15805] = i[573];
  assign o[15804] = i[572];
  assign o[15803] = i[571];
  assign o[15802] = i[570];
  assign o[15801] = i[569];
  assign o[15800] = i[568];
  assign o[15799] = i[567];
  assign o[15798] = i[566];
  assign o[15797] = i[565];
  assign o[15796] = i[564];
  assign o[15795] = i[563];
  assign o[15794] = i[562];
  assign o[15793] = i[561];
  assign o[15792] = i[560];
  assign o[15791] = i[559];
  assign o[15790] = i[558];
  assign o[15789] = i[557];
  assign o[15788] = i[556];
  assign o[15787] = i[555];
  assign o[15786] = i[554];
  assign o[15785] = i[553];
  assign o[15784] = i[552];
  assign o[15783] = i[551];
  assign o[15782] = i[550];
  assign o[15781] = i[549];
  assign o[15780] = i[548];
  assign o[15779] = i[547];
  assign o[15778] = i[546];
  assign o[15777] = i[545];
  assign o[15776] = i[544];
  assign o[15775] = i[543];
  assign o[15774] = i[542];
  assign o[15773] = i[541];
  assign o[15772] = i[540];
  assign o[15771] = i[539];
  assign o[15770] = i[538];
  assign o[15769] = i[537];
  assign o[15768] = i[536];
  assign o[15767] = i[535];
  assign o[15766] = i[534];
  assign o[15765] = i[533];
  assign o[15764] = i[532];
  assign o[15763] = i[531];
  assign o[15762] = i[530];
  assign o[15761] = i[529];
  assign o[15760] = i[528];
  assign o[15759] = i[527];
  assign o[15758] = i[526];
  assign o[15757] = i[525];
  assign o[15756] = i[524];
  assign o[15755] = i[523];
  assign o[15754] = i[522];
  assign o[15753] = i[521];
  assign o[15752] = i[520];
  assign o[15751] = i[519];
  assign o[15750] = i[518];
  assign o[15749] = i[517];
  assign o[15748] = i[516];
  assign o[15747] = i[515];
  assign o[15746] = i[514];
  assign o[15745] = i[513];
  assign o[15744] = i[512];
  assign o[15743] = i[767];
  assign o[15742] = i[766];
  assign o[15741] = i[765];
  assign o[15740] = i[764];
  assign o[15739] = i[763];
  assign o[15738] = i[762];
  assign o[15737] = i[761];
  assign o[15736] = i[760];
  assign o[15735] = i[759];
  assign o[15734] = i[758];
  assign o[15733] = i[757];
  assign o[15732] = i[756];
  assign o[15731] = i[755];
  assign o[15730] = i[754];
  assign o[15729] = i[753];
  assign o[15728] = i[752];
  assign o[15727] = i[751];
  assign o[15726] = i[750];
  assign o[15725] = i[749];
  assign o[15724] = i[748];
  assign o[15723] = i[747];
  assign o[15722] = i[746];
  assign o[15721] = i[745];
  assign o[15720] = i[744];
  assign o[15719] = i[743];
  assign o[15718] = i[742];
  assign o[15717] = i[741];
  assign o[15716] = i[740];
  assign o[15715] = i[739];
  assign o[15714] = i[738];
  assign o[15713] = i[737];
  assign o[15712] = i[736];
  assign o[15711] = i[735];
  assign o[15710] = i[734];
  assign o[15709] = i[733];
  assign o[15708] = i[732];
  assign o[15707] = i[731];
  assign o[15706] = i[730];
  assign o[15705] = i[729];
  assign o[15704] = i[728];
  assign o[15703] = i[727];
  assign o[15702] = i[726];
  assign o[15701] = i[725];
  assign o[15700] = i[724];
  assign o[15699] = i[723];
  assign o[15698] = i[722];
  assign o[15697] = i[721];
  assign o[15696] = i[720];
  assign o[15695] = i[719];
  assign o[15694] = i[718];
  assign o[15693] = i[717];
  assign o[15692] = i[716];
  assign o[15691] = i[715];
  assign o[15690] = i[714];
  assign o[15689] = i[713];
  assign o[15688] = i[712];
  assign o[15687] = i[711];
  assign o[15686] = i[710];
  assign o[15685] = i[709];
  assign o[15684] = i[708];
  assign o[15683] = i[707];
  assign o[15682] = i[706];
  assign o[15681] = i[705];
  assign o[15680] = i[704];
  assign o[15679] = i[703];
  assign o[15678] = i[702];
  assign o[15677] = i[701];
  assign o[15676] = i[700];
  assign o[15675] = i[699];
  assign o[15674] = i[698];
  assign o[15673] = i[697];
  assign o[15672] = i[696];
  assign o[15671] = i[695];
  assign o[15670] = i[694];
  assign o[15669] = i[693];
  assign o[15668] = i[692];
  assign o[15667] = i[691];
  assign o[15666] = i[690];
  assign o[15665] = i[689];
  assign o[15664] = i[688];
  assign o[15663] = i[687];
  assign o[15662] = i[686];
  assign o[15661] = i[685];
  assign o[15660] = i[684];
  assign o[15659] = i[683];
  assign o[15658] = i[682];
  assign o[15657] = i[681];
  assign o[15656] = i[680];
  assign o[15655] = i[679];
  assign o[15654] = i[678];
  assign o[15653] = i[677];
  assign o[15652] = i[676];
  assign o[15651] = i[675];
  assign o[15650] = i[674];
  assign o[15649] = i[673];
  assign o[15648] = i[672];
  assign o[15647] = i[671];
  assign o[15646] = i[670];
  assign o[15645] = i[669];
  assign o[15644] = i[668];
  assign o[15643] = i[667];
  assign o[15642] = i[666];
  assign o[15641] = i[665];
  assign o[15640] = i[664];
  assign o[15639] = i[663];
  assign o[15638] = i[662];
  assign o[15637] = i[661];
  assign o[15636] = i[660];
  assign o[15635] = i[659];
  assign o[15634] = i[658];
  assign o[15633] = i[657];
  assign o[15632] = i[656];
  assign o[15631] = i[655];
  assign o[15630] = i[654];
  assign o[15629] = i[653];
  assign o[15628] = i[652];
  assign o[15627] = i[651];
  assign o[15626] = i[650];
  assign o[15625] = i[649];
  assign o[15624] = i[648];
  assign o[15623] = i[647];
  assign o[15622] = i[646];
  assign o[15621] = i[645];
  assign o[15620] = i[644];
  assign o[15619] = i[643];
  assign o[15618] = i[642];
  assign o[15617] = i[641];
  assign o[15616] = i[640];
  assign o[15615] = i[895];
  assign o[15614] = i[894];
  assign o[15613] = i[893];
  assign o[15612] = i[892];
  assign o[15611] = i[891];
  assign o[15610] = i[890];
  assign o[15609] = i[889];
  assign o[15608] = i[888];
  assign o[15607] = i[887];
  assign o[15606] = i[886];
  assign o[15605] = i[885];
  assign o[15604] = i[884];
  assign o[15603] = i[883];
  assign o[15602] = i[882];
  assign o[15601] = i[881];
  assign o[15600] = i[880];
  assign o[15599] = i[879];
  assign o[15598] = i[878];
  assign o[15597] = i[877];
  assign o[15596] = i[876];
  assign o[15595] = i[875];
  assign o[15594] = i[874];
  assign o[15593] = i[873];
  assign o[15592] = i[872];
  assign o[15591] = i[871];
  assign o[15590] = i[870];
  assign o[15589] = i[869];
  assign o[15588] = i[868];
  assign o[15587] = i[867];
  assign o[15586] = i[866];
  assign o[15585] = i[865];
  assign o[15584] = i[864];
  assign o[15583] = i[863];
  assign o[15582] = i[862];
  assign o[15581] = i[861];
  assign o[15580] = i[860];
  assign o[15579] = i[859];
  assign o[15578] = i[858];
  assign o[15577] = i[857];
  assign o[15576] = i[856];
  assign o[15575] = i[855];
  assign o[15574] = i[854];
  assign o[15573] = i[853];
  assign o[15572] = i[852];
  assign o[15571] = i[851];
  assign o[15570] = i[850];
  assign o[15569] = i[849];
  assign o[15568] = i[848];
  assign o[15567] = i[847];
  assign o[15566] = i[846];
  assign o[15565] = i[845];
  assign o[15564] = i[844];
  assign o[15563] = i[843];
  assign o[15562] = i[842];
  assign o[15561] = i[841];
  assign o[15560] = i[840];
  assign o[15559] = i[839];
  assign o[15558] = i[838];
  assign o[15557] = i[837];
  assign o[15556] = i[836];
  assign o[15555] = i[835];
  assign o[15554] = i[834];
  assign o[15553] = i[833];
  assign o[15552] = i[832];
  assign o[15551] = i[831];
  assign o[15550] = i[830];
  assign o[15549] = i[829];
  assign o[15548] = i[828];
  assign o[15547] = i[827];
  assign o[15546] = i[826];
  assign o[15545] = i[825];
  assign o[15544] = i[824];
  assign o[15543] = i[823];
  assign o[15542] = i[822];
  assign o[15541] = i[821];
  assign o[15540] = i[820];
  assign o[15539] = i[819];
  assign o[15538] = i[818];
  assign o[15537] = i[817];
  assign o[15536] = i[816];
  assign o[15535] = i[815];
  assign o[15534] = i[814];
  assign o[15533] = i[813];
  assign o[15532] = i[812];
  assign o[15531] = i[811];
  assign o[15530] = i[810];
  assign o[15529] = i[809];
  assign o[15528] = i[808];
  assign o[15527] = i[807];
  assign o[15526] = i[806];
  assign o[15525] = i[805];
  assign o[15524] = i[804];
  assign o[15523] = i[803];
  assign o[15522] = i[802];
  assign o[15521] = i[801];
  assign o[15520] = i[800];
  assign o[15519] = i[799];
  assign o[15518] = i[798];
  assign o[15517] = i[797];
  assign o[15516] = i[796];
  assign o[15515] = i[795];
  assign o[15514] = i[794];
  assign o[15513] = i[793];
  assign o[15512] = i[792];
  assign o[15511] = i[791];
  assign o[15510] = i[790];
  assign o[15509] = i[789];
  assign o[15508] = i[788];
  assign o[15507] = i[787];
  assign o[15506] = i[786];
  assign o[15505] = i[785];
  assign o[15504] = i[784];
  assign o[15503] = i[783];
  assign o[15502] = i[782];
  assign o[15501] = i[781];
  assign o[15500] = i[780];
  assign o[15499] = i[779];
  assign o[15498] = i[778];
  assign o[15497] = i[777];
  assign o[15496] = i[776];
  assign o[15495] = i[775];
  assign o[15494] = i[774];
  assign o[15493] = i[773];
  assign o[15492] = i[772];
  assign o[15491] = i[771];
  assign o[15490] = i[770];
  assign o[15489] = i[769];
  assign o[15488] = i[768];
  assign o[15487] = i[1023];
  assign o[15486] = i[1022];
  assign o[15485] = i[1021];
  assign o[15484] = i[1020];
  assign o[15483] = i[1019];
  assign o[15482] = i[1018];
  assign o[15481] = i[1017];
  assign o[15480] = i[1016];
  assign o[15479] = i[1015];
  assign o[15478] = i[1014];
  assign o[15477] = i[1013];
  assign o[15476] = i[1012];
  assign o[15475] = i[1011];
  assign o[15474] = i[1010];
  assign o[15473] = i[1009];
  assign o[15472] = i[1008];
  assign o[15471] = i[1007];
  assign o[15470] = i[1006];
  assign o[15469] = i[1005];
  assign o[15468] = i[1004];
  assign o[15467] = i[1003];
  assign o[15466] = i[1002];
  assign o[15465] = i[1001];
  assign o[15464] = i[1000];
  assign o[15463] = i[999];
  assign o[15462] = i[998];
  assign o[15461] = i[997];
  assign o[15460] = i[996];
  assign o[15459] = i[995];
  assign o[15458] = i[994];
  assign o[15457] = i[993];
  assign o[15456] = i[992];
  assign o[15455] = i[991];
  assign o[15454] = i[990];
  assign o[15453] = i[989];
  assign o[15452] = i[988];
  assign o[15451] = i[987];
  assign o[15450] = i[986];
  assign o[15449] = i[985];
  assign o[15448] = i[984];
  assign o[15447] = i[983];
  assign o[15446] = i[982];
  assign o[15445] = i[981];
  assign o[15444] = i[980];
  assign o[15443] = i[979];
  assign o[15442] = i[978];
  assign o[15441] = i[977];
  assign o[15440] = i[976];
  assign o[15439] = i[975];
  assign o[15438] = i[974];
  assign o[15437] = i[973];
  assign o[15436] = i[972];
  assign o[15435] = i[971];
  assign o[15434] = i[970];
  assign o[15433] = i[969];
  assign o[15432] = i[968];
  assign o[15431] = i[967];
  assign o[15430] = i[966];
  assign o[15429] = i[965];
  assign o[15428] = i[964];
  assign o[15427] = i[963];
  assign o[15426] = i[962];
  assign o[15425] = i[961];
  assign o[15424] = i[960];
  assign o[15423] = i[959];
  assign o[15422] = i[958];
  assign o[15421] = i[957];
  assign o[15420] = i[956];
  assign o[15419] = i[955];
  assign o[15418] = i[954];
  assign o[15417] = i[953];
  assign o[15416] = i[952];
  assign o[15415] = i[951];
  assign o[15414] = i[950];
  assign o[15413] = i[949];
  assign o[15412] = i[948];
  assign o[15411] = i[947];
  assign o[15410] = i[946];
  assign o[15409] = i[945];
  assign o[15408] = i[944];
  assign o[15407] = i[943];
  assign o[15406] = i[942];
  assign o[15405] = i[941];
  assign o[15404] = i[940];
  assign o[15403] = i[939];
  assign o[15402] = i[938];
  assign o[15401] = i[937];
  assign o[15400] = i[936];
  assign o[15399] = i[935];
  assign o[15398] = i[934];
  assign o[15397] = i[933];
  assign o[15396] = i[932];
  assign o[15395] = i[931];
  assign o[15394] = i[930];
  assign o[15393] = i[929];
  assign o[15392] = i[928];
  assign o[15391] = i[927];
  assign o[15390] = i[926];
  assign o[15389] = i[925];
  assign o[15388] = i[924];
  assign o[15387] = i[923];
  assign o[15386] = i[922];
  assign o[15385] = i[921];
  assign o[15384] = i[920];
  assign o[15383] = i[919];
  assign o[15382] = i[918];
  assign o[15381] = i[917];
  assign o[15380] = i[916];
  assign o[15379] = i[915];
  assign o[15378] = i[914];
  assign o[15377] = i[913];
  assign o[15376] = i[912];
  assign o[15375] = i[911];
  assign o[15374] = i[910];
  assign o[15373] = i[909];
  assign o[15372] = i[908];
  assign o[15371] = i[907];
  assign o[15370] = i[906];
  assign o[15369] = i[905];
  assign o[15368] = i[904];
  assign o[15367] = i[903];
  assign o[15366] = i[902];
  assign o[15365] = i[901];
  assign o[15364] = i[900];
  assign o[15363] = i[899];
  assign o[15362] = i[898];
  assign o[15361] = i[897];
  assign o[15360] = i[896];
  assign o[15359] = i[1151];
  assign o[15358] = i[1150];
  assign o[15357] = i[1149];
  assign o[15356] = i[1148];
  assign o[15355] = i[1147];
  assign o[15354] = i[1146];
  assign o[15353] = i[1145];
  assign o[15352] = i[1144];
  assign o[15351] = i[1143];
  assign o[15350] = i[1142];
  assign o[15349] = i[1141];
  assign o[15348] = i[1140];
  assign o[15347] = i[1139];
  assign o[15346] = i[1138];
  assign o[15345] = i[1137];
  assign o[15344] = i[1136];
  assign o[15343] = i[1135];
  assign o[15342] = i[1134];
  assign o[15341] = i[1133];
  assign o[15340] = i[1132];
  assign o[15339] = i[1131];
  assign o[15338] = i[1130];
  assign o[15337] = i[1129];
  assign o[15336] = i[1128];
  assign o[15335] = i[1127];
  assign o[15334] = i[1126];
  assign o[15333] = i[1125];
  assign o[15332] = i[1124];
  assign o[15331] = i[1123];
  assign o[15330] = i[1122];
  assign o[15329] = i[1121];
  assign o[15328] = i[1120];
  assign o[15327] = i[1119];
  assign o[15326] = i[1118];
  assign o[15325] = i[1117];
  assign o[15324] = i[1116];
  assign o[15323] = i[1115];
  assign o[15322] = i[1114];
  assign o[15321] = i[1113];
  assign o[15320] = i[1112];
  assign o[15319] = i[1111];
  assign o[15318] = i[1110];
  assign o[15317] = i[1109];
  assign o[15316] = i[1108];
  assign o[15315] = i[1107];
  assign o[15314] = i[1106];
  assign o[15313] = i[1105];
  assign o[15312] = i[1104];
  assign o[15311] = i[1103];
  assign o[15310] = i[1102];
  assign o[15309] = i[1101];
  assign o[15308] = i[1100];
  assign o[15307] = i[1099];
  assign o[15306] = i[1098];
  assign o[15305] = i[1097];
  assign o[15304] = i[1096];
  assign o[15303] = i[1095];
  assign o[15302] = i[1094];
  assign o[15301] = i[1093];
  assign o[15300] = i[1092];
  assign o[15299] = i[1091];
  assign o[15298] = i[1090];
  assign o[15297] = i[1089];
  assign o[15296] = i[1088];
  assign o[15295] = i[1087];
  assign o[15294] = i[1086];
  assign o[15293] = i[1085];
  assign o[15292] = i[1084];
  assign o[15291] = i[1083];
  assign o[15290] = i[1082];
  assign o[15289] = i[1081];
  assign o[15288] = i[1080];
  assign o[15287] = i[1079];
  assign o[15286] = i[1078];
  assign o[15285] = i[1077];
  assign o[15284] = i[1076];
  assign o[15283] = i[1075];
  assign o[15282] = i[1074];
  assign o[15281] = i[1073];
  assign o[15280] = i[1072];
  assign o[15279] = i[1071];
  assign o[15278] = i[1070];
  assign o[15277] = i[1069];
  assign o[15276] = i[1068];
  assign o[15275] = i[1067];
  assign o[15274] = i[1066];
  assign o[15273] = i[1065];
  assign o[15272] = i[1064];
  assign o[15271] = i[1063];
  assign o[15270] = i[1062];
  assign o[15269] = i[1061];
  assign o[15268] = i[1060];
  assign o[15267] = i[1059];
  assign o[15266] = i[1058];
  assign o[15265] = i[1057];
  assign o[15264] = i[1056];
  assign o[15263] = i[1055];
  assign o[15262] = i[1054];
  assign o[15261] = i[1053];
  assign o[15260] = i[1052];
  assign o[15259] = i[1051];
  assign o[15258] = i[1050];
  assign o[15257] = i[1049];
  assign o[15256] = i[1048];
  assign o[15255] = i[1047];
  assign o[15254] = i[1046];
  assign o[15253] = i[1045];
  assign o[15252] = i[1044];
  assign o[15251] = i[1043];
  assign o[15250] = i[1042];
  assign o[15249] = i[1041];
  assign o[15248] = i[1040];
  assign o[15247] = i[1039];
  assign o[15246] = i[1038];
  assign o[15245] = i[1037];
  assign o[15244] = i[1036];
  assign o[15243] = i[1035];
  assign o[15242] = i[1034];
  assign o[15241] = i[1033];
  assign o[15240] = i[1032];
  assign o[15239] = i[1031];
  assign o[15238] = i[1030];
  assign o[15237] = i[1029];
  assign o[15236] = i[1028];
  assign o[15235] = i[1027];
  assign o[15234] = i[1026];
  assign o[15233] = i[1025];
  assign o[15232] = i[1024];
  assign o[15231] = i[1279];
  assign o[15230] = i[1278];
  assign o[15229] = i[1277];
  assign o[15228] = i[1276];
  assign o[15227] = i[1275];
  assign o[15226] = i[1274];
  assign o[15225] = i[1273];
  assign o[15224] = i[1272];
  assign o[15223] = i[1271];
  assign o[15222] = i[1270];
  assign o[15221] = i[1269];
  assign o[15220] = i[1268];
  assign o[15219] = i[1267];
  assign o[15218] = i[1266];
  assign o[15217] = i[1265];
  assign o[15216] = i[1264];
  assign o[15215] = i[1263];
  assign o[15214] = i[1262];
  assign o[15213] = i[1261];
  assign o[15212] = i[1260];
  assign o[15211] = i[1259];
  assign o[15210] = i[1258];
  assign o[15209] = i[1257];
  assign o[15208] = i[1256];
  assign o[15207] = i[1255];
  assign o[15206] = i[1254];
  assign o[15205] = i[1253];
  assign o[15204] = i[1252];
  assign o[15203] = i[1251];
  assign o[15202] = i[1250];
  assign o[15201] = i[1249];
  assign o[15200] = i[1248];
  assign o[15199] = i[1247];
  assign o[15198] = i[1246];
  assign o[15197] = i[1245];
  assign o[15196] = i[1244];
  assign o[15195] = i[1243];
  assign o[15194] = i[1242];
  assign o[15193] = i[1241];
  assign o[15192] = i[1240];
  assign o[15191] = i[1239];
  assign o[15190] = i[1238];
  assign o[15189] = i[1237];
  assign o[15188] = i[1236];
  assign o[15187] = i[1235];
  assign o[15186] = i[1234];
  assign o[15185] = i[1233];
  assign o[15184] = i[1232];
  assign o[15183] = i[1231];
  assign o[15182] = i[1230];
  assign o[15181] = i[1229];
  assign o[15180] = i[1228];
  assign o[15179] = i[1227];
  assign o[15178] = i[1226];
  assign o[15177] = i[1225];
  assign o[15176] = i[1224];
  assign o[15175] = i[1223];
  assign o[15174] = i[1222];
  assign o[15173] = i[1221];
  assign o[15172] = i[1220];
  assign o[15171] = i[1219];
  assign o[15170] = i[1218];
  assign o[15169] = i[1217];
  assign o[15168] = i[1216];
  assign o[15167] = i[1215];
  assign o[15166] = i[1214];
  assign o[15165] = i[1213];
  assign o[15164] = i[1212];
  assign o[15163] = i[1211];
  assign o[15162] = i[1210];
  assign o[15161] = i[1209];
  assign o[15160] = i[1208];
  assign o[15159] = i[1207];
  assign o[15158] = i[1206];
  assign o[15157] = i[1205];
  assign o[15156] = i[1204];
  assign o[15155] = i[1203];
  assign o[15154] = i[1202];
  assign o[15153] = i[1201];
  assign o[15152] = i[1200];
  assign o[15151] = i[1199];
  assign o[15150] = i[1198];
  assign o[15149] = i[1197];
  assign o[15148] = i[1196];
  assign o[15147] = i[1195];
  assign o[15146] = i[1194];
  assign o[15145] = i[1193];
  assign o[15144] = i[1192];
  assign o[15143] = i[1191];
  assign o[15142] = i[1190];
  assign o[15141] = i[1189];
  assign o[15140] = i[1188];
  assign o[15139] = i[1187];
  assign o[15138] = i[1186];
  assign o[15137] = i[1185];
  assign o[15136] = i[1184];
  assign o[15135] = i[1183];
  assign o[15134] = i[1182];
  assign o[15133] = i[1181];
  assign o[15132] = i[1180];
  assign o[15131] = i[1179];
  assign o[15130] = i[1178];
  assign o[15129] = i[1177];
  assign o[15128] = i[1176];
  assign o[15127] = i[1175];
  assign o[15126] = i[1174];
  assign o[15125] = i[1173];
  assign o[15124] = i[1172];
  assign o[15123] = i[1171];
  assign o[15122] = i[1170];
  assign o[15121] = i[1169];
  assign o[15120] = i[1168];
  assign o[15119] = i[1167];
  assign o[15118] = i[1166];
  assign o[15117] = i[1165];
  assign o[15116] = i[1164];
  assign o[15115] = i[1163];
  assign o[15114] = i[1162];
  assign o[15113] = i[1161];
  assign o[15112] = i[1160];
  assign o[15111] = i[1159];
  assign o[15110] = i[1158];
  assign o[15109] = i[1157];
  assign o[15108] = i[1156];
  assign o[15107] = i[1155];
  assign o[15106] = i[1154];
  assign o[15105] = i[1153];
  assign o[15104] = i[1152];
  assign o[15103] = i[1407];
  assign o[15102] = i[1406];
  assign o[15101] = i[1405];
  assign o[15100] = i[1404];
  assign o[15099] = i[1403];
  assign o[15098] = i[1402];
  assign o[15097] = i[1401];
  assign o[15096] = i[1400];
  assign o[15095] = i[1399];
  assign o[15094] = i[1398];
  assign o[15093] = i[1397];
  assign o[15092] = i[1396];
  assign o[15091] = i[1395];
  assign o[15090] = i[1394];
  assign o[15089] = i[1393];
  assign o[15088] = i[1392];
  assign o[15087] = i[1391];
  assign o[15086] = i[1390];
  assign o[15085] = i[1389];
  assign o[15084] = i[1388];
  assign o[15083] = i[1387];
  assign o[15082] = i[1386];
  assign o[15081] = i[1385];
  assign o[15080] = i[1384];
  assign o[15079] = i[1383];
  assign o[15078] = i[1382];
  assign o[15077] = i[1381];
  assign o[15076] = i[1380];
  assign o[15075] = i[1379];
  assign o[15074] = i[1378];
  assign o[15073] = i[1377];
  assign o[15072] = i[1376];
  assign o[15071] = i[1375];
  assign o[15070] = i[1374];
  assign o[15069] = i[1373];
  assign o[15068] = i[1372];
  assign o[15067] = i[1371];
  assign o[15066] = i[1370];
  assign o[15065] = i[1369];
  assign o[15064] = i[1368];
  assign o[15063] = i[1367];
  assign o[15062] = i[1366];
  assign o[15061] = i[1365];
  assign o[15060] = i[1364];
  assign o[15059] = i[1363];
  assign o[15058] = i[1362];
  assign o[15057] = i[1361];
  assign o[15056] = i[1360];
  assign o[15055] = i[1359];
  assign o[15054] = i[1358];
  assign o[15053] = i[1357];
  assign o[15052] = i[1356];
  assign o[15051] = i[1355];
  assign o[15050] = i[1354];
  assign o[15049] = i[1353];
  assign o[15048] = i[1352];
  assign o[15047] = i[1351];
  assign o[15046] = i[1350];
  assign o[15045] = i[1349];
  assign o[15044] = i[1348];
  assign o[15043] = i[1347];
  assign o[15042] = i[1346];
  assign o[15041] = i[1345];
  assign o[15040] = i[1344];
  assign o[15039] = i[1343];
  assign o[15038] = i[1342];
  assign o[15037] = i[1341];
  assign o[15036] = i[1340];
  assign o[15035] = i[1339];
  assign o[15034] = i[1338];
  assign o[15033] = i[1337];
  assign o[15032] = i[1336];
  assign o[15031] = i[1335];
  assign o[15030] = i[1334];
  assign o[15029] = i[1333];
  assign o[15028] = i[1332];
  assign o[15027] = i[1331];
  assign o[15026] = i[1330];
  assign o[15025] = i[1329];
  assign o[15024] = i[1328];
  assign o[15023] = i[1327];
  assign o[15022] = i[1326];
  assign o[15021] = i[1325];
  assign o[15020] = i[1324];
  assign o[15019] = i[1323];
  assign o[15018] = i[1322];
  assign o[15017] = i[1321];
  assign o[15016] = i[1320];
  assign o[15015] = i[1319];
  assign o[15014] = i[1318];
  assign o[15013] = i[1317];
  assign o[15012] = i[1316];
  assign o[15011] = i[1315];
  assign o[15010] = i[1314];
  assign o[15009] = i[1313];
  assign o[15008] = i[1312];
  assign o[15007] = i[1311];
  assign o[15006] = i[1310];
  assign o[15005] = i[1309];
  assign o[15004] = i[1308];
  assign o[15003] = i[1307];
  assign o[15002] = i[1306];
  assign o[15001] = i[1305];
  assign o[15000] = i[1304];
  assign o[14999] = i[1303];
  assign o[14998] = i[1302];
  assign o[14997] = i[1301];
  assign o[14996] = i[1300];
  assign o[14995] = i[1299];
  assign o[14994] = i[1298];
  assign o[14993] = i[1297];
  assign o[14992] = i[1296];
  assign o[14991] = i[1295];
  assign o[14990] = i[1294];
  assign o[14989] = i[1293];
  assign o[14988] = i[1292];
  assign o[14987] = i[1291];
  assign o[14986] = i[1290];
  assign o[14985] = i[1289];
  assign o[14984] = i[1288];
  assign o[14983] = i[1287];
  assign o[14982] = i[1286];
  assign o[14981] = i[1285];
  assign o[14980] = i[1284];
  assign o[14979] = i[1283];
  assign o[14978] = i[1282];
  assign o[14977] = i[1281];
  assign o[14976] = i[1280];
  assign o[14975] = i[1535];
  assign o[14974] = i[1534];
  assign o[14973] = i[1533];
  assign o[14972] = i[1532];
  assign o[14971] = i[1531];
  assign o[14970] = i[1530];
  assign o[14969] = i[1529];
  assign o[14968] = i[1528];
  assign o[14967] = i[1527];
  assign o[14966] = i[1526];
  assign o[14965] = i[1525];
  assign o[14964] = i[1524];
  assign o[14963] = i[1523];
  assign o[14962] = i[1522];
  assign o[14961] = i[1521];
  assign o[14960] = i[1520];
  assign o[14959] = i[1519];
  assign o[14958] = i[1518];
  assign o[14957] = i[1517];
  assign o[14956] = i[1516];
  assign o[14955] = i[1515];
  assign o[14954] = i[1514];
  assign o[14953] = i[1513];
  assign o[14952] = i[1512];
  assign o[14951] = i[1511];
  assign o[14950] = i[1510];
  assign o[14949] = i[1509];
  assign o[14948] = i[1508];
  assign o[14947] = i[1507];
  assign o[14946] = i[1506];
  assign o[14945] = i[1505];
  assign o[14944] = i[1504];
  assign o[14943] = i[1503];
  assign o[14942] = i[1502];
  assign o[14941] = i[1501];
  assign o[14940] = i[1500];
  assign o[14939] = i[1499];
  assign o[14938] = i[1498];
  assign o[14937] = i[1497];
  assign o[14936] = i[1496];
  assign o[14935] = i[1495];
  assign o[14934] = i[1494];
  assign o[14933] = i[1493];
  assign o[14932] = i[1492];
  assign o[14931] = i[1491];
  assign o[14930] = i[1490];
  assign o[14929] = i[1489];
  assign o[14928] = i[1488];
  assign o[14927] = i[1487];
  assign o[14926] = i[1486];
  assign o[14925] = i[1485];
  assign o[14924] = i[1484];
  assign o[14923] = i[1483];
  assign o[14922] = i[1482];
  assign o[14921] = i[1481];
  assign o[14920] = i[1480];
  assign o[14919] = i[1479];
  assign o[14918] = i[1478];
  assign o[14917] = i[1477];
  assign o[14916] = i[1476];
  assign o[14915] = i[1475];
  assign o[14914] = i[1474];
  assign o[14913] = i[1473];
  assign o[14912] = i[1472];
  assign o[14911] = i[1471];
  assign o[14910] = i[1470];
  assign o[14909] = i[1469];
  assign o[14908] = i[1468];
  assign o[14907] = i[1467];
  assign o[14906] = i[1466];
  assign o[14905] = i[1465];
  assign o[14904] = i[1464];
  assign o[14903] = i[1463];
  assign o[14902] = i[1462];
  assign o[14901] = i[1461];
  assign o[14900] = i[1460];
  assign o[14899] = i[1459];
  assign o[14898] = i[1458];
  assign o[14897] = i[1457];
  assign o[14896] = i[1456];
  assign o[14895] = i[1455];
  assign o[14894] = i[1454];
  assign o[14893] = i[1453];
  assign o[14892] = i[1452];
  assign o[14891] = i[1451];
  assign o[14890] = i[1450];
  assign o[14889] = i[1449];
  assign o[14888] = i[1448];
  assign o[14887] = i[1447];
  assign o[14886] = i[1446];
  assign o[14885] = i[1445];
  assign o[14884] = i[1444];
  assign o[14883] = i[1443];
  assign o[14882] = i[1442];
  assign o[14881] = i[1441];
  assign o[14880] = i[1440];
  assign o[14879] = i[1439];
  assign o[14878] = i[1438];
  assign o[14877] = i[1437];
  assign o[14876] = i[1436];
  assign o[14875] = i[1435];
  assign o[14874] = i[1434];
  assign o[14873] = i[1433];
  assign o[14872] = i[1432];
  assign o[14871] = i[1431];
  assign o[14870] = i[1430];
  assign o[14869] = i[1429];
  assign o[14868] = i[1428];
  assign o[14867] = i[1427];
  assign o[14866] = i[1426];
  assign o[14865] = i[1425];
  assign o[14864] = i[1424];
  assign o[14863] = i[1423];
  assign o[14862] = i[1422];
  assign o[14861] = i[1421];
  assign o[14860] = i[1420];
  assign o[14859] = i[1419];
  assign o[14858] = i[1418];
  assign o[14857] = i[1417];
  assign o[14856] = i[1416];
  assign o[14855] = i[1415];
  assign o[14854] = i[1414];
  assign o[14853] = i[1413];
  assign o[14852] = i[1412];
  assign o[14851] = i[1411];
  assign o[14850] = i[1410];
  assign o[14849] = i[1409];
  assign o[14848] = i[1408];
  assign o[14847] = i[1663];
  assign o[14846] = i[1662];
  assign o[14845] = i[1661];
  assign o[14844] = i[1660];
  assign o[14843] = i[1659];
  assign o[14842] = i[1658];
  assign o[14841] = i[1657];
  assign o[14840] = i[1656];
  assign o[14839] = i[1655];
  assign o[14838] = i[1654];
  assign o[14837] = i[1653];
  assign o[14836] = i[1652];
  assign o[14835] = i[1651];
  assign o[14834] = i[1650];
  assign o[14833] = i[1649];
  assign o[14832] = i[1648];
  assign o[14831] = i[1647];
  assign o[14830] = i[1646];
  assign o[14829] = i[1645];
  assign o[14828] = i[1644];
  assign o[14827] = i[1643];
  assign o[14826] = i[1642];
  assign o[14825] = i[1641];
  assign o[14824] = i[1640];
  assign o[14823] = i[1639];
  assign o[14822] = i[1638];
  assign o[14821] = i[1637];
  assign o[14820] = i[1636];
  assign o[14819] = i[1635];
  assign o[14818] = i[1634];
  assign o[14817] = i[1633];
  assign o[14816] = i[1632];
  assign o[14815] = i[1631];
  assign o[14814] = i[1630];
  assign o[14813] = i[1629];
  assign o[14812] = i[1628];
  assign o[14811] = i[1627];
  assign o[14810] = i[1626];
  assign o[14809] = i[1625];
  assign o[14808] = i[1624];
  assign o[14807] = i[1623];
  assign o[14806] = i[1622];
  assign o[14805] = i[1621];
  assign o[14804] = i[1620];
  assign o[14803] = i[1619];
  assign o[14802] = i[1618];
  assign o[14801] = i[1617];
  assign o[14800] = i[1616];
  assign o[14799] = i[1615];
  assign o[14798] = i[1614];
  assign o[14797] = i[1613];
  assign o[14796] = i[1612];
  assign o[14795] = i[1611];
  assign o[14794] = i[1610];
  assign o[14793] = i[1609];
  assign o[14792] = i[1608];
  assign o[14791] = i[1607];
  assign o[14790] = i[1606];
  assign o[14789] = i[1605];
  assign o[14788] = i[1604];
  assign o[14787] = i[1603];
  assign o[14786] = i[1602];
  assign o[14785] = i[1601];
  assign o[14784] = i[1600];
  assign o[14783] = i[1599];
  assign o[14782] = i[1598];
  assign o[14781] = i[1597];
  assign o[14780] = i[1596];
  assign o[14779] = i[1595];
  assign o[14778] = i[1594];
  assign o[14777] = i[1593];
  assign o[14776] = i[1592];
  assign o[14775] = i[1591];
  assign o[14774] = i[1590];
  assign o[14773] = i[1589];
  assign o[14772] = i[1588];
  assign o[14771] = i[1587];
  assign o[14770] = i[1586];
  assign o[14769] = i[1585];
  assign o[14768] = i[1584];
  assign o[14767] = i[1583];
  assign o[14766] = i[1582];
  assign o[14765] = i[1581];
  assign o[14764] = i[1580];
  assign o[14763] = i[1579];
  assign o[14762] = i[1578];
  assign o[14761] = i[1577];
  assign o[14760] = i[1576];
  assign o[14759] = i[1575];
  assign o[14758] = i[1574];
  assign o[14757] = i[1573];
  assign o[14756] = i[1572];
  assign o[14755] = i[1571];
  assign o[14754] = i[1570];
  assign o[14753] = i[1569];
  assign o[14752] = i[1568];
  assign o[14751] = i[1567];
  assign o[14750] = i[1566];
  assign o[14749] = i[1565];
  assign o[14748] = i[1564];
  assign o[14747] = i[1563];
  assign o[14746] = i[1562];
  assign o[14745] = i[1561];
  assign o[14744] = i[1560];
  assign o[14743] = i[1559];
  assign o[14742] = i[1558];
  assign o[14741] = i[1557];
  assign o[14740] = i[1556];
  assign o[14739] = i[1555];
  assign o[14738] = i[1554];
  assign o[14737] = i[1553];
  assign o[14736] = i[1552];
  assign o[14735] = i[1551];
  assign o[14734] = i[1550];
  assign o[14733] = i[1549];
  assign o[14732] = i[1548];
  assign o[14731] = i[1547];
  assign o[14730] = i[1546];
  assign o[14729] = i[1545];
  assign o[14728] = i[1544];
  assign o[14727] = i[1543];
  assign o[14726] = i[1542];
  assign o[14725] = i[1541];
  assign o[14724] = i[1540];
  assign o[14723] = i[1539];
  assign o[14722] = i[1538];
  assign o[14721] = i[1537];
  assign o[14720] = i[1536];
  assign o[14719] = i[1791];
  assign o[14718] = i[1790];
  assign o[14717] = i[1789];
  assign o[14716] = i[1788];
  assign o[14715] = i[1787];
  assign o[14714] = i[1786];
  assign o[14713] = i[1785];
  assign o[14712] = i[1784];
  assign o[14711] = i[1783];
  assign o[14710] = i[1782];
  assign o[14709] = i[1781];
  assign o[14708] = i[1780];
  assign o[14707] = i[1779];
  assign o[14706] = i[1778];
  assign o[14705] = i[1777];
  assign o[14704] = i[1776];
  assign o[14703] = i[1775];
  assign o[14702] = i[1774];
  assign o[14701] = i[1773];
  assign o[14700] = i[1772];
  assign o[14699] = i[1771];
  assign o[14698] = i[1770];
  assign o[14697] = i[1769];
  assign o[14696] = i[1768];
  assign o[14695] = i[1767];
  assign o[14694] = i[1766];
  assign o[14693] = i[1765];
  assign o[14692] = i[1764];
  assign o[14691] = i[1763];
  assign o[14690] = i[1762];
  assign o[14689] = i[1761];
  assign o[14688] = i[1760];
  assign o[14687] = i[1759];
  assign o[14686] = i[1758];
  assign o[14685] = i[1757];
  assign o[14684] = i[1756];
  assign o[14683] = i[1755];
  assign o[14682] = i[1754];
  assign o[14681] = i[1753];
  assign o[14680] = i[1752];
  assign o[14679] = i[1751];
  assign o[14678] = i[1750];
  assign o[14677] = i[1749];
  assign o[14676] = i[1748];
  assign o[14675] = i[1747];
  assign o[14674] = i[1746];
  assign o[14673] = i[1745];
  assign o[14672] = i[1744];
  assign o[14671] = i[1743];
  assign o[14670] = i[1742];
  assign o[14669] = i[1741];
  assign o[14668] = i[1740];
  assign o[14667] = i[1739];
  assign o[14666] = i[1738];
  assign o[14665] = i[1737];
  assign o[14664] = i[1736];
  assign o[14663] = i[1735];
  assign o[14662] = i[1734];
  assign o[14661] = i[1733];
  assign o[14660] = i[1732];
  assign o[14659] = i[1731];
  assign o[14658] = i[1730];
  assign o[14657] = i[1729];
  assign o[14656] = i[1728];
  assign o[14655] = i[1727];
  assign o[14654] = i[1726];
  assign o[14653] = i[1725];
  assign o[14652] = i[1724];
  assign o[14651] = i[1723];
  assign o[14650] = i[1722];
  assign o[14649] = i[1721];
  assign o[14648] = i[1720];
  assign o[14647] = i[1719];
  assign o[14646] = i[1718];
  assign o[14645] = i[1717];
  assign o[14644] = i[1716];
  assign o[14643] = i[1715];
  assign o[14642] = i[1714];
  assign o[14641] = i[1713];
  assign o[14640] = i[1712];
  assign o[14639] = i[1711];
  assign o[14638] = i[1710];
  assign o[14637] = i[1709];
  assign o[14636] = i[1708];
  assign o[14635] = i[1707];
  assign o[14634] = i[1706];
  assign o[14633] = i[1705];
  assign o[14632] = i[1704];
  assign o[14631] = i[1703];
  assign o[14630] = i[1702];
  assign o[14629] = i[1701];
  assign o[14628] = i[1700];
  assign o[14627] = i[1699];
  assign o[14626] = i[1698];
  assign o[14625] = i[1697];
  assign o[14624] = i[1696];
  assign o[14623] = i[1695];
  assign o[14622] = i[1694];
  assign o[14621] = i[1693];
  assign o[14620] = i[1692];
  assign o[14619] = i[1691];
  assign o[14618] = i[1690];
  assign o[14617] = i[1689];
  assign o[14616] = i[1688];
  assign o[14615] = i[1687];
  assign o[14614] = i[1686];
  assign o[14613] = i[1685];
  assign o[14612] = i[1684];
  assign o[14611] = i[1683];
  assign o[14610] = i[1682];
  assign o[14609] = i[1681];
  assign o[14608] = i[1680];
  assign o[14607] = i[1679];
  assign o[14606] = i[1678];
  assign o[14605] = i[1677];
  assign o[14604] = i[1676];
  assign o[14603] = i[1675];
  assign o[14602] = i[1674];
  assign o[14601] = i[1673];
  assign o[14600] = i[1672];
  assign o[14599] = i[1671];
  assign o[14598] = i[1670];
  assign o[14597] = i[1669];
  assign o[14596] = i[1668];
  assign o[14595] = i[1667];
  assign o[14594] = i[1666];
  assign o[14593] = i[1665];
  assign o[14592] = i[1664];
  assign o[14591] = i[1919];
  assign o[14590] = i[1918];
  assign o[14589] = i[1917];
  assign o[14588] = i[1916];
  assign o[14587] = i[1915];
  assign o[14586] = i[1914];
  assign o[14585] = i[1913];
  assign o[14584] = i[1912];
  assign o[14583] = i[1911];
  assign o[14582] = i[1910];
  assign o[14581] = i[1909];
  assign o[14580] = i[1908];
  assign o[14579] = i[1907];
  assign o[14578] = i[1906];
  assign o[14577] = i[1905];
  assign o[14576] = i[1904];
  assign o[14575] = i[1903];
  assign o[14574] = i[1902];
  assign o[14573] = i[1901];
  assign o[14572] = i[1900];
  assign o[14571] = i[1899];
  assign o[14570] = i[1898];
  assign o[14569] = i[1897];
  assign o[14568] = i[1896];
  assign o[14567] = i[1895];
  assign o[14566] = i[1894];
  assign o[14565] = i[1893];
  assign o[14564] = i[1892];
  assign o[14563] = i[1891];
  assign o[14562] = i[1890];
  assign o[14561] = i[1889];
  assign o[14560] = i[1888];
  assign o[14559] = i[1887];
  assign o[14558] = i[1886];
  assign o[14557] = i[1885];
  assign o[14556] = i[1884];
  assign o[14555] = i[1883];
  assign o[14554] = i[1882];
  assign o[14553] = i[1881];
  assign o[14552] = i[1880];
  assign o[14551] = i[1879];
  assign o[14550] = i[1878];
  assign o[14549] = i[1877];
  assign o[14548] = i[1876];
  assign o[14547] = i[1875];
  assign o[14546] = i[1874];
  assign o[14545] = i[1873];
  assign o[14544] = i[1872];
  assign o[14543] = i[1871];
  assign o[14542] = i[1870];
  assign o[14541] = i[1869];
  assign o[14540] = i[1868];
  assign o[14539] = i[1867];
  assign o[14538] = i[1866];
  assign o[14537] = i[1865];
  assign o[14536] = i[1864];
  assign o[14535] = i[1863];
  assign o[14534] = i[1862];
  assign o[14533] = i[1861];
  assign o[14532] = i[1860];
  assign o[14531] = i[1859];
  assign o[14530] = i[1858];
  assign o[14529] = i[1857];
  assign o[14528] = i[1856];
  assign o[14527] = i[1855];
  assign o[14526] = i[1854];
  assign o[14525] = i[1853];
  assign o[14524] = i[1852];
  assign o[14523] = i[1851];
  assign o[14522] = i[1850];
  assign o[14521] = i[1849];
  assign o[14520] = i[1848];
  assign o[14519] = i[1847];
  assign o[14518] = i[1846];
  assign o[14517] = i[1845];
  assign o[14516] = i[1844];
  assign o[14515] = i[1843];
  assign o[14514] = i[1842];
  assign o[14513] = i[1841];
  assign o[14512] = i[1840];
  assign o[14511] = i[1839];
  assign o[14510] = i[1838];
  assign o[14509] = i[1837];
  assign o[14508] = i[1836];
  assign o[14507] = i[1835];
  assign o[14506] = i[1834];
  assign o[14505] = i[1833];
  assign o[14504] = i[1832];
  assign o[14503] = i[1831];
  assign o[14502] = i[1830];
  assign o[14501] = i[1829];
  assign o[14500] = i[1828];
  assign o[14499] = i[1827];
  assign o[14498] = i[1826];
  assign o[14497] = i[1825];
  assign o[14496] = i[1824];
  assign o[14495] = i[1823];
  assign o[14494] = i[1822];
  assign o[14493] = i[1821];
  assign o[14492] = i[1820];
  assign o[14491] = i[1819];
  assign o[14490] = i[1818];
  assign o[14489] = i[1817];
  assign o[14488] = i[1816];
  assign o[14487] = i[1815];
  assign o[14486] = i[1814];
  assign o[14485] = i[1813];
  assign o[14484] = i[1812];
  assign o[14483] = i[1811];
  assign o[14482] = i[1810];
  assign o[14481] = i[1809];
  assign o[14480] = i[1808];
  assign o[14479] = i[1807];
  assign o[14478] = i[1806];
  assign o[14477] = i[1805];
  assign o[14476] = i[1804];
  assign o[14475] = i[1803];
  assign o[14474] = i[1802];
  assign o[14473] = i[1801];
  assign o[14472] = i[1800];
  assign o[14471] = i[1799];
  assign o[14470] = i[1798];
  assign o[14469] = i[1797];
  assign o[14468] = i[1796];
  assign o[14467] = i[1795];
  assign o[14466] = i[1794];
  assign o[14465] = i[1793];
  assign o[14464] = i[1792];
  assign o[14463] = i[2047];
  assign o[14462] = i[2046];
  assign o[14461] = i[2045];
  assign o[14460] = i[2044];
  assign o[14459] = i[2043];
  assign o[14458] = i[2042];
  assign o[14457] = i[2041];
  assign o[14456] = i[2040];
  assign o[14455] = i[2039];
  assign o[14454] = i[2038];
  assign o[14453] = i[2037];
  assign o[14452] = i[2036];
  assign o[14451] = i[2035];
  assign o[14450] = i[2034];
  assign o[14449] = i[2033];
  assign o[14448] = i[2032];
  assign o[14447] = i[2031];
  assign o[14446] = i[2030];
  assign o[14445] = i[2029];
  assign o[14444] = i[2028];
  assign o[14443] = i[2027];
  assign o[14442] = i[2026];
  assign o[14441] = i[2025];
  assign o[14440] = i[2024];
  assign o[14439] = i[2023];
  assign o[14438] = i[2022];
  assign o[14437] = i[2021];
  assign o[14436] = i[2020];
  assign o[14435] = i[2019];
  assign o[14434] = i[2018];
  assign o[14433] = i[2017];
  assign o[14432] = i[2016];
  assign o[14431] = i[2015];
  assign o[14430] = i[2014];
  assign o[14429] = i[2013];
  assign o[14428] = i[2012];
  assign o[14427] = i[2011];
  assign o[14426] = i[2010];
  assign o[14425] = i[2009];
  assign o[14424] = i[2008];
  assign o[14423] = i[2007];
  assign o[14422] = i[2006];
  assign o[14421] = i[2005];
  assign o[14420] = i[2004];
  assign o[14419] = i[2003];
  assign o[14418] = i[2002];
  assign o[14417] = i[2001];
  assign o[14416] = i[2000];
  assign o[14415] = i[1999];
  assign o[14414] = i[1998];
  assign o[14413] = i[1997];
  assign o[14412] = i[1996];
  assign o[14411] = i[1995];
  assign o[14410] = i[1994];
  assign o[14409] = i[1993];
  assign o[14408] = i[1992];
  assign o[14407] = i[1991];
  assign o[14406] = i[1990];
  assign o[14405] = i[1989];
  assign o[14404] = i[1988];
  assign o[14403] = i[1987];
  assign o[14402] = i[1986];
  assign o[14401] = i[1985];
  assign o[14400] = i[1984];
  assign o[14399] = i[1983];
  assign o[14398] = i[1982];
  assign o[14397] = i[1981];
  assign o[14396] = i[1980];
  assign o[14395] = i[1979];
  assign o[14394] = i[1978];
  assign o[14393] = i[1977];
  assign o[14392] = i[1976];
  assign o[14391] = i[1975];
  assign o[14390] = i[1974];
  assign o[14389] = i[1973];
  assign o[14388] = i[1972];
  assign o[14387] = i[1971];
  assign o[14386] = i[1970];
  assign o[14385] = i[1969];
  assign o[14384] = i[1968];
  assign o[14383] = i[1967];
  assign o[14382] = i[1966];
  assign o[14381] = i[1965];
  assign o[14380] = i[1964];
  assign o[14379] = i[1963];
  assign o[14378] = i[1962];
  assign o[14377] = i[1961];
  assign o[14376] = i[1960];
  assign o[14375] = i[1959];
  assign o[14374] = i[1958];
  assign o[14373] = i[1957];
  assign o[14372] = i[1956];
  assign o[14371] = i[1955];
  assign o[14370] = i[1954];
  assign o[14369] = i[1953];
  assign o[14368] = i[1952];
  assign o[14367] = i[1951];
  assign o[14366] = i[1950];
  assign o[14365] = i[1949];
  assign o[14364] = i[1948];
  assign o[14363] = i[1947];
  assign o[14362] = i[1946];
  assign o[14361] = i[1945];
  assign o[14360] = i[1944];
  assign o[14359] = i[1943];
  assign o[14358] = i[1942];
  assign o[14357] = i[1941];
  assign o[14356] = i[1940];
  assign o[14355] = i[1939];
  assign o[14354] = i[1938];
  assign o[14353] = i[1937];
  assign o[14352] = i[1936];
  assign o[14351] = i[1935];
  assign o[14350] = i[1934];
  assign o[14349] = i[1933];
  assign o[14348] = i[1932];
  assign o[14347] = i[1931];
  assign o[14346] = i[1930];
  assign o[14345] = i[1929];
  assign o[14344] = i[1928];
  assign o[14343] = i[1927];
  assign o[14342] = i[1926];
  assign o[14341] = i[1925];
  assign o[14340] = i[1924];
  assign o[14339] = i[1923];
  assign o[14338] = i[1922];
  assign o[14337] = i[1921];
  assign o[14336] = i[1920];
  assign o[14335] = i[2175];
  assign o[14334] = i[2174];
  assign o[14333] = i[2173];
  assign o[14332] = i[2172];
  assign o[14331] = i[2171];
  assign o[14330] = i[2170];
  assign o[14329] = i[2169];
  assign o[14328] = i[2168];
  assign o[14327] = i[2167];
  assign o[14326] = i[2166];
  assign o[14325] = i[2165];
  assign o[14324] = i[2164];
  assign o[14323] = i[2163];
  assign o[14322] = i[2162];
  assign o[14321] = i[2161];
  assign o[14320] = i[2160];
  assign o[14319] = i[2159];
  assign o[14318] = i[2158];
  assign o[14317] = i[2157];
  assign o[14316] = i[2156];
  assign o[14315] = i[2155];
  assign o[14314] = i[2154];
  assign o[14313] = i[2153];
  assign o[14312] = i[2152];
  assign o[14311] = i[2151];
  assign o[14310] = i[2150];
  assign o[14309] = i[2149];
  assign o[14308] = i[2148];
  assign o[14307] = i[2147];
  assign o[14306] = i[2146];
  assign o[14305] = i[2145];
  assign o[14304] = i[2144];
  assign o[14303] = i[2143];
  assign o[14302] = i[2142];
  assign o[14301] = i[2141];
  assign o[14300] = i[2140];
  assign o[14299] = i[2139];
  assign o[14298] = i[2138];
  assign o[14297] = i[2137];
  assign o[14296] = i[2136];
  assign o[14295] = i[2135];
  assign o[14294] = i[2134];
  assign o[14293] = i[2133];
  assign o[14292] = i[2132];
  assign o[14291] = i[2131];
  assign o[14290] = i[2130];
  assign o[14289] = i[2129];
  assign o[14288] = i[2128];
  assign o[14287] = i[2127];
  assign o[14286] = i[2126];
  assign o[14285] = i[2125];
  assign o[14284] = i[2124];
  assign o[14283] = i[2123];
  assign o[14282] = i[2122];
  assign o[14281] = i[2121];
  assign o[14280] = i[2120];
  assign o[14279] = i[2119];
  assign o[14278] = i[2118];
  assign o[14277] = i[2117];
  assign o[14276] = i[2116];
  assign o[14275] = i[2115];
  assign o[14274] = i[2114];
  assign o[14273] = i[2113];
  assign o[14272] = i[2112];
  assign o[14271] = i[2111];
  assign o[14270] = i[2110];
  assign o[14269] = i[2109];
  assign o[14268] = i[2108];
  assign o[14267] = i[2107];
  assign o[14266] = i[2106];
  assign o[14265] = i[2105];
  assign o[14264] = i[2104];
  assign o[14263] = i[2103];
  assign o[14262] = i[2102];
  assign o[14261] = i[2101];
  assign o[14260] = i[2100];
  assign o[14259] = i[2099];
  assign o[14258] = i[2098];
  assign o[14257] = i[2097];
  assign o[14256] = i[2096];
  assign o[14255] = i[2095];
  assign o[14254] = i[2094];
  assign o[14253] = i[2093];
  assign o[14252] = i[2092];
  assign o[14251] = i[2091];
  assign o[14250] = i[2090];
  assign o[14249] = i[2089];
  assign o[14248] = i[2088];
  assign o[14247] = i[2087];
  assign o[14246] = i[2086];
  assign o[14245] = i[2085];
  assign o[14244] = i[2084];
  assign o[14243] = i[2083];
  assign o[14242] = i[2082];
  assign o[14241] = i[2081];
  assign o[14240] = i[2080];
  assign o[14239] = i[2079];
  assign o[14238] = i[2078];
  assign o[14237] = i[2077];
  assign o[14236] = i[2076];
  assign o[14235] = i[2075];
  assign o[14234] = i[2074];
  assign o[14233] = i[2073];
  assign o[14232] = i[2072];
  assign o[14231] = i[2071];
  assign o[14230] = i[2070];
  assign o[14229] = i[2069];
  assign o[14228] = i[2068];
  assign o[14227] = i[2067];
  assign o[14226] = i[2066];
  assign o[14225] = i[2065];
  assign o[14224] = i[2064];
  assign o[14223] = i[2063];
  assign o[14222] = i[2062];
  assign o[14221] = i[2061];
  assign o[14220] = i[2060];
  assign o[14219] = i[2059];
  assign o[14218] = i[2058];
  assign o[14217] = i[2057];
  assign o[14216] = i[2056];
  assign o[14215] = i[2055];
  assign o[14214] = i[2054];
  assign o[14213] = i[2053];
  assign o[14212] = i[2052];
  assign o[14211] = i[2051];
  assign o[14210] = i[2050];
  assign o[14209] = i[2049];
  assign o[14208] = i[2048];
  assign o[14207] = i[2303];
  assign o[14206] = i[2302];
  assign o[14205] = i[2301];
  assign o[14204] = i[2300];
  assign o[14203] = i[2299];
  assign o[14202] = i[2298];
  assign o[14201] = i[2297];
  assign o[14200] = i[2296];
  assign o[14199] = i[2295];
  assign o[14198] = i[2294];
  assign o[14197] = i[2293];
  assign o[14196] = i[2292];
  assign o[14195] = i[2291];
  assign o[14194] = i[2290];
  assign o[14193] = i[2289];
  assign o[14192] = i[2288];
  assign o[14191] = i[2287];
  assign o[14190] = i[2286];
  assign o[14189] = i[2285];
  assign o[14188] = i[2284];
  assign o[14187] = i[2283];
  assign o[14186] = i[2282];
  assign o[14185] = i[2281];
  assign o[14184] = i[2280];
  assign o[14183] = i[2279];
  assign o[14182] = i[2278];
  assign o[14181] = i[2277];
  assign o[14180] = i[2276];
  assign o[14179] = i[2275];
  assign o[14178] = i[2274];
  assign o[14177] = i[2273];
  assign o[14176] = i[2272];
  assign o[14175] = i[2271];
  assign o[14174] = i[2270];
  assign o[14173] = i[2269];
  assign o[14172] = i[2268];
  assign o[14171] = i[2267];
  assign o[14170] = i[2266];
  assign o[14169] = i[2265];
  assign o[14168] = i[2264];
  assign o[14167] = i[2263];
  assign o[14166] = i[2262];
  assign o[14165] = i[2261];
  assign o[14164] = i[2260];
  assign o[14163] = i[2259];
  assign o[14162] = i[2258];
  assign o[14161] = i[2257];
  assign o[14160] = i[2256];
  assign o[14159] = i[2255];
  assign o[14158] = i[2254];
  assign o[14157] = i[2253];
  assign o[14156] = i[2252];
  assign o[14155] = i[2251];
  assign o[14154] = i[2250];
  assign o[14153] = i[2249];
  assign o[14152] = i[2248];
  assign o[14151] = i[2247];
  assign o[14150] = i[2246];
  assign o[14149] = i[2245];
  assign o[14148] = i[2244];
  assign o[14147] = i[2243];
  assign o[14146] = i[2242];
  assign o[14145] = i[2241];
  assign o[14144] = i[2240];
  assign o[14143] = i[2239];
  assign o[14142] = i[2238];
  assign o[14141] = i[2237];
  assign o[14140] = i[2236];
  assign o[14139] = i[2235];
  assign o[14138] = i[2234];
  assign o[14137] = i[2233];
  assign o[14136] = i[2232];
  assign o[14135] = i[2231];
  assign o[14134] = i[2230];
  assign o[14133] = i[2229];
  assign o[14132] = i[2228];
  assign o[14131] = i[2227];
  assign o[14130] = i[2226];
  assign o[14129] = i[2225];
  assign o[14128] = i[2224];
  assign o[14127] = i[2223];
  assign o[14126] = i[2222];
  assign o[14125] = i[2221];
  assign o[14124] = i[2220];
  assign o[14123] = i[2219];
  assign o[14122] = i[2218];
  assign o[14121] = i[2217];
  assign o[14120] = i[2216];
  assign o[14119] = i[2215];
  assign o[14118] = i[2214];
  assign o[14117] = i[2213];
  assign o[14116] = i[2212];
  assign o[14115] = i[2211];
  assign o[14114] = i[2210];
  assign o[14113] = i[2209];
  assign o[14112] = i[2208];
  assign o[14111] = i[2207];
  assign o[14110] = i[2206];
  assign o[14109] = i[2205];
  assign o[14108] = i[2204];
  assign o[14107] = i[2203];
  assign o[14106] = i[2202];
  assign o[14105] = i[2201];
  assign o[14104] = i[2200];
  assign o[14103] = i[2199];
  assign o[14102] = i[2198];
  assign o[14101] = i[2197];
  assign o[14100] = i[2196];
  assign o[14099] = i[2195];
  assign o[14098] = i[2194];
  assign o[14097] = i[2193];
  assign o[14096] = i[2192];
  assign o[14095] = i[2191];
  assign o[14094] = i[2190];
  assign o[14093] = i[2189];
  assign o[14092] = i[2188];
  assign o[14091] = i[2187];
  assign o[14090] = i[2186];
  assign o[14089] = i[2185];
  assign o[14088] = i[2184];
  assign o[14087] = i[2183];
  assign o[14086] = i[2182];
  assign o[14085] = i[2181];
  assign o[14084] = i[2180];
  assign o[14083] = i[2179];
  assign o[14082] = i[2178];
  assign o[14081] = i[2177];
  assign o[14080] = i[2176];
  assign o[14079] = i[2431];
  assign o[14078] = i[2430];
  assign o[14077] = i[2429];
  assign o[14076] = i[2428];
  assign o[14075] = i[2427];
  assign o[14074] = i[2426];
  assign o[14073] = i[2425];
  assign o[14072] = i[2424];
  assign o[14071] = i[2423];
  assign o[14070] = i[2422];
  assign o[14069] = i[2421];
  assign o[14068] = i[2420];
  assign o[14067] = i[2419];
  assign o[14066] = i[2418];
  assign o[14065] = i[2417];
  assign o[14064] = i[2416];
  assign o[14063] = i[2415];
  assign o[14062] = i[2414];
  assign o[14061] = i[2413];
  assign o[14060] = i[2412];
  assign o[14059] = i[2411];
  assign o[14058] = i[2410];
  assign o[14057] = i[2409];
  assign o[14056] = i[2408];
  assign o[14055] = i[2407];
  assign o[14054] = i[2406];
  assign o[14053] = i[2405];
  assign o[14052] = i[2404];
  assign o[14051] = i[2403];
  assign o[14050] = i[2402];
  assign o[14049] = i[2401];
  assign o[14048] = i[2400];
  assign o[14047] = i[2399];
  assign o[14046] = i[2398];
  assign o[14045] = i[2397];
  assign o[14044] = i[2396];
  assign o[14043] = i[2395];
  assign o[14042] = i[2394];
  assign o[14041] = i[2393];
  assign o[14040] = i[2392];
  assign o[14039] = i[2391];
  assign o[14038] = i[2390];
  assign o[14037] = i[2389];
  assign o[14036] = i[2388];
  assign o[14035] = i[2387];
  assign o[14034] = i[2386];
  assign o[14033] = i[2385];
  assign o[14032] = i[2384];
  assign o[14031] = i[2383];
  assign o[14030] = i[2382];
  assign o[14029] = i[2381];
  assign o[14028] = i[2380];
  assign o[14027] = i[2379];
  assign o[14026] = i[2378];
  assign o[14025] = i[2377];
  assign o[14024] = i[2376];
  assign o[14023] = i[2375];
  assign o[14022] = i[2374];
  assign o[14021] = i[2373];
  assign o[14020] = i[2372];
  assign o[14019] = i[2371];
  assign o[14018] = i[2370];
  assign o[14017] = i[2369];
  assign o[14016] = i[2368];
  assign o[14015] = i[2367];
  assign o[14014] = i[2366];
  assign o[14013] = i[2365];
  assign o[14012] = i[2364];
  assign o[14011] = i[2363];
  assign o[14010] = i[2362];
  assign o[14009] = i[2361];
  assign o[14008] = i[2360];
  assign o[14007] = i[2359];
  assign o[14006] = i[2358];
  assign o[14005] = i[2357];
  assign o[14004] = i[2356];
  assign o[14003] = i[2355];
  assign o[14002] = i[2354];
  assign o[14001] = i[2353];
  assign o[14000] = i[2352];
  assign o[13999] = i[2351];
  assign o[13998] = i[2350];
  assign o[13997] = i[2349];
  assign o[13996] = i[2348];
  assign o[13995] = i[2347];
  assign o[13994] = i[2346];
  assign o[13993] = i[2345];
  assign o[13992] = i[2344];
  assign o[13991] = i[2343];
  assign o[13990] = i[2342];
  assign o[13989] = i[2341];
  assign o[13988] = i[2340];
  assign o[13987] = i[2339];
  assign o[13986] = i[2338];
  assign o[13985] = i[2337];
  assign o[13984] = i[2336];
  assign o[13983] = i[2335];
  assign o[13982] = i[2334];
  assign o[13981] = i[2333];
  assign o[13980] = i[2332];
  assign o[13979] = i[2331];
  assign o[13978] = i[2330];
  assign o[13977] = i[2329];
  assign o[13976] = i[2328];
  assign o[13975] = i[2327];
  assign o[13974] = i[2326];
  assign o[13973] = i[2325];
  assign o[13972] = i[2324];
  assign o[13971] = i[2323];
  assign o[13970] = i[2322];
  assign o[13969] = i[2321];
  assign o[13968] = i[2320];
  assign o[13967] = i[2319];
  assign o[13966] = i[2318];
  assign o[13965] = i[2317];
  assign o[13964] = i[2316];
  assign o[13963] = i[2315];
  assign o[13962] = i[2314];
  assign o[13961] = i[2313];
  assign o[13960] = i[2312];
  assign o[13959] = i[2311];
  assign o[13958] = i[2310];
  assign o[13957] = i[2309];
  assign o[13956] = i[2308];
  assign o[13955] = i[2307];
  assign o[13954] = i[2306];
  assign o[13953] = i[2305];
  assign o[13952] = i[2304];
  assign o[13951] = i[2559];
  assign o[13950] = i[2558];
  assign o[13949] = i[2557];
  assign o[13948] = i[2556];
  assign o[13947] = i[2555];
  assign o[13946] = i[2554];
  assign o[13945] = i[2553];
  assign o[13944] = i[2552];
  assign o[13943] = i[2551];
  assign o[13942] = i[2550];
  assign o[13941] = i[2549];
  assign o[13940] = i[2548];
  assign o[13939] = i[2547];
  assign o[13938] = i[2546];
  assign o[13937] = i[2545];
  assign o[13936] = i[2544];
  assign o[13935] = i[2543];
  assign o[13934] = i[2542];
  assign o[13933] = i[2541];
  assign o[13932] = i[2540];
  assign o[13931] = i[2539];
  assign o[13930] = i[2538];
  assign o[13929] = i[2537];
  assign o[13928] = i[2536];
  assign o[13927] = i[2535];
  assign o[13926] = i[2534];
  assign o[13925] = i[2533];
  assign o[13924] = i[2532];
  assign o[13923] = i[2531];
  assign o[13922] = i[2530];
  assign o[13921] = i[2529];
  assign o[13920] = i[2528];
  assign o[13919] = i[2527];
  assign o[13918] = i[2526];
  assign o[13917] = i[2525];
  assign o[13916] = i[2524];
  assign o[13915] = i[2523];
  assign o[13914] = i[2522];
  assign o[13913] = i[2521];
  assign o[13912] = i[2520];
  assign o[13911] = i[2519];
  assign o[13910] = i[2518];
  assign o[13909] = i[2517];
  assign o[13908] = i[2516];
  assign o[13907] = i[2515];
  assign o[13906] = i[2514];
  assign o[13905] = i[2513];
  assign o[13904] = i[2512];
  assign o[13903] = i[2511];
  assign o[13902] = i[2510];
  assign o[13901] = i[2509];
  assign o[13900] = i[2508];
  assign o[13899] = i[2507];
  assign o[13898] = i[2506];
  assign o[13897] = i[2505];
  assign o[13896] = i[2504];
  assign o[13895] = i[2503];
  assign o[13894] = i[2502];
  assign o[13893] = i[2501];
  assign o[13892] = i[2500];
  assign o[13891] = i[2499];
  assign o[13890] = i[2498];
  assign o[13889] = i[2497];
  assign o[13888] = i[2496];
  assign o[13887] = i[2495];
  assign o[13886] = i[2494];
  assign o[13885] = i[2493];
  assign o[13884] = i[2492];
  assign o[13883] = i[2491];
  assign o[13882] = i[2490];
  assign o[13881] = i[2489];
  assign o[13880] = i[2488];
  assign o[13879] = i[2487];
  assign o[13878] = i[2486];
  assign o[13877] = i[2485];
  assign o[13876] = i[2484];
  assign o[13875] = i[2483];
  assign o[13874] = i[2482];
  assign o[13873] = i[2481];
  assign o[13872] = i[2480];
  assign o[13871] = i[2479];
  assign o[13870] = i[2478];
  assign o[13869] = i[2477];
  assign o[13868] = i[2476];
  assign o[13867] = i[2475];
  assign o[13866] = i[2474];
  assign o[13865] = i[2473];
  assign o[13864] = i[2472];
  assign o[13863] = i[2471];
  assign o[13862] = i[2470];
  assign o[13861] = i[2469];
  assign o[13860] = i[2468];
  assign o[13859] = i[2467];
  assign o[13858] = i[2466];
  assign o[13857] = i[2465];
  assign o[13856] = i[2464];
  assign o[13855] = i[2463];
  assign o[13854] = i[2462];
  assign o[13853] = i[2461];
  assign o[13852] = i[2460];
  assign o[13851] = i[2459];
  assign o[13850] = i[2458];
  assign o[13849] = i[2457];
  assign o[13848] = i[2456];
  assign o[13847] = i[2455];
  assign o[13846] = i[2454];
  assign o[13845] = i[2453];
  assign o[13844] = i[2452];
  assign o[13843] = i[2451];
  assign o[13842] = i[2450];
  assign o[13841] = i[2449];
  assign o[13840] = i[2448];
  assign o[13839] = i[2447];
  assign o[13838] = i[2446];
  assign o[13837] = i[2445];
  assign o[13836] = i[2444];
  assign o[13835] = i[2443];
  assign o[13834] = i[2442];
  assign o[13833] = i[2441];
  assign o[13832] = i[2440];
  assign o[13831] = i[2439];
  assign o[13830] = i[2438];
  assign o[13829] = i[2437];
  assign o[13828] = i[2436];
  assign o[13827] = i[2435];
  assign o[13826] = i[2434];
  assign o[13825] = i[2433];
  assign o[13824] = i[2432];
  assign o[13823] = i[2687];
  assign o[13822] = i[2686];
  assign o[13821] = i[2685];
  assign o[13820] = i[2684];
  assign o[13819] = i[2683];
  assign o[13818] = i[2682];
  assign o[13817] = i[2681];
  assign o[13816] = i[2680];
  assign o[13815] = i[2679];
  assign o[13814] = i[2678];
  assign o[13813] = i[2677];
  assign o[13812] = i[2676];
  assign o[13811] = i[2675];
  assign o[13810] = i[2674];
  assign o[13809] = i[2673];
  assign o[13808] = i[2672];
  assign o[13807] = i[2671];
  assign o[13806] = i[2670];
  assign o[13805] = i[2669];
  assign o[13804] = i[2668];
  assign o[13803] = i[2667];
  assign o[13802] = i[2666];
  assign o[13801] = i[2665];
  assign o[13800] = i[2664];
  assign o[13799] = i[2663];
  assign o[13798] = i[2662];
  assign o[13797] = i[2661];
  assign o[13796] = i[2660];
  assign o[13795] = i[2659];
  assign o[13794] = i[2658];
  assign o[13793] = i[2657];
  assign o[13792] = i[2656];
  assign o[13791] = i[2655];
  assign o[13790] = i[2654];
  assign o[13789] = i[2653];
  assign o[13788] = i[2652];
  assign o[13787] = i[2651];
  assign o[13786] = i[2650];
  assign o[13785] = i[2649];
  assign o[13784] = i[2648];
  assign o[13783] = i[2647];
  assign o[13782] = i[2646];
  assign o[13781] = i[2645];
  assign o[13780] = i[2644];
  assign o[13779] = i[2643];
  assign o[13778] = i[2642];
  assign o[13777] = i[2641];
  assign o[13776] = i[2640];
  assign o[13775] = i[2639];
  assign o[13774] = i[2638];
  assign o[13773] = i[2637];
  assign o[13772] = i[2636];
  assign o[13771] = i[2635];
  assign o[13770] = i[2634];
  assign o[13769] = i[2633];
  assign o[13768] = i[2632];
  assign o[13767] = i[2631];
  assign o[13766] = i[2630];
  assign o[13765] = i[2629];
  assign o[13764] = i[2628];
  assign o[13763] = i[2627];
  assign o[13762] = i[2626];
  assign o[13761] = i[2625];
  assign o[13760] = i[2624];
  assign o[13759] = i[2623];
  assign o[13758] = i[2622];
  assign o[13757] = i[2621];
  assign o[13756] = i[2620];
  assign o[13755] = i[2619];
  assign o[13754] = i[2618];
  assign o[13753] = i[2617];
  assign o[13752] = i[2616];
  assign o[13751] = i[2615];
  assign o[13750] = i[2614];
  assign o[13749] = i[2613];
  assign o[13748] = i[2612];
  assign o[13747] = i[2611];
  assign o[13746] = i[2610];
  assign o[13745] = i[2609];
  assign o[13744] = i[2608];
  assign o[13743] = i[2607];
  assign o[13742] = i[2606];
  assign o[13741] = i[2605];
  assign o[13740] = i[2604];
  assign o[13739] = i[2603];
  assign o[13738] = i[2602];
  assign o[13737] = i[2601];
  assign o[13736] = i[2600];
  assign o[13735] = i[2599];
  assign o[13734] = i[2598];
  assign o[13733] = i[2597];
  assign o[13732] = i[2596];
  assign o[13731] = i[2595];
  assign o[13730] = i[2594];
  assign o[13729] = i[2593];
  assign o[13728] = i[2592];
  assign o[13727] = i[2591];
  assign o[13726] = i[2590];
  assign o[13725] = i[2589];
  assign o[13724] = i[2588];
  assign o[13723] = i[2587];
  assign o[13722] = i[2586];
  assign o[13721] = i[2585];
  assign o[13720] = i[2584];
  assign o[13719] = i[2583];
  assign o[13718] = i[2582];
  assign o[13717] = i[2581];
  assign o[13716] = i[2580];
  assign o[13715] = i[2579];
  assign o[13714] = i[2578];
  assign o[13713] = i[2577];
  assign o[13712] = i[2576];
  assign o[13711] = i[2575];
  assign o[13710] = i[2574];
  assign o[13709] = i[2573];
  assign o[13708] = i[2572];
  assign o[13707] = i[2571];
  assign o[13706] = i[2570];
  assign o[13705] = i[2569];
  assign o[13704] = i[2568];
  assign o[13703] = i[2567];
  assign o[13702] = i[2566];
  assign o[13701] = i[2565];
  assign o[13700] = i[2564];
  assign o[13699] = i[2563];
  assign o[13698] = i[2562];
  assign o[13697] = i[2561];
  assign o[13696] = i[2560];
  assign o[13695] = i[2815];
  assign o[13694] = i[2814];
  assign o[13693] = i[2813];
  assign o[13692] = i[2812];
  assign o[13691] = i[2811];
  assign o[13690] = i[2810];
  assign o[13689] = i[2809];
  assign o[13688] = i[2808];
  assign o[13687] = i[2807];
  assign o[13686] = i[2806];
  assign o[13685] = i[2805];
  assign o[13684] = i[2804];
  assign o[13683] = i[2803];
  assign o[13682] = i[2802];
  assign o[13681] = i[2801];
  assign o[13680] = i[2800];
  assign o[13679] = i[2799];
  assign o[13678] = i[2798];
  assign o[13677] = i[2797];
  assign o[13676] = i[2796];
  assign o[13675] = i[2795];
  assign o[13674] = i[2794];
  assign o[13673] = i[2793];
  assign o[13672] = i[2792];
  assign o[13671] = i[2791];
  assign o[13670] = i[2790];
  assign o[13669] = i[2789];
  assign o[13668] = i[2788];
  assign o[13667] = i[2787];
  assign o[13666] = i[2786];
  assign o[13665] = i[2785];
  assign o[13664] = i[2784];
  assign o[13663] = i[2783];
  assign o[13662] = i[2782];
  assign o[13661] = i[2781];
  assign o[13660] = i[2780];
  assign o[13659] = i[2779];
  assign o[13658] = i[2778];
  assign o[13657] = i[2777];
  assign o[13656] = i[2776];
  assign o[13655] = i[2775];
  assign o[13654] = i[2774];
  assign o[13653] = i[2773];
  assign o[13652] = i[2772];
  assign o[13651] = i[2771];
  assign o[13650] = i[2770];
  assign o[13649] = i[2769];
  assign o[13648] = i[2768];
  assign o[13647] = i[2767];
  assign o[13646] = i[2766];
  assign o[13645] = i[2765];
  assign o[13644] = i[2764];
  assign o[13643] = i[2763];
  assign o[13642] = i[2762];
  assign o[13641] = i[2761];
  assign o[13640] = i[2760];
  assign o[13639] = i[2759];
  assign o[13638] = i[2758];
  assign o[13637] = i[2757];
  assign o[13636] = i[2756];
  assign o[13635] = i[2755];
  assign o[13634] = i[2754];
  assign o[13633] = i[2753];
  assign o[13632] = i[2752];
  assign o[13631] = i[2751];
  assign o[13630] = i[2750];
  assign o[13629] = i[2749];
  assign o[13628] = i[2748];
  assign o[13627] = i[2747];
  assign o[13626] = i[2746];
  assign o[13625] = i[2745];
  assign o[13624] = i[2744];
  assign o[13623] = i[2743];
  assign o[13622] = i[2742];
  assign o[13621] = i[2741];
  assign o[13620] = i[2740];
  assign o[13619] = i[2739];
  assign o[13618] = i[2738];
  assign o[13617] = i[2737];
  assign o[13616] = i[2736];
  assign o[13615] = i[2735];
  assign o[13614] = i[2734];
  assign o[13613] = i[2733];
  assign o[13612] = i[2732];
  assign o[13611] = i[2731];
  assign o[13610] = i[2730];
  assign o[13609] = i[2729];
  assign o[13608] = i[2728];
  assign o[13607] = i[2727];
  assign o[13606] = i[2726];
  assign o[13605] = i[2725];
  assign o[13604] = i[2724];
  assign o[13603] = i[2723];
  assign o[13602] = i[2722];
  assign o[13601] = i[2721];
  assign o[13600] = i[2720];
  assign o[13599] = i[2719];
  assign o[13598] = i[2718];
  assign o[13597] = i[2717];
  assign o[13596] = i[2716];
  assign o[13595] = i[2715];
  assign o[13594] = i[2714];
  assign o[13593] = i[2713];
  assign o[13592] = i[2712];
  assign o[13591] = i[2711];
  assign o[13590] = i[2710];
  assign o[13589] = i[2709];
  assign o[13588] = i[2708];
  assign o[13587] = i[2707];
  assign o[13586] = i[2706];
  assign o[13585] = i[2705];
  assign o[13584] = i[2704];
  assign o[13583] = i[2703];
  assign o[13582] = i[2702];
  assign o[13581] = i[2701];
  assign o[13580] = i[2700];
  assign o[13579] = i[2699];
  assign o[13578] = i[2698];
  assign o[13577] = i[2697];
  assign o[13576] = i[2696];
  assign o[13575] = i[2695];
  assign o[13574] = i[2694];
  assign o[13573] = i[2693];
  assign o[13572] = i[2692];
  assign o[13571] = i[2691];
  assign o[13570] = i[2690];
  assign o[13569] = i[2689];
  assign o[13568] = i[2688];
  assign o[13567] = i[2943];
  assign o[13566] = i[2942];
  assign o[13565] = i[2941];
  assign o[13564] = i[2940];
  assign o[13563] = i[2939];
  assign o[13562] = i[2938];
  assign o[13561] = i[2937];
  assign o[13560] = i[2936];
  assign o[13559] = i[2935];
  assign o[13558] = i[2934];
  assign o[13557] = i[2933];
  assign o[13556] = i[2932];
  assign o[13555] = i[2931];
  assign o[13554] = i[2930];
  assign o[13553] = i[2929];
  assign o[13552] = i[2928];
  assign o[13551] = i[2927];
  assign o[13550] = i[2926];
  assign o[13549] = i[2925];
  assign o[13548] = i[2924];
  assign o[13547] = i[2923];
  assign o[13546] = i[2922];
  assign o[13545] = i[2921];
  assign o[13544] = i[2920];
  assign o[13543] = i[2919];
  assign o[13542] = i[2918];
  assign o[13541] = i[2917];
  assign o[13540] = i[2916];
  assign o[13539] = i[2915];
  assign o[13538] = i[2914];
  assign o[13537] = i[2913];
  assign o[13536] = i[2912];
  assign o[13535] = i[2911];
  assign o[13534] = i[2910];
  assign o[13533] = i[2909];
  assign o[13532] = i[2908];
  assign o[13531] = i[2907];
  assign o[13530] = i[2906];
  assign o[13529] = i[2905];
  assign o[13528] = i[2904];
  assign o[13527] = i[2903];
  assign o[13526] = i[2902];
  assign o[13525] = i[2901];
  assign o[13524] = i[2900];
  assign o[13523] = i[2899];
  assign o[13522] = i[2898];
  assign o[13521] = i[2897];
  assign o[13520] = i[2896];
  assign o[13519] = i[2895];
  assign o[13518] = i[2894];
  assign o[13517] = i[2893];
  assign o[13516] = i[2892];
  assign o[13515] = i[2891];
  assign o[13514] = i[2890];
  assign o[13513] = i[2889];
  assign o[13512] = i[2888];
  assign o[13511] = i[2887];
  assign o[13510] = i[2886];
  assign o[13509] = i[2885];
  assign o[13508] = i[2884];
  assign o[13507] = i[2883];
  assign o[13506] = i[2882];
  assign o[13505] = i[2881];
  assign o[13504] = i[2880];
  assign o[13503] = i[2879];
  assign o[13502] = i[2878];
  assign o[13501] = i[2877];
  assign o[13500] = i[2876];
  assign o[13499] = i[2875];
  assign o[13498] = i[2874];
  assign o[13497] = i[2873];
  assign o[13496] = i[2872];
  assign o[13495] = i[2871];
  assign o[13494] = i[2870];
  assign o[13493] = i[2869];
  assign o[13492] = i[2868];
  assign o[13491] = i[2867];
  assign o[13490] = i[2866];
  assign o[13489] = i[2865];
  assign o[13488] = i[2864];
  assign o[13487] = i[2863];
  assign o[13486] = i[2862];
  assign o[13485] = i[2861];
  assign o[13484] = i[2860];
  assign o[13483] = i[2859];
  assign o[13482] = i[2858];
  assign o[13481] = i[2857];
  assign o[13480] = i[2856];
  assign o[13479] = i[2855];
  assign o[13478] = i[2854];
  assign o[13477] = i[2853];
  assign o[13476] = i[2852];
  assign o[13475] = i[2851];
  assign o[13474] = i[2850];
  assign o[13473] = i[2849];
  assign o[13472] = i[2848];
  assign o[13471] = i[2847];
  assign o[13470] = i[2846];
  assign o[13469] = i[2845];
  assign o[13468] = i[2844];
  assign o[13467] = i[2843];
  assign o[13466] = i[2842];
  assign o[13465] = i[2841];
  assign o[13464] = i[2840];
  assign o[13463] = i[2839];
  assign o[13462] = i[2838];
  assign o[13461] = i[2837];
  assign o[13460] = i[2836];
  assign o[13459] = i[2835];
  assign o[13458] = i[2834];
  assign o[13457] = i[2833];
  assign o[13456] = i[2832];
  assign o[13455] = i[2831];
  assign o[13454] = i[2830];
  assign o[13453] = i[2829];
  assign o[13452] = i[2828];
  assign o[13451] = i[2827];
  assign o[13450] = i[2826];
  assign o[13449] = i[2825];
  assign o[13448] = i[2824];
  assign o[13447] = i[2823];
  assign o[13446] = i[2822];
  assign o[13445] = i[2821];
  assign o[13444] = i[2820];
  assign o[13443] = i[2819];
  assign o[13442] = i[2818];
  assign o[13441] = i[2817];
  assign o[13440] = i[2816];
  assign o[13439] = i[3071];
  assign o[13438] = i[3070];
  assign o[13437] = i[3069];
  assign o[13436] = i[3068];
  assign o[13435] = i[3067];
  assign o[13434] = i[3066];
  assign o[13433] = i[3065];
  assign o[13432] = i[3064];
  assign o[13431] = i[3063];
  assign o[13430] = i[3062];
  assign o[13429] = i[3061];
  assign o[13428] = i[3060];
  assign o[13427] = i[3059];
  assign o[13426] = i[3058];
  assign o[13425] = i[3057];
  assign o[13424] = i[3056];
  assign o[13423] = i[3055];
  assign o[13422] = i[3054];
  assign o[13421] = i[3053];
  assign o[13420] = i[3052];
  assign o[13419] = i[3051];
  assign o[13418] = i[3050];
  assign o[13417] = i[3049];
  assign o[13416] = i[3048];
  assign o[13415] = i[3047];
  assign o[13414] = i[3046];
  assign o[13413] = i[3045];
  assign o[13412] = i[3044];
  assign o[13411] = i[3043];
  assign o[13410] = i[3042];
  assign o[13409] = i[3041];
  assign o[13408] = i[3040];
  assign o[13407] = i[3039];
  assign o[13406] = i[3038];
  assign o[13405] = i[3037];
  assign o[13404] = i[3036];
  assign o[13403] = i[3035];
  assign o[13402] = i[3034];
  assign o[13401] = i[3033];
  assign o[13400] = i[3032];
  assign o[13399] = i[3031];
  assign o[13398] = i[3030];
  assign o[13397] = i[3029];
  assign o[13396] = i[3028];
  assign o[13395] = i[3027];
  assign o[13394] = i[3026];
  assign o[13393] = i[3025];
  assign o[13392] = i[3024];
  assign o[13391] = i[3023];
  assign o[13390] = i[3022];
  assign o[13389] = i[3021];
  assign o[13388] = i[3020];
  assign o[13387] = i[3019];
  assign o[13386] = i[3018];
  assign o[13385] = i[3017];
  assign o[13384] = i[3016];
  assign o[13383] = i[3015];
  assign o[13382] = i[3014];
  assign o[13381] = i[3013];
  assign o[13380] = i[3012];
  assign o[13379] = i[3011];
  assign o[13378] = i[3010];
  assign o[13377] = i[3009];
  assign o[13376] = i[3008];
  assign o[13375] = i[3007];
  assign o[13374] = i[3006];
  assign o[13373] = i[3005];
  assign o[13372] = i[3004];
  assign o[13371] = i[3003];
  assign o[13370] = i[3002];
  assign o[13369] = i[3001];
  assign o[13368] = i[3000];
  assign o[13367] = i[2999];
  assign o[13366] = i[2998];
  assign o[13365] = i[2997];
  assign o[13364] = i[2996];
  assign o[13363] = i[2995];
  assign o[13362] = i[2994];
  assign o[13361] = i[2993];
  assign o[13360] = i[2992];
  assign o[13359] = i[2991];
  assign o[13358] = i[2990];
  assign o[13357] = i[2989];
  assign o[13356] = i[2988];
  assign o[13355] = i[2987];
  assign o[13354] = i[2986];
  assign o[13353] = i[2985];
  assign o[13352] = i[2984];
  assign o[13351] = i[2983];
  assign o[13350] = i[2982];
  assign o[13349] = i[2981];
  assign o[13348] = i[2980];
  assign o[13347] = i[2979];
  assign o[13346] = i[2978];
  assign o[13345] = i[2977];
  assign o[13344] = i[2976];
  assign o[13343] = i[2975];
  assign o[13342] = i[2974];
  assign o[13341] = i[2973];
  assign o[13340] = i[2972];
  assign o[13339] = i[2971];
  assign o[13338] = i[2970];
  assign o[13337] = i[2969];
  assign o[13336] = i[2968];
  assign o[13335] = i[2967];
  assign o[13334] = i[2966];
  assign o[13333] = i[2965];
  assign o[13332] = i[2964];
  assign o[13331] = i[2963];
  assign o[13330] = i[2962];
  assign o[13329] = i[2961];
  assign o[13328] = i[2960];
  assign o[13327] = i[2959];
  assign o[13326] = i[2958];
  assign o[13325] = i[2957];
  assign o[13324] = i[2956];
  assign o[13323] = i[2955];
  assign o[13322] = i[2954];
  assign o[13321] = i[2953];
  assign o[13320] = i[2952];
  assign o[13319] = i[2951];
  assign o[13318] = i[2950];
  assign o[13317] = i[2949];
  assign o[13316] = i[2948];
  assign o[13315] = i[2947];
  assign o[13314] = i[2946];
  assign o[13313] = i[2945];
  assign o[13312] = i[2944];
  assign o[13311] = i[3199];
  assign o[13310] = i[3198];
  assign o[13309] = i[3197];
  assign o[13308] = i[3196];
  assign o[13307] = i[3195];
  assign o[13306] = i[3194];
  assign o[13305] = i[3193];
  assign o[13304] = i[3192];
  assign o[13303] = i[3191];
  assign o[13302] = i[3190];
  assign o[13301] = i[3189];
  assign o[13300] = i[3188];
  assign o[13299] = i[3187];
  assign o[13298] = i[3186];
  assign o[13297] = i[3185];
  assign o[13296] = i[3184];
  assign o[13295] = i[3183];
  assign o[13294] = i[3182];
  assign o[13293] = i[3181];
  assign o[13292] = i[3180];
  assign o[13291] = i[3179];
  assign o[13290] = i[3178];
  assign o[13289] = i[3177];
  assign o[13288] = i[3176];
  assign o[13287] = i[3175];
  assign o[13286] = i[3174];
  assign o[13285] = i[3173];
  assign o[13284] = i[3172];
  assign o[13283] = i[3171];
  assign o[13282] = i[3170];
  assign o[13281] = i[3169];
  assign o[13280] = i[3168];
  assign o[13279] = i[3167];
  assign o[13278] = i[3166];
  assign o[13277] = i[3165];
  assign o[13276] = i[3164];
  assign o[13275] = i[3163];
  assign o[13274] = i[3162];
  assign o[13273] = i[3161];
  assign o[13272] = i[3160];
  assign o[13271] = i[3159];
  assign o[13270] = i[3158];
  assign o[13269] = i[3157];
  assign o[13268] = i[3156];
  assign o[13267] = i[3155];
  assign o[13266] = i[3154];
  assign o[13265] = i[3153];
  assign o[13264] = i[3152];
  assign o[13263] = i[3151];
  assign o[13262] = i[3150];
  assign o[13261] = i[3149];
  assign o[13260] = i[3148];
  assign o[13259] = i[3147];
  assign o[13258] = i[3146];
  assign o[13257] = i[3145];
  assign o[13256] = i[3144];
  assign o[13255] = i[3143];
  assign o[13254] = i[3142];
  assign o[13253] = i[3141];
  assign o[13252] = i[3140];
  assign o[13251] = i[3139];
  assign o[13250] = i[3138];
  assign o[13249] = i[3137];
  assign o[13248] = i[3136];
  assign o[13247] = i[3135];
  assign o[13246] = i[3134];
  assign o[13245] = i[3133];
  assign o[13244] = i[3132];
  assign o[13243] = i[3131];
  assign o[13242] = i[3130];
  assign o[13241] = i[3129];
  assign o[13240] = i[3128];
  assign o[13239] = i[3127];
  assign o[13238] = i[3126];
  assign o[13237] = i[3125];
  assign o[13236] = i[3124];
  assign o[13235] = i[3123];
  assign o[13234] = i[3122];
  assign o[13233] = i[3121];
  assign o[13232] = i[3120];
  assign o[13231] = i[3119];
  assign o[13230] = i[3118];
  assign o[13229] = i[3117];
  assign o[13228] = i[3116];
  assign o[13227] = i[3115];
  assign o[13226] = i[3114];
  assign o[13225] = i[3113];
  assign o[13224] = i[3112];
  assign o[13223] = i[3111];
  assign o[13222] = i[3110];
  assign o[13221] = i[3109];
  assign o[13220] = i[3108];
  assign o[13219] = i[3107];
  assign o[13218] = i[3106];
  assign o[13217] = i[3105];
  assign o[13216] = i[3104];
  assign o[13215] = i[3103];
  assign o[13214] = i[3102];
  assign o[13213] = i[3101];
  assign o[13212] = i[3100];
  assign o[13211] = i[3099];
  assign o[13210] = i[3098];
  assign o[13209] = i[3097];
  assign o[13208] = i[3096];
  assign o[13207] = i[3095];
  assign o[13206] = i[3094];
  assign o[13205] = i[3093];
  assign o[13204] = i[3092];
  assign o[13203] = i[3091];
  assign o[13202] = i[3090];
  assign o[13201] = i[3089];
  assign o[13200] = i[3088];
  assign o[13199] = i[3087];
  assign o[13198] = i[3086];
  assign o[13197] = i[3085];
  assign o[13196] = i[3084];
  assign o[13195] = i[3083];
  assign o[13194] = i[3082];
  assign o[13193] = i[3081];
  assign o[13192] = i[3080];
  assign o[13191] = i[3079];
  assign o[13190] = i[3078];
  assign o[13189] = i[3077];
  assign o[13188] = i[3076];
  assign o[13187] = i[3075];
  assign o[13186] = i[3074];
  assign o[13185] = i[3073];
  assign o[13184] = i[3072];
  assign o[13183] = i[3327];
  assign o[13182] = i[3326];
  assign o[13181] = i[3325];
  assign o[13180] = i[3324];
  assign o[13179] = i[3323];
  assign o[13178] = i[3322];
  assign o[13177] = i[3321];
  assign o[13176] = i[3320];
  assign o[13175] = i[3319];
  assign o[13174] = i[3318];
  assign o[13173] = i[3317];
  assign o[13172] = i[3316];
  assign o[13171] = i[3315];
  assign o[13170] = i[3314];
  assign o[13169] = i[3313];
  assign o[13168] = i[3312];
  assign o[13167] = i[3311];
  assign o[13166] = i[3310];
  assign o[13165] = i[3309];
  assign o[13164] = i[3308];
  assign o[13163] = i[3307];
  assign o[13162] = i[3306];
  assign o[13161] = i[3305];
  assign o[13160] = i[3304];
  assign o[13159] = i[3303];
  assign o[13158] = i[3302];
  assign o[13157] = i[3301];
  assign o[13156] = i[3300];
  assign o[13155] = i[3299];
  assign o[13154] = i[3298];
  assign o[13153] = i[3297];
  assign o[13152] = i[3296];
  assign o[13151] = i[3295];
  assign o[13150] = i[3294];
  assign o[13149] = i[3293];
  assign o[13148] = i[3292];
  assign o[13147] = i[3291];
  assign o[13146] = i[3290];
  assign o[13145] = i[3289];
  assign o[13144] = i[3288];
  assign o[13143] = i[3287];
  assign o[13142] = i[3286];
  assign o[13141] = i[3285];
  assign o[13140] = i[3284];
  assign o[13139] = i[3283];
  assign o[13138] = i[3282];
  assign o[13137] = i[3281];
  assign o[13136] = i[3280];
  assign o[13135] = i[3279];
  assign o[13134] = i[3278];
  assign o[13133] = i[3277];
  assign o[13132] = i[3276];
  assign o[13131] = i[3275];
  assign o[13130] = i[3274];
  assign o[13129] = i[3273];
  assign o[13128] = i[3272];
  assign o[13127] = i[3271];
  assign o[13126] = i[3270];
  assign o[13125] = i[3269];
  assign o[13124] = i[3268];
  assign o[13123] = i[3267];
  assign o[13122] = i[3266];
  assign o[13121] = i[3265];
  assign o[13120] = i[3264];
  assign o[13119] = i[3263];
  assign o[13118] = i[3262];
  assign o[13117] = i[3261];
  assign o[13116] = i[3260];
  assign o[13115] = i[3259];
  assign o[13114] = i[3258];
  assign o[13113] = i[3257];
  assign o[13112] = i[3256];
  assign o[13111] = i[3255];
  assign o[13110] = i[3254];
  assign o[13109] = i[3253];
  assign o[13108] = i[3252];
  assign o[13107] = i[3251];
  assign o[13106] = i[3250];
  assign o[13105] = i[3249];
  assign o[13104] = i[3248];
  assign o[13103] = i[3247];
  assign o[13102] = i[3246];
  assign o[13101] = i[3245];
  assign o[13100] = i[3244];
  assign o[13099] = i[3243];
  assign o[13098] = i[3242];
  assign o[13097] = i[3241];
  assign o[13096] = i[3240];
  assign o[13095] = i[3239];
  assign o[13094] = i[3238];
  assign o[13093] = i[3237];
  assign o[13092] = i[3236];
  assign o[13091] = i[3235];
  assign o[13090] = i[3234];
  assign o[13089] = i[3233];
  assign o[13088] = i[3232];
  assign o[13087] = i[3231];
  assign o[13086] = i[3230];
  assign o[13085] = i[3229];
  assign o[13084] = i[3228];
  assign o[13083] = i[3227];
  assign o[13082] = i[3226];
  assign o[13081] = i[3225];
  assign o[13080] = i[3224];
  assign o[13079] = i[3223];
  assign o[13078] = i[3222];
  assign o[13077] = i[3221];
  assign o[13076] = i[3220];
  assign o[13075] = i[3219];
  assign o[13074] = i[3218];
  assign o[13073] = i[3217];
  assign o[13072] = i[3216];
  assign o[13071] = i[3215];
  assign o[13070] = i[3214];
  assign o[13069] = i[3213];
  assign o[13068] = i[3212];
  assign o[13067] = i[3211];
  assign o[13066] = i[3210];
  assign o[13065] = i[3209];
  assign o[13064] = i[3208];
  assign o[13063] = i[3207];
  assign o[13062] = i[3206];
  assign o[13061] = i[3205];
  assign o[13060] = i[3204];
  assign o[13059] = i[3203];
  assign o[13058] = i[3202];
  assign o[13057] = i[3201];
  assign o[13056] = i[3200];
  assign o[13055] = i[3455];
  assign o[13054] = i[3454];
  assign o[13053] = i[3453];
  assign o[13052] = i[3452];
  assign o[13051] = i[3451];
  assign o[13050] = i[3450];
  assign o[13049] = i[3449];
  assign o[13048] = i[3448];
  assign o[13047] = i[3447];
  assign o[13046] = i[3446];
  assign o[13045] = i[3445];
  assign o[13044] = i[3444];
  assign o[13043] = i[3443];
  assign o[13042] = i[3442];
  assign o[13041] = i[3441];
  assign o[13040] = i[3440];
  assign o[13039] = i[3439];
  assign o[13038] = i[3438];
  assign o[13037] = i[3437];
  assign o[13036] = i[3436];
  assign o[13035] = i[3435];
  assign o[13034] = i[3434];
  assign o[13033] = i[3433];
  assign o[13032] = i[3432];
  assign o[13031] = i[3431];
  assign o[13030] = i[3430];
  assign o[13029] = i[3429];
  assign o[13028] = i[3428];
  assign o[13027] = i[3427];
  assign o[13026] = i[3426];
  assign o[13025] = i[3425];
  assign o[13024] = i[3424];
  assign o[13023] = i[3423];
  assign o[13022] = i[3422];
  assign o[13021] = i[3421];
  assign o[13020] = i[3420];
  assign o[13019] = i[3419];
  assign o[13018] = i[3418];
  assign o[13017] = i[3417];
  assign o[13016] = i[3416];
  assign o[13015] = i[3415];
  assign o[13014] = i[3414];
  assign o[13013] = i[3413];
  assign o[13012] = i[3412];
  assign o[13011] = i[3411];
  assign o[13010] = i[3410];
  assign o[13009] = i[3409];
  assign o[13008] = i[3408];
  assign o[13007] = i[3407];
  assign o[13006] = i[3406];
  assign o[13005] = i[3405];
  assign o[13004] = i[3404];
  assign o[13003] = i[3403];
  assign o[13002] = i[3402];
  assign o[13001] = i[3401];
  assign o[13000] = i[3400];
  assign o[12999] = i[3399];
  assign o[12998] = i[3398];
  assign o[12997] = i[3397];
  assign o[12996] = i[3396];
  assign o[12995] = i[3395];
  assign o[12994] = i[3394];
  assign o[12993] = i[3393];
  assign o[12992] = i[3392];
  assign o[12991] = i[3391];
  assign o[12990] = i[3390];
  assign o[12989] = i[3389];
  assign o[12988] = i[3388];
  assign o[12987] = i[3387];
  assign o[12986] = i[3386];
  assign o[12985] = i[3385];
  assign o[12984] = i[3384];
  assign o[12983] = i[3383];
  assign o[12982] = i[3382];
  assign o[12981] = i[3381];
  assign o[12980] = i[3380];
  assign o[12979] = i[3379];
  assign o[12978] = i[3378];
  assign o[12977] = i[3377];
  assign o[12976] = i[3376];
  assign o[12975] = i[3375];
  assign o[12974] = i[3374];
  assign o[12973] = i[3373];
  assign o[12972] = i[3372];
  assign o[12971] = i[3371];
  assign o[12970] = i[3370];
  assign o[12969] = i[3369];
  assign o[12968] = i[3368];
  assign o[12967] = i[3367];
  assign o[12966] = i[3366];
  assign o[12965] = i[3365];
  assign o[12964] = i[3364];
  assign o[12963] = i[3363];
  assign o[12962] = i[3362];
  assign o[12961] = i[3361];
  assign o[12960] = i[3360];
  assign o[12959] = i[3359];
  assign o[12958] = i[3358];
  assign o[12957] = i[3357];
  assign o[12956] = i[3356];
  assign o[12955] = i[3355];
  assign o[12954] = i[3354];
  assign o[12953] = i[3353];
  assign o[12952] = i[3352];
  assign o[12951] = i[3351];
  assign o[12950] = i[3350];
  assign o[12949] = i[3349];
  assign o[12948] = i[3348];
  assign o[12947] = i[3347];
  assign o[12946] = i[3346];
  assign o[12945] = i[3345];
  assign o[12944] = i[3344];
  assign o[12943] = i[3343];
  assign o[12942] = i[3342];
  assign o[12941] = i[3341];
  assign o[12940] = i[3340];
  assign o[12939] = i[3339];
  assign o[12938] = i[3338];
  assign o[12937] = i[3337];
  assign o[12936] = i[3336];
  assign o[12935] = i[3335];
  assign o[12934] = i[3334];
  assign o[12933] = i[3333];
  assign o[12932] = i[3332];
  assign o[12931] = i[3331];
  assign o[12930] = i[3330];
  assign o[12929] = i[3329];
  assign o[12928] = i[3328];
  assign o[12927] = i[3583];
  assign o[12926] = i[3582];
  assign o[12925] = i[3581];
  assign o[12924] = i[3580];
  assign o[12923] = i[3579];
  assign o[12922] = i[3578];
  assign o[12921] = i[3577];
  assign o[12920] = i[3576];
  assign o[12919] = i[3575];
  assign o[12918] = i[3574];
  assign o[12917] = i[3573];
  assign o[12916] = i[3572];
  assign o[12915] = i[3571];
  assign o[12914] = i[3570];
  assign o[12913] = i[3569];
  assign o[12912] = i[3568];
  assign o[12911] = i[3567];
  assign o[12910] = i[3566];
  assign o[12909] = i[3565];
  assign o[12908] = i[3564];
  assign o[12907] = i[3563];
  assign o[12906] = i[3562];
  assign o[12905] = i[3561];
  assign o[12904] = i[3560];
  assign o[12903] = i[3559];
  assign o[12902] = i[3558];
  assign o[12901] = i[3557];
  assign o[12900] = i[3556];
  assign o[12899] = i[3555];
  assign o[12898] = i[3554];
  assign o[12897] = i[3553];
  assign o[12896] = i[3552];
  assign o[12895] = i[3551];
  assign o[12894] = i[3550];
  assign o[12893] = i[3549];
  assign o[12892] = i[3548];
  assign o[12891] = i[3547];
  assign o[12890] = i[3546];
  assign o[12889] = i[3545];
  assign o[12888] = i[3544];
  assign o[12887] = i[3543];
  assign o[12886] = i[3542];
  assign o[12885] = i[3541];
  assign o[12884] = i[3540];
  assign o[12883] = i[3539];
  assign o[12882] = i[3538];
  assign o[12881] = i[3537];
  assign o[12880] = i[3536];
  assign o[12879] = i[3535];
  assign o[12878] = i[3534];
  assign o[12877] = i[3533];
  assign o[12876] = i[3532];
  assign o[12875] = i[3531];
  assign o[12874] = i[3530];
  assign o[12873] = i[3529];
  assign o[12872] = i[3528];
  assign o[12871] = i[3527];
  assign o[12870] = i[3526];
  assign o[12869] = i[3525];
  assign o[12868] = i[3524];
  assign o[12867] = i[3523];
  assign o[12866] = i[3522];
  assign o[12865] = i[3521];
  assign o[12864] = i[3520];
  assign o[12863] = i[3519];
  assign o[12862] = i[3518];
  assign o[12861] = i[3517];
  assign o[12860] = i[3516];
  assign o[12859] = i[3515];
  assign o[12858] = i[3514];
  assign o[12857] = i[3513];
  assign o[12856] = i[3512];
  assign o[12855] = i[3511];
  assign o[12854] = i[3510];
  assign o[12853] = i[3509];
  assign o[12852] = i[3508];
  assign o[12851] = i[3507];
  assign o[12850] = i[3506];
  assign o[12849] = i[3505];
  assign o[12848] = i[3504];
  assign o[12847] = i[3503];
  assign o[12846] = i[3502];
  assign o[12845] = i[3501];
  assign o[12844] = i[3500];
  assign o[12843] = i[3499];
  assign o[12842] = i[3498];
  assign o[12841] = i[3497];
  assign o[12840] = i[3496];
  assign o[12839] = i[3495];
  assign o[12838] = i[3494];
  assign o[12837] = i[3493];
  assign o[12836] = i[3492];
  assign o[12835] = i[3491];
  assign o[12834] = i[3490];
  assign o[12833] = i[3489];
  assign o[12832] = i[3488];
  assign o[12831] = i[3487];
  assign o[12830] = i[3486];
  assign o[12829] = i[3485];
  assign o[12828] = i[3484];
  assign o[12827] = i[3483];
  assign o[12826] = i[3482];
  assign o[12825] = i[3481];
  assign o[12824] = i[3480];
  assign o[12823] = i[3479];
  assign o[12822] = i[3478];
  assign o[12821] = i[3477];
  assign o[12820] = i[3476];
  assign o[12819] = i[3475];
  assign o[12818] = i[3474];
  assign o[12817] = i[3473];
  assign o[12816] = i[3472];
  assign o[12815] = i[3471];
  assign o[12814] = i[3470];
  assign o[12813] = i[3469];
  assign o[12812] = i[3468];
  assign o[12811] = i[3467];
  assign o[12810] = i[3466];
  assign o[12809] = i[3465];
  assign o[12808] = i[3464];
  assign o[12807] = i[3463];
  assign o[12806] = i[3462];
  assign o[12805] = i[3461];
  assign o[12804] = i[3460];
  assign o[12803] = i[3459];
  assign o[12802] = i[3458];
  assign o[12801] = i[3457];
  assign o[12800] = i[3456];
  assign o[12799] = i[3711];
  assign o[12798] = i[3710];
  assign o[12797] = i[3709];
  assign o[12796] = i[3708];
  assign o[12795] = i[3707];
  assign o[12794] = i[3706];
  assign o[12793] = i[3705];
  assign o[12792] = i[3704];
  assign o[12791] = i[3703];
  assign o[12790] = i[3702];
  assign o[12789] = i[3701];
  assign o[12788] = i[3700];
  assign o[12787] = i[3699];
  assign o[12786] = i[3698];
  assign o[12785] = i[3697];
  assign o[12784] = i[3696];
  assign o[12783] = i[3695];
  assign o[12782] = i[3694];
  assign o[12781] = i[3693];
  assign o[12780] = i[3692];
  assign o[12779] = i[3691];
  assign o[12778] = i[3690];
  assign o[12777] = i[3689];
  assign o[12776] = i[3688];
  assign o[12775] = i[3687];
  assign o[12774] = i[3686];
  assign o[12773] = i[3685];
  assign o[12772] = i[3684];
  assign o[12771] = i[3683];
  assign o[12770] = i[3682];
  assign o[12769] = i[3681];
  assign o[12768] = i[3680];
  assign o[12767] = i[3679];
  assign o[12766] = i[3678];
  assign o[12765] = i[3677];
  assign o[12764] = i[3676];
  assign o[12763] = i[3675];
  assign o[12762] = i[3674];
  assign o[12761] = i[3673];
  assign o[12760] = i[3672];
  assign o[12759] = i[3671];
  assign o[12758] = i[3670];
  assign o[12757] = i[3669];
  assign o[12756] = i[3668];
  assign o[12755] = i[3667];
  assign o[12754] = i[3666];
  assign o[12753] = i[3665];
  assign o[12752] = i[3664];
  assign o[12751] = i[3663];
  assign o[12750] = i[3662];
  assign o[12749] = i[3661];
  assign o[12748] = i[3660];
  assign o[12747] = i[3659];
  assign o[12746] = i[3658];
  assign o[12745] = i[3657];
  assign o[12744] = i[3656];
  assign o[12743] = i[3655];
  assign o[12742] = i[3654];
  assign o[12741] = i[3653];
  assign o[12740] = i[3652];
  assign o[12739] = i[3651];
  assign o[12738] = i[3650];
  assign o[12737] = i[3649];
  assign o[12736] = i[3648];
  assign o[12735] = i[3647];
  assign o[12734] = i[3646];
  assign o[12733] = i[3645];
  assign o[12732] = i[3644];
  assign o[12731] = i[3643];
  assign o[12730] = i[3642];
  assign o[12729] = i[3641];
  assign o[12728] = i[3640];
  assign o[12727] = i[3639];
  assign o[12726] = i[3638];
  assign o[12725] = i[3637];
  assign o[12724] = i[3636];
  assign o[12723] = i[3635];
  assign o[12722] = i[3634];
  assign o[12721] = i[3633];
  assign o[12720] = i[3632];
  assign o[12719] = i[3631];
  assign o[12718] = i[3630];
  assign o[12717] = i[3629];
  assign o[12716] = i[3628];
  assign o[12715] = i[3627];
  assign o[12714] = i[3626];
  assign o[12713] = i[3625];
  assign o[12712] = i[3624];
  assign o[12711] = i[3623];
  assign o[12710] = i[3622];
  assign o[12709] = i[3621];
  assign o[12708] = i[3620];
  assign o[12707] = i[3619];
  assign o[12706] = i[3618];
  assign o[12705] = i[3617];
  assign o[12704] = i[3616];
  assign o[12703] = i[3615];
  assign o[12702] = i[3614];
  assign o[12701] = i[3613];
  assign o[12700] = i[3612];
  assign o[12699] = i[3611];
  assign o[12698] = i[3610];
  assign o[12697] = i[3609];
  assign o[12696] = i[3608];
  assign o[12695] = i[3607];
  assign o[12694] = i[3606];
  assign o[12693] = i[3605];
  assign o[12692] = i[3604];
  assign o[12691] = i[3603];
  assign o[12690] = i[3602];
  assign o[12689] = i[3601];
  assign o[12688] = i[3600];
  assign o[12687] = i[3599];
  assign o[12686] = i[3598];
  assign o[12685] = i[3597];
  assign o[12684] = i[3596];
  assign o[12683] = i[3595];
  assign o[12682] = i[3594];
  assign o[12681] = i[3593];
  assign o[12680] = i[3592];
  assign o[12679] = i[3591];
  assign o[12678] = i[3590];
  assign o[12677] = i[3589];
  assign o[12676] = i[3588];
  assign o[12675] = i[3587];
  assign o[12674] = i[3586];
  assign o[12673] = i[3585];
  assign o[12672] = i[3584];
  assign o[12671] = i[3839];
  assign o[12670] = i[3838];
  assign o[12669] = i[3837];
  assign o[12668] = i[3836];
  assign o[12667] = i[3835];
  assign o[12666] = i[3834];
  assign o[12665] = i[3833];
  assign o[12664] = i[3832];
  assign o[12663] = i[3831];
  assign o[12662] = i[3830];
  assign o[12661] = i[3829];
  assign o[12660] = i[3828];
  assign o[12659] = i[3827];
  assign o[12658] = i[3826];
  assign o[12657] = i[3825];
  assign o[12656] = i[3824];
  assign o[12655] = i[3823];
  assign o[12654] = i[3822];
  assign o[12653] = i[3821];
  assign o[12652] = i[3820];
  assign o[12651] = i[3819];
  assign o[12650] = i[3818];
  assign o[12649] = i[3817];
  assign o[12648] = i[3816];
  assign o[12647] = i[3815];
  assign o[12646] = i[3814];
  assign o[12645] = i[3813];
  assign o[12644] = i[3812];
  assign o[12643] = i[3811];
  assign o[12642] = i[3810];
  assign o[12641] = i[3809];
  assign o[12640] = i[3808];
  assign o[12639] = i[3807];
  assign o[12638] = i[3806];
  assign o[12637] = i[3805];
  assign o[12636] = i[3804];
  assign o[12635] = i[3803];
  assign o[12634] = i[3802];
  assign o[12633] = i[3801];
  assign o[12632] = i[3800];
  assign o[12631] = i[3799];
  assign o[12630] = i[3798];
  assign o[12629] = i[3797];
  assign o[12628] = i[3796];
  assign o[12627] = i[3795];
  assign o[12626] = i[3794];
  assign o[12625] = i[3793];
  assign o[12624] = i[3792];
  assign o[12623] = i[3791];
  assign o[12622] = i[3790];
  assign o[12621] = i[3789];
  assign o[12620] = i[3788];
  assign o[12619] = i[3787];
  assign o[12618] = i[3786];
  assign o[12617] = i[3785];
  assign o[12616] = i[3784];
  assign o[12615] = i[3783];
  assign o[12614] = i[3782];
  assign o[12613] = i[3781];
  assign o[12612] = i[3780];
  assign o[12611] = i[3779];
  assign o[12610] = i[3778];
  assign o[12609] = i[3777];
  assign o[12608] = i[3776];
  assign o[12607] = i[3775];
  assign o[12606] = i[3774];
  assign o[12605] = i[3773];
  assign o[12604] = i[3772];
  assign o[12603] = i[3771];
  assign o[12602] = i[3770];
  assign o[12601] = i[3769];
  assign o[12600] = i[3768];
  assign o[12599] = i[3767];
  assign o[12598] = i[3766];
  assign o[12597] = i[3765];
  assign o[12596] = i[3764];
  assign o[12595] = i[3763];
  assign o[12594] = i[3762];
  assign o[12593] = i[3761];
  assign o[12592] = i[3760];
  assign o[12591] = i[3759];
  assign o[12590] = i[3758];
  assign o[12589] = i[3757];
  assign o[12588] = i[3756];
  assign o[12587] = i[3755];
  assign o[12586] = i[3754];
  assign o[12585] = i[3753];
  assign o[12584] = i[3752];
  assign o[12583] = i[3751];
  assign o[12582] = i[3750];
  assign o[12581] = i[3749];
  assign o[12580] = i[3748];
  assign o[12579] = i[3747];
  assign o[12578] = i[3746];
  assign o[12577] = i[3745];
  assign o[12576] = i[3744];
  assign o[12575] = i[3743];
  assign o[12574] = i[3742];
  assign o[12573] = i[3741];
  assign o[12572] = i[3740];
  assign o[12571] = i[3739];
  assign o[12570] = i[3738];
  assign o[12569] = i[3737];
  assign o[12568] = i[3736];
  assign o[12567] = i[3735];
  assign o[12566] = i[3734];
  assign o[12565] = i[3733];
  assign o[12564] = i[3732];
  assign o[12563] = i[3731];
  assign o[12562] = i[3730];
  assign o[12561] = i[3729];
  assign o[12560] = i[3728];
  assign o[12559] = i[3727];
  assign o[12558] = i[3726];
  assign o[12557] = i[3725];
  assign o[12556] = i[3724];
  assign o[12555] = i[3723];
  assign o[12554] = i[3722];
  assign o[12553] = i[3721];
  assign o[12552] = i[3720];
  assign o[12551] = i[3719];
  assign o[12550] = i[3718];
  assign o[12549] = i[3717];
  assign o[12548] = i[3716];
  assign o[12547] = i[3715];
  assign o[12546] = i[3714];
  assign o[12545] = i[3713];
  assign o[12544] = i[3712];
  assign o[12543] = i[3967];
  assign o[12542] = i[3966];
  assign o[12541] = i[3965];
  assign o[12540] = i[3964];
  assign o[12539] = i[3963];
  assign o[12538] = i[3962];
  assign o[12537] = i[3961];
  assign o[12536] = i[3960];
  assign o[12535] = i[3959];
  assign o[12534] = i[3958];
  assign o[12533] = i[3957];
  assign o[12532] = i[3956];
  assign o[12531] = i[3955];
  assign o[12530] = i[3954];
  assign o[12529] = i[3953];
  assign o[12528] = i[3952];
  assign o[12527] = i[3951];
  assign o[12526] = i[3950];
  assign o[12525] = i[3949];
  assign o[12524] = i[3948];
  assign o[12523] = i[3947];
  assign o[12522] = i[3946];
  assign o[12521] = i[3945];
  assign o[12520] = i[3944];
  assign o[12519] = i[3943];
  assign o[12518] = i[3942];
  assign o[12517] = i[3941];
  assign o[12516] = i[3940];
  assign o[12515] = i[3939];
  assign o[12514] = i[3938];
  assign o[12513] = i[3937];
  assign o[12512] = i[3936];
  assign o[12511] = i[3935];
  assign o[12510] = i[3934];
  assign o[12509] = i[3933];
  assign o[12508] = i[3932];
  assign o[12507] = i[3931];
  assign o[12506] = i[3930];
  assign o[12505] = i[3929];
  assign o[12504] = i[3928];
  assign o[12503] = i[3927];
  assign o[12502] = i[3926];
  assign o[12501] = i[3925];
  assign o[12500] = i[3924];
  assign o[12499] = i[3923];
  assign o[12498] = i[3922];
  assign o[12497] = i[3921];
  assign o[12496] = i[3920];
  assign o[12495] = i[3919];
  assign o[12494] = i[3918];
  assign o[12493] = i[3917];
  assign o[12492] = i[3916];
  assign o[12491] = i[3915];
  assign o[12490] = i[3914];
  assign o[12489] = i[3913];
  assign o[12488] = i[3912];
  assign o[12487] = i[3911];
  assign o[12486] = i[3910];
  assign o[12485] = i[3909];
  assign o[12484] = i[3908];
  assign o[12483] = i[3907];
  assign o[12482] = i[3906];
  assign o[12481] = i[3905];
  assign o[12480] = i[3904];
  assign o[12479] = i[3903];
  assign o[12478] = i[3902];
  assign o[12477] = i[3901];
  assign o[12476] = i[3900];
  assign o[12475] = i[3899];
  assign o[12474] = i[3898];
  assign o[12473] = i[3897];
  assign o[12472] = i[3896];
  assign o[12471] = i[3895];
  assign o[12470] = i[3894];
  assign o[12469] = i[3893];
  assign o[12468] = i[3892];
  assign o[12467] = i[3891];
  assign o[12466] = i[3890];
  assign o[12465] = i[3889];
  assign o[12464] = i[3888];
  assign o[12463] = i[3887];
  assign o[12462] = i[3886];
  assign o[12461] = i[3885];
  assign o[12460] = i[3884];
  assign o[12459] = i[3883];
  assign o[12458] = i[3882];
  assign o[12457] = i[3881];
  assign o[12456] = i[3880];
  assign o[12455] = i[3879];
  assign o[12454] = i[3878];
  assign o[12453] = i[3877];
  assign o[12452] = i[3876];
  assign o[12451] = i[3875];
  assign o[12450] = i[3874];
  assign o[12449] = i[3873];
  assign o[12448] = i[3872];
  assign o[12447] = i[3871];
  assign o[12446] = i[3870];
  assign o[12445] = i[3869];
  assign o[12444] = i[3868];
  assign o[12443] = i[3867];
  assign o[12442] = i[3866];
  assign o[12441] = i[3865];
  assign o[12440] = i[3864];
  assign o[12439] = i[3863];
  assign o[12438] = i[3862];
  assign o[12437] = i[3861];
  assign o[12436] = i[3860];
  assign o[12435] = i[3859];
  assign o[12434] = i[3858];
  assign o[12433] = i[3857];
  assign o[12432] = i[3856];
  assign o[12431] = i[3855];
  assign o[12430] = i[3854];
  assign o[12429] = i[3853];
  assign o[12428] = i[3852];
  assign o[12427] = i[3851];
  assign o[12426] = i[3850];
  assign o[12425] = i[3849];
  assign o[12424] = i[3848];
  assign o[12423] = i[3847];
  assign o[12422] = i[3846];
  assign o[12421] = i[3845];
  assign o[12420] = i[3844];
  assign o[12419] = i[3843];
  assign o[12418] = i[3842];
  assign o[12417] = i[3841];
  assign o[12416] = i[3840];
  assign o[12415] = i[4095];
  assign o[12414] = i[4094];
  assign o[12413] = i[4093];
  assign o[12412] = i[4092];
  assign o[12411] = i[4091];
  assign o[12410] = i[4090];
  assign o[12409] = i[4089];
  assign o[12408] = i[4088];
  assign o[12407] = i[4087];
  assign o[12406] = i[4086];
  assign o[12405] = i[4085];
  assign o[12404] = i[4084];
  assign o[12403] = i[4083];
  assign o[12402] = i[4082];
  assign o[12401] = i[4081];
  assign o[12400] = i[4080];
  assign o[12399] = i[4079];
  assign o[12398] = i[4078];
  assign o[12397] = i[4077];
  assign o[12396] = i[4076];
  assign o[12395] = i[4075];
  assign o[12394] = i[4074];
  assign o[12393] = i[4073];
  assign o[12392] = i[4072];
  assign o[12391] = i[4071];
  assign o[12390] = i[4070];
  assign o[12389] = i[4069];
  assign o[12388] = i[4068];
  assign o[12387] = i[4067];
  assign o[12386] = i[4066];
  assign o[12385] = i[4065];
  assign o[12384] = i[4064];
  assign o[12383] = i[4063];
  assign o[12382] = i[4062];
  assign o[12381] = i[4061];
  assign o[12380] = i[4060];
  assign o[12379] = i[4059];
  assign o[12378] = i[4058];
  assign o[12377] = i[4057];
  assign o[12376] = i[4056];
  assign o[12375] = i[4055];
  assign o[12374] = i[4054];
  assign o[12373] = i[4053];
  assign o[12372] = i[4052];
  assign o[12371] = i[4051];
  assign o[12370] = i[4050];
  assign o[12369] = i[4049];
  assign o[12368] = i[4048];
  assign o[12367] = i[4047];
  assign o[12366] = i[4046];
  assign o[12365] = i[4045];
  assign o[12364] = i[4044];
  assign o[12363] = i[4043];
  assign o[12362] = i[4042];
  assign o[12361] = i[4041];
  assign o[12360] = i[4040];
  assign o[12359] = i[4039];
  assign o[12358] = i[4038];
  assign o[12357] = i[4037];
  assign o[12356] = i[4036];
  assign o[12355] = i[4035];
  assign o[12354] = i[4034];
  assign o[12353] = i[4033];
  assign o[12352] = i[4032];
  assign o[12351] = i[4031];
  assign o[12350] = i[4030];
  assign o[12349] = i[4029];
  assign o[12348] = i[4028];
  assign o[12347] = i[4027];
  assign o[12346] = i[4026];
  assign o[12345] = i[4025];
  assign o[12344] = i[4024];
  assign o[12343] = i[4023];
  assign o[12342] = i[4022];
  assign o[12341] = i[4021];
  assign o[12340] = i[4020];
  assign o[12339] = i[4019];
  assign o[12338] = i[4018];
  assign o[12337] = i[4017];
  assign o[12336] = i[4016];
  assign o[12335] = i[4015];
  assign o[12334] = i[4014];
  assign o[12333] = i[4013];
  assign o[12332] = i[4012];
  assign o[12331] = i[4011];
  assign o[12330] = i[4010];
  assign o[12329] = i[4009];
  assign o[12328] = i[4008];
  assign o[12327] = i[4007];
  assign o[12326] = i[4006];
  assign o[12325] = i[4005];
  assign o[12324] = i[4004];
  assign o[12323] = i[4003];
  assign o[12322] = i[4002];
  assign o[12321] = i[4001];
  assign o[12320] = i[4000];
  assign o[12319] = i[3999];
  assign o[12318] = i[3998];
  assign o[12317] = i[3997];
  assign o[12316] = i[3996];
  assign o[12315] = i[3995];
  assign o[12314] = i[3994];
  assign o[12313] = i[3993];
  assign o[12312] = i[3992];
  assign o[12311] = i[3991];
  assign o[12310] = i[3990];
  assign o[12309] = i[3989];
  assign o[12308] = i[3988];
  assign o[12307] = i[3987];
  assign o[12306] = i[3986];
  assign o[12305] = i[3985];
  assign o[12304] = i[3984];
  assign o[12303] = i[3983];
  assign o[12302] = i[3982];
  assign o[12301] = i[3981];
  assign o[12300] = i[3980];
  assign o[12299] = i[3979];
  assign o[12298] = i[3978];
  assign o[12297] = i[3977];
  assign o[12296] = i[3976];
  assign o[12295] = i[3975];
  assign o[12294] = i[3974];
  assign o[12293] = i[3973];
  assign o[12292] = i[3972];
  assign o[12291] = i[3971];
  assign o[12290] = i[3970];
  assign o[12289] = i[3969];
  assign o[12288] = i[3968];
  assign o[12287] = i[4223];
  assign o[12286] = i[4222];
  assign o[12285] = i[4221];
  assign o[12284] = i[4220];
  assign o[12283] = i[4219];
  assign o[12282] = i[4218];
  assign o[12281] = i[4217];
  assign o[12280] = i[4216];
  assign o[12279] = i[4215];
  assign o[12278] = i[4214];
  assign o[12277] = i[4213];
  assign o[12276] = i[4212];
  assign o[12275] = i[4211];
  assign o[12274] = i[4210];
  assign o[12273] = i[4209];
  assign o[12272] = i[4208];
  assign o[12271] = i[4207];
  assign o[12270] = i[4206];
  assign o[12269] = i[4205];
  assign o[12268] = i[4204];
  assign o[12267] = i[4203];
  assign o[12266] = i[4202];
  assign o[12265] = i[4201];
  assign o[12264] = i[4200];
  assign o[12263] = i[4199];
  assign o[12262] = i[4198];
  assign o[12261] = i[4197];
  assign o[12260] = i[4196];
  assign o[12259] = i[4195];
  assign o[12258] = i[4194];
  assign o[12257] = i[4193];
  assign o[12256] = i[4192];
  assign o[12255] = i[4191];
  assign o[12254] = i[4190];
  assign o[12253] = i[4189];
  assign o[12252] = i[4188];
  assign o[12251] = i[4187];
  assign o[12250] = i[4186];
  assign o[12249] = i[4185];
  assign o[12248] = i[4184];
  assign o[12247] = i[4183];
  assign o[12246] = i[4182];
  assign o[12245] = i[4181];
  assign o[12244] = i[4180];
  assign o[12243] = i[4179];
  assign o[12242] = i[4178];
  assign o[12241] = i[4177];
  assign o[12240] = i[4176];
  assign o[12239] = i[4175];
  assign o[12238] = i[4174];
  assign o[12237] = i[4173];
  assign o[12236] = i[4172];
  assign o[12235] = i[4171];
  assign o[12234] = i[4170];
  assign o[12233] = i[4169];
  assign o[12232] = i[4168];
  assign o[12231] = i[4167];
  assign o[12230] = i[4166];
  assign o[12229] = i[4165];
  assign o[12228] = i[4164];
  assign o[12227] = i[4163];
  assign o[12226] = i[4162];
  assign o[12225] = i[4161];
  assign o[12224] = i[4160];
  assign o[12223] = i[4159];
  assign o[12222] = i[4158];
  assign o[12221] = i[4157];
  assign o[12220] = i[4156];
  assign o[12219] = i[4155];
  assign o[12218] = i[4154];
  assign o[12217] = i[4153];
  assign o[12216] = i[4152];
  assign o[12215] = i[4151];
  assign o[12214] = i[4150];
  assign o[12213] = i[4149];
  assign o[12212] = i[4148];
  assign o[12211] = i[4147];
  assign o[12210] = i[4146];
  assign o[12209] = i[4145];
  assign o[12208] = i[4144];
  assign o[12207] = i[4143];
  assign o[12206] = i[4142];
  assign o[12205] = i[4141];
  assign o[12204] = i[4140];
  assign o[12203] = i[4139];
  assign o[12202] = i[4138];
  assign o[12201] = i[4137];
  assign o[12200] = i[4136];
  assign o[12199] = i[4135];
  assign o[12198] = i[4134];
  assign o[12197] = i[4133];
  assign o[12196] = i[4132];
  assign o[12195] = i[4131];
  assign o[12194] = i[4130];
  assign o[12193] = i[4129];
  assign o[12192] = i[4128];
  assign o[12191] = i[4127];
  assign o[12190] = i[4126];
  assign o[12189] = i[4125];
  assign o[12188] = i[4124];
  assign o[12187] = i[4123];
  assign o[12186] = i[4122];
  assign o[12185] = i[4121];
  assign o[12184] = i[4120];
  assign o[12183] = i[4119];
  assign o[12182] = i[4118];
  assign o[12181] = i[4117];
  assign o[12180] = i[4116];
  assign o[12179] = i[4115];
  assign o[12178] = i[4114];
  assign o[12177] = i[4113];
  assign o[12176] = i[4112];
  assign o[12175] = i[4111];
  assign o[12174] = i[4110];
  assign o[12173] = i[4109];
  assign o[12172] = i[4108];
  assign o[12171] = i[4107];
  assign o[12170] = i[4106];
  assign o[12169] = i[4105];
  assign o[12168] = i[4104];
  assign o[12167] = i[4103];
  assign o[12166] = i[4102];
  assign o[12165] = i[4101];
  assign o[12164] = i[4100];
  assign o[12163] = i[4099];
  assign o[12162] = i[4098];
  assign o[12161] = i[4097];
  assign o[12160] = i[4096];
  assign o[12159] = i[4351];
  assign o[12158] = i[4350];
  assign o[12157] = i[4349];
  assign o[12156] = i[4348];
  assign o[12155] = i[4347];
  assign o[12154] = i[4346];
  assign o[12153] = i[4345];
  assign o[12152] = i[4344];
  assign o[12151] = i[4343];
  assign o[12150] = i[4342];
  assign o[12149] = i[4341];
  assign o[12148] = i[4340];
  assign o[12147] = i[4339];
  assign o[12146] = i[4338];
  assign o[12145] = i[4337];
  assign o[12144] = i[4336];
  assign o[12143] = i[4335];
  assign o[12142] = i[4334];
  assign o[12141] = i[4333];
  assign o[12140] = i[4332];
  assign o[12139] = i[4331];
  assign o[12138] = i[4330];
  assign o[12137] = i[4329];
  assign o[12136] = i[4328];
  assign o[12135] = i[4327];
  assign o[12134] = i[4326];
  assign o[12133] = i[4325];
  assign o[12132] = i[4324];
  assign o[12131] = i[4323];
  assign o[12130] = i[4322];
  assign o[12129] = i[4321];
  assign o[12128] = i[4320];
  assign o[12127] = i[4319];
  assign o[12126] = i[4318];
  assign o[12125] = i[4317];
  assign o[12124] = i[4316];
  assign o[12123] = i[4315];
  assign o[12122] = i[4314];
  assign o[12121] = i[4313];
  assign o[12120] = i[4312];
  assign o[12119] = i[4311];
  assign o[12118] = i[4310];
  assign o[12117] = i[4309];
  assign o[12116] = i[4308];
  assign o[12115] = i[4307];
  assign o[12114] = i[4306];
  assign o[12113] = i[4305];
  assign o[12112] = i[4304];
  assign o[12111] = i[4303];
  assign o[12110] = i[4302];
  assign o[12109] = i[4301];
  assign o[12108] = i[4300];
  assign o[12107] = i[4299];
  assign o[12106] = i[4298];
  assign o[12105] = i[4297];
  assign o[12104] = i[4296];
  assign o[12103] = i[4295];
  assign o[12102] = i[4294];
  assign o[12101] = i[4293];
  assign o[12100] = i[4292];
  assign o[12099] = i[4291];
  assign o[12098] = i[4290];
  assign o[12097] = i[4289];
  assign o[12096] = i[4288];
  assign o[12095] = i[4287];
  assign o[12094] = i[4286];
  assign o[12093] = i[4285];
  assign o[12092] = i[4284];
  assign o[12091] = i[4283];
  assign o[12090] = i[4282];
  assign o[12089] = i[4281];
  assign o[12088] = i[4280];
  assign o[12087] = i[4279];
  assign o[12086] = i[4278];
  assign o[12085] = i[4277];
  assign o[12084] = i[4276];
  assign o[12083] = i[4275];
  assign o[12082] = i[4274];
  assign o[12081] = i[4273];
  assign o[12080] = i[4272];
  assign o[12079] = i[4271];
  assign o[12078] = i[4270];
  assign o[12077] = i[4269];
  assign o[12076] = i[4268];
  assign o[12075] = i[4267];
  assign o[12074] = i[4266];
  assign o[12073] = i[4265];
  assign o[12072] = i[4264];
  assign o[12071] = i[4263];
  assign o[12070] = i[4262];
  assign o[12069] = i[4261];
  assign o[12068] = i[4260];
  assign o[12067] = i[4259];
  assign o[12066] = i[4258];
  assign o[12065] = i[4257];
  assign o[12064] = i[4256];
  assign o[12063] = i[4255];
  assign o[12062] = i[4254];
  assign o[12061] = i[4253];
  assign o[12060] = i[4252];
  assign o[12059] = i[4251];
  assign o[12058] = i[4250];
  assign o[12057] = i[4249];
  assign o[12056] = i[4248];
  assign o[12055] = i[4247];
  assign o[12054] = i[4246];
  assign o[12053] = i[4245];
  assign o[12052] = i[4244];
  assign o[12051] = i[4243];
  assign o[12050] = i[4242];
  assign o[12049] = i[4241];
  assign o[12048] = i[4240];
  assign o[12047] = i[4239];
  assign o[12046] = i[4238];
  assign o[12045] = i[4237];
  assign o[12044] = i[4236];
  assign o[12043] = i[4235];
  assign o[12042] = i[4234];
  assign o[12041] = i[4233];
  assign o[12040] = i[4232];
  assign o[12039] = i[4231];
  assign o[12038] = i[4230];
  assign o[12037] = i[4229];
  assign o[12036] = i[4228];
  assign o[12035] = i[4227];
  assign o[12034] = i[4226];
  assign o[12033] = i[4225];
  assign o[12032] = i[4224];
  assign o[12031] = i[4479];
  assign o[12030] = i[4478];
  assign o[12029] = i[4477];
  assign o[12028] = i[4476];
  assign o[12027] = i[4475];
  assign o[12026] = i[4474];
  assign o[12025] = i[4473];
  assign o[12024] = i[4472];
  assign o[12023] = i[4471];
  assign o[12022] = i[4470];
  assign o[12021] = i[4469];
  assign o[12020] = i[4468];
  assign o[12019] = i[4467];
  assign o[12018] = i[4466];
  assign o[12017] = i[4465];
  assign o[12016] = i[4464];
  assign o[12015] = i[4463];
  assign o[12014] = i[4462];
  assign o[12013] = i[4461];
  assign o[12012] = i[4460];
  assign o[12011] = i[4459];
  assign o[12010] = i[4458];
  assign o[12009] = i[4457];
  assign o[12008] = i[4456];
  assign o[12007] = i[4455];
  assign o[12006] = i[4454];
  assign o[12005] = i[4453];
  assign o[12004] = i[4452];
  assign o[12003] = i[4451];
  assign o[12002] = i[4450];
  assign o[12001] = i[4449];
  assign o[12000] = i[4448];
  assign o[11999] = i[4447];
  assign o[11998] = i[4446];
  assign o[11997] = i[4445];
  assign o[11996] = i[4444];
  assign o[11995] = i[4443];
  assign o[11994] = i[4442];
  assign o[11993] = i[4441];
  assign o[11992] = i[4440];
  assign o[11991] = i[4439];
  assign o[11990] = i[4438];
  assign o[11989] = i[4437];
  assign o[11988] = i[4436];
  assign o[11987] = i[4435];
  assign o[11986] = i[4434];
  assign o[11985] = i[4433];
  assign o[11984] = i[4432];
  assign o[11983] = i[4431];
  assign o[11982] = i[4430];
  assign o[11981] = i[4429];
  assign o[11980] = i[4428];
  assign o[11979] = i[4427];
  assign o[11978] = i[4426];
  assign o[11977] = i[4425];
  assign o[11976] = i[4424];
  assign o[11975] = i[4423];
  assign o[11974] = i[4422];
  assign o[11973] = i[4421];
  assign o[11972] = i[4420];
  assign o[11971] = i[4419];
  assign o[11970] = i[4418];
  assign o[11969] = i[4417];
  assign o[11968] = i[4416];
  assign o[11967] = i[4415];
  assign o[11966] = i[4414];
  assign o[11965] = i[4413];
  assign o[11964] = i[4412];
  assign o[11963] = i[4411];
  assign o[11962] = i[4410];
  assign o[11961] = i[4409];
  assign o[11960] = i[4408];
  assign o[11959] = i[4407];
  assign o[11958] = i[4406];
  assign o[11957] = i[4405];
  assign o[11956] = i[4404];
  assign o[11955] = i[4403];
  assign o[11954] = i[4402];
  assign o[11953] = i[4401];
  assign o[11952] = i[4400];
  assign o[11951] = i[4399];
  assign o[11950] = i[4398];
  assign o[11949] = i[4397];
  assign o[11948] = i[4396];
  assign o[11947] = i[4395];
  assign o[11946] = i[4394];
  assign o[11945] = i[4393];
  assign o[11944] = i[4392];
  assign o[11943] = i[4391];
  assign o[11942] = i[4390];
  assign o[11941] = i[4389];
  assign o[11940] = i[4388];
  assign o[11939] = i[4387];
  assign o[11938] = i[4386];
  assign o[11937] = i[4385];
  assign o[11936] = i[4384];
  assign o[11935] = i[4383];
  assign o[11934] = i[4382];
  assign o[11933] = i[4381];
  assign o[11932] = i[4380];
  assign o[11931] = i[4379];
  assign o[11930] = i[4378];
  assign o[11929] = i[4377];
  assign o[11928] = i[4376];
  assign o[11927] = i[4375];
  assign o[11926] = i[4374];
  assign o[11925] = i[4373];
  assign o[11924] = i[4372];
  assign o[11923] = i[4371];
  assign o[11922] = i[4370];
  assign o[11921] = i[4369];
  assign o[11920] = i[4368];
  assign o[11919] = i[4367];
  assign o[11918] = i[4366];
  assign o[11917] = i[4365];
  assign o[11916] = i[4364];
  assign o[11915] = i[4363];
  assign o[11914] = i[4362];
  assign o[11913] = i[4361];
  assign o[11912] = i[4360];
  assign o[11911] = i[4359];
  assign o[11910] = i[4358];
  assign o[11909] = i[4357];
  assign o[11908] = i[4356];
  assign o[11907] = i[4355];
  assign o[11906] = i[4354];
  assign o[11905] = i[4353];
  assign o[11904] = i[4352];
  assign o[11903] = i[4607];
  assign o[11902] = i[4606];
  assign o[11901] = i[4605];
  assign o[11900] = i[4604];
  assign o[11899] = i[4603];
  assign o[11898] = i[4602];
  assign o[11897] = i[4601];
  assign o[11896] = i[4600];
  assign o[11895] = i[4599];
  assign o[11894] = i[4598];
  assign o[11893] = i[4597];
  assign o[11892] = i[4596];
  assign o[11891] = i[4595];
  assign o[11890] = i[4594];
  assign o[11889] = i[4593];
  assign o[11888] = i[4592];
  assign o[11887] = i[4591];
  assign o[11886] = i[4590];
  assign o[11885] = i[4589];
  assign o[11884] = i[4588];
  assign o[11883] = i[4587];
  assign o[11882] = i[4586];
  assign o[11881] = i[4585];
  assign o[11880] = i[4584];
  assign o[11879] = i[4583];
  assign o[11878] = i[4582];
  assign o[11877] = i[4581];
  assign o[11876] = i[4580];
  assign o[11875] = i[4579];
  assign o[11874] = i[4578];
  assign o[11873] = i[4577];
  assign o[11872] = i[4576];
  assign o[11871] = i[4575];
  assign o[11870] = i[4574];
  assign o[11869] = i[4573];
  assign o[11868] = i[4572];
  assign o[11867] = i[4571];
  assign o[11866] = i[4570];
  assign o[11865] = i[4569];
  assign o[11864] = i[4568];
  assign o[11863] = i[4567];
  assign o[11862] = i[4566];
  assign o[11861] = i[4565];
  assign o[11860] = i[4564];
  assign o[11859] = i[4563];
  assign o[11858] = i[4562];
  assign o[11857] = i[4561];
  assign o[11856] = i[4560];
  assign o[11855] = i[4559];
  assign o[11854] = i[4558];
  assign o[11853] = i[4557];
  assign o[11852] = i[4556];
  assign o[11851] = i[4555];
  assign o[11850] = i[4554];
  assign o[11849] = i[4553];
  assign o[11848] = i[4552];
  assign o[11847] = i[4551];
  assign o[11846] = i[4550];
  assign o[11845] = i[4549];
  assign o[11844] = i[4548];
  assign o[11843] = i[4547];
  assign o[11842] = i[4546];
  assign o[11841] = i[4545];
  assign o[11840] = i[4544];
  assign o[11839] = i[4543];
  assign o[11838] = i[4542];
  assign o[11837] = i[4541];
  assign o[11836] = i[4540];
  assign o[11835] = i[4539];
  assign o[11834] = i[4538];
  assign o[11833] = i[4537];
  assign o[11832] = i[4536];
  assign o[11831] = i[4535];
  assign o[11830] = i[4534];
  assign o[11829] = i[4533];
  assign o[11828] = i[4532];
  assign o[11827] = i[4531];
  assign o[11826] = i[4530];
  assign o[11825] = i[4529];
  assign o[11824] = i[4528];
  assign o[11823] = i[4527];
  assign o[11822] = i[4526];
  assign o[11821] = i[4525];
  assign o[11820] = i[4524];
  assign o[11819] = i[4523];
  assign o[11818] = i[4522];
  assign o[11817] = i[4521];
  assign o[11816] = i[4520];
  assign o[11815] = i[4519];
  assign o[11814] = i[4518];
  assign o[11813] = i[4517];
  assign o[11812] = i[4516];
  assign o[11811] = i[4515];
  assign o[11810] = i[4514];
  assign o[11809] = i[4513];
  assign o[11808] = i[4512];
  assign o[11807] = i[4511];
  assign o[11806] = i[4510];
  assign o[11805] = i[4509];
  assign o[11804] = i[4508];
  assign o[11803] = i[4507];
  assign o[11802] = i[4506];
  assign o[11801] = i[4505];
  assign o[11800] = i[4504];
  assign o[11799] = i[4503];
  assign o[11798] = i[4502];
  assign o[11797] = i[4501];
  assign o[11796] = i[4500];
  assign o[11795] = i[4499];
  assign o[11794] = i[4498];
  assign o[11793] = i[4497];
  assign o[11792] = i[4496];
  assign o[11791] = i[4495];
  assign o[11790] = i[4494];
  assign o[11789] = i[4493];
  assign o[11788] = i[4492];
  assign o[11787] = i[4491];
  assign o[11786] = i[4490];
  assign o[11785] = i[4489];
  assign o[11784] = i[4488];
  assign o[11783] = i[4487];
  assign o[11782] = i[4486];
  assign o[11781] = i[4485];
  assign o[11780] = i[4484];
  assign o[11779] = i[4483];
  assign o[11778] = i[4482];
  assign o[11777] = i[4481];
  assign o[11776] = i[4480];
  assign o[11775] = i[4735];
  assign o[11774] = i[4734];
  assign o[11773] = i[4733];
  assign o[11772] = i[4732];
  assign o[11771] = i[4731];
  assign o[11770] = i[4730];
  assign o[11769] = i[4729];
  assign o[11768] = i[4728];
  assign o[11767] = i[4727];
  assign o[11766] = i[4726];
  assign o[11765] = i[4725];
  assign o[11764] = i[4724];
  assign o[11763] = i[4723];
  assign o[11762] = i[4722];
  assign o[11761] = i[4721];
  assign o[11760] = i[4720];
  assign o[11759] = i[4719];
  assign o[11758] = i[4718];
  assign o[11757] = i[4717];
  assign o[11756] = i[4716];
  assign o[11755] = i[4715];
  assign o[11754] = i[4714];
  assign o[11753] = i[4713];
  assign o[11752] = i[4712];
  assign o[11751] = i[4711];
  assign o[11750] = i[4710];
  assign o[11749] = i[4709];
  assign o[11748] = i[4708];
  assign o[11747] = i[4707];
  assign o[11746] = i[4706];
  assign o[11745] = i[4705];
  assign o[11744] = i[4704];
  assign o[11743] = i[4703];
  assign o[11742] = i[4702];
  assign o[11741] = i[4701];
  assign o[11740] = i[4700];
  assign o[11739] = i[4699];
  assign o[11738] = i[4698];
  assign o[11737] = i[4697];
  assign o[11736] = i[4696];
  assign o[11735] = i[4695];
  assign o[11734] = i[4694];
  assign o[11733] = i[4693];
  assign o[11732] = i[4692];
  assign o[11731] = i[4691];
  assign o[11730] = i[4690];
  assign o[11729] = i[4689];
  assign o[11728] = i[4688];
  assign o[11727] = i[4687];
  assign o[11726] = i[4686];
  assign o[11725] = i[4685];
  assign o[11724] = i[4684];
  assign o[11723] = i[4683];
  assign o[11722] = i[4682];
  assign o[11721] = i[4681];
  assign o[11720] = i[4680];
  assign o[11719] = i[4679];
  assign o[11718] = i[4678];
  assign o[11717] = i[4677];
  assign o[11716] = i[4676];
  assign o[11715] = i[4675];
  assign o[11714] = i[4674];
  assign o[11713] = i[4673];
  assign o[11712] = i[4672];
  assign o[11711] = i[4671];
  assign o[11710] = i[4670];
  assign o[11709] = i[4669];
  assign o[11708] = i[4668];
  assign o[11707] = i[4667];
  assign o[11706] = i[4666];
  assign o[11705] = i[4665];
  assign o[11704] = i[4664];
  assign o[11703] = i[4663];
  assign o[11702] = i[4662];
  assign o[11701] = i[4661];
  assign o[11700] = i[4660];
  assign o[11699] = i[4659];
  assign o[11698] = i[4658];
  assign o[11697] = i[4657];
  assign o[11696] = i[4656];
  assign o[11695] = i[4655];
  assign o[11694] = i[4654];
  assign o[11693] = i[4653];
  assign o[11692] = i[4652];
  assign o[11691] = i[4651];
  assign o[11690] = i[4650];
  assign o[11689] = i[4649];
  assign o[11688] = i[4648];
  assign o[11687] = i[4647];
  assign o[11686] = i[4646];
  assign o[11685] = i[4645];
  assign o[11684] = i[4644];
  assign o[11683] = i[4643];
  assign o[11682] = i[4642];
  assign o[11681] = i[4641];
  assign o[11680] = i[4640];
  assign o[11679] = i[4639];
  assign o[11678] = i[4638];
  assign o[11677] = i[4637];
  assign o[11676] = i[4636];
  assign o[11675] = i[4635];
  assign o[11674] = i[4634];
  assign o[11673] = i[4633];
  assign o[11672] = i[4632];
  assign o[11671] = i[4631];
  assign o[11670] = i[4630];
  assign o[11669] = i[4629];
  assign o[11668] = i[4628];
  assign o[11667] = i[4627];
  assign o[11666] = i[4626];
  assign o[11665] = i[4625];
  assign o[11664] = i[4624];
  assign o[11663] = i[4623];
  assign o[11662] = i[4622];
  assign o[11661] = i[4621];
  assign o[11660] = i[4620];
  assign o[11659] = i[4619];
  assign o[11658] = i[4618];
  assign o[11657] = i[4617];
  assign o[11656] = i[4616];
  assign o[11655] = i[4615];
  assign o[11654] = i[4614];
  assign o[11653] = i[4613];
  assign o[11652] = i[4612];
  assign o[11651] = i[4611];
  assign o[11650] = i[4610];
  assign o[11649] = i[4609];
  assign o[11648] = i[4608];
  assign o[11647] = i[4863];
  assign o[11646] = i[4862];
  assign o[11645] = i[4861];
  assign o[11644] = i[4860];
  assign o[11643] = i[4859];
  assign o[11642] = i[4858];
  assign o[11641] = i[4857];
  assign o[11640] = i[4856];
  assign o[11639] = i[4855];
  assign o[11638] = i[4854];
  assign o[11637] = i[4853];
  assign o[11636] = i[4852];
  assign o[11635] = i[4851];
  assign o[11634] = i[4850];
  assign o[11633] = i[4849];
  assign o[11632] = i[4848];
  assign o[11631] = i[4847];
  assign o[11630] = i[4846];
  assign o[11629] = i[4845];
  assign o[11628] = i[4844];
  assign o[11627] = i[4843];
  assign o[11626] = i[4842];
  assign o[11625] = i[4841];
  assign o[11624] = i[4840];
  assign o[11623] = i[4839];
  assign o[11622] = i[4838];
  assign o[11621] = i[4837];
  assign o[11620] = i[4836];
  assign o[11619] = i[4835];
  assign o[11618] = i[4834];
  assign o[11617] = i[4833];
  assign o[11616] = i[4832];
  assign o[11615] = i[4831];
  assign o[11614] = i[4830];
  assign o[11613] = i[4829];
  assign o[11612] = i[4828];
  assign o[11611] = i[4827];
  assign o[11610] = i[4826];
  assign o[11609] = i[4825];
  assign o[11608] = i[4824];
  assign o[11607] = i[4823];
  assign o[11606] = i[4822];
  assign o[11605] = i[4821];
  assign o[11604] = i[4820];
  assign o[11603] = i[4819];
  assign o[11602] = i[4818];
  assign o[11601] = i[4817];
  assign o[11600] = i[4816];
  assign o[11599] = i[4815];
  assign o[11598] = i[4814];
  assign o[11597] = i[4813];
  assign o[11596] = i[4812];
  assign o[11595] = i[4811];
  assign o[11594] = i[4810];
  assign o[11593] = i[4809];
  assign o[11592] = i[4808];
  assign o[11591] = i[4807];
  assign o[11590] = i[4806];
  assign o[11589] = i[4805];
  assign o[11588] = i[4804];
  assign o[11587] = i[4803];
  assign o[11586] = i[4802];
  assign o[11585] = i[4801];
  assign o[11584] = i[4800];
  assign o[11583] = i[4799];
  assign o[11582] = i[4798];
  assign o[11581] = i[4797];
  assign o[11580] = i[4796];
  assign o[11579] = i[4795];
  assign o[11578] = i[4794];
  assign o[11577] = i[4793];
  assign o[11576] = i[4792];
  assign o[11575] = i[4791];
  assign o[11574] = i[4790];
  assign o[11573] = i[4789];
  assign o[11572] = i[4788];
  assign o[11571] = i[4787];
  assign o[11570] = i[4786];
  assign o[11569] = i[4785];
  assign o[11568] = i[4784];
  assign o[11567] = i[4783];
  assign o[11566] = i[4782];
  assign o[11565] = i[4781];
  assign o[11564] = i[4780];
  assign o[11563] = i[4779];
  assign o[11562] = i[4778];
  assign o[11561] = i[4777];
  assign o[11560] = i[4776];
  assign o[11559] = i[4775];
  assign o[11558] = i[4774];
  assign o[11557] = i[4773];
  assign o[11556] = i[4772];
  assign o[11555] = i[4771];
  assign o[11554] = i[4770];
  assign o[11553] = i[4769];
  assign o[11552] = i[4768];
  assign o[11551] = i[4767];
  assign o[11550] = i[4766];
  assign o[11549] = i[4765];
  assign o[11548] = i[4764];
  assign o[11547] = i[4763];
  assign o[11546] = i[4762];
  assign o[11545] = i[4761];
  assign o[11544] = i[4760];
  assign o[11543] = i[4759];
  assign o[11542] = i[4758];
  assign o[11541] = i[4757];
  assign o[11540] = i[4756];
  assign o[11539] = i[4755];
  assign o[11538] = i[4754];
  assign o[11537] = i[4753];
  assign o[11536] = i[4752];
  assign o[11535] = i[4751];
  assign o[11534] = i[4750];
  assign o[11533] = i[4749];
  assign o[11532] = i[4748];
  assign o[11531] = i[4747];
  assign o[11530] = i[4746];
  assign o[11529] = i[4745];
  assign o[11528] = i[4744];
  assign o[11527] = i[4743];
  assign o[11526] = i[4742];
  assign o[11525] = i[4741];
  assign o[11524] = i[4740];
  assign o[11523] = i[4739];
  assign o[11522] = i[4738];
  assign o[11521] = i[4737];
  assign o[11520] = i[4736];
  assign o[11519] = i[4991];
  assign o[11518] = i[4990];
  assign o[11517] = i[4989];
  assign o[11516] = i[4988];
  assign o[11515] = i[4987];
  assign o[11514] = i[4986];
  assign o[11513] = i[4985];
  assign o[11512] = i[4984];
  assign o[11511] = i[4983];
  assign o[11510] = i[4982];
  assign o[11509] = i[4981];
  assign o[11508] = i[4980];
  assign o[11507] = i[4979];
  assign o[11506] = i[4978];
  assign o[11505] = i[4977];
  assign o[11504] = i[4976];
  assign o[11503] = i[4975];
  assign o[11502] = i[4974];
  assign o[11501] = i[4973];
  assign o[11500] = i[4972];
  assign o[11499] = i[4971];
  assign o[11498] = i[4970];
  assign o[11497] = i[4969];
  assign o[11496] = i[4968];
  assign o[11495] = i[4967];
  assign o[11494] = i[4966];
  assign o[11493] = i[4965];
  assign o[11492] = i[4964];
  assign o[11491] = i[4963];
  assign o[11490] = i[4962];
  assign o[11489] = i[4961];
  assign o[11488] = i[4960];
  assign o[11487] = i[4959];
  assign o[11486] = i[4958];
  assign o[11485] = i[4957];
  assign o[11484] = i[4956];
  assign o[11483] = i[4955];
  assign o[11482] = i[4954];
  assign o[11481] = i[4953];
  assign o[11480] = i[4952];
  assign o[11479] = i[4951];
  assign o[11478] = i[4950];
  assign o[11477] = i[4949];
  assign o[11476] = i[4948];
  assign o[11475] = i[4947];
  assign o[11474] = i[4946];
  assign o[11473] = i[4945];
  assign o[11472] = i[4944];
  assign o[11471] = i[4943];
  assign o[11470] = i[4942];
  assign o[11469] = i[4941];
  assign o[11468] = i[4940];
  assign o[11467] = i[4939];
  assign o[11466] = i[4938];
  assign o[11465] = i[4937];
  assign o[11464] = i[4936];
  assign o[11463] = i[4935];
  assign o[11462] = i[4934];
  assign o[11461] = i[4933];
  assign o[11460] = i[4932];
  assign o[11459] = i[4931];
  assign o[11458] = i[4930];
  assign o[11457] = i[4929];
  assign o[11456] = i[4928];
  assign o[11455] = i[4927];
  assign o[11454] = i[4926];
  assign o[11453] = i[4925];
  assign o[11452] = i[4924];
  assign o[11451] = i[4923];
  assign o[11450] = i[4922];
  assign o[11449] = i[4921];
  assign o[11448] = i[4920];
  assign o[11447] = i[4919];
  assign o[11446] = i[4918];
  assign o[11445] = i[4917];
  assign o[11444] = i[4916];
  assign o[11443] = i[4915];
  assign o[11442] = i[4914];
  assign o[11441] = i[4913];
  assign o[11440] = i[4912];
  assign o[11439] = i[4911];
  assign o[11438] = i[4910];
  assign o[11437] = i[4909];
  assign o[11436] = i[4908];
  assign o[11435] = i[4907];
  assign o[11434] = i[4906];
  assign o[11433] = i[4905];
  assign o[11432] = i[4904];
  assign o[11431] = i[4903];
  assign o[11430] = i[4902];
  assign o[11429] = i[4901];
  assign o[11428] = i[4900];
  assign o[11427] = i[4899];
  assign o[11426] = i[4898];
  assign o[11425] = i[4897];
  assign o[11424] = i[4896];
  assign o[11423] = i[4895];
  assign o[11422] = i[4894];
  assign o[11421] = i[4893];
  assign o[11420] = i[4892];
  assign o[11419] = i[4891];
  assign o[11418] = i[4890];
  assign o[11417] = i[4889];
  assign o[11416] = i[4888];
  assign o[11415] = i[4887];
  assign o[11414] = i[4886];
  assign o[11413] = i[4885];
  assign o[11412] = i[4884];
  assign o[11411] = i[4883];
  assign o[11410] = i[4882];
  assign o[11409] = i[4881];
  assign o[11408] = i[4880];
  assign o[11407] = i[4879];
  assign o[11406] = i[4878];
  assign o[11405] = i[4877];
  assign o[11404] = i[4876];
  assign o[11403] = i[4875];
  assign o[11402] = i[4874];
  assign o[11401] = i[4873];
  assign o[11400] = i[4872];
  assign o[11399] = i[4871];
  assign o[11398] = i[4870];
  assign o[11397] = i[4869];
  assign o[11396] = i[4868];
  assign o[11395] = i[4867];
  assign o[11394] = i[4866];
  assign o[11393] = i[4865];
  assign o[11392] = i[4864];
  assign o[11391] = i[5119];
  assign o[11390] = i[5118];
  assign o[11389] = i[5117];
  assign o[11388] = i[5116];
  assign o[11387] = i[5115];
  assign o[11386] = i[5114];
  assign o[11385] = i[5113];
  assign o[11384] = i[5112];
  assign o[11383] = i[5111];
  assign o[11382] = i[5110];
  assign o[11381] = i[5109];
  assign o[11380] = i[5108];
  assign o[11379] = i[5107];
  assign o[11378] = i[5106];
  assign o[11377] = i[5105];
  assign o[11376] = i[5104];
  assign o[11375] = i[5103];
  assign o[11374] = i[5102];
  assign o[11373] = i[5101];
  assign o[11372] = i[5100];
  assign o[11371] = i[5099];
  assign o[11370] = i[5098];
  assign o[11369] = i[5097];
  assign o[11368] = i[5096];
  assign o[11367] = i[5095];
  assign o[11366] = i[5094];
  assign o[11365] = i[5093];
  assign o[11364] = i[5092];
  assign o[11363] = i[5091];
  assign o[11362] = i[5090];
  assign o[11361] = i[5089];
  assign o[11360] = i[5088];
  assign o[11359] = i[5087];
  assign o[11358] = i[5086];
  assign o[11357] = i[5085];
  assign o[11356] = i[5084];
  assign o[11355] = i[5083];
  assign o[11354] = i[5082];
  assign o[11353] = i[5081];
  assign o[11352] = i[5080];
  assign o[11351] = i[5079];
  assign o[11350] = i[5078];
  assign o[11349] = i[5077];
  assign o[11348] = i[5076];
  assign o[11347] = i[5075];
  assign o[11346] = i[5074];
  assign o[11345] = i[5073];
  assign o[11344] = i[5072];
  assign o[11343] = i[5071];
  assign o[11342] = i[5070];
  assign o[11341] = i[5069];
  assign o[11340] = i[5068];
  assign o[11339] = i[5067];
  assign o[11338] = i[5066];
  assign o[11337] = i[5065];
  assign o[11336] = i[5064];
  assign o[11335] = i[5063];
  assign o[11334] = i[5062];
  assign o[11333] = i[5061];
  assign o[11332] = i[5060];
  assign o[11331] = i[5059];
  assign o[11330] = i[5058];
  assign o[11329] = i[5057];
  assign o[11328] = i[5056];
  assign o[11327] = i[5055];
  assign o[11326] = i[5054];
  assign o[11325] = i[5053];
  assign o[11324] = i[5052];
  assign o[11323] = i[5051];
  assign o[11322] = i[5050];
  assign o[11321] = i[5049];
  assign o[11320] = i[5048];
  assign o[11319] = i[5047];
  assign o[11318] = i[5046];
  assign o[11317] = i[5045];
  assign o[11316] = i[5044];
  assign o[11315] = i[5043];
  assign o[11314] = i[5042];
  assign o[11313] = i[5041];
  assign o[11312] = i[5040];
  assign o[11311] = i[5039];
  assign o[11310] = i[5038];
  assign o[11309] = i[5037];
  assign o[11308] = i[5036];
  assign o[11307] = i[5035];
  assign o[11306] = i[5034];
  assign o[11305] = i[5033];
  assign o[11304] = i[5032];
  assign o[11303] = i[5031];
  assign o[11302] = i[5030];
  assign o[11301] = i[5029];
  assign o[11300] = i[5028];
  assign o[11299] = i[5027];
  assign o[11298] = i[5026];
  assign o[11297] = i[5025];
  assign o[11296] = i[5024];
  assign o[11295] = i[5023];
  assign o[11294] = i[5022];
  assign o[11293] = i[5021];
  assign o[11292] = i[5020];
  assign o[11291] = i[5019];
  assign o[11290] = i[5018];
  assign o[11289] = i[5017];
  assign o[11288] = i[5016];
  assign o[11287] = i[5015];
  assign o[11286] = i[5014];
  assign o[11285] = i[5013];
  assign o[11284] = i[5012];
  assign o[11283] = i[5011];
  assign o[11282] = i[5010];
  assign o[11281] = i[5009];
  assign o[11280] = i[5008];
  assign o[11279] = i[5007];
  assign o[11278] = i[5006];
  assign o[11277] = i[5005];
  assign o[11276] = i[5004];
  assign o[11275] = i[5003];
  assign o[11274] = i[5002];
  assign o[11273] = i[5001];
  assign o[11272] = i[5000];
  assign o[11271] = i[4999];
  assign o[11270] = i[4998];
  assign o[11269] = i[4997];
  assign o[11268] = i[4996];
  assign o[11267] = i[4995];
  assign o[11266] = i[4994];
  assign o[11265] = i[4993];
  assign o[11264] = i[4992];
  assign o[11263] = i[5247];
  assign o[11262] = i[5246];
  assign o[11261] = i[5245];
  assign o[11260] = i[5244];
  assign o[11259] = i[5243];
  assign o[11258] = i[5242];
  assign o[11257] = i[5241];
  assign o[11256] = i[5240];
  assign o[11255] = i[5239];
  assign o[11254] = i[5238];
  assign o[11253] = i[5237];
  assign o[11252] = i[5236];
  assign o[11251] = i[5235];
  assign o[11250] = i[5234];
  assign o[11249] = i[5233];
  assign o[11248] = i[5232];
  assign o[11247] = i[5231];
  assign o[11246] = i[5230];
  assign o[11245] = i[5229];
  assign o[11244] = i[5228];
  assign o[11243] = i[5227];
  assign o[11242] = i[5226];
  assign o[11241] = i[5225];
  assign o[11240] = i[5224];
  assign o[11239] = i[5223];
  assign o[11238] = i[5222];
  assign o[11237] = i[5221];
  assign o[11236] = i[5220];
  assign o[11235] = i[5219];
  assign o[11234] = i[5218];
  assign o[11233] = i[5217];
  assign o[11232] = i[5216];
  assign o[11231] = i[5215];
  assign o[11230] = i[5214];
  assign o[11229] = i[5213];
  assign o[11228] = i[5212];
  assign o[11227] = i[5211];
  assign o[11226] = i[5210];
  assign o[11225] = i[5209];
  assign o[11224] = i[5208];
  assign o[11223] = i[5207];
  assign o[11222] = i[5206];
  assign o[11221] = i[5205];
  assign o[11220] = i[5204];
  assign o[11219] = i[5203];
  assign o[11218] = i[5202];
  assign o[11217] = i[5201];
  assign o[11216] = i[5200];
  assign o[11215] = i[5199];
  assign o[11214] = i[5198];
  assign o[11213] = i[5197];
  assign o[11212] = i[5196];
  assign o[11211] = i[5195];
  assign o[11210] = i[5194];
  assign o[11209] = i[5193];
  assign o[11208] = i[5192];
  assign o[11207] = i[5191];
  assign o[11206] = i[5190];
  assign o[11205] = i[5189];
  assign o[11204] = i[5188];
  assign o[11203] = i[5187];
  assign o[11202] = i[5186];
  assign o[11201] = i[5185];
  assign o[11200] = i[5184];
  assign o[11199] = i[5183];
  assign o[11198] = i[5182];
  assign o[11197] = i[5181];
  assign o[11196] = i[5180];
  assign o[11195] = i[5179];
  assign o[11194] = i[5178];
  assign o[11193] = i[5177];
  assign o[11192] = i[5176];
  assign o[11191] = i[5175];
  assign o[11190] = i[5174];
  assign o[11189] = i[5173];
  assign o[11188] = i[5172];
  assign o[11187] = i[5171];
  assign o[11186] = i[5170];
  assign o[11185] = i[5169];
  assign o[11184] = i[5168];
  assign o[11183] = i[5167];
  assign o[11182] = i[5166];
  assign o[11181] = i[5165];
  assign o[11180] = i[5164];
  assign o[11179] = i[5163];
  assign o[11178] = i[5162];
  assign o[11177] = i[5161];
  assign o[11176] = i[5160];
  assign o[11175] = i[5159];
  assign o[11174] = i[5158];
  assign o[11173] = i[5157];
  assign o[11172] = i[5156];
  assign o[11171] = i[5155];
  assign o[11170] = i[5154];
  assign o[11169] = i[5153];
  assign o[11168] = i[5152];
  assign o[11167] = i[5151];
  assign o[11166] = i[5150];
  assign o[11165] = i[5149];
  assign o[11164] = i[5148];
  assign o[11163] = i[5147];
  assign o[11162] = i[5146];
  assign o[11161] = i[5145];
  assign o[11160] = i[5144];
  assign o[11159] = i[5143];
  assign o[11158] = i[5142];
  assign o[11157] = i[5141];
  assign o[11156] = i[5140];
  assign o[11155] = i[5139];
  assign o[11154] = i[5138];
  assign o[11153] = i[5137];
  assign o[11152] = i[5136];
  assign o[11151] = i[5135];
  assign o[11150] = i[5134];
  assign o[11149] = i[5133];
  assign o[11148] = i[5132];
  assign o[11147] = i[5131];
  assign o[11146] = i[5130];
  assign o[11145] = i[5129];
  assign o[11144] = i[5128];
  assign o[11143] = i[5127];
  assign o[11142] = i[5126];
  assign o[11141] = i[5125];
  assign o[11140] = i[5124];
  assign o[11139] = i[5123];
  assign o[11138] = i[5122];
  assign o[11137] = i[5121];
  assign o[11136] = i[5120];
  assign o[11135] = i[5375];
  assign o[11134] = i[5374];
  assign o[11133] = i[5373];
  assign o[11132] = i[5372];
  assign o[11131] = i[5371];
  assign o[11130] = i[5370];
  assign o[11129] = i[5369];
  assign o[11128] = i[5368];
  assign o[11127] = i[5367];
  assign o[11126] = i[5366];
  assign o[11125] = i[5365];
  assign o[11124] = i[5364];
  assign o[11123] = i[5363];
  assign o[11122] = i[5362];
  assign o[11121] = i[5361];
  assign o[11120] = i[5360];
  assign o[11119] = i[5359];
  assign o[11118] = i[5358];
  assign o[11117] = i[5357];
  assign o[11116] = i[5356];
  assign o[11115] = i[5355];
  assign o[11114] = i[5354];
  assign o[11113] = i[5353];
  assign o[11112] = i[5352];
  assign o[11111] = i[5351];
  assign o[11110] = i[5350];
  assign o[11109] = i[5349];
  assign o[11108] = i[5348];
  assign o[11107] = i[5347];
  assign o[11106] = i[5346];
  assign o[11105] = i[5345];
  assign o[11104] = i[5344];
  assign o[11103] = i[5343];
  assign o[11102] = i[5342];
  assign o[11101] = i[5341];
  assign o[11100] = i[5340];
  assign o[11099] = i[5339];
  assign o[11098] = i[5338];
  assign o[11097] = i[5337];
  assign o[11096] = i[5336];
  assign o[11095] = i[5335];
  assign o[11094] = i[5334];
  assign o[11093] = i[5333];
  assign o[11092] = i[5332];
  assign o[11091] = i[5331];
  assign o[11090] = i[5330];
  assign o[11089] = i[5329];
  assign o[11088] = i[5328];
  assign o[11087] = i[5327];
  assign o[11086] = i[5326];
  assign o[11085] = i[5325];
  assign o[11084] = i[5324];
  assign o[11083] = i[5323];
  assign o[11082] = i[5322];
  assign o[11081] = i[5321];
  assign o[11080] = i[5320];
  assign o[11079] = i[5319];
  assign o[11078] = i[5318];
  assign o[11077] = i[5317];
  assign o[11076] = i[5316];
  assign o[11075] = i[5315];
  assign o[11074] = i[5314];
  assign o[11073] = i[5313];
  assign o[11072] = i[5312];
  assign o[11071] = i[5311];
  assign o[11070] = i[5310];
  assign o[11069] = i[5309];
  assign o[11068] = i[5308];
  assign o[11067] = i[5307];
  assign o[11066] = i[5306];
  assign o[11065] = i[5305];
  assign o[11064] = i[5304];
  assign o[11063] = i[5303];
  assign o[11062] = i[5302];
  assign o[11061] = i[5301];
  assign o[11060] = i[5300];
  assign o[11059] = i[5299];
  assign o[11058] = i[5298];
  assign o[11057] = i[5297];
  assign o[11056] = i[5296];
  assign o[11055] = i[5295];
  assign o[11054] = i[5294];
  assign o[11053] = i[5293];
  assign o[11052] = i[5292];
  assign o[11051] = i[5291];
  assign o[11050] = i[5290];
  assign o[11049] = i[5289];
  assign o[11048] = i[5288];
  assign o[11047] = i[5287];
  assign o[11046] = i[5286];
  assign o[11045] = i[5285];
  assign o[11044] = i[5284];
  assign o[11043] = i[5283];
  assign o[11042] = i[5282];
  assign o[11041] = i[5281];
  assign o[11040] = i[5280];
  assign o[11039] = i[5279];
  assign o[11038] = i[5278];
  assign o[11037] = i[5277];
  assign o[11036] = i[5276];
  assign o[11035] = i[5275];
  assign o[11034] = i[5274];
  assign o[11033] = i[5273];
  assign o[11032] = i[5272];
  assign o[11031] = i[5271];
  assign o[11030] = i[5270];
  assign o[11029] = i[5269];
  assign o[11028] = i[5268];
  assign o[11027] = i[5267];
  assign o[11026] = i[5266];
  assign o[11025] = i[5265];
  assign o[11024] = i[5264];
  assign o[11023] = i[5263];
  assign o[11022] = i[5262];
  assign o[11021] = i[5261];
  assign o[11020] = i[5260];
  assign o[11019] = i[5259];
  assign o[11018] = i[5258];
  assign o[11017] = i[5257];
  assign o[11016] = i[5256];
  assign o[11015] = i[5255];
  assign o[11014] = i[5254];
  assign o[11013] = i[5253];
  assign o[11012] = i[5252];
  assign o[11011] = i[5251];
  assign o[11010] = i[5250];
  assign o[11009] = i[5249];
  assign o[11008] = i[5248];
  assign o[11007] = i[5503];
  assign o[11006] = i[5502];
  assign o[11005] = i[5501];
  assign o[11004] = i[5500];
  assign o[11003] = i[5499];
  assign o[11002] = i[5498];
  assign o[11001] = i[5497];
  assign o[11000] = i[5496];
  assign o[10999] = i[5495];
  assign o[10998] = i[5494];
  assign o[10997] = i[5493];
  assign o[10996] = i[5492];
  assign o[10995] = i[5491];
  assign o[10994] = i[5490];
  assign o[10993] = i[5489];
  assign o[10992] = i[5488];
  assign o[10991] = i[5487];
  assign o[10990] = i[5486];
  assign o[10989] = i[5485];
  assign o[10988] = i[5484];
  assign o[10987] = i[5483];
  assign o[10986] = i[5482];
  assign o[10985] = i[5481];
  assign o[10984] = i[5480];
  assign o[10983] = i[5479];
  assign o[10982] = i[5478];
  assign o[10981] = i[5477];
  assign o[10980] = i[5476];
  assign o[10979] = i[5475];
  assign o[10978] = i[5474];
  assign o[10977] = i[5473];
  assign o[10976] = i[5472];
  assign o[10975] = i[5471];
  assign o[10974] = i[5470];
  assign o[10973] = i[5469];
  assign o[10972] = i[5468];
  assign o[10971] = i[5467];
  assign o[10970] = i[5466];
  assign o[10969] = i[5465];
  assign o[10968] = i[5464];
  assign o[10967] = i[5463];
  assign o[10966] = i[5462];
  assign o[10965] = i[5461];
  assign o[10964] = i[5460];
  assign o[10963] = i[5459];
  assign o[10962] = i[5458];
  assign o[10961] = i[5457];
  assign o[10960] = i[5456];
  assign o[10959] = i[5455];
  assign o[10958] = i[5454];
  assign o[10957] = i[5453];
  assign o[10956] = i[5452];
  assign o[10955] = i[5451];
  assign o[10954] = i[5450];
  assign o[10953] = i[5449];
  assign o[10952] = i[5448];
  assign o[10951] = i[5447];
  assign o[10950] = i[5446];
  assign o[10949] = i[5445];
  assign o[10948] = i[5444];
  assign o[10947] = i[5443];
  assign o[10946] = i[5442];
  assign o[10945] = i[5441];
  assign o[10944] = i[5440];
  assign o[10943] = i[5439];
  assign o[10942] = i[5438];
  assign o[10941] = i[5437];
  assign o[10940] = i[5436];
  assign o[10939] = i[5435];
  assign o[10938] = i[5434];
  assign o[10937] = i[5433];
  assign o[10936] = i[5432];
  assign o[10935] = i[5431];
  assign o[10934] = i[5430];
  assign o[10933] = i[5429];
  assign o[10932] = i[5428];
  assign o[10931] = i[5427];
  assign o[10930] = i[5426];
  assign o[10929] = i[5425];
  assign o[10928] = i[5424];
  assign o[10927] = i[5423];
  assign o[10926] = i[5422];
  assign o[10925] = i[5421];
  assign o[10924] = i[5420];
  assign o[10923] = i[5419];
  assign o[10922] = i[5418];
  assign o[10921] = i[5417];
  assign o[10920] = i[5416];
  assign o[10919] = i[5415];
  assign o[10918] = i[5414];
  assign o[10917] = i[5413];
  assign o[10916] = i[5412];
  assign o[10915] = i[5411];
  assign o[10914] = i[5410];
  assign o[10913] = i[5409];
  assign o[10912] = i[5408];
  assign o[10911] = i[5407];
  assign o[10910] = i[5406];
  assign o[10909] = i[5405];
  assign o[10908] = i[5404];
  assign o[10907] = i[5403];
  assign o[10906] = i[5402];
  assign o[10905] = i[5401];
  assign o[10904] = i[5400];
  assign o[10903] = i[5399];
  assign o[10902] = i[5398];
  assign o[10901] = i[5397];
  assign o[10900] = i[5396];
  assign o[10899] = i[5395];
  assign o[10898] = i[5394];
  assign o[10897] = i[5393];
  assign o[10896] = i[5392];
  assign o[10895] = i[5391];
  assign o[10894] = i[5390];
  assign o[10893] = i[5389];
  assign o[10892] = i[5388];
  assign o[10891] = i[5387];
  assign o[10890] = i[5386];
  assign o[10889] = i[5385];
  assign o[10888] = i[5384];
  assign o[10887] = i[5383];
  assign o[10886] = i[5382];
  assign o[10885] = i[5381];
  assign o[10884] = i[5380];
  assign o[10883] = i[5379];
  assign o[10882] = i[5378];
  assign o[10881] = i[5377];
  assign o[10880] = i[5376];
  assign o[10879] = i[5631];
  assign o[10878] = i[5630];
  assign o[10877] = i[5629];
  assign o[10876] = i[5628];
  assign o[10875] = i[5627];
  assign o[10874] = i[5626];
  assign o[10873] = i[5625];
  assign o[10872] = i[5624];
  assign o[10871] = i[5623];
  assign o[10870] = i[5622];
  assign o[10869] = i[5621];
  assign o[10868] = i[5620];
  assign o[10867] = i[5619];
  assign o[10866] = i[5618];
  assign o[10865] = i[5617];
  assign o[10864] = i[5616];
  assign o[10863] = i[5615];
  assign o[10862] = i[5614];
  assign o[10861] = i[5613];
  assign o[10860] = i[5612];
  assign o[10859] = i[5611];
  assign o[10858] = i[5610];
  assign o[10857] = i[5609];
  assign o[10856] = i[5608];
  assign o[10855] = i[5607];
  assign o[10854] = i[5606];
  assign o[10853] = i[5605];
  assign o[10852] = i[5604];
  assign o[10851] = i[5603];
  assign o[10850] = i[5602];
  assign o[10849] = i[5601];
  assign o[10848] = i[5600];
  assign o[10847] = i[5599];
  assign o[10846] = i[5598];
  assign o[10845] = i[5597];
  assign o[10844] = i[5596];
  assign o[10843] = i[5595];
  assign o[10842] = i[5594];
  assign o[10841] = i[5593];
  assign o[10840] = i[5592];
  assign o[10839] = i[5591];
  assign o[10838] = i[5590];
  assign o[10837] = i[5589];
  assign o[10836] = i[5588];
  assign o[10835] = i[5587];
  assign o[10834] = i[5586];
  assign o[10833] = i[5585];
  assign o[10832] = i[5584];
  assign o[10831] = i[5583];
  assign o[10830] = i[5582];
  assign o[10829] = i[5581];
  assign o[10828] = i[5580];
  assign o[10827] = i[5579];
  assign o[10826] = i[5578];
  assign o[10825] = i[5577];
  assign o[10824] = i[5576];
  assign o[10823] = i[5575];
  assign o[10822] = i[5574];
  assign o[10821] = i[5573];
  assign o[10820] = i[5572];
  assign o[10819] = i[5571];
  assign o[10818] = i[5570];
  assign o[10817] = i[5569];
  assign o[10816] = i[5568];
  assign o[10815] = i[5567];
  assign o[10814] = i[5566];
  assign o[10813] = i[5565];
  assign o[10812] = i[5564];
  assign o[10811] = i[5563];
  assign o[10810] = i[5562];
  assign o[10809] = i[5561];
  assign o[10808] = i[5560];
  assign o[10807] = i[5559];
  assign o[10806] = i[5558];
  assign o[10805] = i[5557];
  assign o[10804] = i[5556];
  assign o[10803] = i[5555];
  assign o[10802] = i[5554];
  assign o[10801] = i[5553];
  assign o[10800] = i[5552];
  assign o[10799] = i[5551];
  assign o[10798] = i[5550];
  assign o[10797] = i[5549];
  assign o[10796] = i[5548];
  assign o[10795] = i[5547];
  assign o[10794] = i[5546];
  assign o[10793] = i[5545];
  assign o[10792] = i[5544];
  assign o[10791] = i[5543];
  assign o[10790] = i[5542];
  assign o[10789] = i[5541];
  assign o[10788] = i[5540];
  assign o[10787] = i[5539];
  assign o[10786] = i[5538];
  assign o[10785] = i[5537];
  assign o[10784] = i[5536];
  assign o[10783] = i[5535];
  assign o[10782] = i[5534];
  assign o[10781] = i[5533];
  assign o[10780] = i[5532];
  assign o[10779] = i[5531];
  assign o[10778] = i[5530];
  assign o[10777] = i[5529];
  assign o[10776] = i[5528];
  assign o[10775] = i[5527];
  assign o[10774] = i[5526];
  assign o[10773] = i[5525];
  assign o[10772] = i[5524];
  assign o[10771] = i[5523];
  assign o[10770] = i[5522];
  assign o[10769] = i[5521];
  assign o[10768] = i[5520];
  assign o[10767] = i[5519];
  assign o[10766] = i[5518];
  assign o[10765] = i[5517];
  assign o[10764] = i[5516];
  assign o[10763] = i[5515];
  assign o[10762] = i[5514];
  assign o[10761] = i[5513];
  assign o[10760] = i[5512];
  assign o[10759] = i[5511];
  assign o[10758] = i[5510];
  assign o[10757] = i[5509];
  assign o[10756] = i[5508];
  assign o[10755] = i[5507];
  assign o[10754] = i[5506];
  assign o[10753] = i[5505];
  assign o[10752] = i[5504];
  assign o[10751] = i[5759];
  assign o[10750] = i[5758];
  assign o[10749] = i[5757];
  assign o[10748] = i[5756];
  assign o[10747] = i[5755];
  assign o[10746] = i[5754];
  assign o[10745] = i[5753];
  assign o[10744] = i[5752];
  assign o[10743] = i[5751];
  assign o[10742] = i[5750];
  assign o[10741] = i[5749];
  assign o[10740] = i[5748];
  assign o[10739] = i[5747];
  assign o[10738] = i[5746];
  assign o[10737] = i[5745];
  assign o[10736] = i[5744];
  assign o[10735] = i[5743];
  assign o[10734] = i[5742];
  assign o[10733] = i[5741];
  assign o[10732] = i[5740];
  assign o[10731] = i[5739];
  assign o[10730] = i[5738];
  assign o[10729] = i[5737];
  assign o[10728] = i[5736];
  assign o[10727] = i[5735];
  assign o[10726] = i[5734];
  assign o[10725] = i[5733];
  assign o[10724] = i[5732];
  assign o[10723] = i[5731];
  assign o[10722] = i[5730];
  assign o[10721] = i[5729];
  assign o[10720] = i[5728];
  assign o[10719] = i[5727];
  assign o[10718] = i[5726];
  assign o[10717] = i[5725];
  assign o[10716] = i[5724];
  assign o[10715] = i[5723];
  assign o[10714] = i[5722];
  assign o[10713] = i[5721];
  assign o[10712] = i[5720];
  assign o[10711] = i[5719];
  assign o[10710] = i[5718];
  assign o[10709] = i[5717];
  assign o[10708] = i[5716];
  assign o[10707] = i[5715];
  assign o[10706] = i[5714];
  assign o[10705] = i[5713];
  assign o[10704] = i[5712];
  assign o[10703] = i[5711];
  assign o[10702] = i[5710];
  assign o[10701] = i[5709];
  assign o[10700] = i[5708];
  assign o[10699] = i[5707];
  assign o[10698] = i[5706];
  assign o[10697] = i[5705];
  assign o[10696] = i[5704];
  assign o[10695] = i[5703];
  assign o[10694] = i[5702];
  assign o[10693] = i[5701];
  assign o[10692] = i[5700];
  assign o[10691] = i[5699];
  assign o[10690] = i[5698];
  assign o[10689] = i[5697];
  assign o[10688] = i[5696];
  assign o[10687] = i[5695];
  assign o[10686] = i[5694];
  assign o[10685] = i[5693];
  assign o[10684] = i[5692];
  assign o[10683] = i[5691];
  assign o[10682] = i[5690];
  assign o[10681] = i[5689];
  assign o[10680] = i[5688];
  assign o[10679] = i[5687];
  assign o[10678] = i[5686];
  assign o[10677] = i[5685];
  assign o[10676] = i[5684];
  assign o[10675] = i[5683];
  assign o[10674] = i[5682];
  assign o[10673] = i[5681];
  assign o[10672] = i[5680];
  assign o[10671] = i[5679];
  assign o[10670] = i[5678];
  assign o[10669] = i[5677];
  assign o[10668] = i[5676];
  assign o[10667] = i[5675];
  assign o[10666] = i[5674];
  assign o[10665] = i[5673];
  assign o[10664] = i[5672];
  assign o[10663] = i[5671];
  assign o[10662] = i[5670];
  assign o[10661] = i[5669];
  assign o[10660] = i[5668];
  assign o[10659] = i[5667];
  assign o[10658] = i[5666];
  assign o[10657] = i[5665];
  assign o[10656] = i[5664];
  assign o[10655] = i[5663];
  assign o[10654] = i[5662];
  assign o[10653] = i[5661];
  assign o[10652] = i[5660];
  assign o[10651] = i[5659];
  assign o[10650] = i[5658];
  assign o[10649] = i[5657];
  assign o[10648] = i[5656];
  assign o[10647] = i[5655];
  assign o[10646] = i[5654];
  assign o[10645] = i[5653];
  assign o[10644] = i[5652];
  assign o[10643] = i[5651];
  assign o[10642] = i[5650];
  assign o[10641] = i[5649];
  assign o[10640] = i[5648];
  assign o[10639] = i[5647];
  assign o[10638] = i[5646];
  assign o[10637] = i[5645];
  assign o[10636] = i[5644];
  assign o[10635] = i[5643];
  assign o[10634] = i[5642];
  assign o[10633] = i[5641];
  assign o[10632] = i[5640];
  assign o[10631] = i[5639];
  assign o[10630] = i[5638];
  assign o[10629] = i[5637];
  assign o[10628] = i[5636];
  assign o[10627] = i[5635];
  assign o[10626] = i[5634];
  assign o[10625] = i[5633];
  assign o[10624] = i[5632];
  assign o[10623] = i[5887];
  assign o[10622] = i[5886];
  assign o[10621] = i[5885];
  assign o[10620] = i[5884];
  assign o[10619] = i[5883];
  assign o[10618] = i[5882];
  assign o[10617] = i[5881];
  assign o[10616] = i[5880];
  assign o[10615] = i[5879];
  assign o[10614] = i[5878];
  assign o[10613] = i[5877];
  assign o[10612] = i[5876];
  assign o[10611] = i[5875];
  assign o[10610] = i[5874];
  assign o[10609] = i[5873];
  assign o[10608] = i[5872];
  assign o[10607] = i[5871];
  assign o[10606] = i[5870];
  assign o[10605] = i[5869];
  assign o[10604] = i[5868];
  assign o[10603] = i[5867];
  assign o[10602] = i[5866];
  assign o[10601] = i[5865];
  assign o[10600] = i[5864];
  assign o[10599] = i[5863];
  assign o[10598] = i[5862];
  assign o[10597] = i[5861];
  assign o[10596] = i[5860];
  assign o[10595] = i[5859];
  assign o[10594] = i[5858];
  assign o[10593] = i[5857];
  assign o[10592] = i[5856];
  assign o[10591] = i[5855];
  assign o[10590] = i[5854];
  assign o[10589] = i[5853];
  assign o[10588] = i[5852];
  assign o[10587] = i[5851];
  assign o[10586] = i[5850];
  assign o[10585] = i[5849];
  assign o[10584] = i[5848];
  assign o[10583] = i[5847];
  assign o[10582] = i[5846];
  assign o[10581] = i[5845];
  assign o[10580] = i[5844];
  assign o[10579] = i[5843];
  assign o[10578] = i[5842];
  assign o[10577] = i[5841];
  assign o[10576] = i[5840];
  assign o[10575] = i[5839];
  assign o[10574] = i[5838];
  assign o[10573] = i[5837];
  assign o[10572] = i[5836];
  assign o[10571] = i[5835];
  assign o[10570] = i[5834];
  assign o[10569] = i[5833];
  assign o[10568] = i[5832];
  assign o[10567] = i[5831];
  assign o[10566] = i[5830];
  assign o[10565] = i[5829];
  assign o[10564] = i[5828];
  assign o[10563] = i[5827];
  assign o[10562] = i[5826];
  assign o[10561] = i[5825];
  assign o[10560] = i[5824];
  assign o[10559] = i[5823];
  assign o[10558] = i[5822];
  assign o[10557] = i[5821];
  assign o[10556] = i[5820];
  assign o[10555] = i[5819];
  assign o[10554] = i[5818];
  assign o[10553] = i[5817];
  assign o[10552] = i[5816];
  assign o[10551] = i[5815];
  assign o[10550] = i[5814];
  assign o[10549] = i[5813];
  assign o[10548] = i[5812];
  assign o[10547] = i[5811];
  assign o[10546] = i[5810];
  assign o[10545] = i[5809];
  assign o[10544] = i[5808];
  assign o[10543] = i[5807];
  assign o[10542] = i[5806];
  assign o[10541] = i[5805];
  assign o[10540] = i[5804];
  assign o[10539] = i[5803];
  assign o[10538] = i[5802];
  assign o[10537] = i[5801];
  assign o[10536] = i[5800];
  assign o[10535] = i[5799];
  assign o[10534] = i[5798];
  assign o[10533] = i[5797];
  assign o[10532] = i[5796];
  assign o[10531] = i[5795];
  assign o[10530] = i[5794];
  assign o[10529] = i[5793];
  assign o[10528] = i[5792];
  assign o[10527] = i[5791];
  assign o[10526] = i[5790];
  assign o[10525] = i[5789];
  assign o[10524] = i[5788];
  assign o[10523] = i[5787];
  assign o[10522] = i[5786];
  assign o[10521] = i[5785];
  assign o[10520] = i[5784];
  assign o[10519] = i[5783];
  assign o[10518] = i[5782];
  assign o[10517] = i[5781];
  assign o[10516] = i[5780];
  assign o[10515] = i[5779];
  assign o[10514] = i[5778];
  assign o[10513] = i[5777];
  assign o[10512] = i[5776];
  assign o[10511] = i[5775];
  assign o[10510] = i[5774];
  assign o[10509] = i[5773];
  assign o[10508] = i[5772];
  assign o[10507] = i[5771];
  assign o[10506] = i[5770];
  assign o[10505] = i[5769];
  assign o[10504] = i[5768];
  assign o[10503] = i[5767];
  assign o[10502] = i[5766];
  assign o[10501] = i[5765];
  assign o[10500] = i[5764];
  assign o[10499] = i[5763];
  assign o[10498] = i[5762];
  assign o[10497] = i[5761];
  assign o[10496] = i[5760];
  assign o[10495] = i[6015];
  assign o[10494] = i[6014];
  assign o[10493] = i[6013];
  assign o[10492] = i[6012];
  assign o[10491] = i[6011];
  assign o[10490] = i[6010];
  assign o[10489] = i[6009];
  assign o[10488] = i[6008];
  assign o[10487] = i[6007];
  assign o[10486] = i[6006];
  assign o[10485] = i[6005];
  assign o[10484] = i[6004];
  assign o[10483] = i[6003];
  assign o[10482] = i[6002];
  assign o[10481] = i[6001];
  assign o[10480] = i[6000];
  assign o[10479] = i[5999];
  assign o[10478] = i[5998];
  assign o[10477] = i[5997];
  assign o[10476] = i[5996];
  assign o[10475] = i[5995];
  assign o[10474] = i[5994];
  assign o[10473] = i[5993];
  assign o[10472] = i[5992];
  assign o[10471] = i[5991];
  assign o[10470] = i[5990];
  assign o[10469] = i[5989];
  assign o[10468] = i[5988];
  assign o[10467] = i[5987];
  assign o[10466] = i[5986];
  assign o[10465] = i[5985];
  assign o[10464] = i[5984];
  assign o[10463] = i[5983];
  assign o[10462] = i[5982];
  assign o[10461] = i[5981];
  assign o[10460] = i[5980];
  assign o[10459] = i[5979];
  assign o[10458] = i[5978];
  assign o[10457] = i[5977];
  assign o[10456] = i[5976];
  assign o[10455] = i[5975];
  assign o[10454] = i[5974];
  assign o[10453] = i[5973];
  assign o[10452] = i[5972];
  assign o[10451] = i[5971];
  assign o[10450] = i[5970];
  assign o[10449] = i[5969];
  assign o[10448] = i[5968];
  assign o[10447] = i[5967];
  assign o[10446] = i[5966];
  assign o[10445] = i[5965];
  assign o[10444] = i[5964];
  assign o[10443] = i[5963];
  assign o[10442] = i[5962];
  assign o[10441] = i[5961];
  assign o[10440] = i[5960];
  assign o[10439] = i[5959];
  assign o[10438] = i[5958];
  assign o[10437] = i[5957];
  assign o[10436] = i[5956];
  assign o[10435] = i[5955];
  assign o[10434] = i[5954];
  assign o[10433] = i[5953];
  assign o[10432] = i[5952];
  assign o[10431] = i[5951];
  assign o[10430] = i[5950];
  assign o[10429] = i[5949];
  assign o[10428] = i[5948];
  assign o[10427] = i[5947];
  assign o[10426] = i[5946];
  assign o[10425] = i[5945];
  assign o[10424] = i[5944];
  assign o[10423] = i[5943];
  assign o[10422] = i[5942];
  assign o[10421] = i[5941];
  assign o[10420] = i[5940];
  assign o[10419] = i[5939];
  assign o[10418] = i[5938];
  assign o[10417] = i[5937];
  assign o[10416] = i[5936];
  assign o[10415] = i[5935];
  assign o[10414] = i[5934];
  assign o[10413] = i[5933];
  assign o[10412] = i[5932];
  assign o[10411] = i[5931];
  assign o[10410] = i[5930];
  assign o[10409] = i[5929];
  assign o[10408] = i[5928];
  assign o[10407] = i[5927];
  assign o[10406] = i[5926];
  assign o[10405] = i[5925];
  assign o[10404] = i[5924];
  assign o[10403] = i[5923];
  assign o[10402] = i[5922];
  assign o[10401] = i[5921];
  assign o[10400] = i[5920];
  assign o[10399] = i[5919];
  assign o[10398] = i[5918];
  assign o[10397] = i[5917];
  assign o[10396] = i[5916];
  assign o[10395] = i[5915];
  assign o[10394] = i[5914];
  assign o[10393] = i[5913];
  assign o[10392] = i[5912];
  assign o[10391] = i[5911];
  assign o[10390] = i[5910];
  assign o[10389] = i[5909];
  assign o[10388] = i[5908];
  assign o[10387] = i[5907];
  assign o[10386] = i[5906];
  assign o[10385] = i[5905];
  assign o[10384] = i[5904];
  assign o[10383] = i[5903];
  assign o[10382] = i[5902];
  assign o[10381] = i[5901];
  assign o[10380] = i[5900];
  assign o[10379] = i[5899];
  assign o[10378] = i[5898];
  assign o[10377] = i[5897];
  assign o[10376] = i[5896];
  assign o[10375] = i[5895];
  assign o[10374] = i[5894];
  assign o[10373] = i[5893];
  assign o[10372] = i[5892];
  assign o[10371] = i[5891];
  assign o[10370] = i[5890];
  assign o[10369] = i[5889];
  assign o[10368] = i[5888];
  assign o[10367] = i[6143];
  assign o[10366] = i[6142];
  assign o[10365] = i[6141];
  assign o[10364] = i[6140];
  assign o[10363] = i[6139];
  assign o[10362] = i[6138];
  assign o[10361] = i[6137];
  assign o[10360] = i[6136];
  assign o[10359] = i[6135];
  assign o[10358] = i[6134];
  assign o[10357] = i[6133];
  assign o[10356] = i[6132];
  assign o[10355] = i[6131];
  assign o[10354] = i[6130];
  assign o[10353] = i[6129];
  assign o[10352] = i[6128];
  assign o[10351] = i[6127];
  assign o[10350] = i[6126];
  assign o[10349] = i[6125];
  assign o[10348] = i[6124];
  assign o[10347] = i[6123];
  assign o[10346] = i[6122];
  assign o[10345] = i[6121];
  assign o[10344] = i[6120];
  assign o[10343] = i[6119];
  assign o[10342] = i[6118];
  assign o[10341] = i[6117];
  assign o[10340] = i[6116];
  assign o[10339] = i[6115];
  assign o[10338] = i[6114];
  assign o[10337] = i[6113];
  assign o[10336] = i[6112];
  assign o[10335] = i[6111];
  assign o[10334] = i[6110];
  assign o[10333] = i[6109];
  assign o[10332] = i[6108];
  assign o[10331] = i[6107];
  assign o[10330] = i[6106];
  assign o[10329] = i[6105];
  assign o[10328] = i[6104];
  assign o[10327] = i[6103];
  assign o[10326] = i[6102];
  assign o[10325] = i[6101];
  assign o[10324] = i[6100];
  assign o[10323] = i[6099];
  assign o[10322] = i[6098];
  assign o[10321] = i[6097];
  assign o[10320] = i[6096];
  assign o[10319] = i[6095];
  assign o[10318] = i[6094];
  assign o[10317] = i[6093];
  assign o[10316] = i[6092];
  assign o[10315] = i[6091];
  assign o[10314] = i[6090];
  assign o[10313] = i[6089];
  assign o[10312] = i[6088];
  assign o[10311] = i[6087];
  assign o[10310] = i[6086];
  assign o[10309] = i[6085];
  assign o[10308] = i[6084];
  assign o[10307] = i[6083];
  assign o[10306] = i[6082];
  assign o[10305] = i[6081];
  assign o[10304] = i[6080];
  assign o[10303] = i[6079];
  assign o[10302] = i[6078];
  assign o[10301] = i[6077];
  assign o[10300] = i[6076];
  assign o[10299] = i[6075];
  assign o[10298] = i[6074];
  assign o[10297] = i[6073];
  assign o[10296] = i[6072];
  assign o[10295] = i[6071];
  assign o[10294] = i[6070];
  assign o[10293] = i[6069];
  assign o[10292] = i[6068];
  assign o[10291] = i[6067];
  assign o[10290] = i[6066];
  assign o[10289] = i[6065];
  assign o[10288] = i[6064];
  assign o[10287] = i[6063];
  assign o[10286] = i[6062];
  assign o[10285] = i[6061];
  assign o[10284] = i[6060];
  assign o[10283] = i[6059];
  assign o[10282] = i[6058];
  assign o[10281] = i[6057];
  assign o[10280] = i[6056];
  assign o[10279] = i[6055];
  assign o[10278] = i[6054];
  assign o[10277] = i[6053];
  assign o[10276] = i[6052];
  assign o[10275] = i[6051];
  assign o[10274] = i[6050];
  assign o[10273] = i[6049];
  assign o[10272] = i[6048];
  assign o[10271] = i[6047];
  assign o[10270] = i[6046];
  assign o[10269] = i[6045];
  assign o[10268] = i[6044];
  assign o[10267] = i[6043];
  assign o[10266] = i[6042];
  assign o[10265] = i[6041];
  assign o[10264] = i[6040];
  assign o[10263] = i[6039];
  assign o[10262] = i[6038];
  assign o[10261] = i[6037];
  assign o[10260] = i[6036];
  assign o[10259] = i[6035];
  assign o[10258] = i[6034];
  assign o[10257] = i[6033];
  assign o[10256] = i[6032];
  assign o[10255] = i[6031];
  assign o[10254] = i[6030];
  assign o[10253] = i[6029];
  assign o[10252] = i[6028];
  assign o[10251] = i[6027];
  assign o[10250] = i[6026];
  assign o[10249] = i[6025];
  assign o[10248] = i[6024];
  assign o[10247] = i[6023];
  assign o[10246] = i[6022];
  assign o[10245] = i[6021];
  assign o[10244] = i[6020];
  assign o[10243] = i[6019];
  assign o[10242] = i[6018];
  assign o[10241] = i[6017];
  assign o[10240] = i[6016];
  assign o[10239] = i[6271];
  assign o[10238] = i[6270];
  assign o[10237] = i[6269];
  assign o[10236] = i[6268];
  assign o[10235] = i[6267];
  assign o[10234] = i[6266];
  assign o[10233] = i[6265];
  assign o[10232] = i[6264];
  assign o[10231] = i[6263];
  assign o[10230] = i[6262];
  assign o[10229] = i[6261];
  assign o[10228] = i[6260];
  assign o[10227] = i[6259];
  assign o[10226] = i[6258];
  assign o[10225] = i[6257];
  assign o[10224] = i[6256];
  assign o[10223] = i[6255];
  assign o[10222] = i[6254];
  assign o[10221] = i[6253];
  assign o[10220] = i[6252];
  assign o[10219] = i[6251];
  assign o[10218] = i[6250];
  assign o[10217] = i[6249];
  assign o[10216] = i[6248];
  assign o[10215] = i[6247];
  assign o[10214] = i[6246];
  assign o[10213] = i[6245];
  assign o[10212] = i[6244];
  assign o[10211] = i[6243];
  assign o[10210] = i[6242];
  assign o[10209] = i[6241];
  assign o[10208] = i[6240];
  assign o[10207] = i[6239];
  assign o[10206] = i[6238];
  assign o[10205] = i[6237];
  assign o[10204] = i[6236];
  assign o[10203] = i[6235];
  assign o[10202] = i[6234];
  assign o[10201] = i[6233];
  assign o[10200] = i[6232];
  assign o[10199] = i[6231];
  assign o[10198] = i[6230];
  assign o[10197] = i[6229];
  assign o[10196] = i[6228];
  assign o[10195] = i[6227];
  assign o[10194] = i[6226];
  assign o[10193] = i[6225];
  assign o[10192] = i[6224];
  assign o[10191] = i[6223];
  assign o[10190] = i[6222];
  assign o[10189] = i[6221];
  assign o[10188] = i[6220];
  assign o[10187] = i[6219];
  assign o[10186] = i[6218];
  assign o[10185] = i[6217];
  assign o[10184] = i[6216];
  assign o[10183] = i[6215];
  assign o[10182] = i[6214];
  assign o[10181] = i[6213];
  assign o[10180] = i[6212];
  assign o[10179] = i[6211];
  assign o[10178] = i[6210];
  assign o[10177] = i[6209];
  assign o[10176] = i[6208];
  assign o[10175] = i[6207];
  assign o[10174] = i[6206];
  assign o[10173] = i[6205];
  assign o[10172] = i[6204];
  assign o[10171] = i[6203];
  assign o[10170] = i[6202];
  assign o[10169] = i[6201];
  assign o[10168] = i[6200];
  assign o[10167] = i[6199];
  assign o[10166] = i[6198];
  assign o[10165] = i[6197];
  assign o[10164] = i[6196];
  assign o[10163] = i[6195];
  assign o[10162] = i[6194];
  assign o[10161] = i[6193];
  assign o[10160] = i[6192];
  assign o[10159] = i[6191];
  assign o[10158] = i[6190];
  assign o[10157] = i[6189];
  assign o[10156] = i[6188];
  assign o[10155] = i[6187];
  assign o[10154] = i[6186];
  assign o[10153] = i[6185];
  assign o[10152] = i[6184];
  assign o[10151] = i[6183];
  assign o[10150] = i[6182];
  assign o[10149] = i[6181];
  assign o[10148] = i[6180];
  assign o[10147] = i[6179];
  assign o[10146] = i[6178];
  assign o[10145] = i[6177];
  assign o[10144] = i[6176];
  assign o[10143] = i[6175];
  assign o[10142] = i[6174];
  assign o[10141] = i[6173];
  assign o[10140] = i[6172];
  assign o[10139] = i[6171];
  assign o[10138] = i[6170];
  assign o[10137] = i[6169];
  assign o[10136] = i[6168];
  assign o[10135] = i[6167];
  assign o[10134] = i[6166];
  assign o[10133] = i[6165];
  assign o[10132] = i[6164];
  assign o[10131] = i[6163];
  assign o[10130] = i[6162];
  assign o[10129] = i[6161];
  assign o[10128] = i[6160];
  assign o[10127] = i[6159];
  assign o[10126] = i[6158];
  assign o[10125] = i[6157];
  assign o[10124] = i[6156];
  assign o[10123] = i[6155];
  assign o[10122] = i[6154];
  assign o[10121] = i[6153];
  assign o[10120] = i[6152];
  assign o[10119] = i[6151];
  assign o[10118] = i[6150];
  assign o[10117] = i[6149];
  assign o[10116] = i[6148];
  assign o[10115] = i[6147];
  assign o[10114] = i[6146];
  assign o[10113] = i[6145];
  assign o[10112] = i[6144];
  assign o[10111] = i[6399];
  assign o[10110] = i[6398];
  assign o[10109] = i[6397];
  assign o[10108] = i[6396];
  assign o[10107] = i[6395];
  assign o[10106] = i[6394];
  assign o[10105] = i[6393];
  assign o[10104] = i[6392];
  assign o[10103] = i[6391];
  assign o[10102] = i[6390];
  assign o[10101] = i[6389];
  assign o[10100] = i[6388];
  assign o[10099] = i[6387];
  assign o[10098] = i[6386];
  assign o[10097] = i[6385];
  assign o[10096] = i[6384];
  assign o[10095] = i[6383];
  assign o[10094] = i[6382];
  assign o[10093] = i[6381];
  assign o[10092] = i[6380];
  assign o[10091] = i[6379];
  assign o[10090] = i[6378];
  assign o[10089] = i[6377];
  assign o[10088] = i[6376];
  assign o[10087] = i[6375];
  assign o[10086] = i[6374];
  assign o[10085] = i[6373];
  assign o[10084] = i[6372];
  assign o[10083] = i[6371];
  assign o[10082] = i[6370];
  assign o[10081] = i[6369];
  assign o[10080] = i[6368];
  assign o[10079] = i[6367];
  assign o[10078] = i[6366];
  assign o[10077] = i[6365];
  assign o[10076] = i[6364];
  assign o[10075] = i[6363];
  assign o[10074] = i[6362];
  assign o[10073] = i[6361];
  assign o[10072] = i[6360];
  assign o[10071] = i[6359];
  assign o[10070] = i[6358];
  assign o[10069] = i[6357];
  assign o[10068] = i[6356];
  assign o[10067] = i[6355];
  assign o[10066] = i[6354];
  assign o[10065] = i[6353];
  assign o[10064] = i[6352];
  assign o[10063] = i[6351];
  assign o[10062] = i[6350];
  assign o[10061] = i[6349];
  assign o[10060] = i[6348];
  assign o[10059] = i[6347];
  assign o[10058] = i[6346];
  assign o[10057] = i[6345];
  assign o[10056] = i[6344];
  assign o[10055] = i[6343];
  assign o[10054] = i[6342];
  assign o[10053] = i[6341];
  assign o[10052] = i[6340];
  assign o[10051] = i[6339];
  assign o[10050] = i[6338];
  assign o[10049] = i[6337];
  assign o[10048] = i[6336];
  assign o[10047] = i[6335];
  assign o[10046] = i[6334];
  assign o[10045] = i[6333];
  assign o[10044] = i[6332];
  assign o[10043] = i[6331];
  assign o[10042] = i[6330];
  assign o[10041] = i[6329];
  assign o[10040] = i[6328];
  assign o[10039] = i[6327];
  assign o[10038] = i[6326];
  assign o[10037] = i[6325];
  assign o[10036] = i[6324];
  assign o[10035] = i[6323];
  assign o[10034] = i[6322];
  assign o[10033] = i[6321];
  assign o[10032] = i[6320];
  assign o[10031] = i[6319];
  assign o[10030] = i[6318];
  assign o[10029] = i[6317];
  assign o[10028] = i[6316];
  assign o[10027] = i[6315];
  assign o[10026] = i[6314];
  assign o[10025] = i[6313];
  assign o[10024] = i[6312];
  assign o[10023] = i[6311];
  assign o[10022] = i[6310];
  assign o[10021] = i[6309];
  assign o[10020] = i[6308];
  assign o[10019] = i[6307];
  assign o[10018] = i[6306];
  assign o[10017] = i[6305];
  assign o[10016] = i[6304];
  assign o[10015] = i[6303];
  assign o[10014] = i[6302];
  assign o[10013] = i[6301];
  assign o[10012] = i[6300];
  assign o[10011] = i[6299];
  assign o[10010] = i[6298];
  assign o[10009] = i[6297];
  assign o[10008] = i[6296];
  assign o[10007] = i[6295];
  assign o[10006] = i[6294];
  assign o[10005] = i[6293];
  assign o[10004] = i[6292];
  assign o[10003] = i[6291];
  assign o[10002] = i[6290];
  assign o[10001] = i[6289];
  assign o[10000] = i[6288];
  assign o[9999] = i[6287];
  assign o[9998] = i[6286];
  assign o[9997] = i[6285];
  assign o[9996] = i[6284];
  assign o[9995] = i[6283];
  assign o[9994] = i[6282];
  assign o[9993] = i[6281];
  assign o[9992] = i[6280];
  assign o[9991] = i[6279];
  assign o[9990] = i[6278];
  assign o[9989] = i[6277];
  assign o[9988] = i[6276];
  assign o[9987] = i[6275];
  assign o[9986] = i[6274];
  assign o[9985] = i[6273];
  assign o[9984] = i[6272];
  assign o[9983] = i[6527];
  assign o[9982] = i[6526];
  assign o[9981] = i[6525];
  assign o[9980] = i[6524];
  assign o[9979] = i[6523];
  assign o[9978] = i[6522];
  assign o[9977] = i[6521];
  assign o[9976] = i[6520];
  assign o[9975] = i[6519];
  assign o[9974] = i[6518];
  assign o[9973] = i[6517];
  assign o[9972] = i[6516];
  assign o[9971] = i[6515];
  assign o[9970] = i[6514];
  assign o[9969] = i[6513];
  assign o[9968] = i[6512];
  assign o[9967] = i[6511];
  assign o[9966] = i[6510];
  assign o[9965] = i[6509];
  assign o[9964] = i[6508];
  assign o[9963] = i[6507];
  assign o[9962] = i[6506];
  assign o[9961] = i[6505];
  assign o[9960] = i[6504];
  assign o[9959] = i[6503];
  assign o[9958] = i[6502];
  assign o[9957] = i[6501];
  assign o[9956] = i[6500];
  assign o[9955] = i[6499];
  assign o[9954] = i[6498];
  assign o[9953] = i[6497];
  assign o[9952] = i[6496];
  assign o[9951] = i[6495];
  assign o[9950] = i[6494];
  assign o[9949] = i[6493];
  assign o[9948] = i[6492];
  assign o[9947] = i[6491];
  assign o[9946] = i[6490];
  assign o[9945] = i[6489];
  assign o[9944] = i[6488];
  assign o[9943] = i[6487];
  assign o[9942] = i[6486];
  assign o[9941] = i[6485];
  assign o[9940] = i[6484];
  assign o[9939] = i[6483];
  assign o[9938] = i[6482];
  assign o[9937] = i[6481];
  assign o[9936] = i[6480];
  assign o[9935] = i[6479];
  assign o[9934] = i[6478];
  assign o[9933] = i[6477];
  assign o[9932] = i[6476];
  assign o[9931] = i[6475];
  assign o[9930] = i[6474];
  assign o[9929] = i[6473];
  assign o[9928] = i[6472];
  assign o[9927] = i[6471];
  assign o[9926] = i[6470];
  assign o[9925] = i[6469];
  assign o[9924] = i[6468];
  assign o[9923] = i[6467];
  assign o[9922] = i[6466];
  assign o[9921] = i[6465];
  assign o[9920] = i[6464];
  assign o[9919] = i[6463];
  assign o[9918] = i[6462];
  assign o[9917] = i[6461];
  assign o[9916] = i[6460];
  assign o[9915] = i[6459];
  assign o[9914] = i[6458];
  assign o[9913] = i[6457];
  assign o[9912] = i[6456];
  assign o[9911] = i[6455];
  assign o[9910] = i[6454];
  assign o[9909] = i[6453];
  assign o[9908] = i[6452];
  assign o[9907] = i[6451];
  assign o[9906] = i[6450];
  assign o[9905] = i[6449];
  assign o[9904] = i[6448];
  assign o[9903] = i[6447];
  assign o[9902] = i[6446];
  assign o[9901] = i[6445];
  assign o[9900] = i[6444];
  assign o[9899] = i[6443];
  assign o[9898] = i[6442];
  assign o[9897] = i[6441];
  assign o[9896] = i[6440];
  assign o[9895] = i[6439];
  assign o[9894] = i[6438];
  assign o[9893] = i[6437];
  assign o[9892] = i[6436];
  assign o[9891] = i[6435];
  assign o[9890] = i[6434];
  assign o[9889] = i[6433];
  assign o[9888] = i[6432];
  assign o[9887] = i[6431];
  assign o[9886] = i[6430];
  assign o[9885] = i[6429];
  assign o[9884] = i[6428];
  assign o[9883] = i[6427];
  assign o[9882] = i[6426];
  assign o[9881] = i[6425];
  assign o[9880] = i[6424];
  assign o[9879] = i[6423];
  assign o[9878] = i[6422];
  assign o[9877] = i[6421];
  assign o[9876] = i[6420];
  assign o[9875] = i[6419];
  assign o[9874] = i[6418];
  assign o[9873] = i[6417];
  assign o[9872] = i[6416];
  assign o[9871] = i[6415];
  assign o[9870] = i[6414];
  assign o[9869] = i[6413];
  assign o[9868] = i[6412];
  assign o[9867] = i[6411];
  assign o[9866] = i[6410];
  assign o[9865] = i[6409];
  assign o[9864] = i[6408];
  assign o[9863] = i[6407];
  assign o[9862] = i[6406];
  assign o[9861] = i[6405];
  assign o[9860] = i[6404];
  assign o[9859] = i[6403];
  assign o[9858] = i[6402];
  assign o[9857] = i[6401];
  assign o[9856] = i[6400];
  assign o[9855] = i[6655];
  assign o[9854] = i[6654];
  assign o[9853] = i[6653];
  assign o[9852] = i[6652];
  assign o[9851] = i[6651];
  assign o[9850] = i[6650];
  assign o[9849] = i[6649];
  assign o[9848] = i[6648];
  assign o[9847] = i[6647];
  assign o[9846] = i[6646];
  assign o[9845] = i[6645];
  assign o[9844] = i[6644];
  assign o[9843] = i[6643];
  assign o[9842] = i[6642];
  assign o[9841] = i[6641];
  assign o[9840] = i[6640];
  assign o[9839] = i[6639];
  assign o[9838] = i[6638];
  assign o[9837] = i[6637];
  assign o[9836] = i[6636];
  assign o[9835] = i[6635];
  assign o[9834] = i[6634];
  assign o[9833] = i[6633];
  assign o[9832] = i[6632];
  assign o[9831] = i[6631];
  assign o[9830] = i[6630];
  assign o[9829] = i[6629];
  assign o[9828] = i[6628];
  assign o[9827] = i[6627];
  assign o[9826] = i[6626];
  assign o[9825] = i[6625];
  assign o[9824] = i[6624];
  assign o[9823] = i[6623];
  assign o[9822] = i[6622];
  assign o[9821] = i[6621];
  assign o[9820] = i[6620];
  assign o[9819] = i[6619];
  assign o[9818] = i[6618];
  assign o[9817] = i[6617];
  assign o[9816] = i[6616];
  assign o[9815] = i[6615];
  assign o[9814] = i[6614];
  assign o[9813] = i[6613];
  assign o[9812] = i[6612];
  assign o[9811] = i[6611];
  assign o[9810] = i[6610];
  assign o[9809] = i[6609];
  assign o[9808] = i[6608];
  assign o[9807] = i[6607];
  assign o[9806] = i[6606];
  assign o[9805] = i[6605];
  assign o[9804] = i[6604];
  assign o[9803] = i[6603];
  assign o[9802] = i[6602];
  assign o[9801] = i[6601];
  assign o[9800] = i[6600];
  assign o[9799] = i[6599];
  assign o[9798] = i[6598];
  assign o[9797] = i[6597];
  assign o[9796] = i[6596];
  assign o[9795] = i[6595];
  assign o[9794] = i[6594];
  assign o[9793] = i[6593];
  assign o[9792] = i[6592];
  assign o[9791] = i[6591];
  assign o[9790] = i[6590];
  assign o[9789] = i[6589];
  assign o[9788] = i[6588];
  assign o[9787] = i[6587];
  assign o[9786] = i[6586];
  assign o[9785] = i[6585];
  assign o[9784] = i[6584];
  assign o[9783] = i[6583];
  assign o[9782] = i[6582];
  assign o[9781] = i[6581];
  assign o[9780] = i[6580];
  assign o[9779] = i[6579];
  assign o[9778] = i[6578];
  assign o[9777] = i[6577];
  assign o[9776] = i[6576];
  assign o[9775] = i[6575];
  assign o[9774] = i[6574];
  assign o[9773] = i[6573];
  assign o[9772] = i[6572];
  assign o[9771] = i[6571];
  assign o[9770] = i[6570];
  assign o[9769] = i[6569];
  assign o[9768] = i[6568];
  assign o[9767] = i[6567];
  assign o[9766] = i[6566];
  assign o[9765] = i[6565];
  assign o[9764] = i[6564];
  assign o[9763] = i[6563];
  assign o[9762] = i[6562];
  assign o[9761] = i[6561];
  assign o[9760] = i[6560];
  assign o[9759] = i[6559];
  assign o[9758] = i[6558];
  assign o[9757] = i[6557];
  assign o[9756] = i[6556];
  assign o[9755] = i[6555];
  assign o[9754] = i[6554];
  assign o[9753] = i[6553];
  assign o[9752] = i[6552];
  assign o[9751] = i[6551];
  assign o[9750] = i[6550];
  assign o[9749] = i[6549];
  assign o[9748] = i[6548];
  assign o[9747] = i[6547];
  assign o[9746] = i[6546];
  assign o[9745] = i[6545];
  assign o[9744] = i[6544];
  assign o[9743] = i[6543];
  assign o[9742] = i[6542];
  assign o[9741] = i[6541];
  assign o[9740] = i[6540];
  assign o[9739] = i[6539];
  assign o[9738] = i[6538];
  assign o[9737] = i[6537];
  assign o[9736] = i[6536];
  assign o[9735] = i[6535];
  assign o[9734] = i[6534];
  assign o[9733] = i[6533];
  assign o[9732] = i[6532];
  assign o[9731] = i[6531];
  assign o[9730] = i[6530];
  assign o[9729] = i[6529];
  assign o[9728] = i[6528];
  assign o[9727] = i[6783];
  assign o[9726] = i[6782];
  assign o[9725] = i[6781];
  assign o[9724] = i[6780];
  assign o[9723] = i[6779];
  assign o[9722] = i[6778];
  assign o[9721] = i[6777];
  assign o[9720] = i[6776];
  assign o[9719] = i[6775];
  assign o[9718] = i[6774];
  assign o[9717] = i[6773];
  assign o[9716] = i[6772];
  assign o[9715] = i[6771];
  assign o[9714] = i[6770];
  assign o[9713] = i[6769];
  assign o[9712] = i[6768];
  assign o[9711] = i[6767];
  assign o[9710] = i[6766];
  assign o[9709] = i[6765];
  assign o[9708] = i[6764];
  assign o[9707] = i[6763];
  assign o[9706] = i[6762];
  assign o[9705] = i[6761];
  assign o[9704] = i[6760];
  assign o[9703] = i[6759];
  assign o[9702] = i[6758];
  assign o[9701] = i[6757];
  assign o[9700] = i[6756];
  assign o[9699] = i[6755];
  assign o[9698] = i[6754];
  assign o[9697] = i[6753];
  assign o[9696] = i[6752];
  assign o[9695] = i[6751];
  assign o[9694] = i[6750];
  assign o[9693] = i[6749];
  assign o[9692] = i[6748];
  assign o[9691] = i[6747];
  assign o[9690] = i[6746];
  assign o[9689] = i[6745];
  assign o[9688] = i[6744];
  assign o[9687] = i[6743];
  assign o[9686] = i[6742];
  assign o[9685] = i[6741];
  assign o[9684] = i[6740];
  assign o[9683] = i[6739];
  assign o[9682] = i[6738];
  assign o[9681] = i[6737];
  assign o[9680] = i[6736];
  assign o[9679] = i[6735];
  assign o[9678] = i[6734];
  assign o[9677] = i[6733];
  assign o[9676] = i[6732];
  assign o[9675] = i[6731];
  assign o[9674] = i[6730];
  assign o[9673] = i[6729];
  assign o[9672] = i[6728];
  assign o[9671] = i[6727];
  assign o[9670] = i[6726];
  assign o[9669] = i[6725];
  assign o[9668] = i[6724];
  assign o[9667] = i[6723];
  assign o[9666] = i[6722];
  assign o[9665] = i[6721];
  assign o[9664] = i[6720];
  assign o[9663] = i[6719];
  assign o[9662] = i[6718];
  assign o[9661] = i[6717];
  assign o[9660] = i[6716];
  assign o[9659] = i[6715];
  assign o[9658] = i[6714];
  assign o[9657] = i[6713];
  assign o[9656] = i[6712];
  assign o[9655] = i[6711];
  assign o[9654] = i[6710];
  assign o[9653] = i[6709];
  assign o[9652] = i[6708];
  assign o[9651] = i[6707];
  assign o[9650] = i[6706];
  assign o[9649] = i[6705];
  assign o[9648] = i[6704];
  assign o[9647] = i[6703];
  assign o[9646] = i[6702];
  assign o[9645] = i[6701];
  assign o[9644] = i[6700];
  assign o[9643] = i[6699];
  assign o[9642] = i[6698];
  assign o[9641] = i[6697];
  assign o[9640] = i[6696];
  assign o[9639] = i[6695];
  assign o[9638] = i[6694];
  assign o[9637] = i[6693];
  assign o[9636] = i[6692];
  assign o[9635] = i[6691];
  assign o[9634] = i[6690];
  assign o[9633] = i[6689];
  assign o[9632] = i[6688];
  assign o[9631] = i[6687];
  assign o[9630] = i[6686];
  assign o[9629] = i[6685];
  assign o[9628] = i[6684];
  assign o[9627] = i[6683];
  assign o[9626] = i[6682];
  assign o[9625] = i[6681];
  assign o[9624] = i[6680];
  assign o[9623] = i[6679];
  assign o[9622] = i[6678];
  assign o[9621] = i[6677];
  assign o[9620] = i[6676];
  assign o[9619] = i[6675];
  assign o[9618] = i[6674];
  assign o[9617] = i[6673];
  assign o[9616] = i[6672];
  assign o[9615] = i[6671];
  assign o[9614] = i[6670];
  assign o[9613] = i[6669];
  assign o[9612] = i[6668];
  assign o[9611] = i[6667];
  assign o[9610] = i[6666];
  assign o[9609] = i[6665];
  assign o[9608] = i[6664];
  assign o[9607] = i[6663];
  assign o[9606] = i[6662];
  assign o[9605] = i[6661];
  assign o[9604] = i[6660];
  assign o[9603] = i[6659];
  assign o[9602] = i[6658];
  assign o[9601] = i[6657];
  assign o[9600] = i[6656];
  assign o[9599] = i[6911];
  assign o[9598] = i[6910];
  assign o[9597] = i[6909];
  assign o[9596] = i[6908];
  assign o[9595] = i[6907];
  assign o[9594] = i[6906];
  assign o[9593] = i[6905];
  assign o[9592] = i[6904];
  assign o[9591] = i[6903];
  assign o[9590] = i[6902];
  assign o[9589] = i[6901];
  assign o[9588] = i[6900];
  assign o[9587] = i[6899];
  assign o[9586] = i[6898];
  assign o[9585] = i[6897];
  assign o[9584] = i[6896];
  assign o[9583] = i[6895];
  assign o[9582] = i[6894];
  assign o[9581] = i[6893];
  assign o[9580] = i[6892];
  assign o[9579] = i[6891];
  assign o[9578] = i[6890];
  assign o[9577] = i[6889];
  assign o[9576] = i[6888];
  assign o[9575] = i[6887];
  assign o[9574] = i[6886];
  assign o[9573] = i[6885];
  assign o[9572] = i[6884];
  assign o[9571] = i[6883];
  assign o[9570] = i[6882];
  assign o[9569] = i[6881];
  assign o[9568] = i[6880];
  assign o[9567] = i[6879];
  assign o[9566] = i[6878];
  assign o[9565] = i[6877];
  assign o[9564] = i[6876];
  assign o[9563] = i[6875];
  assign o[9562] = i[6874];
  assign o[9561] = i[6873];
  assign o[9560] = i[6872];
  assign o[9559] = i[6871];
  assign o[9558] = i[6870];
  assign o[9557] = i[6869];
  assign o[9556] = i[6868];
  assign o[9555] = i[6867];
  assign o[9554] = i[6866];
  assign o[9553] = i[6865];
  assign o[9552] = i[6864];
  assign o[9551] = i[6863];
  assign o[9550] = i[6862];
  assign o[9549] = i[6861];
  assign o[9548] = i[6860];
  assign o[9547] = i[6859];
  assign o[9546] = i[6858];
  assign o[9545] = i[6857];
  assign o[9544] = i[6856];
  assign o[9543] = i[6855];
  assign o[9542] = i[6854];
  assign o[9541] = i[6853];
  assign o[9540] = i[6852];
  assign o[9539] = i[6851];
  assign o[9538] = i[6850];
  assign o[9537] = i[6849];
  assign o[9536] = i[6848];
  assign o[9535] = i[6847];
  assign o[9534] = i[6846];
  assign o[9533] = i[6845];
  assign o[9532] = i[6844];
  assign o[9531] = i[6843];
  assign o[9530] = i[6842];
  assign o[9529] = i[6841];
  assign o[9528] = i[6840];
  assign o[9527] = i[6839];
  assign o[9526] = i[6838];
  assign o[9525] = i[6837];
  assign o[9524] = i[6836];
  assign o[9523] = i[6835];
  assign o[9522] = i[6834];
  assign o[9521] = i[6833];
  assign o[9520] = i[6832];
  assign o[9519] = i[6831];
  assign o[9518] = i[6830];
  assign o[9517] = i[6829];
  assign o[9516] = i[6828];
  assign o[9515] = i[6827];
  assign o[9514] = i[6826];
  assign o[9513] = i[6825];
  assign o[9512] = i[6824];
  assign o[9511] = i[6823];
  assign o[9510] = i[6822];
  assign o[9509] = i[6821];
  assign o[9508] = i[6820];
  assign o[9507] = i[6819];
  assign o[9506] = i[6818];
  assign o[9505] = i[6817];
  assign o[9504] = i[6816];
  assign o[9503] = i[6815];
  assign o[9502] = i[6814];
  assign o[9501] = i[6813];
  assign o[9500] = i[6812];
  assign o[9499] = i[6811];
  assign o[9498] = i[6810];
  assign o[9497] = i[6809];
  assign o[9496] = i[6808];
  assign o[9495] = i[6807];
  assign o[9494] = i[6806];
  assign o[9493] = i[6805];
  assign o[9492] = i[6804];
  assign o[9491] = i[6803];
  assign o[9490] = i[6802];
  assign o[9489] = i[6801];
  assign o[9488] = i[6800];
  assign o[9487] = i[6799];
  assign o[9486] = i[6798];
  assign o[9485] = i[6797];
  assign o[9484] = i[6796];
  assign o[9483] = i[6795];
  assign o[9482] = i[6794];
  assign o[9481] = i[6793];
  assign o[9480] = i[6792];
  assign o[9479] = i[6791];
  assign o[9478] = i[6790];
  assign o[9477] = i[6789];
  assign o[9476] = i[6788];
  assign o[9475] = i[6787];
  assign o[9474] = i[6786];
  assign o[9473] = i[6785];
  assign o[9472] = i[6784];
  assign o[9471] = i[7039];
  assign o[9470] = i[7038];
  assign o[9469] = i[7037];
  assign o[9468] = i[7036];
  assign o[9467] = i[7035];
  assign o[9466] = i[7034];
  assign o[9465] = i[7033];
  assign o[9464] = i[7032];
  assign o[9463] = i[7031];
  assign o[9462] = i[7030];
  assign o[9461] = i[7029];
  assign o[9460] = i[7028];
  assign o[9459] = i[7027];
  assign o[9458] = i[7026];
  assign o[9457] = i[7025];
  assign o[9456] = i[7024];
  assign o[9455] = i[7023];
  assign o[9454] = i[7022];
  assign o[9453] = i[7021];
  assign o[9452] = i[7020];
  assign o[9451] = i[7019];
  assign o[9450] = i[7018];
  assign o[9449] = i[7017];
  assign o[9448] = i[7016];
  assign o[9447] = i[7015];
  assign o[9446] = i[7014];
  assign o[9445] = i[7013];
  assign o[9444] = i[7012];
  assign o[9443] = i[7011];
  assign o[9442] = i[7010];
  assign o[9441] = i[7009];
  assign o[9440] = i[7008];
  assign o[9439] = i[7007];
  assign o[9438] = i[7006];
  assign o[9437] = i[7005];
  assign o[9436] = i[7004];
  assign o[9435] = i[7003];
  assign o[9434] = i[7002];
  assign o[9433] = i[7001];
  assign o[9432] = i[7000];
  assign o[9431] = i[6999];
  assign o[9430] = i[6998];
  assign o[9429] = i[6997];
  assign o[9428] = i[6996];
  assign o[9427] = i[6995];
  assign o[9426] = i[6994];
  assign o[9425] = i[6993];
  assign o[9424] = i[6992];
  assign o[9423] = i[6991];
  assign o[9422] = i[6990];
  assign o[9421] = i[6989];
  assign o[9420] = i[6988];
  assign o[9419] = i[6987];
  assign o[9418] = i[6986];
  assign o[9417] = i[6985];
  assign o[9416] = i[6984];
  assign o[9415] = i[6983];
  assign o[9414] = i[6982];
  assign o[9413] = i[6981];
  assign o[9412] = i[6980];
  assign o[9411] = i[6979];
  assign o[9410] = i[6978];
  assign o[9409] = i[6977];
  assign o[9408] = i[6976];
  assign o[9407] = i[6975];
  assign o[9406] = i[6974];
  assign o[9405] = i[6973];
  assign o[9404] = i[6972];
  assign o[9403] = i[6971];
  assign o[9402] = i[6970];
  assign o[9401] = i[6969];
  assign o[9400] = i[6968];
  assign o[9399] = i[6967];
  assign o[9398] = i[6966];
  assign o[9397] = i[6965];
  assign o[9396] = i[6964];
  assign o[9395] = i[6963];
  assign o[9394] = i[6962];
  assign o[9393] = i[6961];
  assign o[9392] = i[6960];
  assign o[9391] = i[6959];
  assign o[9390] = i[6958];
  assign o[9389] = i[6957];
  assign o[9388] = i[6956];
  assign o[9387] = i[6955];
  assign o[9386] = i[6954];
  assign o[9385] = i[6953];
  assign o[9384] = i[6952];
  assign o[9383] = i[6951];
  assign o[9382] = i[6950];
  assign o[9381] = i[6949];
  assign o[9380] = i[6948];
  assign o[9379] = i[6947];
  assign o[9378] = i[6946];
  assign o[9377] = i[6945];
  assign o[9376] = i[6944];
  assign o[9375] = i[6943];
  assign o[9374] = i[6942];
  assign o[9373] = i[6941];
  assign o[9372] = i[6940];
  assign o[9371] = i[6939];
  assign o[9370] = i[6938];
  assign o[9369] = i[6937];
  assign o[9368] = i[6936];
  assign o[9367] = i[6935];
  assign o[9366] = i[6934];
  assign o[9365] = i[6933];
  assign o[9364] = i[6932];
  assign o[9363] = i[6931];
  assign o[9362] = i[6930];
  assign o[9361] = i[6929];
  assign o[9360] = i[6928];
  assign o[9359] = i[6927];
  assign o[9358] = i[6926];
  assign o[9357] = i[6925];
  assign o[9356] = i[6924];
  assign o[9355] = i[6923];
  assign o[9354] = i[6922];
  assign o[9353] = i[6921];
  assign o[9352] = i[6920];
  assign o[9351] = i[6919];
  assign o[9350] = i[6918];
  assign o[9349] = i[6917];
  assign o[9348] = i[6916];
  assign o[9347] = i[6915];
  assign o[9346] = i[6914];
  assign o[9345] = i[6913];
  assign o[9344] = i[6912];
  assign o[9343] = i[7167];
  assign o[9342] = i[7166];
  assign o[9341] = i[7165];
  assign o[9340] = i[7164];
  assign o[9339] = i[7163];
  assign o[9338] = i[7162];
  assign o[9337] = i[7161];
  assign o[9336] = i[7160];
  assign o[9335] = i[7159];
  assign o[9334] = i[7158];
  assign o[9333] = i[7157];
  assign o[9332] = i[7156];
  assign o[9331] = i[7155];
  assign o[9330] = i[7154];
  assign o[9329] = i[7153];
  assign o[9328] = i[7152];
  assign o[9327] = i[7151];
  assign o[9326] = i[7150];
  assign o[9325] = i[7149];
  assign o[9324] = i[7148];
  assign o[9323] = i[7147];
  assign o[9322] = i[7146];
  assign o[9321] = i[7145];
  assign o[9320] = i[7144];
  assign o[9319] = i[7143];
  assign o[9318] = i[7142];
  assign o[9317] = i[7141];
  assign o[9316] = i[7140];
  assign o[9315] = i[7139];
  assign o[9314] = i[7138];
  assign o[9313] = i[7137];
  assign o[9312] = i[7136];
  assign o[9311] = i[7135];
  assign o[9310] = i[7134];
  assign o[9309] = i[7133];
  assign o[9308] = i[7132];
  assign o[9307] = i[7131];
  assign o[9306] = i[7130];
  assign o[9305] = i[7129];
  assign o[9304] = i[7128];
  assign o[9303] = i[7127];
  assign o[9302] = i[7126];
  assign o[9301] = i[7125];
  assign o[9300] = i[7124];
  assign o[9299] = i[7123];
  assign o[9298] = i[7122];
  assign o[9297] = i[7121];
  assign o[9296] = i[7120];
  assign o[9295] = i[7119];
  assign o[9294] = i[7118];
  assign o[9293] = i[7117];
  assign o[9292] = i[7116];
  assign o[9291] = i[7115];
  assign o[9290] = i[7114];
  assign o[9289] = i[7113];
  assign o[9288] = i[7112];
  assign o[9287] = i[7111];
  assign o[9286] = i[7110];
  assign o[9285] = i[7109];
  assign o[9284] = i[7108];
  assign o[9283] = i[7107];
  assign o[9282] = i[7106];
  assign o[9281] = i[7105];
  assign o[9280] = i[7104];
  assign o[9279] = i[7103];
  assign o[9278] = i[7102];
  assign o[9277] = i[7101];
  assign o[9276] = i[7100];
  assign o[9275] = i[7099];
  assign o[9274] = i[7098];
  assign o[9273] = i[7097];
  assign o[9272] = i[7096];
  assign o[9271] = i[7095];
  assign o[9270] = i[7094];
  assign o[9269] = i[7093];
  assign o[9268] = i[7092];
  assign o[9267] = i[7091];
  assign o[9266] = i[7090];
  assign o[9265] = i[7089];
  assign o[9264] = i[7088];
  assign o[9263] = i[7087];
  assign o[9262] = i[7086];
  assign o[9261] = i[7085];
  assign o[9260] = i[7084];
  assign o[9259] = i[7083];
  assign o[9258] = i[7082];
  assign o[9257] = i[7081];
  assign o[9256] = i[7080];
  assign o[9255] = i[7079];
  assign o[9254] = i[7078];
  assign o[9253] = i[7077];
  assign o[9252] = i[7076];
  assign o[9251] = i[7075];
  assign o[9250] = i[7074];
  assign o[9249] = i[7073];
  assign o[9248] = i[7072];
  assign o[9247] = i[7071];
  assign o[9246] = i[7070];
  assign o[9245] = i[7069];
  assign o[9244] = i[7068];
  assign o[9243] = i[7067];
  assign o[9242] = i[7066];
  assign o[9241] = i[7065];
  assign o[9240] = i[7064];
  assign o[9239] = i[7063];
  assign o[9238] = i[7062];
  assign o[9237] = i[7061];
  assign o[9236] = i[7060];
  assign o[9235] = i[7059];
  assign o[9234] = i[7058];
  assign o[9233] = i[7057];
  assign o[9232] = i[7056];
  assign o[9231] = i[7055];
  assign o[9230] = i[7054];
  assign o[9229] = i[7053];
  assign o[9228] = i[7052];
  assign o[9227] = i[7051];
  assign o[9226] = i[7050];
  assign o[9225] = i[7049];
  assign o[9224] = i[7048];
  assign o[9223] = i[7047];
  assign o[9222] = i[7046];
  assign o[9221] = i[7045];
  assign o[9220] = i[7044];
  assign o[9219] = i[7043];
  assign o[9218] = i[7042];
  assign o[9217] = i[7041];
  assign o[9216] = i[7040];
  assign o[9215] = i[7295];
  assign o[9214] = i[7294];
  assign o[9213] = i[7293];
  assign o[9212] = i[7292];
  assign o[9211] = i[7291];
  assign o[9210] = i[7290];
  assign o[9209] = i[7289];
  assign o[9208] = i[7288];
  assign o[9207] = i[7287];
  assign o[9206] = i[7286];
  assign o[9205] = i[7285];
  assign o[9204] = i[7284];
  assign o[9203] = i[7283];
  assign o[9202] = i[7282];
  assign o[9201] = i[7281];
  assign o[9200] = i[7280];
  assign o[9199] = i[7279];
  assign o[9198] = i[7278];
  assign o[9197] = i[7277];
  assign o[9196] = i[7276];
  assign o[9195] = i[7275];
  assign o[9194] = i[7274];
  assign o[9193] = i[7273];
  assign o[9192] = i[7272];
  assign o[9191] = i[7271];
  assign o[9190] = i[7270];
  assign o[9189] = i[7269];
  assign o[9188] = i[7268];
  assign o[9187] = i[7267];
  assign o[9186] = i[7266];
  assign o[9185] = i[7265];
  assign o[9184] = i[7264];
  assign o[9183] = i[7263];
  assign o[9182] = i[7262];
  assign o[9181] = i[7261];
  assign o[9180] = i[7260];
  assign o[9179] = i[7259];
  assign o[9178] = i[7258];
  assign o[9177] = i[7257];
  assign o[9176] = i[7256];
  assign o[9175] = i[7255];
  assign o[9174] = i[7254];
  assign o[9173] = i[7253];
  assign o[9172] = i[7252];
  assign o[9171] = i[7251];
  assign o[9170] = i[7250];
  assign o[9169] = i[7249];
  assign o[9168] = i[7248];
  assign o[9167] = i[7247];
  assign o[9166] = i[7246];
  assign o[9165] = i[7245];
  assign o[9164] = i[7244];
  assign o[9163] = i[7243];
  assign o[9162] = i[7242];
  assign o[9161] = i[7241];
  assign o[9160] = i[7240];
  assign o[9159] = i[7239];
  assign o[9158] = i[7238];
  assign o[9157] = i[7237];
  assign o[9156] = i[7236];
  assign o[9155] = i[7235];
  assign o[9154] = i[7234];
  assign o[9153] = i[7233];
  assign o[9152] = i[7232];
  assign o[9151] = i[7231];
  assign o[9150] = i[7230];
  assign o[9149] = i[7229];
  assign o[9148] = i[7228];
  assign o[9147] = i[7227];
  assign o[9146] = i[7226];
  assign o[9145] = i[7225];
  assign o[9144] = i[7224];
  assign o[9143] = i[7223];
  assign o[9142] = i[7222];
  assign o[9141] = i[7221];
  assign o[9140] = i[7220];
  assign o[9139] = i[7219];
  assign o[9138] = i[7218];
  assign o[9137] = i[7217];
  assign o[9136] = i[7216];
  assign o[9135] = i[7215];
  assign o[9134] = i[7214];
  assign o[9133] = i[7213];
  assign o[9132] = i[7212];
  assign o[9131] = i[7211];
  assign o[9130] = i[7210];
  assign o[9129] = i[7209];
  assign o[9128] = i[7208];
  assign o[9127] = i[7207];
  assign o[9126] = i[7206];
  assign o[9125] = i[7205];
  assign o[9124] = i[7204];
  assign o[9123] = i[7203];
  assign o[9122] = i[7202];
  assign o[9121] = i[7201];
  assign o[9120] = i[7200];
  assign o[9119] = i[7199];
  assign o[9118] = i[7198];
  assign o[9117] = i[7197];
  assign o[9116] = i[7196];
  assign o[9115] = i[7195];
  assign o[9114] = i[7194];
  assign o[9113] = i[7193];
  assign o[9112] = i[7192];
  assign o[9111] = i[7191];
  assign o[9110] = i[7190];
  assign o[9109] = i[7189];
  assign o[9108] = i[7188];
  assign o[9107] = i[7187];
  assign o[9106] = i[7186];
  assign o[9105] = i[7185];
  assign o[9104] = i[7184];
  assign o[9103] = i[7183];
  assign o[9102] = i[7182];
  assign o[9101] = i[7181];
  assign o[9100] = i[7180];
  assign o[9099] = i[7179];
  assign o[9098] = i[7178];
  assign o[9097] = i[7177];
  assign o[9096] = i[7176];
  assign o[9095] = i[7175];
  assign o[9094] = i[7174];
  assign o[9093] = i[7173];
  assign o[9092] = i[7172];
  assign o[9091] = i[7171];
  assign o[9090] = i[7170];
  assign o[9089] = i[7169];
  assign o[9088] = i[7168];
  assign o[9087] = i[7423];
  assign o[9086] = i[7422];
  assign o[9085] = i[7421];
  assign o[9084] = i[7420];
  assign o[9083] = i[7419];
  assign o[9082] = i[7418];
  assign o[9081] = i[7417];
  assign o[9080] = i[7416];
  assign o[9079] = i[7415];
  assign o[9078] = i[7414];
  assign o[9077] = i[7413];
  assign o[9076] = i[7412];
  assign o[9075] = i[7411];
  assign o[9074] = i[7410];
  assign o[9073] = i[7409];
  assign o[9072] = i[7408];
  assign o[9071] = i[7407];
  assign o[9070] = i[7406];
  assign o[9069] = i[7405];
  assign o[9068] = i[7404];
  assign o[9067] = i[7403];
  assign o[9066] = i[7402];
  assign o[9065] = i[7401];
  assign o[9064] = i[7400];
  assign o[9063] = i[7399];
  assign o[9062] = i[7398];
  assign o[9061] = i[7397];
  assign o[9060] = i[7396];
  assign o[9059] = i[7395];
  assign o[9058] = i[7394];
  assign o[9057] = i[7393];
  assign o[9056] = i[7392];
  assign o[9055] = i[7391];
  assign o[9054] = i[7390];
  assign o[9053] = i[7389];
  assign o[9052] = i[7388];
  assign o[9051] = i[7387];
  assign o[9050] = i[7386];
  assign o[9049] = i[7385];
  assign o[9048] = i[7384];
  assign o[9047] = i[7383];
  assign o[9046] = i[7382];
  assign o[9045] = i[7381];
  assign o[9044] = i[7380];
  assign o[9043] = i[7379];
  assign o[9042] = i[7378];
  assign o[9041] = i[7377];
  assign o[9040] = i[7376];
  assign o[9039] = i[7375];
  assign o[9038] = i[7374];
  assign o[9037] = i[7373];
  assign o[9036] = i[7372];
  assign o[9035] = i[7371];
  assign o[9034] = i[7370];
  assign o[9033] = i[7369];
  assign o[9032] = i[7368];
  assign o[9031] = i[7367];
  assign o[9030] = i[7366];
  assign o[9029] = i[7365];
  assign o[9028] = i[7364];
  assign o[9027] = i[7363];
  assign o[9026] = i[7362];
  assign o[9025] = i[7361];
  assign o[9024] = i[7360];
  assign o[9023] = i[7359];
  assign o[9022] = i[7358];
  assign o[9021] = i[7357];
  assign o[9020] = i[7356];
  assign o[9019] = i[7355];
  assign o[9018] = i[7354];
  assign o[9017] = i[7353];
  assign o[9016] = i[7352];
  assign o[9015] = i[7351];
  assign o[9014] = i[7350];
  assign o[9013] = i[7349];
  assign o[9012] = i[7348];
  assign o[9011] = i[7347];
  assign o[9010] = i[7346];
  assign o[9009] = i[7345];
  assign o[9008] = i[7344];
  assign o[9007] = i[7343];
  assign o[9006] = i[7342];
  assign o[9005] = i[7341];
  assign o[9004] = i[7340];
  assign o[9003] = i[7339];
  assign o[9002] = i[7338];
  assign o[9001] = i[7337];
  assign o[9000] = i[7336];
  assign o[8999] = i[7335];
  assign o[8998] = i[7334];
  assign o[8997] = i[7333];
  assign o[8996] = i[7332];
  assign o[8995] = i[7331];
  assign o[8994] = i[7330];
  assign o[8993] = i[7329];
  assign o[8992] = i[7328];
  assign o[8991] = i[7327];
  assign o[8990] = i[7326];
  assign o[8989] = i[7325];
  assign o[8988] = i[7324];
  assign o[8987] = i[7323];
  assign o[8986] = i[7322];
  assign o[8985] = i[7321];
  assign o[8984] = i[7320];
  assign o[8983] = i[7319];
  assign o[8982] = i[7318];
  assign o[8981] = i[7317];
  assign o[8980] = i[7316];
  assign o[8979] = i[7315];
  assign o[8978] = i[7314];
  assign o[8977] = i[7313];
  assign o[8976] = i[7312];
  assign o[8975] = i[7311];
  assign o[8974] = i[7310];
  assign o[8973] = i[7309];
  assign o[8972] = i[7308];
  assign o[8971] = i[7307];
  assign o[8970] = i[7306];
  assign o[8969] = i[7305];
  assign o[8968] = i[7304];
  assign o[8967] = i[7303];
  assign o[8966] = i[7302];
  assign o[8965] = i[7301];
  assign o[8964] = i[7300];
  assign o[8963] = i[7299];
  assign o[8962] = i[7298];
  assign o[8961] = i[7297];
  assign o[8960] = i[7296];
  assign o[8959] = i[7551];
  assign o[8958] = i[7550];
  assign o[8957] = i[7549];
  assign o[8956] = i[7548];
  assign o[8955] = i[7547];
  assign o[8954] = i[7546];
  assign o[8953] = i[7545];
  assign o[8952] = i[7544];
  assign o[8951] = i[7543];
  assign o[8950] = i[7542];
  assign o[8949] = i[7541];
  assign o[8948] = i[7540];
  assign o[8947] = i[7539];
  assign o[8946] = i[7538];
  assign o[8945] = i[7537];
  assign o[8944] = i[7536];
  assign o[8943] = i[7535];
  assign o[8942] = i[7534];
  assign o[8941] = i[7533];
  assign o[8940] = i[7532];
  assign o[8939] = i[7531];
  assign o[8938] = i[7530];
  assign o[8937] = i[7529];
  assign o[8936] = i[7528];
  assign o[8935] = i[7527];
  assign o[8934] = i[7526];
  assign o[8933] = i[7525];
  assign o[8932] = i[7524];
  assign o[8931] = i[7523];
  assign o[8930] = i[7522];
  assign o[8929] = i[7521];
  assign o[8928] = i[7520];
  assign o[8927] = i[7519];
  assign o[8926] = i[7518];
  assign o[8925] = i[7517];
  assign o[8924] = i[7516];
  assign o[8923] = i[7515];
  assign o[8922] = i[7514];
  assign o[8921] = i[7513];
  assign o[8920] = i[7512];
  assign o[8919] = i[7511];
  assign o[8918] = i[7510];
  assign o[8917] = i[7509];
  assign o[8916] = i[7508];
  assign o[8915] = i[7507];
  assign o[8914] = i[7506];
  assign o[8913] = i[7505];
  assign o[8912] = i[7504];
  assign o[8911] = i[7503];
  assign o[8910] = i[7502];
  assign o[8909] = i[7501];
  assign o[8908] = i[7500];
  assign o[8907] = i[7499];
  assign o[8906] = i[7498];
  assign o[8905] = i[7497];
  assign o[8904] = i[7496];
  assign o[8903] = i[7495];
  assign o[8902] = i[7494];
  assign o[8901] = i[7493];
  assign o[8900] = i[7492];
  assign o[8899] = i[7491];
  assign o[8898] = i[7490];
  assign o[8897] = i[7489];
  assign o[8896] = i[7488];
  assign o[8895] = i[7487];
  assign o[8894] = i[7486];
  assign o[8893] = i[7485];
  assign o[8892] = i[7484];
  assign o[8891] = i[7483];
  assign o[8890] = i[7482];
  assign o[8889] = i[7481];
  assign o[8888] = i[7480];
  assign o[8887] = i[7479];
  assign o[8886] = i[7478];
  assign o[8885] = i[7477];
  assign o[8884] = i[7476];
  assign o[8883] = i[7475];
  assign o[8882] = i[7474];
  assign o[8881] = i[7473];
  assign o[8880] = i[7472];
  assign o[8879] = i[7471];
  assign o[8878] = i[7470];
  assign o[8877] = i[7469];
  assign o[8876] = i[7468];
  assign o[8875] = i[7467];
  assign o[8874] = i[7466];
  assign o[8873] = i[7465];
  assign o[8872] = i[7464];
  assign o[8871] = i[7463];
  assign o[8870] = i[7462];
  assign o[8869] = i[7461];
  assign o[8868] = i[7460];
  assign o[8867] = i[7459];
  assign o[8866] = i[7458];
  assign o[8865] = i[7457];
  assign o[8864] = i[7456];
  assign o[8863] = i[7455];
  assign o[8862] = i[7454];
  assign o[8861] = i[7453];
  assign o[8860] = i[7452];
  assign o[8859] = i[7451];
  assign o[8858] = i[7450];
  assign o[8857] = i[7449];
  assign o[8856] = i[7448];
  assign o[8855] = i[7447];
  assign o[8854] = i[7446];
  assign o[8853] = i[7445];
  assign o[8852] = i[7444];
  assign o[8851] = i[7443];
  assign o[8850] = i[7442];
  assign o[8849] = i[7441];
  assign o[8848] = i[7440];
  assign o[8847] = i[7439];
  assign o[8846] = i[7438];
  assign o[8845] = i[7437];
  assign o[8844] = i[7436];
  assign o[8843] = i[7435];
  assign o[8842] = i[7434];
  assign o[8841] = i[7433];
  assign o[8840] = i[7432];
  assign o[8839] = i[7431];
  assign o[8838] = i[7430];
  assign o[8837] = i[7429];
  assign o[8836] = i[7428];
  assign o[8835] = i[7427];
  assign o[8834] = i[7426];
  assign o[8833] = i[7425];
  assign o[8832] = i[7424];
  assign o[8831] = i[7679];
  assign o[8830] = i[7678];
  assign o[8829] = i[7677];
  assign o[8828] = i[7676];
  assign o[8827] = i[7675];
  assign o[8826] = i[7674];
  assign o[8825] = i[7673];
  assign o[8824] = i[7672];
  assign o[8823] = i[7671];
  assign o[8822] = i[7670];
  assign o[8821] = i[7669];
  assign o[8820] = i[7668];
  assign o[8819] = i[7667];
  assign o[8818] = i[7666];
  assign o[8817] = i[7665];
  assign o[8816] = i[7664];
  assign o[8815] = i[7663];
  assign o[8814] = i[7662];
  assign o[8813] = i[7661];
  assign o[8812] = i[7660];
  assign o[8811] = i[7659];
  assign o[8810] = i[7658];
  assign o[8809] = i[7657];
  assign o[8808] = i[7656];
  assign o[8807] = i[7655];
  assign o[8806] = i[7654];
  assign o[8805] = i[7653];
  assign o[8804] = i[7652];
  assign o[8803] = i[7651];
  assign o[8802] = i[7650];
  assign o[8801] = i[7649];
  assign o[8800] = i[7648];
  assign o[8799] = i[7647];
  assign o[8798] = i[7646];
  assign o[8797] = i[7645];
  assign o[8796] = i[7644];
  assign o[8795] = i[7643];
  assign o[8794] = i[7642];
  assign o[8793] = i[7641];
  assign o[8792] = i[7640];
  assign o[8791] = i[7639];
  assign o[8790] = i[7638];
  assign o[8789] = i[7637];
  assign o[8788] = i[7636];
  assign o[8787] = i[7635];
  assign o[8786] = i[7634];
  assign o[8785] = i[7633];
  assign o[8784] = i[7632];
  assign o[8783] = i[7631];
  assign o[8782] = i[7630];
  assign o[8781] = i[7629];
  assign o[8780] = i[7628];
  assign o[8779] = i[7627];
  assign o[8778] = i[7626];
  assign o[8777] = i[7625];
  assign o[8776] = i[7624];
  assign o[8775] = i[7623];
  assign o[8774] = i[7622];
  assign o[8773] = i[7621];
  assign o[8772] = i[7620];
  assign o[8771] = i[7619];
  assign o[8770] = i[7618];
  assign o[8769] = i[7617];
  assign o[8768] = i[7616];
  assign o[8767] = i[7615];
  assign o[8766] = i[7614];
  assign o[8765] = i[7613];
  assign o[8764] = i[7612];
  assign o[8763] = i[7611];
  assign o[8762] = i[7610];
  assign o[8761] = i[7609];
  assign o[8760] = i[7608];
  assign o[8759] = i[7607];
  assign o[8758] = i[7606];
  assign o[8757] = i[7605];
  assign o[8756] = i[7604];
  assign o[8755] = i[7603];
  assign o[8754] = i[7602];
  assign o[8753] = i[7601];
  assign o[8752] = i[7600];
  assign o[8751] = i[7599];
  assign o[8750] = i[7598];
  assign o[8749] = i[7597];
  assign o[8748] = i[7596];
  assign o[8747] = i[7595];
  assign o[8746] = i[7594];
  assign o[8745] = i[7593];
  assign o[8744] = i[7592];
  assign o[8743] = i[7591];
  assign o[8742] = i[7590];
  assign o[8741] = i[7589];
  assign o[8740] = i[7588];
  assign o[8739] = i[7587];
  assign o[8738] = i[7586];
  assign o[8737] = i[7585];
  assign o[8736] = i[7584];
  assign o[8735] = i[7583];
  assign o[8734] = i[7582];
  assign o[8733] = i[7581];
  assign o[8732] = i[7580];
  assign o[8731] = i[7579];
  assign o[8730] = i[7578];
  assign o[8729] = i[7577];
  assign o[8728] = i[7576];
  assign o[8727] = i[7575];
  assign o[8726] = i[7574];
  assign o[8725] = i[7573];
  assign o[8724] = i[7572];
  assign o[8723] = i[7571];
  assign o[8722] = i[7570];
  assign o[8721] = i[7569];
  assign o[8720] = i[7568];
  assign o[8719] = i[7567];
  assign o[8718] = i[7566];
  assign o[8717] = i[7565];
  assign o[8716] = i[7564];
  assign o[8715] = i[7563];
  assign o[8714] = i[7562];
  assign o[8713] = i[7561];
  assign o[8712] = i[7560];
  assign o[8711] = i[7559];
  assign o[8710] = i[7558];
  assign o[8709] = i[7557];
  assign o[8708] = i[7556];
  assign o[8707] = i[7555];
  assign o[8706] = i[7554];
  assign o[8705] = i[7553];
  assign o[8704] = i[7552];
  assign o[8703] = i[7807];
  assign o[8702] = i[7806];
  assign o[8701] = i[7805];
  assign o[8700] = i[7804];
  assign o[8699] = i[7803];
  assign o[8698] = i[7802];
  assign o[8697] = i[7801];
  assign o[8696] = i[7800];
  assign o[8695] = i[7799];
  assign o[8694] = i[7798];
  assign o[8693] = i[7797];
  assign o[8692] = i[7796];
  assign o[8691] = i[7795];
  assign o[8690] = i[7794];
  assign o[8689] = i[7793];
  assign o[8688] = i[7792];
  assign o[8687] = i[7791];
  assign o[8686] = i[7790];
  assign o[8685] = i[7789];
  assign o[8684] = i[7788];
  assign o[8683] = i[7787];
  assign o[8682] = i[7786];
  assign o[8681] = i[7785];
  assign o[8680] = i[7784];
  assign o[8679] = i[7783];
  assign o[8678] = i[7782];
  assign o[8677] = i[7781];
  assign o[8676] = i[7780];
  assign o[8675] = i[7779];
  assign o[8674] = i[7778];
  assign o[8673] = i[7777];
  assign o[8672] = i[7776];
  assign o[8671] = i[7775];
  assign o[8670] = i[7774];
  assign o[8669] = i[7773];
  assign o[8668] = i[7772];
  assign o[8667] = i[7771];
  assign o[8666] = i[7770];
  assign o[8665] = i[7769];
  assign o[8664] = i[7768];
  assign o[8663] = i[7767];
  assign o[8662] = i[7766];
  assign o[8661] = i[7765];
  assign o[8660] = i[7764];
  assign o[8659] = i[7763];
  assign o[8658] = i[7762];
  assign o[8657] = i[7761];
  assign o[8656] = i[7760];
  assign o[8655] = i[7759];
  assign o[8654] = i[7758];
  assign o[8653] = i[7757];
  assign o[8652] = i[7756];
  assign o[8651] = i[7755];
  assign o[8650] = i[7754];
  assign o[8649] = i[7753];
  assign o[8648] = i[7752];
  assign o[8647] = i[7751];
  assign o[8646] = i[7750];
  assign o[8645] = i[7749];
  assign o[8644] = i[7748];
  assign o[8643] = i[7747];
  assign o[8642] = i[7746];
  assign o[8641] = i[7745];
  assign o[8640] = i[7744];
  assign o[8639] = i[7743];
  assign o[8638] = i[7742];
  assign o[8637] = i[7741];
  assign o[8636] = i[7740];
  assign o[8635] = i[7739];
  assign o[8634] = i[7738];
  assign o[8633] = i[7737];
  assign o[8632] = i[7736];
  assign o[8631] = i[7735];
  assign o[8630] = i[7734];
  assign o[8629] = i[7733];
  assign o[8628] = i[7732];
  assign o[8627] = i[7731];
  assign o[8626] = i[7730];
  assign o[8625] = i[7729];
  assign o[8624] = i[7728];
  assign o[8623] = i[7727];
  assign o[8622] = i[7726];
  assign o[8621] = i[7725];
  assign o[8620] = i[7724];
  assign o[8619] = i[7723];
  assign o[8618] = i[7722];
  assign o[8617] = i[7721];
  assign o[8616] = i[7720];
  assign o[8615] = i[7719];
  assign o[8614] = i[7718];
  assign o[8613] = i[7717];
  assign o[8612] = i[7716];
  assign o[8611] = i[7715];
  assign o[8610] = i[7714];
  assign o[8609] = i[7713];
  assign o[8608] = i[7712];
  assign o[8607] = i[7711];
  assign o[8606] = i[7710];
  assign o[8605] = i[7709];
  assign o[8604] = i[7708];
  assign o[8603] = i[7707];
  assign o[8602] = i[7706];
  assign o[8601] = i[7705];
  assign o[8600] = i[7704];
  assign o[8599] = i[7703];
  assign o[8598] = i[7702];
  assign o[8597] = i[7701];
  assign o[8596] = i[7700];
  assign o[8595] = i[7699];
  assign o[8594] = i[7698];
  assign o[8593] = i[7697];
  assign o[8592] = i[7696];
  assign o[8591] = i[7695];
  assign o[8590] = i[7694];
  assign o[8589] = i[7693];
  assign o[8588] = i[7692];
  assign o[8587] = i[7691];
  assign o[8586] = i[7690];
  assign o[8585] = i[7689];
  assign o[8584] = i[7688];
  assign o[8583] = i[7687];
  assign o[8582] = i[7686];
  assign o[8581] = i[7685];
  assign o[8580] = i[7684];
  assign o[8579] = i[7683];
  assign o[8578] = i[7682];
  assign o[8577] = i[7681];
  assign o[8576] = i[7680];
  assign o[8575] = i[7935];
  assign o[8574] = i[7934];
  assign o[8573] = i[7933];
  assign o[8572] = i[7932];
  assign o[8571] = i[7931];
  assign o[8570] = i[7930];
  assign o[8569] = i[7929];
  assign o[8568] = i[7928];
  assign o[8567] = i[7927];
  assign o[8566] = i[7926];
  assign o[8565] = i[7925];
  assign o[8564] = i[7924];
  assign o[8563] = i[7923];
  assign o[8562] = i[7922];
  assign o[8561] = i[7921];
  assign o[8560] = i[7920];
  assign o[8559] = i[7919];
  assign o[8558] = i[7918];
  assign o[8557] = i[7917];
  assign o[8556] = i[7916];
  assign o[8555] = i[7915];
  assign o[8554] = i[7914];
  assign o[8553] = i[7913];
  assign o[8552] = i[7912];
  assign o[8551] = i[7911];
  assign o[8550] = i[7910];
  assign o[8549] = i[7909];
  assign o[8548] = i[7908];
  assign o[8547] = i[7907];
  assign o[8546] = i[7906];
  assign o[8545] = i[7905];
  assign o[8544] = i[7904];
  assign o[8543] = i[7903];
  assign o[8542] = i[7902];
  assign o[8541] = i[7901];
  assign o[8540] = i[7900];
  assign o[8539] = i[7899];
  assign o[8538] = i[7898];
  assign o[8537] = i[7897];
  assign o[8536] = i[7896];
  assign o[8535] = i[7895];
  assign o[8534] = i[7894];
  assign o[8533] = i[7893];
  assign o[8532] = i[7892];
  assign o[8531] = i[7891];
  assign o[8530] = i[7890];
  assign o[8529] = i[7889];
  assign o[8528] = i[7888];
  assign o[8527] = i[7887];
  assign o[8526] = i[7886];
  assign o[8525] = i[7885];
  assign o[8524] = i[7884];
  assign o[8523] = i[7883];
  assign o[8522] = i[7882];
  assign o[8521] = i[7881];
  assign o[8520] = i[7880];
  assign o[8519] = i[7879];
  assign o[8518] = i[7878];
  assign o[8517] = i[7877];
  assign o[8516] = i[7876];
  assign o[8515] = i[7875];
  assign o[8514] = i[7874];
  assign o[8513] = i[7873];
  assign o[8512] = i[7872];
  assign o[8511] = i[7871];
  assign o[8510] = i[7870];
  assign o[8509] = i[7869];
  assign o[8508] = i[7868];
  assign o[8507] = i[7867];
  assign o[8506] = i[7866];
  assign o[8505] = i[7865];
  assign o[8504] = i[7864];
  assign o[8503] = i[7863];
  assign o[8502] = i[7862];
  assign o[8501] = i[7861];
  assign o[8500] = i[7860];
  assign o[8499] = i[7859];
  assign o[8498] = i[7858];
  assign o[8497] = i[7857];
  assign o[8496] = i[7856];
  assign o[8495] = i[7855];
  assign o[8494] = i[7854];
  assign o[8493] = i[7853];
  assign o[8492] = i[7852];
  assign o[8491] = i[7851];
  assign o[8490] = i[7850];
  assign o[8489] = i[7849];
  assign o[8488] = i[7848];
  assign o[8487] = i[7847];
  assign o[8486] = i[7846];
  assign o[8485] = i[7845];
  assign o[8484] = i[7844];
  assign o[8483] = i[7843];
  assign o[8482] = i[7842];
  assign o[8481] = i[7841];
  assign o[8480] = i[7840];
  assign o[8479] = i[7839];
  assign o[8478] = i[7838];
  assign o[8477] = i[7837];
  assign o[8476] = i[7836];
  assign o[8475] = i[7835];
  assign o[8474] = i[7834];
  assign o[8473] = i[7833];
  assign o[8472] = i[7832];
  assign o[8471] = i[7831];
  assign o[8470] = i[7830];
  assign o[8469] = i[7829];
  assign o[8468] = i[7828];
  assign o[8467] = i[7827];
  assign o[8466] = i[7826];
  assign o[8465] = i[7825];
  assign o[8464] = i[7824];
  assign o[8463] = i[7823];
  assign o[8462] = i[7822];
  assign o[8461] = i[7821];
  assign o[8460] = i[7820];
  assign o[8459] = i[7819];
  assign o[8458] = i[7818];
  assign o[8457] = i[7817];
  assign o[8456] = i[7816];
  assign o[8455] = i[7815];
  assign o[8454] = i[7814];
  assign o[8453] = i[7813];
  assign o[8452] = i[7812];
  assign o[8451] = i[7811];
  assign o[8450] = i[7810];
  assign o[8449] = i[7809];
  assign o[8448] = i[7808];
  assign o[8447] = i[8063];
  assign o[8446] = i[8062];
  assign o[8445] = i[8061];
  assign o[8444] = i[8060];
  assign o[8443] = i[8059];
  assign o[8442] = i[8058];
  assign o[8441] = i[8057];
  assign o[8440] = i[8056];
  assign o[8439] = i[8055];
  assign o[8438] = i[8054];
  assign o[8437] = i[8053];
  assign o[8436] = i[8052];
  assign o[8435] = i[8051];
  assign o[8434] = i[8050];
  assign o[8433] = i[8049];
  assign o[8432] = i[8048];
  assign o[8431] = i[8047];
  assign o[8430] = i[8046];
  assign o[8429] = i[8045];
  assign o[8428] = i[8044];
  assign o[8427] = i[8043];
  assign o[8426] = i[8042];
  assign o[8425] = i[8041];
  assign o[8424] = i[8040];
  assign o[8423] = i[8039];
  assign o[8422] = i[8038];
  assign o[8421] = i[8037];
  assign o[8420] = i[8036];
  assign o[8419] = i[8035];
  assign o[8418] = i[8034];
  assign o[8417] = i[8033];
  assign o[8416] = i[8032];
  assign o[8415] = i[8031];
  assign o[8414] = i[8030];
  assign o[8413] = i[8029];
  assign o[8412] = i[8028];
  assign o[8411] = i[8027];
  assign o[8410] = i[8026];
  assign o[8409] = i[8025];
  assign o[8408] = i[8024];
  assign o[8407] = i[8023];
  assign o[8406] = i[8022];
  assign o[8405] = i[8021];
  assign o[8404] = i[8020];
  assign o[8403] = i[8019];
  assign o[8402] = i[8018];
  assign o[8401] = i[8017];
  assign o[8400] = i[8016];
  assign o[8399] = i[8015];
  assign o[8398] = i[8014];
  assign o[8397] = i[8013];
  assign o[8396] = i[8012];
  assign o[8395] = i[8011];
  assign o[8394] = i[8010];
  assign o[8393] = i[8009];
  assign o[8392] = i[8008];
  assign o[8391] = i[8007];
  assign o[8390] = i[8006];
  assign o[8389] = i[8005];
  assign o[8388] = i[8004];
  assign o[8387] = i[8003];
  assign o[8386] = i[8002];
  assign o[8385] = i[8001];
  assign o[8384] = i[8000];
  assign o[8383] = i[7999];
  assign o[8382] = i[7998];
  assign o[8381] = i[7997];
  assign o[8380] = i[7996];
  assign o[8379] = i[7995];
  assign o[8378] = i[7994];
  assign o[8377] = i[7993];
  assign o[8376] = i[7992];
  assign o[8375] = i[7991];
  assign o[8374] = i[7990];
  assign o[8373] = i[7989];
  assign o[8372] = i[7988];
  assign o[8371] = i[7987];
  assign o[8370] = i[7986];
  assign o[8369] = i[7985];
  assign o[8368] = i[7984];
  assign o[8367] = i[7983];
  assign o[8366] = i[7982];
  assign o[8365] = i[7981];
  assign o[8364] = i[7980];
  assign o[8363] = i[7979];
  assign o[8362] = i[7978];
  assign o[8361] = i[7977];
  assign o[8360] = i[7976];
  assign o[8359] = i[7975];
  assign o[8358] = i[7974];
  assign o[8357] = i[7973];
  assign o[8356] = i[7972];
  assign o[8355] = i[7971];
  assign o[8354] = i[7970];
  assign o[8353] = i[7969];
  assign o[8352] = i[7968];
  assign o[8351] = i[7967];
  assign o[8350] = i[7966];
  assign o[8349] = i[7965];
  assign o[8348] = i[7964];
  assign o[8347] = i[7963];
  assign o[8346] = i[7962];
  assign o[8345] = i[7961];
  assign o[8344] = i[7960];
  assign o[8343] = i[7959];
  assign o[8342] = i[7958];
  assign o[8341] = i[7957];
  assign o[8340] = i[7956];
  assign o[8339] = i[7955];
  assign o[8338] = i[7954];
  assign o[8337] = i[7953];
  assign o[8336] = i[7952];
  assign o[8335] = i[7951];
  assign o[8334] = i[7950];
  assign o[8333] = i[7949];
  assign o[8332] = i[7948];
  assign o[8331] = i[7947];
  assign o[8330] = i[7946];
  assign o[8329] = i[7945];
  assign o[8328] = i[7944];
  assign o[8327] = i[7943];
  assign o[8326] = i[7942];
  assign o[8325] = i[7941];
  assign o[8324] = i[7940];
  assign o[8323] = i[7939];
  assign o[8322] = i[7938];
  assign o[8321] = i[7937];
  assign o[8320] = i[7936];
  assign o[8319] = i[8191];
  assign o[8318] = i[8190];
  assign o[8317] = i[8189];
  assign o[8316] = i[8188];
  assign o[8315] = i[8187];
  assign o[8314] = i[8186];
  assign o[8313] = i[8185];
  assign o[8312] = i[8184];
  assign o[8311] = i[8183];
  assign o[8310] = i[8182];
  assign o[8309] = i[8181];
  assign o[8308] = i[8180];
  assign o[8307] = i[8179];
  assign o[8306] = i[8178];
  assign o[8305] = i[8177];
  assign o[8304] = i[8176];
  assign o[8303] = i[8175];
  assign o[8302] = i[8174];
  assign o[8301] = i[8173];
  assign o[8300] = i[8172];
  assign o[8299] = i[8171];
  assign o[8298] = i[8170];
  assign o[8297] = i[8169];
  assign o[8296] = i[8168];
  assign o[8295] = i[8167];
  assign o[8294] = i[8166];
  assign o[8293] = i[8165];
  assign o[8292] = i[8164];
  assign o[8291] = i[8163];
  assign o[8290] = i[8162];
  assign o[8289] = i[8161];
  assign o[8288] = i[8160];
  assign o[8287] = i[8159];
  assign o[8286] = i[8158];
  assign o[8285] = i[8157];
  assign o[8284] = i[8156];
  assign o[8283] = i[8155];
  assign o[8282] = i[8154];
  assign o[8281] = i[8153];
  assign o[8280] = i[8152];
  assign o[8279] = i[8151];
  assign o[8278] = i[8150];
  assign o[8277] = i[8149];
  assign o[8276] = i[8148];
  assign o[8275] = i[8147];
  assign o[8274] = i[8146];
  assign o[8273] = i[8145];
  assign o[8272] = i[8144];
  assign o[8271] = i[8143];
  assign o[8270] = i[8142];
  assign o[8269] = i[8141];
  assign o[8268] = i[8140];
  assign o[8267] = i[8139];
  assign o[8266] = i[8138];
  assign o[8265] = i[8137];
  assign o[8264] = i[8136];
  assign o[8263] = i[8135];
  assign o[8262] = i[8134];
  assign o[8261] = i[8133];
  assign o[8260] = i[8132];
  assign o[8259] = i[8131];
  assign o[8258] = i[8130];
  assign o[8257] = i[8129];
  assign o[8256] = i[8128];
  assign o[8255] = i[8127];
  assign o[8254] = i[8126];
  assign o[8253] = i[8125];
  assign o[8252] = i[8124];
  assign o[8251] = i[8123];
  assign o[8250] = i[8122];
  assign o[8249] = i[8121];
  assign o[8248] = i[8120];
  assign o[8247] = i[8119];
  assign o[8246] = i[8118];
  assign o[8245] = i[8117];
  assign o[8244] = i[8116];
  assign o[8243] = i[8115];
  assign o[8242] = i[8114];
  assign o[8241] = i[8113];
  assign o[8240] = i[8112];
  assign o[8239] = i[8111];
  assign o[8238] = i[8110];
  assign o[8237] = i[8109];
  assign o[8236] = i[8108];
  assign o[8235] = i[8107];
  assign o[8234] = i[8106];
  assign o[8233] = i[8105];
  assign o[8232] = i[8104];
  assign o[8231] = i[8103];
  assign o[8230] = i[8102];
  assign o[8229] = i[8101];
  assign o[8228] = i[8100];
  assign o[8227] = i[8099];
  assign o[8226] = i[8098];
  assign o[8225] = i[8097];
  assign o[8224] = i[8096];
  assign o[8223] = i[8095];
  assign o[8222] = i[8094];
  assign o[8221] = i[8093];
  assign o[8220] = i[8092];
  assign o[8219] = i[8091];
  assign o[8218] = i[8090];
  assign o[8217] = i[8089];
  assign o[8216] = i[8088];
  assign o[8215] = i[8087];
  assign o[8214] = i[8086];
  assign o[8213] = i[8085];
  assign o[8212] = i[8084];
  assign o[8211] = i[8083];
  assign o[8210] = i[8082];
  assign o[8209] = i[8081];
  assign o[8208] = i[8080];
  assign o[8207] = i[8079];
  assign o[8206] = i[8078];
  assign o[8205] = i[8077];
  assign o[8204] = i[8076];
  assign o[8203] = i[8075];
  assign o[8202] = i[8074];
  assign o[8201] = i[8073];
  assign o[8200] = i[8072];
  assign o[8199] = i[8071];
  assign o[8198] = i[8070];
  assign o[8197] = i[8069];
  assign o[8196] = i[8068];
  assign o[8195] = i[8067];
  assign o[8194] = i[8066];
  assign o[8193] = i[8065];
  assign o[8192] = i[8064];
  assign o[8191] = i[8319];
  assign o[8190] = i[8318];
  assign o[8189] = i[8317];
  assign o[8188] = i[8316];
  assign o[8187] = i[8315];
  assign o[8186] = i[8314];
  assign o[8185] = i[8313];
  assign o[8184] = i[8312];
  assign o[8183] = i[8311];
  assign o[8182] = i[8310];
  assign o[8181] = i[8309];
  assign o[8180] = i[8308];
  assign o[8179] = i[8307];
  assign o[8178] = i[8306];
  assign o[8177] = i[8305];
  assign o[8176] = i[8304];
  assign o[8175] = i[8303];
  assign o[8174] = i[8302];
  assign o[8173] = i[8301];
  assign o[8172] = i[8300];
  assign o[8171] = i[8299];
  assign o[8170] = i[8298];
  assign o[8169] = i[8297];
  assign o[8168] = i[8296];
  assign o[8167] = i[8295];
  assign o[8166] = i[8294];
  assign o[8165] = i[8293];
  assign o[8164] = i[8292];
  assign o[8163] = i[8291];
  assign o[8162] = i[8290];
  assign o[8161] = i[8289];
  assign o[8160] = i[8288];
  assign o[8159] = i[8287];
  assign o[8158] = i[8286];
  assign o[8157] = i[8285];
  assign o[8156] = i[8284];
  assign o[8155] = i[8283];
  assign o[8154] = i[8282];
  assign o[8153] = i[8281];
  assign o[8152] = i[8280];
  assign o[8151] = i[8279];
  assign o[8150] = i[8278];
  assign o[8149] = i[8277];
  assign o[8148] = i[8276];
  assign o[8147] = i[8275];
  assign o[8146] = i[8274];
  assign o[8145] = i[8273];
  assign o[8144] = i[8272];
  assign o[8143] = i[8271];
  assign o[8142] = i[8270];
  assign o[8141] = i[8269];
  assign o[8140] = i[8268];
  assign o[8139] = i[8267];
  assign o[8138] = i[8266];
  assign o[8137] = i[8265];
  assign o[8136] = i[8264];
  assign o[8135] = i[8263];
  assign o[8134] = i[8262];
  assign o[8133] = i[8261];
  assign o[8132] = i[8260];
  assign o[8131] = i[8259];
  assign o[8130] = i[8258];
  assign o[8129] = i[8257];
  assign o[8128] = i[8256];
  assign o[8127] = i[8255];
  assign o[8126] = i[8254];
  assign o[8125] = i[8253];
  assign o[8124] = i[8252];
  assign o[8123] = i[8251];
  assign o[8122] = i[8250];
  assign o[8121] = i[8249];
  assign o[8120] = i[8248];
  assign o[8119] = i[8247];
  assign o[8118] = i[8246];
  assign o[8117] = i[8245];
  assign o[8116] = i[8244];
  assign o[8115] = i[8243];
  assign o[8114] = i[8242];
  assign o[8113] = i[8241];
  assign o[8112] = i[8240];
  assign o[8111] = i[8239];
  assign o[8110] = i[8238];
  assign o[8109] = i[8237];
  assign o[8108] = i[8236];
  assign o[8107] = i[8235];
  assign o[8106] = i[8234];
  assign o[8105] = i[8233];
  assign o[8104] = i[8232];
  assign o[8103] = i[8231];
  assign o[8102] = i[8230];
  assign o[8101] = i[8229];
  assign o[8100] = i[8228];
  assign o[8099] = i[8227];
  assign o[8098] = i[8226];
  assign o[8097] = i[8225];
  assign o[8096] = i[8224];
  assign o[8095] = i[8223];
  assign o[8094] = i[8222];
  assign o[8093] = i[8221];
  assign o[8092] = i[8220];
  assign o[8091] = i[8219];
  assign o[8090] = i[8218];
  assign o[8089] = i[8217];
  assign o[8088] = i[8216];
  assign o[8087] = i[8215];
  assign o[8086] = i[8214];
  assign o[8085] = i[8213];
  assign o[8084] = i[8212];
  assign o[8083] = i[8211];
  assign o[8082] = i[8210];
  assign o[8081] = i[8209];
  assign o[8080] = i[8208];
  assign o[8079] = i[8207];
  assign o[8078] = i[8206];
  assign o[8077] = i[8205];
  assign o[8076] = i[8204];
  assign o[8075] = i[8203];
  assign o[8074] = i[8202];
  assign o[8073] = i[8201];
  assign o[8072] = i[8200];
  assign o[8071] = i[8199];
  assign o[8070] = i[8198];
  assign o[8069] = i[8197];
  assign o[8068] = i[8196];
  assign o[8067] = i[8195];
  assign o[8066] = i[8194];
  assign o[8065] = i[8193];
  assign o[8064] = i[8192];
  assign o[8063] = i[8447];
  assign o[8062] = i[8446];
  assign o[8061] = i[8445];
  assign o[8060] = i[8444];
  assign o[8059] = i[8443];
  assign o[8058] = i[8442];
  assign o[8057] = i[8441];
  assign o[8056] = i[8440];
  assign o[8055] = i[8439];
  assign o[8054] = i[8438];
  assign o[8053] = i[8437];
  assign o[8052] = i[8436];
  assign o[8051] = i[8435];
  assign o[8050] = i[8434];
  assign o[8049] = i[8433];
  assign o[8048] = i[8432];
  assign o[8047] = i[8431];
  assign o[8046] = i[8430];
  assign o[8045] = i[8429];
  assign o[8044] = i[8428];
  assign o[8043] = i[8427];
  assign o[8042] = i[8426];
  assign o[8041] = i[8425];
  assign o[8040] = i[8424];
  assign o[8039] = i[8423];
  assign o[8038] = i[8422];
  assign o[8037] = i[8421];
  assign o[8036] = i[8420];
  assign o[8035] = i[8419];
  assign o[8034] = i[8418];
  assign o[8033] = i[8417];
  assign o[8032] = i[8416];
  assign o[8031] = i[8415];
  assign o[8030] = i[8414];
  assign o[8029] = i[8413];
  assign o[8028] = i[8412];
  assign o[8027] = i[8411];
  assign o[8026] = i[8410];
  assign o[8025] = i[8409];
  assign o[8024] = i[8408];
  assign o[8023] = i[8407];
  assign o[8022] = i[8406];
  assign o[8021] = i[8405];
  assign o[8020] = i[8404];
  assign o[8019] = i[8403];
  assign o[8018] = i[8402];
  assign o[8017] = i[8401];
  assign o[8016] = i[8400];
  assign o[8015] = i[8399];
  assign o[8014] = i[8398];
  assign o[8013] = i[8397];
  assign o[8012] = i[8396];
  assign o[8011] = i[8395];
  assign o[8010] = i[8394];
  assign o[8009] = i[8393];
  assign o[8008] = i[8392];
  assign o[8007] = i[8391];
  assign o[8006] = i[8390];
  assign o[8005] = i[8389];
  assign o[8004] = i[8388];
  assign o[8003] = i[8387];
  assign o[8002] = i[8386];
  assign o[8001] = i[8385];
  assign o[8000] = i[8384];
  assign o[7999] = i[8383];
  assign o[7998] = i[8382];
  assign o[7997] = i[8381];
  assign o[7996] = i[8380];
  assign o[7995] = i[8379];
  assign o[7994] = i[8378];
  assign o[7993] = i[8377];
  assign o[7992] = i[8376];
  assign o[7991] = i[8375];
  assign o[7990] = i[8374];
  assign o[7989] = i[8373];
  assign o[7988] = i[8372];
  assign o[7987] = i[8371];
  assign o[7986] = i[8370];
  assign o[7985] = i[8369];
  assign o[7984] = i[8368];
  assign o[7983] = i[8367];
  assign o[7982] = i[8366];
  assign o[7981] = i[8365];
  assign o[7980] = i[8364];
  assign o[7979] = i[8363];
  assign o[7978] = i[8362];
  assign o[7977] = i[8361];
  assign o[7976] = i[8360];
  assign o[7975] = i[8359];
  assign o[7974] = i[8358];
  assign o[7973] = i[8357];
  assign o[7972] = i[8356];
  assign o[7971] = i[8355];
  assign o[7970] = i[8354];
  assign o[7969] = i[8353];
  assign o[7968] = i[8352];
  assign o[7967] = i[8351];
  assign o[7966] = i[8350];
  assign o[7965] = i[8349];
  assign o[7964] = i[8348];
  assign o[7963] = i[8347];
  assign o[7962] = i[8346];
  assign o[7961] = i[8345];
  assign o[7960] = i[8344];
  assign o[7959] = i[8343];
  assign o[7958] = i[8342];
  assign o[7957] = i[8341];
  assign o[7956] = i[8340];
  assign o[7955] = i[8339];
  assign o[7954] = i[8338];
  assign o[7953] = i[8337];
  assign o[7952] = i[8336];
  assign o[7951] = i[8335];
  assign o[7950] = i[8334];
  assign o[7949] = i[8333];
  assign o[7948] = i[8332];
  assign o[7947] = i[8331];
  assign o[7946] = i[8330];
  assign o[7945] = i[8329];
  assign o[7944] = i[8328];
  assign o[7943] = i[8327];
  assign o[7942] = i[8326];
  assign o[7941] = i[8325];
  assign o[7940] = i[8324];
  assign o[7939] = i[8323];
  assign o[7938] = i[8322];
  assign o[7937] = i[8321];
  assign o[7936] = i[8320];
  assign o[7935] = i[8575];
  assign o[7934] = i[8574];
  assign o[7933] = i[8573];
  assign o[7932] = i[8572];
  assign o[7931] = i[8571];
  assign o[7930] = i[8570];
  assign o[7929] = i[8569];
  assign o[7928] = i[8568];
  assign o[7927] = i[8567];
  assign o[7926] = i[8566];
  assign o[7925] = i[8565];
  assign o[7924] = i[8564];
  assign o[7923] = i[8563];
  assign o[7922] = i[8562];
  assign o[7921] = i[8561];
  assign o[7920] = i[8560];
  assign o[7919] = i[8559];
  assign o[7918] = i[8558];
  assign o[7917] = i[8557];
  assign o[7916] = i[8556];
  assign o[7915] = i[8555];
  assign o[7914] = i[8554];
  assign o[7913] = i[8553];
  assign o[7912] = i[8552];
  assign o[7911] = i[8551];
  assign o[7910] = i[8550];
  assign o[7909] = i[8549];
  assign o[7908] = i[8548];
  assign o[7907] = i[8547];
  assign o[7906] = i[8546];
  assign o[7905] = i[8545];
  assign o[7904] = i[8544];
  assign o[7903] = i[8543];
  assign o[7902] = i[8542];
  assign o[7901] = i[8541];
  assign o[7900] = i[8540];
  assign o[7899] = i[8539];
  assign o[7898] = i[8538];
  assign o[7897] = i[8537];
  assign o[7896] = i[8536];
  assign o[7895] = i[8535];
  assign o[7894] = i[8534];
  assign o[7893] = i[8533];
  assign o[7892] = i[8532];
  assign o[7891] = i[8531];
  assign o[7890] = i[8530];
  assign o[7889] = i[8529];
  assign o[7888] = i[8528];
  assign o[7887] = i[8527];
  assign o[7886] = i[8526];
  assign o[7885] = i[8525];
  assign o[7884] = i[8524];
  assign o[7883] = i[8523];
  assign o[7882] = i[8522];
  assign o[7881] = i[8521];
  assign o[7880] = i[8520];
  assign o[7879] = i[8519];
  assign o[7878] = i[8518];
  assign o[7877] = i[8517];
  assign o[7876] = i[8516];
  assign o[7875] = i[8515];
  assign o[7874] = i[8514];
  assign o[7873] = i[8513];
  assign o[7872] = i[8512];
  assign o[7871] = i[8511];
  assign o[7870] = i[8510];
  assign o[7869] = i[8509];
  assign o[7868] = i[8508];
  assign o[7867] = i[8507];
  assign o[7866] = i[8506];
  assign o[7865] = i[8505];
  assign o[7864] = i[8504];
  assign o[7863] = i[8503];
  assign o[7862] = i[8502];
  assign o[7861] = i[8501];
  assign o[7860] = i[8500];
  assign o[7859] = i[8499];
  assign o[7858] = i[8498];
  assign o[7857] = i[8497];
  assign o[7856] = i[8496];
  assign o[7855] = i[8495];
  assign o[7854] = i[8494];
  assign o[7853] = i[8493];
  assign o[7852] = i[8492];
  assign o[7851] = i[8491];
  assign o[7850] = i[8490];
  assign o[7849] = i[8489];
  assign o[7848] = i[8488];
  assign o[7847] = i[8487];
  assign o[7846] = i[8486];
  assign o[7845] = i[8485];
  assign o[7844] = i[8484];
  assign o[7843] = i[8483];
  assign o[7842] = i[8482];
  assign o[7841] = i[8481];
  assign o[7840] = i[8480];
  assign o[7839] = i[8479];
  assign o[7838] = i[8478];
  assign o[7837] = i[8477];
  assign o[7836] = i[8476];
  assign o[7835] = i[8475];
  assign o[7834] = i[8474];
  assign o[7833] = i[8473];
  assign o[7832] = i[8472];
  assign o[7831] = i[8471];
  assign o[7830] = i[8470];
  assign o[7829] = i[8469];
  assign o[7828] = i[8468];
  assign o[7827] = i[8467];
  assign o[7826] = i[8466];
  assign o[7825] = i[8465];
  assign o[7824] = i[8464];
  assign o[7823] = i[8463];
  assign o[7822] = i[8462];
  assign o[7821] = i[8461];
  assign o[7820] = i[8460];
  assign o[7819] = i[8459];
  assign o[7818] = i[8458];
  assign o[7817] = i[8457];
  assign o[7816] = i[8456];
  assign o[7815] = i[8455];
  assign o[7814] = i[8454];
  assign o[7813] = i[8453];
  assign o[7812] = i[8452];
  assign o[7811] = i[8451];
  assign o[7810] = i[8450];
  assign o[7809] = i[8449];
  assign o[7808] = i[8448];
  assign o[7807] = i[8703];
  assign o[7806] = i[8702];
  assign o[7805] = i[8701];
  assign o[7804] = i[8700];
  assign o[7803] = i[8699];
  assign o[7802] = i[8698];
  assign o[7801] = i[8697];
  assign o[7800] = i[8696];
  assign o[7799] = i[8695];
  assign o[7798] = i[8694];
  assign o[7797] = i[8693];
  assign o[7796] = i[8692];
  assign o[7795] = i[8691];
  assign o[7794] = i[8690];
  assign o[7793] = i[8689];
  assign o[7792] = i[8688];
  assign o[7791] = i[8687];
  assign o[7790] = i[8686];
  assign o[7789] = i[8685];
  assign o[7788] = i[8684];
  assign o[7787] = i[8683];
  assign o[7786] = i[8682];
  assign o[7785] = i[8681];
  assign o[7784] = i[8680];
  assign o[7783] = i[8679];
  assign o[7782] = i[8678];
  assign o[7781] = i[8677];
  assign o[7780] = i[8676];
  assign o[7779] = i[8675];
  assign o[7778] = i[8674];
  assign o[7777] = i[8673];
  assign o[7776] = i[8672];
  assign o[7775] = i[8671];
  assign o[7774] = i[8670];
  assign o[7773] = i[8669];
  assign o[7772] = i[8668];
  assign o[7771] = i[8667];
  assign o[7770] = i[8666];
  assign o[7769] = i[8665];
  assign o[7768] = i[8664];
  assign o[7767] = i[8663];
  assign o[7766] = i[8662];
  assign o[7765] = i[8661];
  assign o[7764] = i[8660];
  assign o[7763] = i[8659];
  assign o[7762] = i[8658];
  assign o[7761] = i[8657];
  assign o[7760] = i[8656];
  assign o[7759] = i[8655];
  assign o[7758] = i[8654];
  assign o[7757] = i[8653];
  assign o[7756] = i[8652];
  assign o[7755] = i[8651];
  assign o[7754] = i[8650];
  assign o[7753] = i[8649];
  assign o[7752] = i[8648];
  assign o[7751] = i[8647];
  assign o[7750] = i[8646];
  assign o[7749] = i[8645];
  assign o[7748] = i[8644];
  assign o[7747] = i[8643];
  assign o[7746] = i[8642];
  assign o[7745] = i[8641];
  assign o[7744] = i[8640];
  assign o[7743] = i[8639];
  assign o[7742] = i[8638];
  assign o[7741] = i[8637];
  assign o[7740] = i[8636];
  assign o[7739] = i[8635];
  assign o[7738] = i[8634];
  assign o[7737] = i[8633];
  assign o[7736] = i[8632];
  assign o[7735] = i[8631];
  assign o[7734] = i[8630];
  assign o[7733] = i[8629];
  assign o[7732] = i[8628];
  assign o[7731] = i[8627];
  assign o[7730] = i[8626];
  assign o[7729] = i[8625];
  assign o[7728] = i[8624];
  assign o[7727] = i[8623];
  assign o[7726] = i[8622];
  assign o[7725] = i[8621];
  assign o[7724] = i[8620];
  assign o[7723] = i[8619];
  assign o[7722] = i[8618];
  assign o[7721] = i[8617];
  assign o[7720] = i[8616];
  assign o[7719] = i[8615];
  assign o[7718] = i[8614];
  assign o[7717] = i[8613];
  assign o[7716] = i[8612];
  assign o[7715] = i[8611];
  assign o[7714] = i[8610];
  assign o[7713] = i[8609];
  assign o[7712] = i[8608];
  assign o[7711] = i[8607];
  assign o[7710] = i[8606];
  assign o[7709] = i[8605];
  assign o[7708] = i[8604];
  assign o[7707] = i[8603];
  assign o[7706] = i[8602];
  assign o[7705] = i[8601];
  assign o[7704] = i[8600];
  assign o[7703] = i[8599];
  assign o[7702] = i[8598];
  assign o[7701] = i[8597];
  assign o[7700] = i[8596];
  assign o[7699] = i[8595];
  assign o[7698] = i[8594];
  assign o[7697] = i[8593];
  assign o[7696] = i[8592];
  assign o[7695] = i[8591];
  assign o[7694] = i[8590];
  assign o[7693] = i[8589];
  assign o[7692] = i[8588];
  assign o[7691] = i[8587];
  assign o[7690] = i[8586];
  assign o[7689] = i[8585];
  assign o[7688] = i[8584];
  assign o[7687] = i[8583];
  assign o[7686] = i[8582];
  assign o[7685] = i[8581];
  assign o[7684] = i[8580];
  assign o[7683] = i[8579];
  assign o[7682] = i[8578];
  assign o[7681] = i[8577];
  assign o[7680] = i[8576];
  assign o[7679] = i[8831];
  assign o[7678] = i[8830];
  assign o[7677] = i[8829];
  assign o[7676] = i[8828];
  assign o[7675] = i[8827];
  assign o[7674] = i[8826];
  assign o[7673] = i[8825];
  assign o[7672] = i[8824];
  assign o[7671] = i[8823];
  assign o[7670] = i[8822];
  assign o[7669] = i[8821];
  assign o[7668] = i[8820];
  assign o[7667] = i[8819];
  assign o[7666] = i[8818];
  assign o[7665] = i[8817];
  assign o[7664] = i[8816];
  assign o[7663] = i[8815];
  assign o[7662] = i[8814];
  assign o[7661] = i[8813];
  assign o[7660] = i[8812];
  assign o[7659] = i[8811];
  assign o[7658] = i[8810];
  assign o[7657] = i[8809];
  assign o[7656] = i[8808];
  assign o[7655] = i[8807];
  assign o[7654] = i[8806];
  assign o[7653] = i[8805];
  assign o[7652] = i[8804];
  assign o[7651] = i[8803];
  assign o[7650] = i[8802];
  assign o[7649] = i[8801];
  assign o[7648] = i[8800];
  assign o[7647] = i[8799];
  assign o[7646] = i[8798];
  assign o[7645] = i[8797];
  assign o[7644] = i[8796];
  assign o[7643] = i[8795];
  assign o[7642] = i[8794];
  assign o[7641] = i[8793];
  assign o[7640] = i[8792];
  assign o[7639] = i[8791];
  assign o[7638] = i[8790];
  assign o[7637] = i[8789];
  assign o[7636] = i[8788];
  assign o[7635] = i[8787];
  assign o[7634] = i[8786];
  assign o[7633] = i[8785];
  assign o[7632] = i[8784];
  assign o[7631] = i[8783];
  assign o[7630] = i[8782];
  assign o[7629] = i[8781];
  assign o[7628] = i[8780];
  assign o[7627] = i[8779];
  assign o[7626] = i[8778];
  assign o[7625] = i[8777];
  assign o[7624] = i[8776];
  assign o[7623] = i[8775];
  assign o[7622] = i[8774];
  assign o[7621] = i[8773];
  assign o[7620] = i[8772];
  assign o[7619] = i[8771];
  assign o[7618] = i[8770];
  assign o[7617] = i[8769];
  assign o[7616] = i[8768];
  assign o[7615] = i[8767];
  assign o[7614] = i[8766];
  assign o[7613] = i[8765];
  assign o[7612] = i[8764];
  assign o[7611] = i[8763];
  assign o[7610] = i[8762];
  assign o[7609] = i[8761];
  assign o[7608] = i[8760];
  assign o[7607] = i[8759];
  assign o[7606] = i[8758];
  assign o[7605] = i[8757];
  assign o[7604] = i[8756];
  assign o[7603] = i[8755];
  assign o[7602] = i[8754];
  assign o[7601] = i[8753];
  assign o[7600] = i[8752];
  assign o[7599] = i[8751];
  assign o[7598] = i[8750];
  assign o[7597] = i[8749];
  assign o[7596] = i[8748];
  assign o[7595] = i[8747];
  assign o[7594] = i[8746];
  assign o[7593] = i[8745];
  assign o[7592] = i[8744];
  assign o[7591] = i[8743];
  assign o[7590] = i[8742];
  assign o[7589] = i[8741];
  assign o[7588] = i[8740];
  assign o[7587] = i[8739];
  assign o[7586] = i[8738];
  assign o[7585] = i[8737];
  assign o[7584] = i[8736];
  assign o[7583] = i[8735];
  assign o[7582] = i[8734];
  assign o[7581] = i[8733];
  assign o[7580] = i[8732];
  assign o[7579] = i[8731];
  assign o[7578] = i[8730];
  assign o[7577] = i[8729];
  assign o[7576] = i[8728];
  assign o[7575] = i[8727];
  assign o[7574] = i[8726];
  assign o[7573] = i[8725];
  assign o[7572] = i[8724];
  assign o[7571] = i[8723];
  assign o[7570] = i[8722];
  assign o[7569] = i[8721];
  assign o[7568] = i[8720];
  assign o[7567] = i[8719];
  assign o[7566] = i[8718];
  assign o[7565] = i[8717];
  assign o[7564] = i[8716];
  assign o[7563] = i[8715];
  assign o[7562] = i[8714];
  assign o[7561] = i[8713];
  assign o[7560] = i[8712];
  assign o[7559] = i[8711];
  assign o[7558] = i[8710];
  assign o[7557] = i[8709];
  assign o[7556] = i[8708];
  assign o[7555] = i[8707];
  assign o[7554] = i[8706];
  assign o[7553] = i[8705];
  assign o[7552] = i[8704];
  assign o[7551] = i[8959];
  assign o[7550] = i[8958];
  assign o[7549] = i[8957];
  assign o[7548] = i[8956];
  assign o[7547] = i[8955];
  assign o[7546] = i[8954];
  assign o[7545] = i[8953];
  assign o[7544] = i[8952];
  assign o[7543] = i[8951];
  assign o[7542] = i[8950];
  assign o[7541] = i[8949];
  assign o[7540] = i[8948];
  assign o[7539] = i[8947];
  assign o[7538] = i[8946];
  assign o[7537] = i[8945];
  assign o[7536] = i[8944];
  assign o[7535] = i[8943];
  assign o[7534] = i[8942];
  assign o[7533] = i[8941];
  assign o[7532] = i[8940];
  assign o[7531] = i[8939];
  assign o[7530] = i[8938];
  assign o[7529] = i[8937];
  assign o[7528] = i[8936];
  assign o[7527] = i[8935];
  assign o[7526] = i[8934];
  assign o[7525] = i[8933];
  assign o[7524] = i[8932];
  assign o[7523] = i[8931];
  assign o[7522] = i[8930];
  assign o[7521] = i[8929];
  assign o[7520] = i[8928];
  assign o[7519] = i[8927];
  assign o[7518] = i[8926];
  assign o[7517] = i[8925];
  assign o[7516] = i[8924];
  assign o[7515] = i[8923];
  assign o[7514] = i[8922];
  assign o[7513] = i[8921];
  assign o[7512] = i[8920];
  assign o[7511] = i[8919];
  assign o[7510] = i[8918];
  assign o[7509] = i[8917];
  assign o[7508] = i[8916];
  assign o[7507] = i[8915];
  assign o[7506] = i[8914];
  assign o[7505] = i[8913];
  assign o[7504] = i[8912];
  assign o[7503] = i[8911];
  assign o[7502] = i[8910];
  assign o[7501] = i[8909];
  assign o[7500] = i[8908];
  assign o[7499] = i[8907];
  assign o[7498] = i[8906];
  assign o[7497] = i[8905];
  assign o[7496] = i[8904];
  assign o[7495] = i[8903];
  assign o[7494] = i[8902];
  assign o[7493] = i[8901];
  assign o[7492] = i[8900];
  assign o[7491] = i[8899];
  assign o[7490] = i[8898];
  assign o[7489] = i[8897];
  assign o[7488] = i[8896];
  assign o[7487] = i[8895];
  assign o[7486] = i[8894];
  assign o[7485] = i[8893];
  assign o[7484] = i[8892];
  assign o[7483] = i[8891];
  assign o[7482] = i[8890];
  assign o[7481] = i[8889];
  assign o[7480] = i[8888];
  assign o[7479] = i[8887];
  assign o[7478] = i[8886];
  assign o[7477] = i[8885];
  assign o[7476] = i[8884];
  assign o[7475] = i[8883];
  assign o[7474] = i[8882];
  assign o[7473] = i[8881];
  assign o[7472] = i[8880];
  assign o[7471] = i[8879];
  assign o[7470] = i[8878];
  assign o[7469] = i[8877];
  assign o[7468] = i[8876];
  assign o[7467] = i[8875];
  assign o[7466] = i[8874];
  assign o[7465] = i[8873];
  assign o[7464] = i[8872];
  assign o[7463] = i[8871];
  assign o[7462] = i[8870];
  assign o[7461] = i[8869];
  assign o[7460] = i[8868];
  assign o[7459] = i[8867];
  assign o[7458] = i[8866];
  assign o[7457] = i[8865];
  assign o[7456] = i[8864];
  assign o[7455] = i[8863];
  assign o[7454] = i[8862];
  assign o[7453] = i[8861];
  assign o[7452] = i[8860];
  assign o[7451] = i[8859];
  assign o[7450] = i[8858];
  assign o[7449] = i[8857];
  assign o[7448] = i[8856];
  assign o[7447] = i[8855];
  assign o[7446] = i[8854];
  assign o[7445] = i[8853];
  assign o[7444] = i[8852];
  assign o[7443] = i[8851];
  assign o[7442] = i[8850];
  assign o[7441] = i[8849];
  assign o[7440] = i[8848];
  assign o[7439] = i[8847];
  assign o[7438] = i[8846];
  assign o[7437] = i[8845];
  assign o[7436] = i[8844];
  assign o[7435] = i[8843];
  assign o[7434] = i[8842];
  assign o[7433] = i[8841];
  assign o[7432] = i[8840];
  assign o[7431] = i[8839];
  assign o[7430] = i[8838];
  assign o[7429] = i[8837];
  assign o[7428] = i[8836];
  assign o[7427] = i[8835];
  assign o[7426] = i[8834];
  assign o[7425] = i[8833];
  assign o[7424] = i[8832];
  assign o[7423] = i[9087];
  assign o[7422] = i[9086];
  assign o[7421] = i[9085];
  assign o[7420] = i[9084];
  assign o[7419] = i[9083];
  assign o[7418] = i[9082];
  assign o[7417] = i[9081];
  assign o[7416] = i[9080];
  assign o[7415] = i[9079];
  assign o[7414] = i[9078];
  assign o[7413] = i[9077];
  assign o[7412] = i[9076];
  assign o[7411] = i[9075];
  assign o[7410] = i[9074];
  assign o[7409] = i[9073];
  assign o[7408] = i[9072];
  assign o[7407] = i[9071];
  assign o[7406] = i[9070];
  assign o[7405] = i[9069];
  assign o[7404] = i[9068];
  assign o[7403] = i[9067];
  assign o[7402] = i[9066];
  assign o[7401] = i[9065];
  assign o[7400] = i[9064];
  assign o[7399] = i[9063];
  assign o[7398] = i[9062];
  assign o[7397] = i[9061];
  assign o[7396] = i[9060];
  assign o[7395] = i[9059];
  assign o[7394] = i[9058];
  assign o[7393] = i[9057];
  assign o[7392] = i[9056];
  assign o[7391] = i[9055];
  assign o[7390] = i[9054];
  assign o[7389] = i[9053];
  assign o[7388] = i[9052];
  assign o[7387] = i[9051];
  assign o[7386] = i[9050];
  assign o[7385] = i[9049];
  assign o[7384] = i[9048];
  assign o[7383] = i[9047];
  assign o[7382] = i[9046];
  assign o[7381] = i[9045];
  assign o[7380] = i[9044];
  assign o[7379] = i[9043];
  assign o[7378] = i[9042];
  assign o[7377] = i[9041];
  assign o[7376] = i[9040];
  assign o[7375] = i[9039];
  assign o[7374] = i[9038];
  assign o[7373] = i[9037];
  assign o[7372] = i[9036];
  assign o[7371] = i[9035];
  assign o[7370] = i[9034];
  assign o[7369] = i[9033];
  assign o[7368] = i[9032];
  assign o[7367] = i[9031];
  assign o[7366] = i[9030];
  assign o[7365] = i[9029];
  assign o[7364] = i[9028];
  assign o[7363] = i[9027];
  assign o[7362] = i[9026];
  assign o[7361] = i[9025];
  assign o[7360] = i[9024];
  assign o[7359] = i[9023];
  assign o[7358] = i[9022];
  assign o[7357] = i[9021];
  assign o[7356] = i[9020];
  assign o[7355] = i[9019];
  assign o[7354] = i[9018];
  assign o[7353] = i[9017];
  assign o[7352] = i[9016];
  assign o[7351] = i[9015];
  assign o[7350] = i[9014];
  assign o[7349] = i[9013];
  assign o[7348] = i[9012];
  assign o[7347] = i[9011];
  assign o[7346] = i[9010];
  assign o[7345] = i[9009];
  assign o[7344] = i[9008];
  assign o[7343] = i[9007];
  assign o[7342] = i[9006];
  assign o[7341] = i[9005];
  assign o[7340] = i[9004];
  assign o[7339] = i[9003];
  assign o[7338] = i[9002];
  assign o[7337] = i[9001];
  assign o[7336] = i[9000];
  assign o[7335] = i[8999];
  assign o[7334] = i[8998];
  assign o[7333] = i[8997];
  assign o[7332] = i[8996];
  assign o[7331] = i[8995];
  assign o[7330] = i[8994];
  assign o[7329] = i[8993];
  assign o[7328] = i[8992];
  assign o[7327] = i[8991];
  assign o[7326] = i[8990];
  assign o[7325] = i[8989];
  assign o[7324] = i[8988];
  assign o[7323] = i[8987];
  assign o[7322] = i[8986];
  assign o[7321] = i[8985];
  assign o[7320] = i[8984];
  assign o[7319] = i[8983];
  assign o[7318] = i[8982];
  assign o[7317] = i[8981];
  assign o[7316] = i[8980];
  assign o[7315] = i[8979];
  assign o[7314] = i[8978];
  assign o[7313] = i[8977];
  assign o[7312] = i[8976];
  assign o[7311] = i[8975];
  assign o[7310] = i[8974];
  assign o[7309] = i[8973];
  assign o[7308] = i[8972];
  assign o[7307] = i[8971];
  assign o[7306] = i[8970];
  assign o[7305] = i[8969];
  assign o[7304] = i[8968];
  assign o[7303] = i[8967];
  assign o[7302] = i[8966];
  assign o[7301] = i[8965];
  assign o[7300] = i[8964];
  assign o[7299] = i[8963];
  assign o[7298] = i[8962];
  assign o[7297] = i[8961];
  assign o[7296] = i[8960];
  assign o[7295] = i[9215];
  assign o[7294] = i[9214];
  assign o[7293] = i[9213];
  assign o[7292] = i[9212];
  assign o[7291] = i[9211];
  assign o[7290] = i[9210];
  assign o[7289] = i[9209];
  assign o[7288] = i[9208];
  assign o[7287] = i[9207];
  assign o[7286] = i[9206];
  assign o[7285] = i[9205];
  assign o[7284] = i[9204];
  assign o[7283] = i[9203];
  assign o[7282] = i[9202];
  assign o[7281] = i[9201];
  assign o[7280] = i[9200];
  assign o[7279] = i[9199];
  assign o[7278] = i[9198];
  assign o[7277] = i[9197];
  assign o[7276] = i[9196];
  assign o[7275] = i[9195];
  assign o[7274] = i[9194];
  assign o[7273] = i[9193];
  assign o[7272] = i[9192];
  assign o[7271] = i[9191];
  assign o[7270] = i[9190];
  assign o[7269] = i[9189];
  assign o[7268] = i[9188];
  assign o[7267] = i[9187];
  assign o[7266] = i[9186];
  assign o[7265] = i[9185];
  assign o[7264] = i[9184];
  assign o[7263] = i[9183];
  assign o[7262] = i[9182];
  assign o[7261] = i[9181];
  assign o[7260] = i[9180];
  assign o[7259] = i[9179];
  assign o[7258] = i[9178];
  assign o[7257] = i[9177];
  assign o[7256] = i[9176];
  assign o[7255] = i[9175];
  assign o[7254] = i[9174];
  assign o[7253] = i[9173];
  assign o[7252] = i[9172];
  assign o[7251] = i[9171];
  assign o[7250] = i[9170];
  assign o[7249] = i[9169];
  assign o[7248] = i[9168];
  assign o[7247] = i[9167];
  assign o[7246] = i[9166];
  assign o[7245] = i[9165];
  assign o[7244] = i[9164];
  assign o[7243] = i[9163];
  assign o[7242] = i[9162];
  assign o[7241] = i[9161];
  assign o[7240] = i[9160];
  assign o[7239] = i[9159];
  assign o[7238] = i[9158];
  assign o[7237] = i[9157];
  assign o[7236] = i[9156];
  assign o[7235] = i[9155];
  assign o[7234] = i[9154];
  assign o[7233] = i[9153];
  assign o[7232] = i[9152];
  assign o[7231] = i[9151];
  assign o[7230] = i[9150];
  assign o[7229] = i[9149];
  assign o[7228] = i[9148];
  assign o[7227] = i[9147];
  assign o[7226] = i[9146];
  assign o[7225] = i[9145];
  assign o[7224] = i[9144];
  assign o[7223] = i[9143];
  assign o[7222] = i[9142];
  assign o[7221] = i[9141];
  assign o[7220] = i[9140];
  assign o[7219] = i[9139];
  assign o[7218] = i[9138];
  assign o[7217] = i[9137];
  assign o[7216] = i[9136];
  assign o[7215] = i[9135];
  assign o[7214] = i[9134];
  assign o[7213] = i[9133];
  assign o[7212] = i[9132];
  assign o[7211] = i[9131];
  assign o[7210] = i[9130];
  assign o[7209] = i[9129];
  assign o[7208] = i[9128];
  assign o[7207] = i[9127];
  assign o[7206] = i[9126];
  assign o[7205] = i[9125];
  assign o[7204] = i[9124];
  assign o[7203] = i[9123];
  assign o[7202] = i[9122];
  assign o[7201] = i[9121];
  assign o[7200] = i[9120];
  assign o[7199] = i[9119];
  assign o[7198] = i[9118];
  assign o[7197] = i[9117];
  assign o[7196] = i[9116];
  assign o[7195] = i[9115];
  assign o[7194] = i[9114];
  assign o[7193] = i[9113];
  assign o[7192] = i[9112];
  assign o[7191] = i[9111];
  assign o[7190] = i[9110];
  assign o[7189] = i[9109];
  assign o[7188] = i[9108];
  assign o[7187] = i[9107];
  assign o[7186] = i[9106];
  assign o[7185] = i[9105];
  assign o[7184] = i[9104];
  assign o[7183] = i[9103];
  assign o[7182] = i[9102];
  assign o[7181] = i[9101];
  assign o[7180] = i[9100];
  assign o[7179] = i[9099];
  assign o[7178] = i[9098];
  assign o[7177] = i[9097];
  assign o[7176] = i[9096];
  assign o[7175] = i[9095];
  assign o[7174] = i[9094];
  assign o[7173] = i[9093];
  assign o[7172] = i[9092];
  assign o[7171] = i[9091];
  assign o[7170] = i[9090];
  assign o[7169] = i[9089];
  assign o[7168] = i[9088];
  assign o[7167] = i[9343];
  assign o[7166] = i[9342];
  assign o[7165] = i[9341];
  assign o[7164] = i[9340];
  assign o[7163] = i[9339];
  assign o[7162] = i[9338];
  assign o[7161] = i[9337];
  assign o[7160] = i[9336];
  assign o[7159] = i[9335];
  assign o[7158] = i[9334];
  assign o[7157] = i[9333];
  assign o[7156] = i[9332];
  assign o[7155] = i[9331];
  assign o[7154] = i[9330];
  assign o[7153] = i[9329];
  assign o[7152] = i[9328];
  assign o[7151] = i[9327];
  assign o[7150] = i[9326];
  assign o[7149] = i[9325];
  assign o[7148] = i[9324];
  assign o[7147] = i[9323];
  assign o[7146] = i[9322];
  assign o[7145] = i[9321];
  assign o[7144] = i[9320];
  assign o[7143] = i[9319];
  assign o[7142] = i[9318];
  assign o[7141] = i[9317];
  assign o[7140] = i[9316];
  assign o[7139] = i[9315];
  assign o[7138] = i[9314];
  assign o[7137] = i[9313];
  assign o[7136] = i[9312];
  assign o[7135] = i[9311];
  assign o[7134] = i[9310];
  assign o[7133] = i[9309];
  assign o[7132] = i[9308];
  assign o[7131] = i[9307];
  assign o[7130] = i[9306];
  assign o[7129] = i[9305];
  assign o[7128] = i[9304];
  assign o[7127] = i[9303];
  assign o[7126] = i[9302];
  assign o[7125] = i[9301];
  assign o[7124] = i[9300];
  assign o[7123] = i[9299];
  assign o[7122] = i[9298];
  assign o[7121] = i[9297];
  assign o[7120] = i[9296];
  assign o[7119] = i[9295];
  assign o[7118] = i[9294];
  assign o[7117] = i[9293];
  assign o[7116] = i[9292];
  assign o[7115] = i[9291];
  assign o[7114] = i[9290];
  assign o[7113] = i[9289];
  assign o[7112] = i[9288];
  assign o[7111] = i[9287];
  assign o[7110] = i[9286];
  assign o[7109] = i[9285];
  assign o[7108] = i[9284];
  assign o[7107] = i[9283];
  assign o[7106] = i[9282];
  assign o[7105] = i[9281];
  assign o[7104] = i[9280];
  assign o[7103] = i[9279];
  assign o[7102] = i[9278];
  assign o[7101] = i[9277];
  assign o[7100] = i[9276];
  assign o[7099] = i[9275];
  assign o[7098] = i[9274];
  assign o[7097] = i[9273];
  assign o[7096] = i[9272];
  assign o[7095] = i[9271];
  assign o[7094] = i[9270];
  assign o[7093] = i[9269];
  assign o[7092] = i[9268];
  assign o[7091] = i[9267];
  assign o[7090] = i[9266];
  assign o[7089] = i[9265];
  assign o[7088] = i[9264];
  assign o[7087] = i[9263];
  assign o[7086] = i[9262];
  assign o[7085] = i[9261];
  assign o[7084] = i[9260];
  assign o[7083] = i[9259];
  assign o[7082] = i[9258];
  assign o[7081] = i[9257];
  assign o[7080] = i[9256];
  assign o[7079] = i[9255];
  assign o[7078] = i[9254];
  assign o[7077] = i[9253];
  assign o[7076] = i[9252];
  assign o[7075] = i[9251];
  assign o[7074] = i[9250];
  assign o[7073] = i[9249];
  assign o[7072] = i[9248];
  assign o[7071] = i[9247];
  assign o[7070] = i[9246];
  assign o[7069] = i[9245];
  assign o[7068] = i[9244];
  assign o[7067] = i[9243];
  assign o[7066] = i[9242];
  assign o[7065] = i[9241];
  assign o[7064] = i[9240];
  assign o[7063] = i[9239];
  assign o[7062] = i[9238];
  assign o[7061] = i[9237];
  assign o[7060] = i[9236];
  assign o[7059] = i[9235];
  assign o[7058] = i[9234];
  assign o[7057] = i[9233];
  assign o[7056] = i[9232];
  assign o[7055] = i[9231];
  assign o[7054] = i[9230];
  assign o[7053] = i[9229];
  assign o[7052] = i[9228];
  assign o[7051] = i[9227];
  assign o[7050] = i[9226];
  assign o[7049] = i[9225];
  assign o[7048] = i[9224];
  assign o[7047] = i[9223];
  assign o[7046] = i[9222];
  assign o[7045] = i[9221];
  assign o[7044] = i[9220];
  assign o[7043] = i[9219];
  assign o[7042] = i[9218];
  assign o[7041] = i[9217];
  assign o[7040] = i[9216];
  assign o[7039] = i[9471];
  assign o[7038] = i[9470];
  assign o[7037] = i[9469];
  assign o[7036] = i[9468];
  assign o[7035] = i[9467];
  assign o[7034] = i[9466];
  assign o[7033] = i[9465];
  assign o[7032] = i[9464];
  assign o[7031] = i[9463];
  assign o[7030] = i[9462];
  assign o[7029] = i[9461];
  assign o[7028] = i[9460];
  assign o[7027] = i[9459];
  assign o[7026] = i[9458];
  assign o[7025] = i[9457];
  assign o[7024] = i[9456];
  assign o[7023] = i[9455];
  assign o[7022] = i[9454];
  assign o[7021] = i[9453];
  assign o[7020] = i[9452];
  assign o[7019] = i[9451];
  assign o[7018] = i[9450];
  assign o[7017] = i[9449];
  assign o[7016] = i[9448];
  assign o[7015] = i[9447];
  assign o[7014] = i[9446];
  assign o[7013] = i[9445];
  assign o[7012] = i[9444];
  assign o[7011] = i[9443];
  assign o[7010] = i[9442];
  assign o[7009] = i[9441];
  assign o[7008] = i[9440];
  assign o[7007] = i[9439];
  assign o[7006] = i[9438];
  assign o[7005] = i[9437];
  assign o[7004] = i[9436];
  assign o[7003] = i[9435];
  assign o[7002] = i[9434];
  assign o[7001] = i[9433];
  assign o[7000] = i[9432];
  assign o[6999] = i[9431];
  assign o[6998] = i[9430];
  assign o[6997] = i[9429];
  assign o[6996] = i[9428];
  assign o[6995] = i[9427];
  assign o[6994] = i[9426];
  assign o[6993] = i[9425];
  assign o[6992] = i[9424];
  assign o[6991] = i[9423];
  assign o[6990] = i[9422];
  assign o[6989] = i[9421];
  assign o[6988] = i[9420];
  assign o[6987] = i[9419];
  assign o[6986] = i[9418];
  assign o[6985] = i[9417];
  assign o[6984] = i[9416];
  assign o[6983] = i[9415];
  assign o[6982] = i[9414];
  assign o[6981] = i[9413];
  assign o[6980] = i[9412];
  assign o[6979] = i[9411];
  assign o[6978] = i[9410];
  assign o[6977] = i[9409];
  assign o[6976] = i[9408];
  assign o[6975] = i[9407];
  assign o[6974] = i[9406];
  assign o[6973] = i[9405];
  assign o[6972] = i[9404];
  assign o[6971] = i[9403];
  assign o[6970] = i[9402];
  assign o[6969] = i[9401];
  assign o[6968] = i[9400];
  assign o[6967] = i[9399];
  assign o[6966] = i[9398];
  assign o[6965] = i[9397];
  assign o[6964] = i[9396];
  assign o[6963] = i[9395];
  assign o[6962] = i[9394];
  assign o[6961] = i[9393];
  assign o[6960] = i[9392];
  assign o[6959] = i[9391];
  assign o[6958] = i[9390];
  assign o[6957] = i[9389];
  assign o[6956] = i[9388];
  assign o[6955] = i[9387];
  assign o[6954] = i[9386];
  assign o[6953] = i[9385];
  assign o[6952] = i[9384];
  assign o[6951] = i[9383];
  assign o[6950] = i[9382];
  assign o[6949] = i[9381];
  assign o[6948] = i[9380];
  assign o[6947] = i[9379];
  assign o[6946] = i[9378];
  assign o[6945] = i[9377];
  assign o[6944] = i[9376];
  assign o[6943] = i[9375];
  assign o[6942] = i[9374];
  assign o[6941] = i[9373];
  assign o[6940] = i[9372];
  assign o[6939] = i[9371];
  assign o[6938] = i[9370];
  assign o[6937] = i[9369];
  assign o[6936] = i[9368];
  assign o[6935] = i[9367];
  assign o[6934] = i[9366];
  assign o[6933] = i[9365];
  assign o[6932] = i[9364];
  assign o[6931] = i[9363];
  assign o[6930] = i[9362];
  assign o[6929] = i[9361];
  assign o[6928] = i[9360];
  assign o[6927] = i[9359];
  assign o[6926] = i[9358];
  assign o[6925] = i[9357];
  assign o[6924] = i[9356];
  assign o[6923] = i[9355];
  assign o[6922] = i[9354];
  assign o[6921] = i[9353];
  assign o[6920] = i[9352];
  assign o[6919] = i[9351];
  assign o[6918] = i[9350];
  assign o[6917] = i[9349];
  assign o[6916] = i[9348];
  assign o[6915] = i[9347];
  assign o[6914] = i[9346];
  assign o[6913] = i[9345];
  assign o[6912] = i[9344];
  assign o[6911] = i[9599];
  assign o[6910] = i[9598];
  assign o[6909] = i[9597];
  assign o[6908] = i[9596];
  assign o[6907] = i[9595];
  assign o[6906] = i[9594];
  assign o[6905] = i[9593];
  assign o[6904] = i[9592];
  assign o[6903] = i[9591];
  assign o[6902] = i[9590];
  assign o[6901] = i[9589];
  assign o[6900] = i[9588];
  assign o[6899] = i[9587];
  assign o[6898] = i[9586];
  assign o[6897] = i[9585];
  assign o[6896] = i[9584];
  assign o[6895] = i[9583];
  assign o[6894] = i[9582];
  assign o[6893] = i[9581];
  assign o[6892] = i[9580];
  assign o[6891] = i[9579];
  assign o[6890] = i[9578];
  assign o[6889] = i[9577];
  assign o[6888] = i[9576];
  assign o[6887] = i[9575];
  assign o[6886] = i[9574];
  assign o[6885] = i[9573];
  assign o[6884] = i[9572];
  assign o[6883] = i[9571];
  assign o[6882] = i[9570];
  assign o[6881] = i[9569];
  assign o[6880] = i[9568];
  assign o[6879] = i[9567];
  assign o[6878] = i[9566];
  assign o[6877] = i[9565];
  assign o[6876] = i[9564];
  assign o[6875] = i[9563];
  assign o[6874] = i[9562];
  assign o[6873] = i[9561];
  assign o[6872] = i[9560];
  assign o[6871] = i[9559];
  assign o[6870] = i[9558];
  assign o[6869] = i[9557];
  assign o[6868] = i[9556];
  assign o[6867] = i[9555];
  assign o[6866] = i[9554];
  assign o[6865] = i[9553];
  assign o[6864] = i[9552];
  assign o[6863] = i[9551];
  assign o[6862] = i[9550];
  assign o[6861] = i[9549];
  assign o[6860] = i[9548];
  assign o[6859] = i[9547];
  assign o[6858] = i[9546];
  assign o[6857] = i[9545];
  assign o[6856] = i[9544];
  assign o[6855] = i[9543];
  assign o[6854] = i[9542];
  assign o[6853] = i[9541];
  assign o[6852] = i[9540];
  assign o[6851] = i[9539];
  assign o[6850] = i[9538];
  assign o[6849] = i[9537];
  assign o[6848] = i[9536];
  assign o[6847] = i[9535];
  assign o[6846] = i[9534];
  assign o[6845] = i[9533];
  assign o[6844] = i[9532];
  assign o[6843] = i[9531];
  assign o[6842] = i[9530];
  assign o[6841] = i[9529];
  assign o[6840] = i[9528];
  assign o[6839] = i[9527];
  assign o[6838] = i[9526];
  assign o[6837] = i[9525];
  assign o[6836] = i[9524];
  assign o[6835] = i[9523];
  assign o[6834] = i[9522];
  assign o[6833] = i[9521];
  assign o[6832] = i[9520];
  assign o[6831] = i[9519];
  assign o[6830] = i[9518];
  assign o[6829] = i[9517];
  assign o[6828] = i[9516];
  assign o[6827] = i[9515];
  assign o[6826] = i[9514];
  assign o[6825] = i[9513];
  assign o[6824] = i[9512];
  assign o[6823] = i[9511];
  assign o[6822] = i[9510];
  assign o[6821] = i[9509];
  assign o[6820] = i[9508];
  assign o[6819] = i[9507];
  assign o[6818] = i[9506];
  assign o[6817] = i[9505];
  assign o[6816] = i[9504];
  assign o[6815] = i[9503];
  assign o[6814] = i[9502];
  assign o[6813] = i[9501];
  assign o[6812] = i[9500];
  assign o[6811] = i[9499];
  assign o[6810] = i[9498];
  assign o[6809] = i[9497];
  assign o[6808] = i[9496];
  assign o[6807] = i[9495];
  assign o[6806] = i[9494];
  assign o[6805] = i[9493];
  assign o[6804] = i[9492];
  assign o[6803] = i[9491];
  assign o[6802] = i[9490];
  assign o[6801] = i[9489];
  assign o[6800] = i[9488];
  assign o[6799] = i[9487];
  assign o[6798] = i[9486];
  assign o[6797] = i[9485];
  assign o[6796] = i[9484];
  assign o[6795] = i[9483];
  assign o[6794] = i[9482];
  assign o[6793] = i[9481];
  assign o[6792] = i[9480];
  assign o[6791] = i[9479];
  assign o[6790] = i[9478];
  assign o[6789] = i[9477];
  assign o[6788] = i[9476];
  assign o[6787] = i[9475];
  assign o[6786] = i[9474];
  assign o[6785] = i[9473];
  assign o[6784] = i[9472];
  assign o[6783] = i[9727];
  assign o[6782] = i[9726];
  assign o[6781] = i[9725];
  assign o[6780] = i[9724];
  assign o[6779] = i[9723];
  assign o[6778] = i[9722];
  assign o[6777] = i[9721];
  assign o[6776] = i[9720];
  assign o[6775] = i[9719];
  assign o[6774] = i[9718];
  assign o[6773] = i[9717];
  assign o[6772] = i[9716];
  assign o[6771] = i[9715];
  assign o[6770] = i[9714];
  assign o[6769] = i[9713];
  assign o[6768] = i[9712];
  assign o[6767] = i[9711];
  assign o[6766] = i[9710];
  assign o[6765] = i[9709];
  assign o[6764] = i[9708];
  assign o[6763] = i[9707];
  assign o[6762] = i[9706];
  assign o[6761] = i[9705];
  assign o[6760] = i[9704];
  assign o[6759] = i[9703];
  assign o[6758] = i[9702];
  assign o[6757] = i[9701];
  assign o[6756] = i[9700];
  assign o[6755] = i[9699];
  assign o[6754] = i[9698];
  assign o[6753] = i[9697];
  assign o[6752] = i[9696];
  assign o[6751] = i[9695];
  assign o[6750] = i[9694];
  assign o[6749] = i[9693];
  assign o[6748] = i[9692];
  assign o[6747] = i[9691];
  assign o[6746] = i[9690];
  assign o[6745] = i[9689];
  assign o[6744] = i[9688];
  assign o[6743] = i[9687];
  assign o[6742] = i[9686];
  assign o[6741] = i[9685];
  assign o[6740] = i[9684];
  assign o[6739] = i[9683];
  assign o[6738] = i[9682];
  assign o[6737] = i[9681];
  assign o[6736] = i[9680];
  assign o[6735] = i[9679];
  assign o[6734] = i[9678];
  assign o[6733] = i[9677];
  assign o[6732] = i[9676];
  assign o[6731] = i[9675];
  assign o[6730] = i[9674];
  assign o[6729] = i[9673];
  assign o[6728] = i[9672];
  assign o[6727] = i[9671];
  assign o[6726] = i[9670];
  assign o[6725] = i[9669];
  assign o[6724] = i[9668];
  assign o[6723] = i[9667];
  assign o[6722] = i[9666];
  assign o[6721] = i[9665];
  assign o[6720] = i[9664];
  assign o[6719] = i[9663];
  assign o[6718] = i[9662];
  assign o[6717] = i[9661];
  assign o[6716] = i[9660];
  assign o[6715] = i[9659];
  assign o[6714] = i[9658];
  assign o[6713] = i[9657];
  assign o[6712] = i[9656];
  assign o[6711] = i[9655];
  assign o[6710] = i[9654];
  assign o[6709] = i[9653];
  assign o[6708] = i[9652];
  assign o[6707] = i[9651];
  assign o[6706] = i[9650];
  assign o[6705] = i[9649];
  assign o[6704] = i[9648];
  assign o[6703] = i[9647];
  assign o[6702] = i[9646];
  assign o[6701] = i[9645];
  assign o[6700] = i[9644];
  assign o[6699] = i[9643];
  assign o[6698] = i[9642];
  assign o[6697] = i[9641];
  assign o[6696] = i[9640];
  assign o[6695] = i[9639];
  assign o[6694] = i[9638];
  assign o[6693] = i[9637];
  assign o[6692] = i[9636];
  assign o[6691] = i[9635];
  assign o[6690] = i[9634];
  assign o[6689] = i[9633];
  assign o[6688] = i[9632];
  assign o[6687] = i[9631];
  assign o[6686] = i[9630];
  assign o[6685] = i[9629];
  assign o[6684] = i[9628];
  assign o[6683] = i[9627];
  assign o[6682] = i[9626];
  assign o[6681] = i[9625];
  assign o[6680] = i[9624];
  assign o[6679] = i[9623];
  assign o[6678] = i[9622];
  assign o[6677] = i[9621];
  assign o[6676] = i[9620];
  assign o[6675] = i[9619];
  assign o[6674] = i[9618];
  assign o[6673] = i[9617];
  assign o[6672] = i[9616];
  assign o[6671] = i[9615];
  assign o[6670] = i[9614];
  assign o[6669] = i[9613];
  assign o[6668] = i[9612];
  assign o[6667] = i[9611];
  assign o[6666] = i[9610];
  assign o[6665] = i[9609];
  assign o[6664] = i[9608];
  assign o[6663] = i[9607];
  assign o[6662] = i[9606];
  assign o[6661] = i[9605];
  assign o[6660] = i[9604];
  assign o[6659] = i[9603];
  assign o[6658] = i[9602];
  assign o[6657] = i[9601];
  assign o[6656] = i[9600];
  assign o[6655] = i[9855];
  assign o[6654] = i[9854];
  assign o[6653] = i[9853];
  assign o[6652] = i[9852];
  assign o[6651] = i[9851];
  assign o[6650] = i[9850];
  assign o[6649] = i[9849];
  assign o[6648] = i[9848];
  assign o[6647] = i[9847];
  assign o[6646] = i[9846];
  assign o[6645] = i[9845];
  assign o[6644] = i[9844];
  assign o[6643] = i[9843];
  assign o[6642] = i[9842];
  assign o[6641] = i[9841];
  assign o[6640] = i[9840];
  assign o[6639] = i[9839];
  assign o[6638] = i[9838];
  assign o[6637] = i[9837];
  assign o[6636] = i[9836];
  assign o[6635] = i[9835];
  assign o[6634] = i[9834];
  assign o[6633] = i[9833];
  assign o[6632] = i[9832];
  assign o[6631] = i[9831];
  assign o[6630] = i[9830];
  assign o[6629] = i[9829];
  assign o[6628] = i[9828];
  assign o[6627] = i[9827];
  assign o[6626] = i[9826];
  assign o[6625] = i[9825];
  assign o[6624] = i[9824];
  assign o[6623] = i[9823];
  assign o[6622] = i[9822];
  assign o[6621] = i[9821];
  assign o[6620] = i[9820];
  assign o[6619] = i[9819];
  assign o[6618] = i[9818];
  assign o[6617] = i[9817];
  assign o[6616] = i[9816];
  assign o[6615] = i[9815];
  assign o[6614] = i[9814];
  assign o[6613] = i[9813];
  assign o[6612] = i[9812];
  assign o[6611] = i[9811];
  assign o[6610] = i[9810];
  assign o[6609] = i[9809];
  assign o[6608] = i[9808];
  assign o[6607] = i[9807];
  assign o[6606] = i[9806];
  assign o[6605] = i[9805];
  assign o[6604] = i[9804];
  assign o[6603] = i[9803];
  assign o[6602] = i[9802];
  assign o[6601] = i[9801];
  assign o[6600] = i[9800];
  assign o[6599] = i[9799];
  assign o[6598] = i[9798];
  assign o[6597] = i[9797];
  assign o[6596] = i[9796];
  assign o[6595] = i[9795];
  assign o[6594] = i[9794];
  assign o[6593] = i[9793];
  assign o[6592] = i[9792];
  assign o[6591] = i[9791];
  assign o[6590] = i[9790];
  assign o[6589] = i[9789];
  assign o[6588] = i[9788];
  assign o[6587] = i[9787];
  assign o[6586] = i[9786];
  assign o[6585] = i[9785];
  assign o[6584] = i[9784];
  assign o[6583] = i[9783];
  assign o[6582] = i[9782];
  assign o[6581] = i[9781];
  assign o[6580] = i[9780];
  assign o[6579] = i[9779];
  assign o[6578] = i[9778];
  assign o[6577] = i[9777];
  assign o[6576] = i[9776];
  assign o[6575] = i[9775];
  assign o[6574] = i[9774];
  assign o[6573] = i[9773];
  assign o[6572] = i[9772];
  assign o[6571] = i[9771];
  assign o[6570] = i[9770];
  assign o[6569] = i[9769];
  assign o[6568] = i[9768];
  assign o[6567] = i[9767];
  assign o[6566] = i[9766];
  assign o[6565] = i[9765];
  assign o[6564] = i[9764];
  assign o[6563] = i[9763];
  assign o[6562] = i[9762];
  assign o[6561] = i[9761];
  assign o[6560] = i[9760];
  assign o[6559] = i[9759];
  assign o[6558] = i[9758];
  assign o[6557] = i[9757];
  assign o[6556] = i[9756];
  assign o[6555] = i[9755];
  assign o[6554] = i[9754];
  assign o[6553] = i[9753];
  assign o[6552] = i[9752];
  assign o[6551] = i[9751];
  assign o[6550] = i[9750];
  assign o[6549] = i[9749];
  assign o[6548] = i[9748];
  assign o[6547] = i[9747];
  assign o[6546] = i[9746];
  assign o[6545] = i[9745];
  assign o[6544] = i[9744];
  assign o[6543] = i[9743];
  assign o[6542] = i[9742];
  assign o[6541] = i[9741];
  assign o[6540] = i[9740];
  assign o[6539] = i[9739];
  assign o[6538] = i[9738];
  assign o[6537] = i[9737];
  assign o[6536] = i[9736];
  assign o[6535] = i[9735];
  assign o[6534] = i[9734];
  assign o[6533] = i[9733];
  assign o[6532] = i[9732];
  assign o[6531] = i[9731];
  assign o[6530] = i[9730];
  assign o[6529] = i[9729];
  assign o[6528] = i[9728];
  assign o[6527] = i[9983];
  assign o[6526] = i[9982];
  assign o[6525] = i[9981];
  assign o[6524] = i[9980];
  assign o[6523] = i[9979];
  assign o[6522] = i[9978];
  assign o[6521] = i[9977];
  assign o[6520] = i[9976];
  assign o[6519] = i[9975];
  assign o[6518] = i[9974];
  assign o[6517] = i[9973];
  assign o[6516] = i[9972];
  assign o[6515] = i[9971];
  assign o[6514] = i[9970];
  assign o[6513] = i[9969];
  assign o[6512] = i[9968];
  assign o[6511] = i[9967];
  assign o[6510] = i[9966];
  assign o[6509] = i[9965];
  assign o[6508] = i[9964];
  assign o[6507] = i[9963];
  assign o[6506] = i[9962];
  assign o[6505] = i[9961];
  assign o[6504] = i[9960];
  assign o[6503] = i[9959];
  assign o[6502] = i[9958];
  assign o[6501] = i[9957];
  assign o[6500] = i[9956];
  assign o[6499] = i[9955];
  assign o[6498] = i[9954];
  assign o[6497] = i[9953];
  assign o[6496] = i[9952];
  assign o[6495] = i[9951];
  assign o[6494] = i[9950];
  assign o[6493] = i[9949];
  assign o[6492] = i[9948];
  assign o[6491] = i[9947];
  assign o[6490] = i[9946];
  assign o[6489] = i[9945];
  assign o[6488] = i[9944];
  assign o[6487] = i[9943];
  assign o[6486] = i[9942];
  assign o[6485] = i[9941];
  assign o[6484] = i[9940];
  assign o[6483] = i[9939];
  assign o[6482] = i[9938];
  assign o[6481] = i[9937];
  assign o[6480] = i[9936];
  assign o[6479] = i[9935];
  assign o[6478] = i[9934];
  assign o[6477] = i[9933];
  assign o[6476] = i[9932];
  assign o[6475] = i[9931];
  assign o[6474] = i[9930];
  assign o[6473] = i[9929];
  assign o[6472] = i[9928];
  assign o[6471] = i[9927];
  assign o[6470] = i[9926];
  assign o[6469] = i[9925];
  assign o[6468] = i[9924];
  assign o[6467] = i[9923];
  assign o[6466] = i[9922];
  assign o[6465] = i[9921];
  assign o[6464] = i[9920];
  assign o[6463] = i[9919];
  assign o[6462] = i[9918];
  assign o[6461] = i[9917];
  assign o[6460] = i[9916];
  assign o[6459] = i[9915];
  assign o[6458] = i[9914];
  assign o[6457] = i[9913];
  assign o[6456] = i[9912];
  assign o[6455] = i[9911];
  assign o[6454] = i[9910];
  assign o[6453] = i[9909];
  assign o[6452] = i[9908];
  assign o[6451] = i[9907];
  assign o[6450] = i[9906];
  assign o[6449] = i[9905];
  assign o[6448] = i[9904];
  assign o[6447] = i[9903];
  assign o[6446] = i[9902];
  assign o[6445] = i[9901];
  assign o[6444] = i[9900];
  assign o[6443] = i[9899];
  assign o[6442] = i[9898];
  assign o[6441] = i[9897];
  assign o[6440] = i[9896];
  assign o[6439] = i[9895];
  assign o[6438] = i[9894];
  assign o[6437] = i[9893];
  assign o[6436] = i[9892];
  assign o[6435] = i[9891];
  assign o[6434] = i[9890];
  assign o[6433] = i[9889];
  assign o[6432] = i[9888];
  assign o[6431] = i[9887];
  assign o[6430] = i[9886];
  assign o[6429] = i[9885];
  assign o[6428] = i[9884];
  assign o[6427] = i[9883];
  assign o[6426] = i[9882];
  assign o[6425] = i[9881];
  assign o[6424] = i[9880];
  assign o[6423] = i[9879];
  assign o[6422] = i[9878];
  assign o[6421] = i[9877];
  assign o[6420] = i[9876];
  assign o[6419] = i[9875];
  assign o[6418] = i[9874];
  assign o[6417] = i[9873];
  assign o[6416] = i[9872];
  assign o[6415] = i[9871];
  assign o[6414] = i[9870];
  assign o[6413] = i[9869];
  assign o[6412] = i[9868];
  assign o[6411] = i[9867];
  assign o[6410] = i[9866];
  assign o[6409] = i[9865];
  assign o[6408] = i[9864];
  assign o[6407] = i[9863];
  assign o[6406] = i[9862];
  assign o[6405] = i[9861];
  assign o[6404] = i[9860];
  assign o[6403] = i[9859];
  assign o[6402] = i[9858];
  assign o[6401] = i[9857];
  assign o[6400] = i[9856];
  assign o[6399] = i[10111];
  assign o[6398] = i[10110];
  assign o[6397] = i[10109];
  assign o[6396] = i[10108];
  assign o[6395] = i[10107];
  assign o[6394] = i[10106];
  assign o[6393] = i[10105];
  assign o[6392] = i[10104];
  assign o[6391] = i[10103];
  assign o[6390] = i[10102];
  assign o[6389] = i[10101];
  assign o[6388] = i[10100];
  assign o[6387] = i[10099];
  assign o[6386] = i[10098];
  assign o[6385] = i[10097];
  assign o[6384] = i[10096];
  assign o[6383] = i[10095];
  assign o[6382] = i[10094];
  assign o[6381] = i[10093];
  assign o[6380] = i[10092];
  assign o[6379] = i[10091];
  assign o[6378] = i[10090];
  assign o[6377] = i[10089];
  assign o[6376] = i[10088];
  assign o[6375] = i[10087];
  assign o[6374] = i[10086];
  assign o[6373] = i[10085];
  assign o[6372] = i[10084];
  assign o[6371] = i[10083];
  assign o[6370] = i[10082];
  assign o[6369] = i[10081];
  assign o[6368] = i[10080];
  assign o[6367] = i[10079];
  assign o[6366] = i[10078];
  assign o[6365] = i[10077];
  assign o[6364] = i[10076];
  assign o[6363] = i[10075];
  assign o[6362] = i[10074];
  assign o[6361] = i[10073];
  assign o[6360] = i[10072];
  assign o[6359] = i[10071];
  assign o[6358] = i[10070];
  assign o[6357] = i[10069];
  assign o[6356] = i[10068];
  assign o[6355] = i[10067];
  assign o[6354] = i[10066];
  assign o[6353] = i[10065];
  assign o[6352] = i[10064];
  assign o[6351] = i[10063];
  assign o[6350] = i[10062];
  assign o[6349] = i[10061];
  assign o[6348] = i[10060];
  assign o[6347] = i[10059];
  assign o[6346] = i[10058];
  assign o[6345] = i[10057];
  assign o[6344] = i[10056];
  assign o[6343] = i[10055];
  assign o[6342] = i[10054];
  assign o[6341] = i[10053];
  assign o[6340] = i[10052];
  assign o[6339] = i[10051];
  assign o[6338] = i[10050];
  assign o[6337] = i[10049];
  assign o[6336] = i[10048];
  assign o[6335] = i[10047];
  assign o[6334] = i[10046];
  assign o[6333] = i[10045];
  assign o[6332] = i[10044];
  assign o[6331] = i[10043];
  assign o[6330] = i[10042];
  assign o[6329] = i[10041];
  assign o[6328] = i[10040];
  assign o[6327] = i[10039];
  assign o[6326] = i[10038];
  assign o[6325] = i[10037];
  assign o[6324] = i[10036];
  assign o[6323] = i[10035];
  assign o[6322] = i[10034];
  assign o[6321] = i[10033];
  assign o[6320] = i[10032];
  assign o[6319] = i[10031];
  assign o[6318] = i[10030];
  assign o[6317] = i[10029];
  assign o[6316] = i[10028];
  assign o[6315] = i[10027];
  assign o[6314] = i[10026];
  assign o[6313] = i[10025];
  assign o[6312] = i[10024];
  assign o[6311] = i[10023];
  assign o[6310] = i[10022];
  assign o[6309] = i[10021];
  assign o[6308] = i[10020];
  assign o[6307] = i[10019];
  assign o[6306] = i[10018];
  assign o[6305] = i[10017];
  assign o[6304] = i[10016];
  assign o[6303] = i[10015];
  assign o[6302] = i[10014];
  assign o[6301] = i[10013];
  assign o[6300] = i[10012];
  assign o[6299] = i[10011];
  assign o[6298] = i[10010];
  assign o[6297] = i[10009];
  assign o[6296] = i[10008];
  assign o[6295] = i[10007];
  assign o[6294] = i[10006];
  assign o[6293] = i[10005];
  assign o[6292] = i[10004];
  assign o[6291] = i[10003];
  assign o[6290] = i[10002];
  assign o[6289] = i[10001];
  assign o[6288] = i[10000];
  assign o[6287] = i[9999];
  assign o[6286] = i[9998];
  assign o[6285] = i[9997];
  assign o[6284] = i[9996];
  assign o[6283] = i[9995];
  assign o[6282] = i[9994];
  assign o[6281] = i[9993];
  assign o[6280] = i[9992];
  assign o[6279] = i[9991];
  assign o[6278] = i[9990];
  assign o[6277] = i[9989];
  assign o[6276] = i[9988];
  assign o[6275] = i[9987];
  assign o[6274] = i[9986];
  assign o[6273] = i[9985];
  assign o[6272] = i[9984];
  assign o[6271] = i[10239];
  assign o[6270] = i[10238];
  assign o[6269] = i[10237];
  assign o[6268] = i[10236];
  assign o[6267] = i[10235];
  assign o[6266] = i[10234];
  assign o[6265] = i[10233];
  assign o[6264] = i[10232];
  assign o[6263] = i[10231];
  assign o[6262] = i[10230];
  assign o[6261] = i[10229];
  assign o[6260] = i[10228];
  assign o[6259] = i[10227];
  assign o[6258] = i[10226];
  assign o[6257] = i[10225];
  assign o[6256] = i[10224];
  assign o[6255] = i[10223];
  assign o[6254] = i[10222];
  assign o[6253] = i[10221];
  assign o[6252] = i[10220];
  assign o[6251] = i[10219];
  assign o[6250] = i[10218];
  assign o[6249] = i[10217];
  assign o[6248] = i[10216];
  assign o[6247] = i[10215];
  assign o[6246] = i[10214];
  assign o[6245] = i[10213];
  assign o[6244] = i[10212];
  assign o[6243] = i[10211];
  assign o[6242] = i[10210];
  assign o[6241] = i[10209];
  assign o[6240] = i[10208];
  assign o[6239] = i[10207];
  assign o[6238] = i[10206];
  assign o[6237] = i[10205];
  assign o[6236] = i[10204];
  assign o[6235] = i[10203];
  assign o[6234] = i[10202];
  assign o[6233] = i[10201];
  assign o[6232] = i[10200];
  assign o[6231] = i[10199];
  assign o[6230] = i[10198];
  assign o[6229] = i[10197];
  assign o[6228] = i[10196];
  assign o[6227] = i[10195];
  assign o[6226] = i[10194];
  assign o[6225] = i[10193];
  assign o[6224] = i[10192];
  assign o[6223] = i[10191];
  assign o[6222] = i[10190];
  assign o[6221] = i[10189];
  assign o[6220] = i[10188];
  assign o[6219] = i[10187];
  assign o[6218] = i[10186];
  assign o[6217] = i[10185];
  assign o[6216] = i[10184];
  assign o[6215] = i[10183];
  assign o[6214] = i[10182];
  assign o[6213] = i[10181];
  assign o[6212] = i[10180];
  assign o[6211] = i[10179];
  assign o[6210] = i[10178];
  assign o[6209] = i[10177];
  assign o[6208] = i[10176];
  assign o[6207] = i[10175];
  assign o[6206] = i[10174];
  assign o[6205] = i[10173];
  assign o[6204] = i[10172];
  assign o[6203] = i[10171];
  assign o[6202] = i[10170];
  assign o[6201] = i[10169];
  assign o[6200] = i[10168];
  assign o[6199] = i[10167];
  assign o[6198] = i[10166];
  assign o[6197] = i[10165];
  assign o[6196] = i[10164];
  assign o[6195] = i[10163];
  assign o[6194] = i[10162];
  assign o[6193] = i[10161];
  assign o[6192] = i[10160];
  assign o[6191] = i[10159];
  assign o[6190] = i[10158];
  assign o[6189] = i[10157];
  assign o[6188] = i[10156];
  assign o[6187] = i[10155];
  assign o[6186] = i[10154];
  assign o[6185] = i[10153];
  assign o[6184] = i[10152];
  assign o[6183] = i[10151];
  assign o[6182] = i[10150];
  assign o[6181] = i[10149];
  assign o[6180] = i[10148];
  assign o[6179] = i[10147];
  assign o[6178] = i[10146];
  assign o[6177] = i[10145];
  assign o[6176] = i[10144];
  assign o[6175] = i[10143];
  assign o[6174] = i[10142];
  assign o[6173] = i[10141];
  assign o[6172] = i[10140];
  assign o[6171] = i[10139];
  assign o[6170] = i[10138];
  assign o[6169] = i[10137];
  assign o[6168] = i[10136];
  assign o[6167] = i[10135];
  assign o[6166] = i[10134];
  assign o[6165] = i[10133];
  assign o[6164] = i[10132];
  assign o[6163] = i[10131];
  assign o[6162] = i[10130];
  assign o[6161] = i[10129];
  assign o[6160] = i[10128];
  assign o[6159] = i[10127];
  assign o[6158] = i[10126];
  assign o[6157] = i[10125];
  assign o[6156] = i[10124];
  assign o[6155] = i[10123];
  assign o[6154] = i[10122];
  assign o[6153] = i[10121];
  assign o[6152] = i[10120];
  assign o[6151] = i[10119];
  assign o[6150] = i[10118];
  assign o[6149] = i[10117];
  assign o[6148] = i[10116];
  assign o[6147] = i[10115];
  assign o[6146] = i[10114];
  assign o[6145] = i[10113];
  assign o[6144] = i[10112];
  assign o[6143] = i[10367];
  assign o[6142] = i[10366];
  assign o[6141] = i[10365];
  assign o[6140] = i[10364];
  assign o[6139] = i[10363];
  assign o[6138] = i[10362];
  assign o[6137] = i[10361];
  assign o[6136] = i[10360];
  assign o[6135] = i[10359];
  assign o[6134] = i[10358];
  assign o[6133] = i[10357];
  assign o[6132] = i[10356];
  assign o[6131] = i[10355];
  assign o[6130] = i[10354];
  assign o[6129] = i[10353];
  assign o[6128] = i[10352];
  assign o[6127] = i[10351];
  assign o[6126] = i[10350];
  assign o[6125] = i[10349];
  assign o[6124] = i[10348];
  assign o[6123] = i[10347];
  assign o[6122] = i[10346];
  assign o[6121] = i[10345];
  assign o[6120] = i[10344];
  assign o[6119] = i[10343];
  assign o[6118] = i[10342];
  assign o[6117] = i[10341];
  assign o[6116] = i[10340];
  assign o[6115] = i[10339];
  assign o[6114] = i[10338];
  assign o[6113] = i[10337];
  assign o[6112] = i[10336];
  assign o[6111] = i[10335];
  assign o[6110] = i[10334];
  assign o[6109] = i[10333];
  assign o[6108] = i[10332];
  assign o[6107] = i[10331];
  assign o[6106] = i[10330];
  assign o[6105] = i[10329];
  assign o[6104] = i[10328];
  assign o[6103] = i[10327];
  assign o[6102] = i[10326];
  assign o[6101] = i[10325];
  assign o[6100] = i[10324];
  assign o[6099] = i[10323];
  assign o[6098] = i[10322];
  assign o[6097] = i[10321];
  assign o[6096] = i[10320];
  assign o[6095] = i[10319];
  assign o[6094] = i[10318];
  assign o[6093] = i[10317];
  assign o[6092] = i[10316];
  assign o[6091] = i[10315];
  assign o[6090] = i[10314];
  assign o[6089] = i[10313];
  assign o[6088] = i[10312];
  assign o[6087] = i[10311];
  assign o[6086] = i[10310];
  assign o[6085] = i[10309];
  assign o[6084] = i[10308];
  assign o[6083] = i[10307];
  assign o[6082] = i[10306];
  assign o[6081] = i[10305];
  assign o[6080] = i[10304];
  assign o[6079] = i[10303];
  assign o[6078] = i[10302];
  assign o[6077] = i[10301];
  assign o[6076] = i[10300];
  assign o[6075] = i[10299];
  assign o[6074] = i[10298];
  assign o[6073] = i[10297];
  assign o[6072] = i[10296];
  assign o[6071] = i[10295];
  assign o[6070] = i[10294];
  assign o[6069] = i[10293];
  assign o[6068] = i[10292];
  assign o[6067] = i[10291];
  assign o[6066] = i[10290];
  assign o[6065] = i[10289];
  assign o[6064] = i[10288];
  assign o[6063] = i[10287];
  assign o[6062] = i[10286];
  assign o[6061] = i[10285];
  assign o[6060] = i[10284];
  assign o[6059] = i[10283];
  assign o[6058] = i[10282];
  assign o[6057] = i[10281];
  assign o[6056] = i[10280];
  assign o[6055] = i[10279];
  assign o[6054] = i[10278];
  assign o[6053] = i[10277];
  assign o[6052] = i[10276];
  assign o[6051] = i[10275];
  assign o[6050] = i[10274];
  assign o[6049] = i[10273];
  assign o[6048] = i[10272];
  assign o[6047] = i[10271];
  assign o[6046] = i[10270];
  assign o[6045] = i[10269];
  assign o[6044] = i[10268];
  assign o[6043] = i[10267];
  assign o[6042] = i[10266];
  assign o[6041] = i[10265];
  assign o[6040] = i[10264];
  assign o[6039] = i[10263];
  assign o[6038] = i[10262];
  assign o[6037] = i[10261];
  assign o[6036] = i[10260];
  assign o[6035] = i[10259];
  assign o[6034] = i[10258];
  assign o[6033] = i[10257];
  assign o[6032] = i[10256];
  assign o[6031] = i[10255];
  assign o[6030] = i[10254];
  assign o[6029] = i[10253];
  assign o[6028] = i[10252];
  assign o[6027] = i[10251];
  assign o[6026] = i[10250];
  assign o[6025] = i[10249];
  assign o[6024] = i[10248];
  assign o[6023] = i[10247];
  assign o[6022] = i[10246];
  assign o[6021] = i[10245];
  assign o[6020] = i[10244];
  assign o[6019] = i[10243];
  assign o[6018] = i[10242];
  assign o[6017] = i[10241];
  assign o[6016] = i[10240];
  assign o[6015] = i[10495];
  assign o[6014] = i[10494];
  assign o[6013] = i[10493];
  assign o[6012] = i[10492];
  assign o[6011] = i[10491];
  assign o[6010] = i[10490];
  assign o[6009] = i[10489];
  assign o[6008] = i[10488];
  assign o[6007] = i[10487];
  assign o[6006] = i[10486];
  assign o[6005] = i[10485];
  assign o[6004] = i[10484];
  assign o[6003] = i[10483];
  assign o[6002] = i[10482];
  assign o[6001] = i[10481];
  assign o[6000] = i[10480];
  assign o[5999] = i[10479];
  assign o[5998] = i[10478];
  assign o[5997] = i[10477];
  assign o[5996] = i[10476];
  assign o[5995] = i[10475];
  assign o[5994] = i[10474];
  assign o[5993] = i[10473];
  assign o[5992] = i[10472];
  assign o[5991] = i[10471];
  assign o[5990] = i[10470];
  assign o[5989] = i[10469];
  assign o[5988] = i[10468];
  assign o[5987] = i[10467];
  assign o[5986] = i[10466];
  assign o[5985] = i[10465];
  assign o[5984] = i[10464];
  assign o[5983] = i[10463];
  assign o[5982] = i[10462];
  assign o[5981] = i[10461];
  assign o[5980] = i[10460];
  assign o[5979] = i[10459];
  assign o[5978] = i[10458];
  assign o[5977] = i[10457];
  assign o[5976] = i[10456];
  assign o[5975] = i[10455];
  assign o[5974] = i[10454];
  assign o[5973] = i[10453];
  assign o[5972] = i[10452];
  assign o[5971] = i[10451];
  assign o[5970] = i[10450];
  assign o[5969] = i[10449];
  assign o[5968] = i[10448];
  assign o[5967] = i[10447];
  assign o[5966] = i[10446];
  assign o[5965] = i[10445];
  assign o[5964] = i[10444];
  assign o[5963] = i[10443];
  assign o[5962] = i[10442];
  assign o[5961] = i[10441];
  assign o[5960] = i[10440];
  assign o[5959] = i[10439];
  assign o[5958] = i[10438];
  assign o[5957] = i[10437];
  assign o[5956] = i[10436];
  assign o[5955] = i[10435];
  assign o[5954] = i[10434];
  assign o[5953] = i[10433];
  assign o[5952] = i[10432];
  assign o[5951] = i[10431];
  assign o[5950] = i[10430];
  assign o[5949] = i[10429];
  assign o[5948] = i[10428];
  assign o[5947] = i[10427];
  assign o[5946] = i[10426];
  assign o[5945] = i[10425];
  assign o[5944] = i[10424];
  assign o[5943] = i[10423];
  assign o[5942] = i[10422];
  assign o[5941] = i[10421];
  assign o[5940] = i[10420];
  assign o[5939] = i[10419];
  assign o[5938] = i[10418];
  assign o[5937] = i[10417];
  assign o[5936] = i[10416];
  assign o[5935] = i[10415];
  assign o[5934] = i[10414];
  assign o[5933] = i[10413];
  assign o[5932] = i[10412];
  assign o[5931] = i[10411];
  assign o[5930] = i[10410];
  assign o[5929] = i[10409];
  assign o[5928] = i[10408];
  assign o[5927] = i[10407];
  assign o[5926] = i[10406];
  assign o[5925] = i[10405];
  assign o[5924] = i[10404];
  assign o[5923] = i[10403];
  assign o[5922] = i[10402];
  assign o[5921] = i[10401];
  assign o[5920] = i[10400];
  assign o[5919] = i[10399];
  assign o[5918] = i[10398];
  assign o[5917] = i[10397];
  assign o[5916] = i[10396];
  assign o[5915] = i[10395];
  assign o[5914] = i[10394];
  assign o[5913] = i[10393];
  assign o[5912] = i[10392];
  assign o[5911] = i[10391];
  assign o[5910] = i[10390];
  assign o[5909] = i[10389];
  assign o[5908] = i[10388];
  assign o[5907] = i[10387];
  assign o[5906] = i[10386];
  assign o[5905] = i[10385];
  assign o[5904] = i[10384];
  assign o[5903] = i[10383];
  assign o[5902] = i[10382];
  assign o[5901] = i[10381];
  assign o[5900] = i[10380];
  assign o[5899] = i[10379];
  assign o[5898] = i[10378];
  assign o[5897] = i[10377];
  assign o[5896] = i[10376];
  assign o[5895] = i[10375];
  assign o[5894] = i[10374];
  assign o[5893] = i[10373];
  assign o[5892] = i[10372];
  assign o[5891] = i[10371];
  assign o[5890] = i[10370];
  assign o[5889] = i[10369];
  assign o[5888] = i[10368];
  assign o[5887] = i[10623];
  assign o[5886] = i[10622];
  assign o[5885] = i[10621];
  assign o[5884] = i[10620];
  assign o[5883] = i[10619];
  assign o[5882] = i[10618];
  assign o[5881] = i[10617];
  assign o[5880] = i[10616];
  assign o[5879] = i[10615];
  assign o[5878] = i[10614];
  assign o[5877] = i[10613];
  assign o[5876] = i[10612];
  assign o[5875] = i[10611];
  assign o[5874] = i[10610];
  assign o[5873] = i[10609];
  assign o[5872] = i[10608];
  assign o[5871] = i[10607];
  assign o[5870] = i[10606];
  assign o[5869] = i[10605];
  assign o[5868] = i[10604];
  assign o[5867] = i[10603];
  assign o[5866] = i[10602];
  assign o[5865] = i[10601];
  assign o[5864] = i[10600];
  assign o[5863] = i[10599];
  assign o[5862] = i[10598];
  assign o[5861] = i[10597];
  assign o[5860] = i[10596];
  assign o[5859] = i[10595];
  assign o[5858] = i[10594];
  assign o[5857] = i[10593];
  assign o[5856] = i[10592];
  assign o[5855] = i[10591];
  assign o[5854] = i[10590];
  assign o[5853] = i[10589];
  assign o[5852] = i[10588];
  assign o[5851] = i[10587];
  assign o[5850] = i[10586];
  assign o[5849] = i[10585];
  assign o[5848] = i[10584];
  assign o[5847] = i[10583];
  assign o[5846] = i[10582];
  assign o[5845] = i[10581];
  assign o[5844] = i[10580];
  assign o[5843] = i[10579];
  assign o[5842] = i[10578];
  assign o[5841] = i[10577];
  assign o[5840] = i[10576];
  assign o[5839] = i[10575];
  assign o[5838] = i[10574];
  assign o[5837] = i[10573];
  assign o[5836] = i[10572];
  assign o[5835] = i[10571];
  assign o[5834] = i[10570];
  assign o[5833] = i[10569];
  assign o[5832] = i[10568];
  assign o[5831] = i[10567];
  assign o[5830] = i[10566];
  assign o[5829] = i[10565];
  assign o[5828] = i[10564];
  assign o[5827] = i[10563];
  assign o[5826] = i[10562];
  assign o[5825] = i[10561];
  assign o[5824] = i[10560];
  assign o[5823] = i[10559];
  assign o[5822] = i[10558];
  assign o[5821] = i[10557];
  assign o[5820] = i[10556];
  assign o[5819] = i[10555];
  assign o[5818] = i[10554];
  assign o[5817] = i[10553];
  assign o[5816] = i[10552];
  assign o[5815] = i[10551];
  assign o[5814] = i[10550];
  assign o[5813] = i[10549];
  assign o[5812] = i[10548];
  assign o[5811] = i[10547];
  assign o[5810] = i[10546];
  assign o[5809] = i[10545];
  assign o[5808] = i[10544];
  assign o[5807] = i[10543];
  assign o[5806] = i[10542];
  assign o[5805] = i[10541];
  assign o[5804] = i[10540];
  assign o[5803] = i[10539];
  assign o[5802] = i[10538];
  assign o[5801] = i[10537];
  assign o[5800] = i[10536];
  assign o[5799] = i[10535];
  assign o[5798] = i[10534];
  assign o[5797] = i[10533];
  assign o[5796] = i[10532];
  assign o[5795] = i[10531];
  assign o[5794] = i[10530];
  assign o[5793] = i[10529];
  assign o[5792] = i[10528];
  assign o[5791] = i[10527];
  assign o[5790] = i[10526];
  assign o[5789] = i[10525];
  assign o[5788] = i[10524];
  assign o[5787] = i[10523];
  assign o[5786] = i[10522];
  assign o[5785] = i[10521];
  assign o[5784] = i[10520];
  assign o[5783] = i[10519];
  assign o[5782] = i[10518];
  assign o[5781] = i[10517];
  assign o[5780] = i[10516];
  assign o[5779] = i[10515];
  assign o[5778] = i[10514];
  assign o[5777] = i[10513];
  assign o[5776] = i[10512];
  assign o[5775] = i[10511];
  assign o[5774] = i[10510];
  assign o[5773] = i[10509];
  assign o[5772] = i[10508];
  assign o[5771] = i[10507];
  assign o[5770] = i[10506];
  assign o[5769] = i[10505];
  assign o[5768] = i[10504];
  assign o[5767] = i[10503];
  assign o[5766] = i[10502];
  assign o[5765] = i[10501];
  assign o[5764] = i[10500];
  assign o[5763] = i[10499];
  assign o[5762] = i[10498];
  assign o[5761] = i[10497];
  assign o[5760] = i[10496];
  assign o[5759] = i[10751];
  assign o[5758] = i[10750];
  assign o[5757] = i[10749];
  assign o[5756] = i[10748];
  assign o[5755] = i[10747];
  assign o[5754] = i[10746];
  assign o[5753] = i[10745];
  assign o[5752] = i[10744];
  assign o[5751] = i[10743];
  assign o[5750] = i[10742];
  assign o[5749] = i[10741];
  assign o[5748] = i[10740];
  assign o[5747] = i[10739];
  assign o[5746] = i[10738];
  assign o[5745] = i[10737];
  assign o[5744] = i[10736];
  assign o[5743] = i[10735];
  assign o[5742] = i[10734];
  assign o[5741] = i[10733];
  assign o[5740] = i[10732];
  assign o[5739] = i[10731];
  assign o[5738] = i[10730];
  assign o[5737] = i[10729];
  assign o[5736] = i[10728];
  assign o[5735] = i[10727];
  assign o[5734] = i[10726];
  assign o[5733] = i[10725];
  assign o[5732] = i[10724];
  assign o[5731] = i[10723];
  assign o[5730] = i[10722];
  assign o[5729] = i[10721];
  assign o[5728] = i[10720];
  assign o[5727] = i[10719];
  assign o[5726] = i[10718];
  assign o[5725] = i[10717];
  assign o[5724] = i[10716];
  assign o[5723] = i[10715];
  assign o[5722] = i[10714];
  assign o[5721] = i[10713];
  assign o[5720] = i[10712];
  assign o[5719] = i[10711];
  assign o[5718] = i[10710];
  assign o[5717] = i[10709];
  assign o[5716] = i[10708];
  assign o[5715] = i[10707];
  assign o[5714] = i[10706];
  assign o[5713] = i[10705];
  assign o[5712] = i[10704];
  assign o[5711] = i[10703];
  assign o[5710] = i[10702];
  assign o[5709] = i[10701];
  assign o[5708] = i[10700];
  assign o[5707] = i[10699];
  assign o[5706] = i[10698];
  assign o[5705] = i[10697];
  assign o[5704] = i[10696];
  assign o[5703] = i[10695];
  assign o[5702] = i[10694];
  assign o[5701] = i[10693];
  assign o[5700] = i[10692];
  assign o[5699] = i[10691];
  assign o[5698] = i[10690];
  assign o[5697] = i[10689];
  assign o[5696] = i[10688];
  assign o[5695] = i[10687];
  assign o[5694] = i[10686];
  assign o[5693] = i[10685];
  assign o[5692] = i[10684];
  assign o[5691] = i[10683];
  assign o[5690] = i[10682];
  assign o[5689] = i[10681];
  assign o[5688] = i[10680];
  assign o[5687] = i[10679];
  assign o[5686] = i[10678];
  assign o[5685] = i[10677];
  assign o[5684] = i[10676];
  assign o[5683] = i[10675];
  assign o[5682] = i[10674];
  assign o[5681] = i[10673];
  assign o[5680] = i[10672];
  assign o[5679] = i[10671];
  assign o[5678] = i[10670];
  assign o[5677] = i[10669];
  assign o[5676] = i[10668];
  assign o[5675] = i[10667];
  assign o[5674] = i[10666];
  assign o[5673] = i[10665];
  assign o[5672] = i[10664];
  assign o[5671] = i[10663];
  assign o[5670] = i[10662];
  assign o[5669] = i[10661];
  assign o[5668] = i[10660];
  assign o[5667] = i[10659];
  assign o[5666] = i[10658];
  assign o[5665] = i[10657];
  assign o[5664] = i[10656];
  assign o[5663] = i[10655];
  assign o[5662] = i[10654];
  assign o[5661] = i[10653];
  assign o[5660] = i[10652];
  assign o[5659] = i[10651];
  assign o[5658] = i[10650];
  assign o[5657] = i[10649];
  assign o[5656] = i[10648];
  assign o[5655] = i[10647];
  assign o[5654] = i[10646];
  assign o[5653] = i[10645];
  assign o[5652] = i[10644];
  assign o[5651] = i[10643];
  assign o[5650] = i[10642];
  assign o[5649] = i[10641];
  assign o[5648] = i[10640];
  assign o[5647] = i[10639];
  assign o[5646] = i[10638];
  assign o[5645] = i[10637];
  assign o[5644] = i[10636];
  assign o[5643] = i[10635];
  assign o[5642] = i[10634];
  assign o[5641] = i[10633];
  assign o[5640] = i[10632];
  assign o[5639] = i[10631];
  assign o[5638] = i[10630];
  assign o[5637] = i[10629];
  assign o[5636] = i[10628];
  assign o[5635] = i[10627];
  assign o[5634] = i[10626];
  assign o[5633] = i[10625];
  assign o[5632] = i[10624];
  assign o[5631] = i[10879];
  assign o[5630] = i[10878];
  assign o[5629] = i[10877];
  assign o[5628] = i[10876];
  assign o[5627] = i[10875];
  assign o[5626] = i[10874];
  assign o[5625] = i[10873];
  assign o[5624] = i[10872];
  assign o[5623] = i[10871];
  assign o[5622] = i[10870];
  assign o[5621] = i[10869];
  assign o[5620] = i[10868];
  assign o[5619] = i[10867];
  assign o[5618] = i[10866];
  assign o[5617] = i[10865];
  assign o[5616] = i[10864];
  assign o[5615] = i[10863];
  assign o[5614] = i[10862];
  assign o[5613] = i[10861];
  assign o[5612] = i[10860];
  assign o[5611] = i[10859];
  assign o[5610] = i[10858];
  assign o[5609] = i[10857];
  assign o[5608] = i[10856];
  assign o[5607] = i[10855];
  assign o[5606] = i[10854];
  assign o[5605] = i[10853];
  assign o[5604] = i[10852];
  assign o[5603] = i[10851];
  assign o[5602] = i[10850];
  assign o[5601] = i[10849];
  assign o[5600] = i[10848];
  assign o[5599] = i[10847];
  assign o[5598] = i[10846];
  assign o[5597] = i[10845];
  assign o[5596] = i[10844];
  assign o[5595] = i[10843];
  assign o[5594] = i[10842];
  assign o[5593] = i[10841];
  assign o[5592] = i[10840];
  assign o[5591] = i[10839];
  assign o[5590] = i[10838];
  assign o[5589] = i[10837];
  assign o[5588] = i[10836];
  assign o[5587] = i[10835];
  assign o[5586] = i[10834];
  assign o[5585] = i[10833];
  assign o[5584] = i[10832];
  assign o[5583] = i[10831];
  assign o[5582] = i[10830];
  assign o[5581] = i[10829];
  assign o[5580] = i[10828];
  assign o[5579] = i[10827];
  assign o[5578] = i[10826];
  assign o[5577] = i[10825];
  assign o[5576] = i[10824];
  assign o[5575] = i[10823];
  assign o[5574] = i[10822];
  assign o[5573] = i[10821];
  assign o[5572] = i[10820];
  assign o[5571] = i[10819];
  assign o[5570] = i[10818];
  assign o[5569] = i[10817];
  assign o[5568] = i[10816];
  assign o[5567] = i[10815];
  assign o[5566] = i[10814];
  assign o[5565] = i[10813];
  assign o[5564] = i[10812];
  assign o[5563] = i[10811];
  assign o[5562] = i[10810];
  assign o[5561] = i[10809];
  assign o[5560] = i[10808];
  assign o[5559] = i[10807];
  assign o[5558] = i[10806];
  assign o[5557] = i[10805];
  assign o[5556] = i[10804];
  assign o[5555] = i[10803];
  assign o[5554] = i[10802];
  assign o[5553] = i[10801];
  assign o[5552] = i[10800];
  assign o[5551] = i[10799];
  assign o[5550] = i[10798];
  assign o[5549] = i[10797];
  assign o[5548] = i[10796];
  assign o[5547] = i[10795];
  assign o[5546] = i[10794];
  assign o[5545] = i[10793];
  assign o[5544] = i[10792];
  assign o[5543] = i[10791];
  assign o[5542] = i[10790];
  assign o[5541] = i[10789];
  assign o[5540] = i[10788];
  assign o[5539] = i[10787];
  assign o[5538] = i[10786];
  assign o[5537] = i[10785];
  assign o[5536] = i[10784];
  assign o[5535] = i[10783];
  assign o[5534] = i[10782];
  assign o[5533] = i[10781];
  assign o[5532] = i[10780];
  assign o[5531] = i[10779];
  assign o[5530] = i[10778];
  assign o[5529] = i[10777];
  assign o[5528] = i[10776];
  assign o[5527] = i[10775];
  assign o[5526] = i[10774];
  assign o[5525] = i[10773];
  assign o[5524] = i[10772];
  assign o[5523] = i[10771];
  assign o[5522] = i[10770];
  assign o[5521] = i[10769];
  assign o[5520] = i[10768];
  assign o[5519] = i[10767];
  assign o[5518] = i[10766];
  assign o[5517] = i[10765];
  assign o[5516] = i[10764];
  assign o[5515] = i[10763];
  assign o[5514] = i[10762];
  assign o[5513] = i[10761];
  assign o[5512] = i[10760];
  assign o[5511] = i[10759];
  assign o[5510] = i[10758];
  assign o[5509] = i[10757];
  assign o[5508] = i[10756];
  assign o[5507] = i[10755];
  assign o[5506] = i[10754];
  assign o[5505] = i[10753];
  assign o[5504] = i[10752];
  assign o[5503] = i[11007];
  assign o[5502] = i[11006];
  assign o[5501] = i[11005];
  assign o[5500] = i[11004];
  assign o[5499] = i[11003];
  assign o[5498] = i[11002];
  assign o[5497] = i[11001];
  assign o[5496] = i[11000];
  assign o[5495] = i[10999];
  assign o[5494] = i[10998];
  assign o[5493] = i[10997];
  assign o[5492] = i[10996];
  assign o[5491] = i[10995];
  assign o[5490] = i[10994];
  assign o[5489] = i[10993];
  assign o[5488] = i[10992];
  assign o[5487] = i[10991];
  assign o[5486] = i[10990];
  assign o[5485] = i[10989];
  assign o[5484] = i[10988];
  assign o[5483] = i[10987];
  assign o[5482] = i[10986];
  assign o[5481] = i[10985];
  assign o[5480] = i[10984];
  assign o[5479] = i[10983];
  assign o[5478] = i[10982];
  assign o[5477] = i[10981];
  assign o[5476] = i[10980];
  assign o[5475] = i[10979];
  assign o[5474] = i[10978];
  assign o[5473] = i[10977];
  assign o[5472] = i[10976];
  assign o[5471] = i[10975];
  assign o[5470] = i[10974];
  assign o[5469] = i[10973];
  assign o[5468] = i[10972];
  assign o[5467] = i[10971];
  assign o[5466] = i[10970];
  assign o[5465] = i[10969];
  assign o[5464] = i[10968];
  assign o[5463] = i[10967];
  assign o[5462] = i[10966];
  assign o[5461] = i[10965];
  assign o[5460] = i[10964];
  assign o[5459] = i[10963];
  assign o[5458] = i[10962];
  assign o[5457] = i[10961];
  assign o[5456] = i[10960];
  assign o[5455] = i[10959];
  assign o[5454] = i[10958];
  assign o[5453] = i[10957];
  assign o[5452] = i[10956];
  assign o[5451] = i[10955];
  assign o[5450] = i[10954];
  assign o[5449] = i[10953];
  assign o[5448] = i[10952];
  assign o[5447] = i[10951];
  assign o[5446] = i[10950];
  assign o[5445] = i[10949];
  assign o[5444] = i[10948];
  assign o[5443] = i[10947];
  assign o[5442] = i[10946];
  assign o[5441] = i[10945];
  assign o[5440] = i[10944];
  assign o[5439] = i[10943];
  assign o[5438] = i[10942];
  assign o[5437] = i[10941];
  assign o[5436] = i[10940];
  assign o[5435] = i[10939];
  assign o[5434] = i[10938];
  assign o[5433] = i[10937];
  assign o[5432] = i[10936];
  assign o[5431] = i[10935];
  assign o[5430] = i[10934];
  assign o[5429] = i[10933];
  assign o[5428] = i[10932];
  assign o[5427] = i[10931];
  assign o[5426] = i[10930];
  assign o[5425] = i[10929];
  assign o[5424] = i[10928];
  assign o[5423] = i[10927];
  assign o[5422] = i[10926];
  assign o[5421] = i[10925];
  assign o[5420] = i[10924];
  assign o[5419] = i[10923];
  assign o[5418] = i[10922];
  assign o[5417] = i[10921];
  assign o[5416] = i[10920];
  assign o[5415] = i[10919];
  assign o[5414] = i[10918];
  assign o[5413] = i[10917];
  assign o[5412] = i[10916];
  assign o[5411] = i[10915];
  assign o[5410] = i[10914];
  assign o[5409] = i[10913];
  assign o[5408] = i[10912];
  assign o[5407] = i[10911];
  assign o[5406] = i[10910];
  assign o[5405] = i[10909];
  assign o[5404] = i[10908];
  assign o[5403] = i[10907];
  assign o[5402] = i[10906];
  assign o[5401] = i[10905];
  assign o[5400] = i[10904];
  assign o[5399] = i[10903];
  assign o[5398] = i[10902];
  assign o[5397] = i[10901];
  assign o[5396] = i[10900];
  assign o[5395] = i[10899];
  assign o[5394] = i[10898];
  assign o[5393] = i[10897];
  assign o[5392] = i[10896];
  assign o[5391] = i[10895];
  assign o[5390] = i[10894];
  assign o[5389] = i[10893];
  assign o[5388] = i[10892];
  assign o[5387] = i[10891];
  assign o[5386] = i[10890];
  assign o[5385] = i[10889];
  assign o[5384] = i[10888];
  assign o[5383] = i[10887];
  assign o[5382] = i[10886];
  assign o[5381] = i[10885];
  assign o[5380] = i[10884];
  assign o[5379] = i[10883];
  assign o[5378] = i[10882];
  assign o[5377] = i[10881];
  assign o[5376] = i[10880];
  assign o[5375] = i[11135];
  assign o[5374] = i[11134];
  assign o[5373] = i[11133];
  assign o[5372] = i[11132];
  assign o[5371] = i[11131];
  assign o[5370] = i[11130];
  assign o[5369] = i[11129];
  assign o[5368] = i[11128];
  assign o[5367] = i[11127];
  assign o[5366] = i[11126];
  assign o[5365] = i[11125];
  assign o[5364] = i[11124];
  assign o[5363] = i[11123];
  assign o[5362] = i[11122];
  assign o[5361] = i[11121];
  assign o[5360] = i[11120];
  assign o[5359] = i[11119];
  assign o[5358] = i[11118];
  assign o[5357] = i[11117];
  assign o[5356] = i[11116];
  assign o[5355] = i[11115];
  assign o[5354] = i[11114];
  assign o[5353] = i[11113];
  assign o[5352] = i[11112];
  assign o[5351] = i[11111];
  assign o[5350] = i[11110];
  assign o[5349] = i[11109];
  assign o[5348] = i[11108];
  assign o[5347] = i[11107];
  assign o[5346] = i[11106];
  assign o[5345] = i[11105];
  assign o[5344] = i[11104];
  assign o[5343] = i[11103];
  assign o[5342] = i[11102];
  assign o[5341] = i[11101];
  assign o[5340] = i[11100];
  assign o[5339] = i[11099];
  assign o[5338] = i[11098];
  assign o[5337] = i[11097];
  assign o[5336] = i[11096];
  assign o[5335] = i[11095];
  assign o[5334] = i[11094];
  assign o[5333] = i[11093];
  assign o[5332] = i[11092];
  assign o[5331] = i[11091];
  assign o[5330] = i[11090];
  assign o[5329] = i[11089];
  assign o[5328] = i[11088];
  assign o[5327] = i[11087];
  assign o[5326] = i[11086];
  assign o[5325] = i[11085];
  assign o[5324] = i[11084];
  assign o[5323] = i[11083];
  assign o[5322] = i[11082];
  assign o[5321] = i[11081];
  assign o[5320] = i[11080];
  assign o[5319] = i[11079];
  assign o[5318] = i[11078];
  assign o[5317] = i[11077];
  assign o[5316] = i[11076];
  assign o[5315] = i[11075];
  assign o[5314] = i[11074];
  assign o[5313] = i[11073];
  assign o[5312] = i[11072];
  assign o[5311] = i[11071];
  assign o[5310] = i[11070];
  assign o[5309] = i[11069];
  assign o[5308] = i[11068];
  assign o[5307] = i[11067];
  assign o[5306] = i[11066];
  assign o[5305] = i[11065];
  assign o[5304] = i[11064];
  assign o[5303] = i[11063];
  assign o[5302] = i[11062];
  assign o[5301] = i[11061];
  assign o[5300] = i[11060];
  assign o[5299] = i[11059];
  assign o[5298] = i[11058];
  assign o[5297] = i[11057];
  assign o[5296] = i[11056];
  assign o[5295] = i[11055];
  assign o[5294] = i[11054];
  assign o[5293] = i[11053];
  assign o[5292] = i[11052];
  assign o[5291] = i[11051];
  assign o[5290] = i[11050];
  assign o[5289] = i[11049];
  assign o[5288] = i[11048];
  assign o[5287] = i[11047];
  assign o[5286] = i[11046];
  assign o[5285] = i[11045];
  assign o[5284] = i[11044];
  assign o[5283] = i[11043];
  assign o[5282] = i[11042];
  assign o[5281] = i[11041];
  assign o[5280] = i[11040];
  assign o[5279] = i[11039];
  assign o[5278] = i[11038];
  assign o[5277] = i[11037];
  assign o[5276] = i[11036];
  assign o[5275] = i[11035];
  assign o[5274] = i[11034];
  assign o[5273] = i[11033];
  assign o[5272] = i[11032];
  assign o[5271] = i[11031];
  assign o[5270] = i[11030];
  assign o[5269] = i[11029];
  assign o[5268] = i[11028];
  assign o[5267] = i[11027];
  assign o[5266] = i[11026];
  assign o[5265] = i[11025];
  assign o[5264] = i[11024];
  assign o[5263] = i[11023];
  assign o[5262] = i[11022];
  assign o[5261] = i[11021];
  assign o[5260] = i[11020];
  assign o[5259] = i[11019];
  assign o[5258] = i[11018];
  assign o[5257] = i[11017];
  assign o[5256] = i[11016];
  assign o[5255] = i[11015];
  assign o[5254] = i[11014];
  assign o[5253] = i[11013];
  assign o[5252] = i[11012];
  assign o[5251] = i[11011];
  assign o[5250] = i[11010];
  assign o[5249] = i[11009];
  assign o[5248] = i[11008];
  assign o[5247] = i[11263];
  assign o[5246] = i[11262];
  assign o[5245] = i[11261];
  assign o[5244] = i[11260];
  assign o[5243] = i[11259];
  assign o[5242] = i[11258];
  assign o[5241] = i[11257];
  assign o[5240] = i[11256];
  assign o[5239] = i[11255];
  assign o[5238] = i[11254];
  assign o[5237] = i[11253];
  assign o[5236] = i[11252];
  assign o[5235] = i[11251];
  assign o[5234] = i[11250];
  assign o[5233] = i[11249];
  assign o[5232] = i[11248];
  assign o[5231] = i[11247];
  assign o[5230] = i[11246];
  assign o[5229] = i[11245];
  assign o[5228] = i[11244];
  assign o[5227] = i[11243];
  assign o[5226] = i[11242];
  assign o[5225] = i[11241];
  assign o[5224] = i[11240];
  assign o[5223] = i[11239];
  assign o[5222] = i[11238];
  assign o[5221] = i[11237];
  assign o[5220] = i[11236];
  assign o[5219] = i[11235];
  assign o[5218] = i[11234];
  assign o[5217] = i[11233];
  assign o[5216] = i[11232];
  assign o[5215] = i[11231];
  assign o[5214] = i[11230];
  assign o[5213] = i[11229];
  assign o[5212] = i[11228];
  assign o[5211] = i[11227];
  assign o[5210] = i[11226];
  assign o[5209] = i[11225];
  assign o[5208] = i[11224];
  assign o[5207] = i[11223];
  assign o[5206] = i[11222];
  assign o[5205] = i[11221];
  assign o[5204] = i[11220];
  assign o[5203] = i[11219];
  assign o[5202] = i[11218];
  assign o[5201] = i[11217];
  assign o[5200] = i[11216];
  assign o[5199] = i[11215];
  assign o[5198] = i[11214];
  assign o[5197] = i[11213];
  assign o[5196] = i[11212];
  assign o[5195] = i[11211];
  assign o[5194] = i[11210];
  assign o[5193] = i[11209];
  assign o[5192] = i[11208];
  assign o[5191] = i[11207];
  assign o[5190] = i[11206];
  assign o[5189] = i[11205];
  assign o[5188] = i[11204];
  assign o[5187] = i[11203];
  assign o[5186] = i[11202];
  assign o[5185] = i[11201];
  assign o[5184] = i[11200];
  assign o[5183] = i[11199];
  assign o[5182] = i[11198];
  assign o[5181] = i[11197];
  assign o[5180] = i[11196];
  assign o[5179] = i[11195];
  assign o[5178] = i[11194];
  assign o[5177] = i[11193];
  assign o[5176] = i[11192];
  assign o[5175] = i[11191];
  assign o[5174] = i[11190];
  assign o[5173] = i[11189];
  assign o[5172] = i[11188];
  assign o[5171] = i[11187];
  assign o[5170] = i[11186];
  assign o[5169] = i[11185];
  assign o[5168] = i[11184];
  assign o[5167] = i[11183];
  assign o[5166] = i[11182];
  assign o[5165] = i[11181];
  assign o[5164] = i[11180];
  assign o[5163] = i[11179];
  assign o[5162] = i[11178];
  assign o[5161] = i[11177];
  assign o[5160] = i[11176];
  assign o[5159] = i[11175];
  assign o[5158] = i[11174];
  assign o[5157] = i[11173];
  assign o[5156] = i[11172];
  assign o[5155] = i[11171];
  assign o[5154] = i[11170];
  assign o[5153] = i[11169];
  assign o[5152] = i[11168];
  assign o[5151] = i[11167];
  assign o[5150] = i[11166];
  assign o[5149] = i[11165];
  assign o[5148] = i[11164];
  assign o[5147] = i[11163];
  assign o[5146] = i[11162];
  assign o[5145] = i[11161];
  assign o[5144] = i[11160];
  assign o[5143] = i[11159];
  assign o[5142] = i[11158];
  assign o[5141] = i[11157];
  assign o[5140] = i[11156];
  assign o[5139] = i[11155];
  assign o[5138] = i[11154];
  assign o[5137] = i[11153];
  assign o[5136] = i[11152];
  assign o[5135] = i[11151];
  assign o[5134] = i[11150];
  assign o[5133] = i[11149];
  assign o[5132] = i[11148];
  assign o[5131] = i[11147];
  assign o[5130] = i[11146];
  assign o[5129] = i[11145];
  assign o[5128] = i[11144];
  assign o[5127] = i[11143];
  assign o[5126] = i[11142];
  assign o[5125] = i[11141];
  assign o[5124] = i[11140];
  assign o[5123] = i[11139];
  assign o[5122] = i[11138];
  assign o[5121] = i[11137];
  assign o[5120] = i[11136];
  assign o[5119] = i[11391];
  assign o[5118] = i[11390];
  assign o[5117] = i[11389];
  assign o[5116] = i[11388];
  assign o[5115] = i[11387];
  assign o[5114] = i[11386];
  assign o[5113] = i[11385];
  assign o[5112] = i[11384];
  assign o[5111] = i[11383];
  assign o[5110] = i[11382];
  assign o[5109] = i[11381];
  assign o[5108] = i[11380];
  assign o[5107] = i[11379];
  assign o[5106] = i[11378];
  assign o[5105] = i[11377];
  assign o[5104] = i[11376];
  assign o[5103] = i[11375];
  assign o[5102] = i[11374];
  assign o[5101] = i[11373];
  assign o[5100] = i[11372];
  assign o[5099] = i[11371];
  assign o[5098] = i[11370];
  assign o[5097] = i[11369];
  assign o[5096] = i[11368];
  assign o[5095] = i[11367];
  assign o[5094] = i[11366];
  assign o[5093] = i[11365];
  assign o[5092] = i[11364];
  assign o[5091] = i[11363];
  assign o[5090] = i[11362];
  assign o[5089] = i[11361];
  assign o[5088] = i[11360];
  assign o[5087] = i[11359];
  assign o[5086] = i[11358];
  assign o[5085] = i[11357];
  assign o[5084] = i[11356];
  assign o[5083] = i[11355];
  assign o[5082] = i[11354];
  assign o[5081] = i[11353];
  assign o[5080] = i[11352];
  assign o[5079] = i[11351];
  assign o[5078] = i[11350];
  assign o[5077] = i[11349];
  assign o[5076] = i[11348];
  assign o[5075] = i[11347];
  assign o[5074] = i[11346];
  assign o[5073] = i[11345];
  assign o[5072] = i[11344];
  assign o[5071] = i[11343];
  assign o[5070] = i[11342];
  assign o[5069] = i[11341];
  assign o[5068] = i[11340];
  assign o[5067] = i[11339];
  assign o[5066] = i[11338];
  assign o[5065] = i[11337];
  assign o[5064] = i[11336];
  assign o[5063] = i[11335];
  assign o[5062] = i[11334];
  assign o[5061] = i[11333];
  assign o[5060] = i[11332];
  assign o[5059] = i[11331];
  assign o[5058] = i[11330];
  assign o[5057] = i[11329];
  assign o[5056] = i[11328];
  assign o[5055] = i[11327];
  assign o[5054] = i[11326];
  assign o[5053] = i[11325];
  assign o[5052] = i[11324];
  assign o[5051] = i[11323];
  assign o[5050] = i[11322];
  assign o[5049] = i[11321];
  assign o[5048] = i[11320];
  assign o[5047] = i[11319];
  assign o[5046] = i[11318];
  assign o[5045] = i[11317];
  assign o[5044] = i[11316];
  assign o[5043] = i[11315];
  assign o[5042] = i[11314];
  assign o[5041] = i[11313];
  assign o[5040] = i[11312];
  assign o[5039] = i[11311];
  assign o[5038] = i[11310];
  assign o[5037] = i[11309];
  assign o[5036] = i[11308];
  assign o[5035] = i[11307];
  assign o[5034] = i[11306];
  assign o[5033] = i[11305];
  assign o[5032] = i[11304];
  assign o[5031] = i[11303];
  assign o[5030] = i[11302];
  assign o[5029] = i[11301];
  assign o[5028] = i[11300];
  assign o[5027] = i[11299];
  assign o[5026] = i[11298];
  assign o[5025] = i[11297];
  assign o[5024] = i[11296];
  assign o[5023] = i[11295];
  assign o[5022] = i[11294];
  assign o[5021] = i[11293];
  assign o[5020] = i[11292];
  assign o[5019] = i[11291];
  assign o[5018] = i[11290];
  assign o[5017] = i[11289];
  assign o[5016] = i[11288];
  assign o[5015] = i[11287];
  assign o[5014] = i[11286];
  assign o[5013] = i[11285];
  assign o[5012] = i[11284];
  assign o[5011] = i[11283];
  assign o[5010] = i[11282];
  assign o[5009] = i[11281];
  assign o[5008] = i[11280];
  assign o[5007] = i[11279];
  assign o[5006] = i[11278];
  assign o[5005] = i[11277];
  assign o[5004] = i[11276];
  assign o[5003] = i[11275];
  assign o[5002] = i[11274];
  assign o[5001] = i[11273];
  assign o[5000] = i[11272];
  assign o[4999] = i[11271];
  assign o[4998] = i[11270];
  assign o[4997] = i[11269];
  assign o[4996] = i[11268];
  assign o[4995] = i[11267];
  assign o[4994] = i[11266];
  assign o[4993] = i[11265];
  assign o[4992] = i[11264];
  assign o[4991] = i[11519];
  assign o[4990] = i[11518];
  assign o[4989] = i[11517];
  assign o[4988] = i[11516];
  assign o[4987] = i[11515];
  assign o[4986] = i[11514];
  assign o[4985] = i[11513];
  assign o[4984] = i[11512];
  assign o[4983] = i[11511];
  assign o[4982] = i[11510];
  assign o[4981] = i[11509];
  assign o[4980] = i[11508];
  assign o[4979] = i[11507];
  assign o[4978] = i[11506];
  assign o[4977] = i[11505];
  assign o[4976] = i[11504];
  assign o[4975] = i[11503];
  assign o[4974] = i[11502];
  assign o[4973] = i[11501];
  assign o[4972] = i[11500];
  assign o[4971] = i[11499];
  assign o[4970] = i[11498];
  assign o[4969] = i[11497];
  assign o[4968] = i[11496];
  assign o[4967] = i[11495];
  assign o[4966] = i[11494];
  assign o[4965] = i[11493];
  assign o[4964] = i[11492];
  assign o[4963] = i[11491];
  assign o[4962] = i[11490];
  assign o[4961] = i[11489];
  assign o[4960] = i[11488];
  assign o[4959] = i[11487];
  assign o[4958] = i[11486];
  assign o[4957] = i[11485];
  assign o[4956] = i[11484];
  assign o[4955] = i[11483];
  assign o[4954] = i[11482];
  assign o[4953] = i[11481];
  assign o[4952] = i[11480];
  assign o[4951] = i[11479];
  assign o[4950] = i[11478];
  assign o[4949] = i[11477];
  assign o[4948] = i[11476];
  assign o[4947] = i[11475];
  assign o[4946] = i[11474];
  assign o[4945] = i[11473];
  assign o[4944] = i[11472];
  assign o[4943] = i[11471];
  assign o[4942] = i[11470];
  assign o[4941] = i[11469];
  assign o[4940] = i[11468];
  assign o[4939] = i[11467];
  assign o[4938] = i[11466];
  assign o[4937] = i[11465];
  assign o[4936] = i[11464];
  assign o[4935] = i[11463];
  assign o[4934] = i[11462];
  assign o[4933] = i[11461];
  assign o[4932] = i[11460];
  assign o[4931] = i[11459];
  assign o[4930] = i[11458];
  assign o[4929] = i[11457];
  assign o[4928] = i[11456];
  assign o[4927] = i[11455];
  assign o[4926] = i[11454];
  assign o[4925] = i[11453];
  assign o[4924] = i[11452];
  assign o[4923] = i[11451];
  assign o[4922] = i[11450];
  assign o[4921] = i[11449];
  assign o[4920] = i[11448];
  assign o[4919] = i[11447];
  assign o[4918] = i[11446];
  assign o[4917] = i[11445];
  assign o[4916] = i[11444];
  assign o[4915] = i[11443];
  assign o[4914] = i[11442];
  assign o[4913] = i[11441];
  assign o[4912] = i[11440];
  assign o[4911] = i[11439];
  assign o[4910] = i[11438];
  assign o[4909] = i[11437];
  assign o[4908] = i[11436];
  assign o[4907] = i[11435];
  assign o[4906] = i[11434];
  assign o[4905] = i[11433];
  assign o[4904] = i[11432];
  assign o[4903] = i[11431];
  assign o[4902] = i[11430];
  assign o[4901] = i[11429];
  assign o[4900] = i[11428];
  assign o[4899] = i[11427];
  assign o[4898] = i[11426];
  assign o[4897] = i[11425];
  assign o[4896] = i[11424];
  assign o[4895] = i[11423];
  assign o[4894] = i[11422];
  assign o[4893] = i[11421];
  assign o[4892] = i[11420];
  assign o[4891] = i[11419];
  assign o[4890] = i[11418];
  assign o[4889] = i[11417];
  assign o[4888] = i[11416];
  assign o[4887] = i[11415];
  assign o[4886] = i[11414];
  assign o[4885] = i[11413];
  assign o[4884] = i[11412];
  assign o[4883] = i[11411];
  assign o[4882] = i[11410];
  assign o[4881] = i[11409];
  assign o[4880] = i[11408];
  assign o[4879] = i[11407];
  assign o[4878] = i[11406];
  assign o[4877] = i[11405];
  assign o[4876] = i[11404];
  assign o[4875] = i[11403];
  assign o[4874] = i[11402];
  assign o[4873] = i[11401];
  assign o[4872] = i[11400];
  assign o[4871] = i[11399];
  assign o[4870] = i[11398];
  assign o[4869] = i[11397];
  assign o[4868] = i[11396];
  assign o[4867] = i[11395];
  assign o[4866] = i[11394];
  assign o[4865] = i[11393];
  assign o[4864] = i[11392];
  assign o[4863] = i[11647];
  assign o[4862] = i[11646];
  assign o[4861] = i[11645];
  assign o[4860] = i[11644];
  assign o[4859] = i[11643];
  assign o[4858] = i[11642];
  assign o[4857] = i[11641];
  assign o[4856] = i[11640];
  assign o[4855] = i[11639];
  assign o[4854] = i[11638];
  assign o[4853] = i[11637];
  assign o[4852] = i[11636];
  assign o[4851] = i[11635];
  assign o[4850] = i[11634];
  assign o[4849] = i[11633];
  assign o[4848] = i[11632];
  assign o[4847] = i[11631];
  assign o[4846] = i[11630];
  assign o[4845] = i[11629];
  assign o[4844] = i[11628];
  assign o[4843] = i[11627];
  assign o[4842] = i[11626];
  assign o[4841] = i[11625];
  assign o[4840] = i[11624];
  assign o[4839] = i[11623];
  assign o[4838] = i[11622];
  assign o[4837] = i[11621];
  assign o[4836] = i[11620];
  assign o[4835] = i[11619];
  assign o[4834] = i[11618];
  assign o[4833] = i[11617];
  assign o[4832] = i[11616];
  assign o[4831] = i[11615];
  assign o[4830] = i[11614];
  assign o[4829] = i[11613];
  assign o[4828] = i[11612];
  assign o[4827] = i[11611];
  assign o[4826] = i[11610];
  assign o[4825] = i[11609];
  assign o[4824] = i[11608];
  assign o[4823] = i[11607];
  assign o[4822] = i[11606];
  assign o[4821] = i[11605];
  assign o[4820] = i[11604];
  assign o[4819] = i[11603];
  assign o[4818] = i[11602];
  assign o[4817] = i[11601];
  assign o[4816] = i[11600];
  assign o[4815] = i[11599];
  assign o[4814] = i[11598];
  assign o[4813] = i[11597];
  assign o[4812] = i[11596];
  assign o[4811] = i[11595];
  assign o[4810] = i[11594];
  assign o[4809] = i[11593];
  assign o[4808] = i[11592];
  assign o[4807] = i[11591];
  assign o[4806] = i[11590];
  assign o[4805] = i[11589];
  assign o[4804] = i[11588];
  assign o[4803] = i[11587];
  assign o[4802] = i[11586];
  assign o[4801] = i[11585];
  assign o[4800] = i[11584];
  assign o[4799] = i[11583];
  assign o[4798] = i[11582];
  assign o[4797] = i[11581];
  assign o[4796] = i[11580];
  assign o[4795] = i[11579];
  assign o[4794] = i[11578];
  assign o[4793] = i[11577];
  assign o[4792] = i[11576];
  assign o[4791] = i[11575];
  assign o[4790] = i[11574];
  assign o[4789] = i[11573];
  assign o[4788] = i[11572];
  assign o[4787] = i[11571];
  assign o[4786] = i[11570];
  assign o[4785] = i[11569];
  assign o[4784] = i[11568];
  assign o[4783] = i[11567];
  assign o[4782] = i[11566];
  assign o[4781] = i[11565];
  assign o[4780] = i[11564];
  assign o[4779] = i[11563];
  assign o[4778] = i[11562];
  assign o[4777] = i[11561];
  assign o[4776] = i[11560];
  assign o[4775] = i[11559];
  assign o[4774] = i[11558];
  assign o[4773] = i[11557];
  assign o[4772] = i[11556];
  assign o[4771] = i[11555];
  assign o[4770] = i[11554];
  assign o[4769] = i[11553];
  assign o[4768] = i[11552];
  assign o[4767] = i[11551];
  assign o[4766] = i[11550];
  assign o[4765] = i[11549];
  assign o[4764] = i[11548];
  assign o[4763] = i[11547];
  assign o[4762] = i[11546];
  assign o[4761] = i[11545];
  assign o[4760] = i[11544];
  assign o[4759] = i[11543];
  assign o[4758] = i[11542];
  assign o[4757] = i[11541];
  assign o[4756] = i[11540];
  assign o[4755] = i[11539];
  assign o[4754] = i[11538];
  assign o[4753] = i[11537];
  assign o[4752] = i[11536];
  assign o[4751] = i[11535];
  assign o[4750] = i[11534];
  assign o[4749] = i[11533];
  assign o[4748] = i[11532];
  assign o[4747] = i[11531];
  assign o[4746] = i[11530];
  assign o[4745] = i[11529];
  assign o[4744] = i[11528];
  assign o[4743] = i[11527];
  assign o[4742] = i[11526];
  assign o[4741] = i[11525];
  assign o[4740] = i[11524];
  assign o[4739] = i[11523];
  assign o[4738] = i[11522];
  assign o[4737] = i[11521];
  assign o[4736] = i[11520];
  assign o[4735] = i[11775];
  assign o[4734] = i[11774];
  assign o[4733] = i[11773];
  assign o[4732] = i[11772];
  assign o[4731] = i[11771];
  assign o[4730] = i[11770];
  assign o[4729] = i[11769];
  assign o[4728] = i[11768];
  assign o[4727] = i[11767];
  assign o[4726] = i[11766];
  assign o[4725] = i[11765];
  assign o[4724] = i[11764];
  assign o[4723] = i[11763];
  assign o[4722] = i[11762];
  assign o[4721] = i[11761];
  assign o[4720] = i[11760];
  assign o[4719] = i[11759];
  assign o[4718] = i[11758];
  assign o[4717] = i[11757];
  assign o[4716] = i[11756];
  assign o[4715] = i[11755];
  assign o[4714] = i[11754];
  assign o[4713] = i[11753];
  assign o[4712] = i[11752];
  assign o[4711] = i[11751];
  assign o[4710] = i[11750];
  assign o[4709] = i[11749];
  assign o[4708] = i[11748];
  assign o[4707] = i[11747];
  assign o[4706] = i[11746];
  assign o[4705] = i[11745];
  assign o[4704] = i[11744];
  assign o[4703] = i[11743];
  assign o[4702] = i[11742];
  assign o[4701] = i[11741];
  assign o[4700] = i[11740];
  assign o[4699] = i[11739];
  assign o[4698] = i[11738];
  assign o[4697] = i[11737];
  assign o[4696] = i[11736];
  assign o[4695] = i[11735];
  assign o[4694] = i[11734];
  assign o[4693] = i[11733];
  assign o[4692] = i[11732];
  assign o[4691] = i[11731];
  assign o[4690] = i[11730];
  assign o[4689] = i[11729];
  assign o[4688] = i[11728];
  assign o[4687] = i[11727];
  assign o[4686] = i[11726];
  assign o[4685] = i[11725];
  assign o[4684] = i[11724];
  assign o[4683] = i[11723];
  assign o[4682] = i[11722];
  assign o[4681] = i[11721];
  assign o[4680] = i[11720];
  assign o[4679] = i[11719];
  assign o[4678] = i[11718];
  assign o[4677] = i[11717];
  assign o[4676] = i[11716];
  assign o[4675] = i[11715];
  assign o[4674] = i[11714];
  assign o[4673] = i[11713];
  assign o[4672] = i[11712];
  assign o[4671] = i[11711];
  assign o[4670] = i[11710];
  assign o[4669] = i[11709];
  assign o[4668] = i[11708];
  assign o[4667] = i[11707];
  assign o[4666] = i[11706];
  assign o[4665] = i[11705];
  assign o[4664] = i[11704];
  assign o[4663] = i[11703];
  assign o[4662] = i[11702];
  assign o[4661] = i[11701];
  assign o[4660] = i[11700];
  assign o[4659] = i[11699];
  assign o[4658] = i[11698];
  assign o[4657] = i[11697];
  assign o[4656] = i[11696];
  assign o[4655] = i[11695];
  assign o[4654] = i[11694];
  assign o[4653] = i[11693];
  assign o[4652] = i[11692];
  assign o[4651] = i[11691];
  assign o[4650] = i[11690];
  assign o[4649] = i[11689];
  assign o[4648] = i[11688];
  assign o[4647] = i[11687];
  assign o[4646] = i[11686];
  assign o[4645] = i[11685];
  assign o[4644] = i[11684];
  assign o[4643] = i[11683];
  assign o[4642] = i[11682];
  assign o[4641] = i[11681];
  assign o[4640] = i[11680];
  assign o[4639] = i[11679];
  assign o[4638] = i[11678];
  assign o[4637] = i[11677];
  assign o[4636] = i[11676];
  assign o[4635] = i[11675];
  assign o[4634] = i[11674];
  assign o[4633] = i[11673];
  assign o[4632] = i[11672];
  assign o[4631] = i[11671];
  assign o[4630] = i[11670];
  assign o[4629] = i[11669];
  assign o[4628] = i[11668];
  assign o[4627] = i[11667];
  assign o[4626] = i[11666];
  assign o[4625] = i[11665];
  assign o[4624] = i[11664];
  assign o[4623] = i[11663];
  assign o[4622] = i[11662];
  assign o[4621] = i[11661];
  assign o[4620] = i[11660];
  assign o[4619] = i[11659];
  assign o[4618] = i[11658];
  assign o[4617] = i[11657];
  assign o[4616] = i[11656];
  assign o[4615] = i[11655];
  assign o[4614] = i[11654];
  assign o[4613] = i[11653];
  assign o[4612] = i[11652];
  assign o[4611] = i[11651];
  assign o[4610] = i[11650];
  assign o[4609] = i[11649];
  assign o[4608] = i[11648];
  assign o[4607] = i[11903];
  assign o[4606] = i[11902];
  assign o[4605] = i[11901];
  assign o[4604] = i[11900];
  assign o[4603] = i[11899];
  assign o[4602] = i[11898];
  assign o[4601] = i[11897];
  assign o[4600] = i[11896];
  assign o[4599] = i[11895];
  assign o[4598] = i[11894];
  assign o[4597] = i[11893];
  assign o[4596] = i[11892];
  assign o[4595] = i[11891];
  assign o[4594] = i[11890];
  assign o[4593] = i[11889];
  assign o[4592] = i[11888];
  assign o[4591] = i[11887];
  assign o[4590] = i[11886];
  assign o[4589] = i[11885];
  assign o[4588] = i[11884];
  assign o[4587] = i[11883];
  assign o[4586] = i[11882];
  assign o[4585] = i[11881];
  assign o[4584] = i[11880];
  assign o[4583] = i[11879];
  assign o[4582] = i[11878];
  assign o[4581] = i[11877];
  assign o[4580] = i[11876];
  assign o[4579] = i[11875];
  assign o[4578] = i[11874];
  assign o[4577] = i[11873];
  assign o[4576] = i[11872];
  assign o[4575] = i[11871];
  assign o[4574] = i[11870];
  assign o[4573] = i[11869];
  assign o[4572] = i[11868];
  assign o[4571] = i[11867];
  assign o[4570] = i[11866];
  assign o[4569] = i[11865];
  assign o[4568] = i[11864];
  assign o[4567] = i[11863];
  assign o[4566] = i[11862];
  assign o[4565] = i[11861];
  assign o[4564] = i[11860];
  assign o[4563] = i[11859];
  assign o[4562] = i[11858];
  assign o[4561] = i[11857];
  assign o[4560] = i[11856];
  assign o[4559] = i[11855];
  assign o[4558] = i[11854];
  assign o[4557] = i[11853];
  assign o[4556] = i[11852];
  assign o[4555] = i[11851];
  assign o[4554] = i[11850];
  assign o[4553] = i[11849];
  assign o[4552] = i[11848];
  assign o[4551] = i[11847];
  assign o[4550] = i[11846];
  assign o[4549] = i[11845];
  assign o[4548] = i[11844];
  assign o[4547] = i[11843];
  assign o[4546] = i[11842];
  assign o[4545] = i[11841];
  assign o[4544] = i[11840];
  assign o[4543] = i[11839];
  assign o[4542] = i[11838];
  assign o[4541] = i[11837];
  assign o[4540] = i[11836];
  assign o[4539] = i[11835];
  assign o[4538] = i[11834];
  assign o[4537] = i[11833];
  assign o[4536] = i[11832];
  assign o[4535] = i[11831];
  assign o[4534] = i[11830];
  assign o[4533] = i[11829];
  assign o[4532] = i[11828];
  assign o[4531] = i[11827];
  assign o[4530] = i[11826];
  assign o[4529] = i[11825];
  assign o[4528] = i[11824];
  assign o[4527] = i[11823];
  assign o[4526] = i[11822];
  assign o[4525] = i[11821];
  assign o[4524] = i[11820];
  assign o[4523] = i[11819];
  assign o[4522] = i[11818];
  assign o[4521] = i[11817];
  assign o[4520] = i[11816];
  assign o[4519] = i[11815];
  assign o[4518] = i[11814];
  assign o[4517] = i[11813];
  assign o[4516] = i[11812];
  assign o[4515] = i[11811];
  assign o[4514] = i[11810];
  assign o[4513] = i[11809];
  assign o[4512] = i[11808];
  assign o[4511] = i[11807];
  assign o[4510] = i[11806];
  assign o[4509] = i[11805];
  assign o[4508] = i[11804];
  assign o[4507] = i[11803];
  assign o[4506] = i[11802];
  assign o[4505] = i[11801];
  assign o[4504] = i[11800];
  assign o[4503] = i[11799];
  assign o[4502] = i[11798];
  assign o[4501] = i[11797];
  assign o[4500] = i[11796];
  assign o[4499] = i[11795];
  assign o[4498] = i[11794];
  assign o[4497] = i[11793];
  assign o[4496] = i[11792];
  assign o[4495] = i[11791];
  assign o[4494] = i[11790];
  assign o[4493] = i[11789];
  assign o[4492] = i[11788];
  assign o[4491] = i[11787];
  assign o[4490] = i[11786];
  assign o[4489] = i[11785];
  assign o[4488] = i[11784];
  assign o[4487] = i[11783];
  assign o[4486] = i[11782];
  assign o[4485] = i[11781];
  assign o[4484] = i[11780];
  assign o[4483] = i[11779];
  assign o[4482] = i[11778];
  assign o[4481] = i[11777];
  assign o[4480] = i[11776];
  assign o[4479] = i[12031];
  assign o[4478] = i[12030];
  assign o[4477] = i[12029];
  assign o[4476] = i[12028];
  assign o[4475] = i[12027];
  assign o[4474] = i[12026];
  assign o[4473] = i[12025];
  assign o[4472] = i[12024];
  assign o[4471] = i[12023];
  assign o[4470] = i[12022];
  assign o[4469] = i[12021];
  assign o[4468] = i[12020];
  assign o[4467] = i[12019];
  assign o[4466] = i[12018];
  assign o[4465] = i[12017];
  assign o[4464] = i[12016];
  assign o[4463] = i[12015];
  assign o[4462] = i[12014];
  assign o[4461] = i[12013];
  assign o[4460] = i[12012];
  assign o[4459] = i[12011];
  assign o[4458] = i[12010];
  assign o[4457] = i[12009];
  assign o[4456] = i[12008];
  assign o[4455] = i[12007];
  assign o[4454] = i[12006];
  assign o[4453] = i[12005];
  assign o[4452] = i[12004];
  assign o[4451] = i[12003];
  assign o[4450] = i[12002];
  assign o[4449] = i[12001];
  assign o[4448] = i[12000];
  assign o[4447] = i[11999];
  assign o[4446] = i[11998];
  assign o[4445] = i[11997];
  assign o[4444] = i[11996];
  assign o[4443] = i[11995];
  assign o[4442] = i[11994];
  assign o[4441] = i[11993];
  assign o[4440] = i[11992];
  assign o[4439] = i[11991];
  assign o[4438] = i[11990];
  assign o[4437] = i[11989];
  assign o[4436] = i[11988];
  assign o[4435] = i[11987];
  assign o[4434] = i[11986];
  assign o[4433] = i[11985];
  assign o[4432] = i[11984];
  assign o[4431] = i[11983];
  assign o[4430] = i[11982];
  assign o[4429] = i[11981];
  assign o[4428] = i[11980];
  assign o[4427] = i[11979];
  assign o[4426] = i[11978];
  assign o[4425] = i[11977];
  assign o[4424] = i[11976];
  assign o[4423] = i[11975];
  assign o[4422] = i[11974];
  assign o[4421] = i[11973];
  assign o[4420] = i[11972];
  assign o[4419] = i[11971];
  assign o[4418] = i[11970];
  assign o[4417] = i[11969];
  assign o[4416] = i[11968];
  assign o[4415] = i[11967];
  assign o[4414] = i[11966];
  assign o[4413] = i[11965];
  assign o[4412] = i[11964];
  assign o[4411] = i[11963];
  assign o[4410] = i[11962];
  assign o[4409] = i[11961];
  assign o[4408] = i[11960];
  assign o[4407] = i[11959];
  assign o[4406] = i[11958];
  assign o[4405] = i[11957];
  assign o[4404] = i[11956];
  assign o[4403] = i[11955];
  assign o[4402] = i[11954];
  assign o[4401] = i[11953];
  assign o[4400] = i[11952];
  assign o[4399] = i[11951];
  assign o[4398] = i[11950];
  assign o[4397] = i[11949];
  assign o[4396] = i[11948];
  assign o[4395] = i[11947];
  assign o[4394] = i[11946];
  assign o[4393] = i[11945];
  assign o[4392] = i[11944];
  assign o[4391] = i[11943];
  assign o[4390] = i[11942];
  assign o[4389] = i[11941];
  assign o[4388] = i[11940];
  assign o[4387] = i[11939];
  assign o[4386] = i[11938];
  assign o[4385] = i[11937];
  assign o[4384] = i[11936];
  assign o[4383] = i[11935];
  assign o[4382] = i[11934];
  assign o[4381] = i[11933];
  assign o[4380] = i[11932];
  assign o[4379] = i[11931];
  assign o[4378] = i[11930];
  assign o[4377] = i[11929];
  assign o[4376] = i[11928];
  assign o[4375] = i[11927];
  assign o[4374] = i[11926];
  assign o[4373] = i[11925];
  assign o[4372] = i[11924];
  assign o[4371] = i[11923];
  assign o[4370] = i[11922];
  assign o[4369] = i[11921];
  assign o[4368] = i[11920];
  assign o[4367] = i[11919];
  assign o[4366] = i[11918];
  assign o[4365] = i[11917];
  assign o[4364] = i[11916];
  assign o[4363] = i[11915];
  assign o[4362] = i[11914];
  assign o[4361] = i[11913];
  assign o[4360] = i[11912];
  assign o[4359] = i[11911];
  assign o[4358] = i[11910];
  assign o[4357] = i[11909];
  assign o[4356] = i[11908];
  assign o[4355] = i[11907];
  assign o[4354] = i[11906];
  assign o[4353] = i[11905];
  assign o[4352] = i[11904];
  assign o[4351] = i[12159];
  assign o[4350] = i[12158];
  assign o[4349] = i[12157];
  assign o[4348] = i[12156];
  assign o[4347] = i[12155];
  assign o[4346] = i[12154];
  assign o[4345] = i[12153];
  assign o[4344] = i[12152];
  assign o[4343] = i[12151];
  assign o[4342] = i[12150];
  assign o[4341] = i[12149];
  assign o[4340] = i[12148];
  assign o[4339] = i[12147];
  assign o[4338] = i[12146];
  assign o[4337] = i[12145];
  assign o[4336] = i[12144];
  assign o[4335] = i[12143];
  assign o[4334] = i[12142];
  assign o[4333] = i[12141];
  assign o[4332] = i[12140];
  assign o[4331] = i[12139];
  assign o[4330] = i[12138];
  assign o[4329] = i[12137];
  assign o[4328] = i[12136];
  assign o[4327] = i[12135];
  assign o[4326] = i[12134];
  assign o[4325] = i[12133];
  assign o[4324] = i[12132];
  assign o[4323] = i[12131];
  assign o[4322] = i[12130];
  assign o[4321] = i[12129];
  assign o[4320] = i[12128];
  assign o[4319] = i[12127];
  assign o[4318] = i[12126];
  assign o[4317] = i[12125];
  assign o[4316] = i[12124];
  assign o[4315] = i[12123];
  assign o[4314] = i[12122];
  assign o[4313] = i[12121];
  assign o[4312] = i[12120];
  assign o[4311] = i[12119];
  assign o[4310] = i[12118];
  assign o[4309] = i[12117];
  assign o[4308] = i[12116];
  assign o[4307] = i[12115];
  assign o[4306] = i[12114];
  assign o[4305] = i[12113];
  assign o[4304] = i[12112];
  assign o[4303] = i[12111];
  assign o[4302] = i[12110];
  assign o[4301] = i[12109];
  assign o[4300] = i[12108];
  assign o[4299] = i[12107];
  assign o[4298] = i[12106];
  assign o[4297] = i[12105];
  assign o[4296] = i[12104];
  assign o[4295] = i[12103];
  assign o[4294] = i[12102];
  assign o[4293] = i[12101];
  assign o[4292] = i[12100];
  assign o[4291] = i[12099];
  assign o[4290] = i[12098];
  assign o[4289] = i[12097];
  assign o[4288] = i[12096];
  assign o[4287] = i[12095];
  assign o[4286] = i[12094];
  assign o[4285] = i[12093];
  assign o[4284] = i[12092];
  assign o[4283] = i[12091];
  assign o[4282] = i[12090];
  assign o[4281] = i[12089];
  assign o[4280] = i[12088];
  assign o[4279] = i[12087];
  assign o[4278] = i[12086];
  assign o[4277] = i[12085];
  assign o[4276] = i[12084];
  assign o[4275] = i[12083];
  assign o[4274] = i[12082];
  assign o[4273] = i[12081];
  assign o[4272] = i[12080];
  assign o[4271] = i[12079];
  assign o[4270] = i[12078];
  assign o[4269] = i[12077];
  assign o[4268] = i[12076];
  assign o[4267] = i[12075];
  assign o[4266] = i[12074];
  assign o[4265] = i[12073];
  assign o[4264] = i[12072];
  assign o[4263] = i[12071];
  assign o[4262] = i[12070];
  assign o[4261] = i[12069];
  assign o[4260] = i[12068];
  assign o[4259] = i[12067];
  assign o[4258] = i[12066];
  assign o[4257] = i[12065];
  assign o[4256] = i[12064];
  assign o[4255] = i[12063];
  assign o[4254] = i[12062];
  assign o[4253] = i[12061];
  assign o[4252] = i[12060];
  assign o[4251] = i[12059];
  assign o[4250] = i[12058];
  assign o[4249] = i[12057];
  assign o[4248] = i[12056];
  assign o[4247] = i[12055];
  assign o[4246] = i[12054];
  assign o[4245] = i[12053];
  assign o[4244] = i[12052];
  assign o[4243] = i[12051];
  assign o[4242] = i[12050];
  assign o[4241] = i[12049];
  assign o[4240] = i[12048];
  assign o[4239] = i[12047];
  assign o[4238] = i[12046];
  assign o[4237] = i[12045];
  assign o[4236] = i[12044];
  assign o[4235] = i[12043];
  assign o[4234] = i[12042];
  assign o[4233] = i[12041];
  assign o[4232] = i[12040];
  assign o[4231] = i[12039];
  assign o[4230] = i[12038];
  assign o[4229] = i[12037];
  assign o[4228] = i[12036];
  assign o[4227] = i[12035];
  assign o[4226] = i[12034];
  assign o[4225] = i[12033];
  assign o[4224] = i[12032];
  assign o[4223] = i[12287];
  assign o[4222] = i[12286];
  assign o[4221] = i[12285];
  assign o[4220] = i[12284];
  assign o[4219] = i[12283];
  assign o[4218] = i[12282];
  assign o[4217] = i[12281];
  assign o[4216] = i[12280];
  assign o[4215] = i[12279];
  assign o[4214] = i[12278];
  assign o[4213] = i[12277];
  assign o[4212] = i[12276];
  assign o[4211] = i[12275];
  assign o[4210] = i[12274];
  assign o[4209] = i[12273];
  assign o[4208] = i[12272];
  assign o[4207] = i[12271];
  assign o[4206] = i[12270];
  assign o[4205] = i[12269];
  assign o[4204] = i[12268];
  assign o[4203] = i[12267];
  assign o[4202] = i[12266];
  assign o[4201] = i[12265];
  assign o[4200] = i[12264];
  assign o[4199] = i[12263];
  assign o[4198] = i[12262];
  assign o[4197] = i[12261];
  assign o[4196] = i[12260];
  assign o[4195] = i[12259];
  assign o[4194] = i[12258];
  assign o[4193] = i[12257];
  assign o[4192] = i[12256];
  assign o[4191] = i[12255];
  assign o[4190] = i[12254];
  assign o[4189] = i[12253];
  assign o[4188] = i[12252];
  assign o[4187] = i[12251];
  assign o[4186] = i[12250];
  assign o[4185] = i[12249];
  assign o[4184] = i[12248];
  assign o[4183] = i[12247];
  assign o[4182] = i[12246];
  assign o[4181] = i[12245];
  assign o[4180] = i[12244];
  assign o[4179] = i[12243];
  assign o[4178] = i[12242];
  assign o[4177] = i[12241];
  assign o[4176] = i[12240];
  assign o[4175] = i[12239];
  assign o[4174] = i[12238];
  assign o[4173] = i[12237];
  assign o[4172] = i[12236];
  assign o[4171] = i[12235];
  assign o[4170] = i[12234];
  assign o[4169] = i[12233];
  assign o[4168] = i[12232];
  assign o[4167] = i[12231];
  assign o[4166] = i[12230];
  assign o[4165] = i[12229];
  assign o[4164] = i[12228];
  assign o[4163] = i[12227];
  assign o[4162] = i[12226];
  assign o[4161] = i[12225];
  assign o[4160] = i[12224];
  assign o[4159] = i[12223];
  assign o[4158] = i[12222];
  assign o[4157] = i[12221];
  assign o[4156] = i[12220];
  assign o[4155] = i[12219];
  assign o[4154] = i[12218];
  assign o[4153] = i[12217];
  assign o[4152] = i[12216];
  assign o[4151] = i[12215];
  assign o[4150] = i[12214];
  assign o[4149] = i[12213];
  assign o[4148] = i[12212];
  assign o[4147] = i[12211];
  assign o[4146] = i[12210];
  assign o[4145] = i[12209];
  assign o[4144] = i[12208];
  assign o[4143] = i[12207];
  assign o[4142] = i[12206];
  assign o[4141] = i[12205];
  assign o[4140] = i[12204];
  assign o[4139] = i[12203];
  assign o[4138] = i[12202];
  assign o[4137] = i[12201];
  assign o[4136] = i[12200];
  assign o[4135] = i[12199];
  assign o[4134] = i[12198];
  assign o[4133] = i[12197];
  assign o[4132] = i[12196];
  assign o[4131] = i[12195];
  assign o[4130] = i[12194];
  assign o[4129] = i[12193];
  assign o[4128] = i[12192];
  assign o[4127] = i[12191];
  assign o[4126] = i[12190];
  assign o[4125] = i[12189];
  assign o[4124] = i[12188];
  assign o[4123] = i[12187];
  assign o[4122] = i[12186];
  assign o[4121] = i[12185];
  assign o[4120] = i[12184];
  assign o[4119] = i[12183];
  assign o[4118] = i[12182];
  assign o[4117] = i[12181];
  assign o[4116] = i[12180];
  assign o[4115] = i[12179];
  assign o[4114] = i[12178];
  assign o[4113] = i[12177];
  assign o[4112] = i[12176];
  assign o[4111] = i[12175];
  assign o[4110] = i[12174];
  assign o[4109] = i[12173];
  assign o[4108] = i[12172];
  assign o[4107] = i[12171];
  assign o[4106] = i[12170];
  assign o[4105] = i[12169];
  assign o[4104] = i[12168];
  assign o[4103] = i[12167];
  assign o[4102] = i[12166];
  assign o[4101] = i[12165];
  assign o[4100] = i[12164];
  assign o[4099] = i[12163];
  assign o[4098] = i[12162];
  assign o[4097] = i[12161];
  assign o[4096] = i[12160];
  assign o[4095] = i[12415];
  assign o[4094] = i[12414];
  assign o[4093] = i[12413];
  assign o[4092] = i[12412];
  assign o[4091] = i[12411];
  assign o[4090] = i[12410];
  assign o[4089] = i[12409];
  assign o[4088] = i[12408];
  assign o[4087] = i[12407];
  assign o[4086] = i[12406];
  assign o[4085] = i[12405];
  assign o[4084] = i[12404];
  assign o[4083] = i[12403];
  assign o[4082] = i[12402];
  assign o[4081] = i[12401];
  assign o[4080] = i[12400];
  assign o[4079] = i[12399];
  assign o[4078] = i[12398];
  assign o[4077] = i[12397];
  assign o[4076] = i[12396];
  assign o[4075] = i[12395];
  assign o[4074] = i[12394];
  assign o[4073] = i[12393];
  assign o[4072] = i[12392];
  assign o[4071] = i[12391];
  assign o[4070] = i[12390];
  assign o[4069] = i[12389];
  assign o[4068] = i[12388];
  assign o[4067] = i[12387];
  assign o[4066] = i[12386];
  assign o[4065] = i[12385];
  assign o[4064] = i[12384];
  assign o[4063] = i[12383];
  assign o[4062] = i[12382];
  assign o[4061] = i[12381];
  assign o[4060] = i[12380];
  assign o[4059] = i[12379];
  assign o[4058] = i[12378];
  assign o[4057] = i[12377];
  assign o[4056] = i[12376];
  assign o[4055] = i[12375];
  assign o[4054] = i[12374];
  assign o[4053] = i[12373];
  assign o[4052] = i[12372];
  assign o[4051] = i[12371];
  assign o[4050] = i[12370];
  assign o[4049] = i[12369];
  assign o[4048] = i[12368];
  assign o[4047] = i[12367];
  assign o[4046] = i[12366];
  assign o[4045] = i[12365];
  assign o[4044] = i[12364];
  assign o[4043] = i[12363];
  assign o[4042] = i[12362];
  assign o[4041] = i[12361];
  assign o[4040] = i[12360];
  assign o[4039] = i[12359];
  assign o[4038] = i[12358];
  assign o[4037] = i[12357];
  assign o[4036] = i[12356];
  assign o[4035] = i[12355];
  assign o[4034] = i[12354];
  assign o[4033] = i[12353];
  assign o[4032] = i[12352];
  assign o[4031] = i[12351];
  assign o[4030] = i[12350];
  assign o[4029] = i[12349];
  assign o[4028] = i[12348];
  assign o[4027] = i[12347];
  assign o[4026] = i[12346];
  assign o[4025] = i[12345];
  assign o[4024] = i[12344];
  assign o[4023] = i[12343];
  assign o[4022] = i[12342];
  assign o[4021] = i[12341];
  assign o[4020] = i[12340];
  assign o[4019] = i[12339];
  assign o[4018] = i[12338];
  assign o[4017] = i[12337];
  assign o[4016] = i[12336];
  assign o[4015] = i[12335];
  assign o[4014] = i[12334];
  assign o[4013] = i[12333];
  assign o[4012] = i[12332];
  assign o[4011] = i[12331];
  assign o[4010] = i[12330];
  assign o[4009] = i[12329];
  assign o[4008] = i[12328];
  assign o[4007] = i[12327];
  assign o[4006] = i[12326];
  assign o[4005] = i[12325];
  assign o[4004] = i[12324];
  assign o[4003] = i[12323];
  assign o[4002] = i[12322];
  assign o[4001] = i[12321];
  assign o[4000] = i[12320];
  assign o[3999] = i[12319];
  assign o[3998] = i[12318];
  assign o[3997] = i[12317];
  assign o[3996] = i[12316];
  assign o[3995] = i[12315];
  assign o[3994] = i[12314];
  assign o[3993] = i[12313];
  assign o[3992] = i[12312];
  assign o[3991] = i[12311];
  assign o[3990] = i[12310];
  assign o[3989] = i[12309];
  assign o[3988] = i[12308];
  assign o[3987] = i[12307];
  assign o[3986] = i[12306];
  assign o[3985] = i[12305];
  assign o[3984] = i[12304];
  assign o[3983] = i[12303];
  assign o[3982] = i[12302];
  assign o[3981] = i[12301];
  assign o[3980] = i[12300];
  assign o[3979] = i[12299];
  assign o[3978] = i[12298];
  assign o[3977] = i[12297];
  assign o[3976] = i[12296];
  assign o[3975] = i[12295];
  assign o[3974] = i[12294];
  assign o[3973] = i[12293];
  assign o[3972] = i[12292];
  assign o[3971] = i[12291];
  assign o[3970] = i[12290];
  assign o[3969] = i[12289];
  assign o[3968] = i[12288];
  assign o[3967] = i[12543];
  assign o[3966] = i[12542];
  assign o[3965] = i[12541];
  assign o[3964] = i[12540];
  assign o[3963] = i[12539];
  assign o[3962] = i[12538];
  assign o[3961] = i[12537];
  assign o[3960] = i[12536];
  assign o[3959] = i[12535];
  assign o[3958] = i[12534];
  assign o[3957] = i[12533];
  assign o[3956] = i[12532];
  assign o[3955] = i[12531];
  assign o[3954] = i[12530];
  assign o[3953] = i[12529];
  assign o[3952] = i[12528];
  assign o[3951] = i[12527];
  assign o[3950] = i[12526];
  assign o[3949] = i[12525];
  assign o[3948] = i[12524];
  assign o[3947] = i[12523];
  assign o[3946] = i[12522];
  assign o[3945] = i[12521];
  assign o[3944] = i[12520];
  assign o[3943] = i[12519];
  assign o[3942] = i[12518];
  assign o[3941] = i[12517];
  assign o[3940] = i[12516];
  assign o[3939] = i[12515];
  assign o[3938] = i[12514];
  assign o[3937] = i[12513];
  assign o[3936] = i[12512];
  assign o[3935] = i[12511];
  assign o[3934] = i[12510];
  assign o[3933] = i[12509];
  assign o[3932] = i[12508];
  assign o[3931] = i[12507];
  assign o[3930] = i[12506];
  assign o[3929] = i[12505];
  assign o[3928] = i[12504];
  assign o[3927] = i[12503];
  assign o[3926] = i[12502];
  assign o[3925] = i[12501];
  assign o[3924] = i[12500];
  assign o[3923] = i[12499];
  assign o[3922] = i[12498];
  assign o[3921] = i[12497];
  assign o[3920] = i[12496];
  assign o[3919] = i[12495];
  assign o[3918] = i[12494];
  assign o[3917] = i[12493];
  assign o[3916] = i[12492];
  assign o[3915] = i[12491];
  assign o[3914] = i[12490];
  assign o[3913] = i[12489];
  assign o[3912] = i[12488];
  assign o[3911] = i[12487];
  assign o[3910] = i[12486];
  assign o[3909] = i[12485];
  assign o[3908] = i[12484];
  assign o[3907] = i[12483];
  assign o[3906] = i[12482];
  assign o[3905] = i[12481];
  assign o[3904] = i[12480];
  assign o[3903] = i[12479];
  assign o[3902] = i[12478];
  assign o[3901] = i[12477];
  assign o[3900] = i[12476];
  assign o[3899] = i[12475];
  assign o[3898] = i[12474];
  assign o[3897] = i[12473];
  assign o[3896] = i[12472];
  assign o[3895] = i[12471];
  assign o[3894] = i[12470];
  assign o[3893] = i[12469];
  assign o[3892] = i[12468];
  assign o[3891] = i[12467];
  assign o[3890] = i[12466];
  assign o[3889] = i[12465];
  assign o[3888] = i[12464];
  assign o[3887] = i[12463];
  assign o[3886] = i[12462];
  assign o[3885] = i[12461];
  assign o[3884] = i[12460];
  assign o[3883] = i[12459];
  assign o[3882] = i[12458];
  assign o[3881] = i[12457];
  assign o[3880] = i[12456];
  assign o[3879] = i[12455];
  assign o[3878] = i[12454];
  assign o[3877] = i[12453];
  assign o[3876] = i[12452];
  assign o[3875] = i[12451];
  assign o[3874] = i[12450];
  assign o[3873] = i[12449];
  assign o[3872] = i[12448];
  assign o[3871] = i[12447];
  assign o[3870] = i[12446];
  assign o[3869] = i[12445];
  assign o[3868] = i[12444];
  assign o[3867] = i[12443];
  assign o[3866] = i[12442];
  assign o[3865] = i[12441];
  assign o[3864] = i[12440];
  assign o[3863] = i[12439];
  assign o[3862] = i[12438];
  assign o[3861] = i[12437];
  assign o[3860] = i[12436];
  assign o[3859] = i[12435];
  assign o[3858] = i[12434];
  assign o[3857] = i[12433];
  assign o[3856] = i[12432];
  assign o[3855] = i[12431];
  assign o[3854] = i[12430];
  assign o[3853] = i[12429];
  assign o[3852] = i[12428];
  assign o[3851] = i[12427];
  assign o[3850] = i[12426];
  assign o[3849] = i[12425];
  assign o[3848] = i[12424];
  assign o[3847] = i[12423];
  assign o[3846] = i[12422];
  assign o[3845] = i[12421];
  assign o[3844] = i[12420];
  assign o[3843] = i[12419];
  assign o[3842] = i[12418];
  assign o[3841] = i[12417];
  assign o[3840] = i[12416];
  assign o[3839] = i[12671];
  assign o[3838] = i[12670];
  assign o[3837] = i[12669];
  assign o[3836] = i[12668];
  assign o[3835] = i[12667];
  assign o[3834] = i[12666];
  assign o[3833] = i[12665];
  assign o[3832] = i[12664];
  assign o[3831] = i[12663];
  assign o[3830] = i[12662];
  assign o[3829] = i[12661];
  assign o[3828] = i[12660];
  assign o[3827] = i[12659];
  assign o[3826] = i[12658];
  assign o[3825] = i[12657];
  assign o[3824] = i[12656];
  assign o[3823] = i[12655];
  assign o[3822] = i[12654];
  assign o[3821] = i[12653];
  assign o[3820] = i[12652];
  assign o[3819] = i[12651];
  assign o[3818] = i[12650];
  assign o[3817] = i[12649];
  assign o[3816] = i[12648];
  assign o[3815] = i[12647];
  assign o[3814] = i[12646];
  assign o[3813] = i[12645];
  assign o[3812] = i[12644];
  assign o[3811] = i[12643];
  assign o[3810] = i[12642];
  assign o[3809] = i[12641];
  assign o[3808] = i[12640];
  assign o[3807] = i[12639];
  assign o[3806] = i[12638];
  assign o[3805] = i[12637];
  assign o[3804] = i[12636];
  assign o[3803] = i[12635];
  assign o[3802] = i[12634];
  assign o[3801] = i[12633];
  assign o[3800] = i[12632];
  assign o[3799] = i[12631];
  assign o[3798] = i[12630];
  assign o[3797] = i[12629];
  assign o[3796] = i[12628];
  assign o[3795] = i[12627];
  assign o[3794] = i[12626];
  assign o[3793] = i[12625];
  assign o[3792] = i[12624];
  assign o[3791] = i[12623];
  assign o[3790] = i[12622];
  assign o[3789] = i[12621];
  assign o[3788] = i[12620];
  assign o[3787] = i[12619];
  assign o[3786] = i[12618];
  assign o[3785] = i[12617];
  assign o[3784] = i[12616];
  assign o[3783] = i[12615];
  assign o[3782] = i[12614];
  assign o[3781] = i[12613];
  assign o[3780] = i[12612];
  assign o[3779] = i[12611];
  assign o[3778] = i[12610];
  assign o[3777] = i[12609];
  assign o[3776] = i[12608];
  assign o[3775] = i[12607];
  assign o[3774] = i[12606];
  assign o[3773] = i[12605];
  assign o[3772] = i[12604];
  assign o[3771] = i[12603];
  assign o[3770] = i[12602];
  assign o[3769] = i[12601];
  assign o[3768] = i[12600];
  assign o[3767] = i[12599];
  assign o[3766] = i[12598];
  assign o[3765] = i[12597];
  assign o[3764] = i[12596];
  assign o[3763] = i[12595];
  assign o[3762] = i[12594];
  assign o[3761] = i[12593];
  assign o[3760] = i[12592];
  assign o[3759] = i[12591];
  assign o[3758] = i[12590];
  assign o[3757] = i[12589];
  assign o[3756] = i[12588];
  assign o[3755] = i[12587];
  assign o[3754] = i[12586];
  assign o[3753] = i[12585];
  assign o[3752] = i[12584];
  assign o[3751] = i[12583];
  assign o[3750] = i[12582];
  assign o[3749] = i[12581];
  assign o[3748] = i[12580];
  assign o[3747] = i[12579];
  assign o[3746] = i[12578];
  assign o[3745] = i[12577];
  assign o[3744] = i[12576];
  assign o[3743] = i[12575];
  assign o[3742] = i[12574];
  assign o[3741] = i[12573];
  assign o[3740] = i[12572];
  assign o[3739] = i[12571];
  assign o[3738] = i[12570];
  assign o[3737] = i[12569];
  assign o[3736] = i[12568];
  assign o[3735] = i[12567];
  assign o[3734] = i[12566];
  assign o[3733] = i[12565];
  assign o[3732] = i[12564];
  assign o[3731] = i[12563];
  assign o[3730] = i[12562];
  assign o[3729] = i[12561];
  assign o[3728] = i[12560];
  assign o[3727] = i[12559];
  assign o[3726] = i[12558];
  assign o[3725] = i[12557];
  assign o[3724] = i[12556];
  assign o[3723] = i[12555];
  assign o[3722] = i[12554];
  assign o[3721] = i[12553];
  assign o[3720] = i[12552];
  assign o[3719] = i[12551];
  assign o[3718] = i[12550];
  assign o[3717] = i[12549];
  assign o[3716] = i[12548];
  assign o[3715] = i[12547];
  assign o[3714] = i[12546];
  assign o[3713] = i[12545];
  assign o[3712] = i[12544];
  assign o[3711] = i[12799];
  assign o[3710] = i[12798];
  assign o[3709] = i[12797];
  assign o[3708] = i[12796];
  assign o[3707] = i[12795];
  assign o[3706] = i[12794];
  assign o[3705] = i[12793];
  assign o[3704] = i[12792];
  assign o[3703] = i[12791];
  assign o[3702] = i[12790];
  assign o[3701] = i[12789];
  assign o[3700] = i[12788];
  assign o[3699] = i[12787];
  assign o[3698] = i[12786];
  assign o[3697] = i[12785];
  assign o[3696] = i[12784];
  assign o[3695] = i[12783];
  assign o[3694] = i[12782];
  assign o[3693] = i[12781];
  assign o[3692] = i[12780];
  assign o[3691] = i[12779];
  assign o[3690] = i[12778];
  assign o[3689] = i[12777];
  assign o[3688] = i[12776];
  assign o[3687] = i[12775];
  assign o[3686] = i[12774];
  assign o[3685] = i[12773];
  assign o[3684] = i[12772];
  assign o[3683] = i[12771];
  assign o[3682] = i[12770];
  assign o[3681] = i[12769];
  assign o[3680] = i[12768];
  assign o[3679] = i[12767];
  assign o[3678] = i[12766];
  assign o[3677] = i[12765];
  assign o[3676] = i[12764];
  assign o[3675] = i[12763];
  assign o[3674] = i[12762];
  assign o[3673] = i[12761];
  assign o[3672] = i[12760];
  assign o[3671] = i[12759];
  assign o[3670] = i[12758];
  assign o[3669] = i[12757];
  assign o[3668] = i[12756];
  assign o[3667] = i[12755];
  assign o[3666] = i[12754];
  assign o[3665] = i[12753];
  assign o[3664] = i[12752];
  assign o[3663] = i[12751];
  assign o[3662] = i[12750];
  assign o[3661] = i[12749];
  assign o[3660] = i[12748];
  assign o[3659] = i[12747];
  assign o[3658] = i[12746];
  assign o[3657] = i[12745];
  assign o[3656] = i[12744];
  assign o[3655] = i[12743];
  assign o[3654] = i[12742];
  assign o[3653] = i[12741];
  assign o[3652] = i[12740];
  assign o[3651] = i[12739];
  assign o[3650] = i[12738];
  assign o[3649] = i[12737];
  assign o[3648] = i[12736];
  assign o[3647] = i[12735];
  assign o[3646] = i[12734];
  assign o[3645] = i[12733];
  assign o[3644] = i[12732];
  assign o[3643] = i[12731];
  assign o[3642] = i[12730];
  assign o[3641] = i[12729];
  assign o[3640] = i[12728];
  assign o[3639] = i[12727];
  assign o[3638] = i[12726];
  assign o[3637] = i[12725];
  assign o[3636] = i[12724];
  assign o[3635] = i[12723];
  assign o[3634] = i[12722];
  assign o[3633] = i[12721];
  assign o[3632] = i[12720];
  assign o[3631] = i[12719];
  assign o[3630] = i[12718];
  assign o[3629] = i[12717];
  assign o[3628] = i[12716];
  assign o[3627] = i[12715];
  assign o[3626] = i[12714];
  assign o[3625] = i[12713];
  assign o[3624] = i[12712];
  assign o[3623] = i[12711];
  assign o[3622] = i[12710];
  assign o[3621] = i[12709];
  assign o[3620] = i[12708];
  assign o[3619] = i[12707];
  assign o[3618] = i[12706];
  assign o[3617] = i[12705];
  assign o[3616] = i[12704];
  assign o[3615] = i[12703];
  assign o[3614] = i[12702];
  assign o[3613] = i[12701];
  assign o[3612] = i[12700];
  assign o[3611] = i[12699];
  assign o[3610] = i[12698];
  assign o[3609] = i[12697];
  assign o[3608] = i[12696];
  assign o[3607] = i[12695];
  assign o[3606] = i[12694];
  assign o[3605] = i[12693];
  assign o[3604] = i[12692];
  assign o[3603] = i[12691];
  assign o[3602] = i[12690];
  assign o[3601] = i[12689];
  assign o[3600] = i[12688];
  assign o[3599] = i[12687];
  assign o[3598] = i[12686];
  assign o[3597] = i[12685];
  assign o[3596] = i[12684];
  assign o[3595] = i[12683];
  assign o[3594] = i[12682];
  assign o[3593] = i[12681];
  assign o[3592] = i[12680];
  assign o[3591] = i[12679];
  assign o[3590] = i[12678];
  assign o[3589] = i[12677];
  assign o[3588] = i[12676];
  assign o[3587] = i[12675];
  assign o[3586] = i[12674];
  assign o[3585] = i[12673];
  assign o[3584] = i[12672];
  assign o[3583] = i[12927];
  assign o[3582] = i[12926];
  assign o[3581] = i[12925];
  assign o[3580] = i[12924];
  assign o[3579] = i[12923];
  assign o[3578] = i[12922];
  assign o[3577] = i[12921];
  assign o[3576] = i[12920];
  assign o[3575] = i[12919];
  assign o[3574] = i[12918];
  assign o[3573] = i[12917];
  assign o[3572] = i[12916];
  assign o[3571] = i[12915];
  assign o[3570] = i[12914];
  assign o[3569] = i[12913];
  assign o[3568] = i[12912];
  assign o[3567] = i[12911];
  assign o[3566] = i[12910];
  assign o[3565] = i[12909];
  assign o[3564] = i[12908];
  assign o[3563] = i[12907];
  assign o[3562] = i[12906];
  assign o[3561] = i[12905];
  assign o[3560] = i[12904];
  assign o[3559] = i[12903];
  assign o[3558] = i[12902];
  assign o[3557] = i[12901];
  assign o[3556] = i[12900];
  assign o[3555] = i[12899];
  assign o[3554] = i[12898];
  assign o[3553] = i[12897];
  assign o[3552] = i[12896];
  assign o[3551] = i[12895];
  assign o[3550] = i[12894];
  assign o[3549] = i[12893];
  assign o[3548] = i[12892];
  assign o[3547] = i[12891];
  assign o[3546] = i[12890];
  assign o[3545] = i[12889];
  assign o[3544] = i[12888];
  assign o[3543] = i[12887];
  assign o[3542] = i[12886];
  assign o[3541] = i[12885];
  assign o[3540] = i[12884];
  assign o[3539] = i[12883];
  assign o[3538] = i[12882];
  assign o[3537] = i[12881];
  assign o[3536] = i[12880];
  assign o[3535] = i[12879];
  assign o[3534] = i[12878];
  assign o[3533] = i[12877];
  assign o[3532] = i[12876];
  assign o[3531] = i[12875];
  assign o[3530] = i[12874];
  assign o[3529] = i[12873];
  assign o[3528] = i[12872];
  assign o[3527] = i[12871];
  assign o[3526] = i[12870];
  assign o[3525] = i[12869];
  assign o[3524] = i[12868];
  assign o[3523] = i[12867];
  assign o[3522] = i[12866];
  assign o[3521] = i[12865];
  assign o[3520] = i[12864];
  assign o[3519] = i[12863];
  assign o[3518] = i[12862];
  assign o[3517] = i[12861];
  assign o[3516] = i[12860];
  assign o[3515] = i[12859];
  assign o[3514] = i[12858];
  assign o[3513] = i[12857];
  assign o[3512] = i[12856];
  assign o[3511] = i[12855];
  assign o[3510] = i[12854];
  assign o[3509] = i[12853];
  assign o[3508] = i[12852];
  assign o[3507] = i[12851];
  assign o[3506] = i[12850];
  assign o[3505] = i[12849];
  assign o[3504] = i[12848];
  assign o[3503] = i[12847];
  assign o[3502] = i[12846];
  assign o[3501] = i[12845];
  assign o[3500] = i[12844];
  assign o[3499] = i[12843];
  assign o[3498] = i[12842];
  assign o[3497] = i[12841];
  assign o[3496] = i[12840];
  assign o[3495] = i[12839];
  assign o[3494] = i[12838];
  assign o[3493] = i[12837];
  assign o[3492] = i[12836];
  assign o[3491] = i[12835];
  assign o[3490] = i[12834];
  assign o[3489] = i[12833];
  assign o[3488] = i[12832];
  assign o[3487] = i[12831];
  assign o[3486] = i[12830];
  assign o[3485] = i[12829];
  assign o[3484] = i[12828];
  assign o[3483] = i[12827];
  assign o[3482] = i[12826];
  assign o[3481] = i[12825];
  assign o[3480] = i[12824];
  assign o[3479] = i[12823];
  assign o[3478] = i[12822];
  assign o[3477] = i[12821];
  assign o[3476] = i[12820];
  assign o[3475] = i[12819];
  assign o[3474] = i[12818];
  assign o[3473] = i[12817];
  assign o[3472] = i[12816];
  assign o[3471] = i[12815];
  assign o[3470] = i[12814];
  assign o[3469] = i[12813];
  assign o[3468] = i[12812];
  assign o[3467] = i[12811];
  assign o[3466] = i[12810];
  assign o[3465] = i[12809];
  assign o[3464] = i[12808];
  assign o[3463] = i[12807];
  assign o[3462] = i[12806];
  assign o[3461] = i[12805];
  assign o[3460] = i[12804];
  assign o[3459] = i[12803];
  assign o[3458] = i[12802];
  assign o[3457] = i[12801];
  assign o[3456] = i[12800];
  assign o[3455] = i[13055];
  assign o[3454] = i[13054];
  assign o[3453] = i[13053];
  assign o[3452] = i[13052];
  assign o[3451] = i[13051];
  assign o[3450] = i[13050];
  assign o[3449] = i[13049];
  assign o[3448] = i[13048];
  assign o[3447] = i[13047];
  assign o[3446] = i[13046];
  assign o[3445] = i[13045];
  assign o[3444] = i[13044];
  assign o[3443] = i[13043];
  assign o[3442] = i[13042];
  assign o[3441] = i[13041];
  assign o[3440] = i[13040];
  assign o[3439] = i[13039];
  assign o[3438] = i[13038];
  assign o[3437] = i[13037];
  assign o[3436] = i[13036];
  assign o[3435] = i[13035];
  assign o[3434] = i[13034];
  assign o[3433] = i[13033];
  assign o[3432] = i[13032];
  assign o[3431] = i[13031];
  assign o[3430] = i[13030];
  assign o[3429] = i[13029];
  assign o[3428] = i[13028];
  assign o[3427] = i[13027];
  assign o[3426] = i[13026];
  assign o[3425] = i[13025];
  assign o[3424] = i[13024];
  assign o[3423] = i[13023];
  assign o[3422] = i[13022];
  assign o[3421] = i[13021];
  assign o[3420] = i[13020];
  assign o[3419] = i[13019];
  assign o[3418] = i[13018];
  assign o[3417] = i[13017];
  assign o[3416] = i[13016];
  assign o[3415] = i[13015];
  assign o[3414] = i[13014];
  assign o[3413] = i[13013];
  assign o[3412] = i[13012];
  assign o[3411] = i[13011];
  assign o[3410] = i[13010];
  assign o[3409] = i[13009];
  assign o[3408] = i[13008];
  assign o[3407] = i[13007];
  assign o[3406] = i[13006];
  assign o[3405] = i[13005];
  assign o[3404] = i[13004];
  assign o[3403] = i[13003];
  assign o[3402] = i[13002];
  assign o[3401] = i[13001];
  assign o[3400] = i[13000];
  assign o[3399] = i[12999];
  assign o[3398] = i[12998];
  assign o[3397] = i[12997];
  assign o[3396] = i[12996];
  assign o[3395] = i[12995];
  assign o[3394] = i[12994];
  assign o[3393] = i[12993];
  assign o[3392] = i[12992];
  assign o[3391] = i[12991];
  assign o[3390] = i[12990];
  assign o[3389] = i[12989];
  assign o[3388] = i[12988];
  assign o[3387] = i[12987];
  assign o[3386] = i[12986];
  assign o[3385] = i[12985];
  assign o[3384] = i[12984];
  assign o[3383] = i[12983];
  assign o[3382] = i[12982];
  assign o[3381] = i[12981];
  assign o[3380] = i[12980];
  assign o[3379] = i[12979];
  assign o[3378] = i[12978];
  assign o[3377] = i[12977];
  assign o[3376] = i[12976];
  assign o[3375] = i[12975];
  assign o[3374] = i[12974];
  assign o[3373] = i[12973];
  assign o[3372] = i[12972];
  assign o[3371] = i[12971];
  assign o[3370] = i[12970];
  assign o[3369] = i[12969];
  assign o[3368] = i[12968];
  assign o[3367] = i[12967];
  assign o[3366] = i[12966];
  assign o[3365] = i[12965];
  assign o[3364] = i[12964];
  assign o[3363] = i[12963];
  assign o[3362] = i[12962];
  assign o[3361] = i[12961];
  assign o[3360] = i[12960];
  assign o[3359] = i[12959];
  assign o[3358] = i[12958];
  assign o[3357] = i[12957];
  assign o[3356] = i[12956];
  assign o[3355] = i[12955];
  assign o[3354] = i[12954];
  assign o[3353] = i[12953];
  assign o[3352] = i[12952];
  assign o[3351] = i[12951];
  assign o[3350] = i[12950];
  assign o[3349] = i[12949];
  assign o[3348] = i[12948];
  assign o[3347] = i[12947];
  assign o[3346] = i[12946];
  assign o[3345] = i[12945];
  assign o[3344] = i[12944];
  assign o[3343] = i[12943];
  assign o[3342] = i[12942];
  assign o[3341] = i[12941];
  assign o[3340] = i[12940];
  assign o[3339] = i[12939];
  assign o[3338] = i[12938];
  assign o[3337] = i[12937];
  assign o[3336] = i[12936];
  assign o[3335] = i[12935];
  assign o[3334] = i[12934];
  assign o[3333] = i[12933];
  assign o[3332] = i[12932];
  assign o[3331] = i[12931];
  assign o[3330] = i[12930];
  assign o[3329] = i[12929];
  assign o[3328] = i[12928];
  assign o[3327] = i[13183];
  assign o[3326] = i[13182];
  assign o[3325] = i[13181];
  assign o[3324] = i[13180];
  assign o[3323] = i[13179];
  assign o[3322] = i[13178];
  assign o[3321] = i[13177];
  assign o[3320] = i[13176];
  assign o[3319] = i[13175];
  assign o[3318] = i[13174];
  assign o[3317] = i[13173];
  assign o[3316] = i[13172];
  assign o[3315] = i[13171];
  assign o[3314] = i[13170];
  assign o[3313] = i[13169];
  assign o[3312] = i[13168];
  assign o[3311] = i[13167];
  assign o[3310] = i[13166];
  assign o[3309] = i[13165];
  assign o[3308] = i[13164];
  assign o[3307] = i[13163];
  assign o[3306] = i[13162];
  assign o[3305] = i[13161];
  assign o[3304] = i[13160];
  assign o[3303] = i[13159];
  assign o[3302] = i[13158];
  assign o[3301] = i[13157];
  assign o[3300] = i[13156];
  assign o[3299] = i[13155];
  assign o[3298] = i[13154];
  assign o[3297] = i[13153];
  assign o[3296] = i[13152];
  assign o[3295] = i[13151];
  assign o[3294] = i[13150];
  assign o[3293] = i[13149];
  assign o[3292] = i[13148];
  assign o[3291] = i[13147];
  assign o[3290] = i[13146];
  assign o[3289] = i[13145];
  assign o[3288] = i[13144];
  assign o[3287] = i[13143];
  assign o[3286] = i[13142];
  assign o[3285] = i[13141];
  assign o[3284] = i[13140];
  assign o[3283] = i[13139];
  assign o[3282] = i[13138];
  assign o[3281] = i[13137];
  assign o[3280] = i[13136];
  assign o[3279] = i[13135];
  assign o[3278] = i[13134];
  assign o[3277] = i[13133];
  assign o[3276] = i[13132];
  assign o[3275] = i[13131];
  assign o[3274] = i[13130];
  assign o[3273] = i[13129];
  assign o[3272] = i[13128];
  assign o[3271] = i[13127];
  assign o[3270] = i[13126];
  assign o[3269] = i[13125];
  assign o[3268] = i[13124];
  assign o[3267] = i[13123];
  assign o[3266] = i[13122];
  assign o[3265] = i[13121];
  assign o[3264] = i[13120];
  assign o[3263] = i[13119];
  assign o[3262] = i[13118];
  assign o[3261] = i[13117];
  assign o[3260] = i[13116];
  assign o[3259] = i[13115];
  assign o[3258] = i[13114];
  assign o[3257] = i[13113];
  assign o[3256] = i[13112];
  assign o[3255] = i[13111];
  assign o[3254] = i[13110];
  assign o[3253] = i[13109];
  assign o[3252] = i[13108];
  assign o[3251] = i[13107];
  assign o[3250] = i[13106];
  assign o[3249] = i[13105];
  assign o[3248] = i[13104];
  assign o[3247] = i[13103];
  assign o[3246] = i[13102];
  assign o[3245] = i[13101];
  assign o[3244] = i[13100];
  assign o[3243] = i[13099];
  assign o[3242] = i[13098];
  assign o[3241] = i[13097];
  assign o[3240] = i[13096];
  assign o[3239] = i[13095];
  assign o[3238] = i[13094];
  assign o[3237] = i[13093];
  assign o[3236] = i[13092];
  assign o[3235] = i[13091];
  assign o[3234] = i[13090];
  assign o[3233] = i[13089];
  assign o[3232] = i[13088];
  assign o[3231] = i[13087];
  assign o[3230] = i[13086];
  assign o[3229] = i[13085];
  assign o[3228] = i[13084];
  assign o[3227] = i[13083];
  assign o[3226] = i[13082];
  assign o[3225] = i[13081];
  assign o[3224] = i[13080];
  assign o[3223] = i[13079];
  assign o[3222] = i[13078];
  assign o[3221] = i[13077];
  assign o[3220] = i[13076];
  assign o[3219] = i[13075];
  assign o[3218] = i[13074];
  assign o[3217] = i[13073];
  assign o[3216] = i[13072];
  assign o[3215] = i[13071];
  assign o[3214] = i[13070];
  assign o[3213] = i[13069];
  assign o[3212] = i[13068];
  assign o[3211] = i[13067];
  assign o[3210] = i[13066];
  assign o[3209] = i[13065];
  assign o[3208] = i[13064];
  assign o[3207] = i[13063];
  assign o[3206] = i[13062];
  assign o[3205] = i[13061];
  assign o[3204] = i[13060];
  assign o[3203] = i[13059];
  assign o[3202] = i[13058];
  assign o[3201] = i[13057];
  assign o[3200] = i[13056];
  assign o[3199] = i[13311];
  assign o[3198] = i[13310];
  assign o[3197] = i[13309];
  assign o[3196] = i[13308];
  assign o[3195] = i[13307];
  assign o[3194] = i[13306];
  assign o[3193] = i[13305];
  assign o[3192] = i[13304];
  assign o[3191] = i[13303];
  assign o[3190] = i[13302];
  assign o[3189] = i[13301];
  assign o[3188] = i[13300];
  assign o[3187] = i[13299];
  assign o[3186] = i[13298];
  assign o[3185] = i[13297];
  assign o[3184] = i[13296];
  assign o[3183] = i[13295];
  assign o[3182] = i[13294];
  assign o[3181] = i[13293];
  assign o[3180] = i[13292];
  assign o[3179] = i[13291];
  assign o[3178] = i[13290];
  assign o[3177] = i[13289];
  assign o[3176] = i[13288];
  assign o[3175] = i[13287];
  assign o[3174] = i[13286];
  assign o[3173] = i[13285];
  assign o[3172] = i[13284];
  assign o[3171] = i[13283];
  assign o[3170] = i[13282];
  assign o[3169] = i[13281];
  assign o[3168] = i[13280];
  assign o[3167] = i[13279];
  assign o[3166] = i[13278];
  assign o[3165] = i[13277];
  assign o[3164] = i[13276];
  assign o[3163] = i[13275];
  assign o[3162] = i[13274];
  assign o[3161] = i[13273];
  assign o[3160] = i[13272];
  assign o[3159] = i[13271];
  assign o[3158] = i[13270];
  assign o[3157] = i[13269];
  assign o[3156] = i[13268];
  assign o[3155] = i[13267];
  assign o[3154] = i[13266];
  assign o[3153] = i[13265];
  assign o[3152] = i[13264];
  assign o[3151] = i[13263];
  assign o[3150] = i[13262];
  assign o[3149] = i[13261];
  assign o[3148] = i[13260];
  assign o[3147] = i[13259];
  assign o[3146] = i[13258];
  assign o[3145] = i[13257];
  assign o[3144] = i[13256];
  assign o[3143] = i[13255];
  assign o[3142] = i[13254];
  assign o[3141] = i[13253];
  assign o[3140] = i[13252];
  assign o[3139] = i[13251];
  assign o[3138] = i[13250];
  assign o[3137] = i[13249];
  assign o[3136] = i[13248];
  assign o[3135] = i[13247];
  assign o[3134] = i[13246];
  assign o[3133] = i[13245];
  assign o[3132] = i[13244];
  assign o[3131] = i[13243];
  assign o[3130] = i[13242];
  assign o[3129] = i[13241];
  assign o[3128] = i[13240];
  assign o[3127] = i[13239];
  assign o[3126] = i[13238];
  assign o[3125] = i[13237];
  assign o[3124] = i[13236];
  assign o[3123] = i[13235];
  assign o[3122] = i[13234];
  assign o[3121] = i[13233];
  assign o[3120] = i[13232];
  assign o[3119] = i[13231];
  assign o[3118] = i[13230];
  assign o[3117] = i[13229];
  assign o[3116] = i[13228];
  assign o[3115] = i[13227];
  assign o[3114] = i[13226];
  assign o[3113] = i[13225];
  assign o[3112] = i[13224];
  assign o[3111] = i[13223];
  assign o[3110] = i[13222];
  assign o[3109] = i[13221];
  assign o[3108] = i[13220];
  assign o[3107] = i[13219];
  assign o[3106] = i[13218];
  assign o[3105] = i[13217];
  assign o[3104] = i[13216];
  assign o[3103] = i[13215];
  assign o[3102] = i[13214];
  assign o[3101] = i[13213];
  assign o[3100] = i[13212];
  assign o[3099] = i[13211];
  assign o[3098] = i[13210];
  assign o[3097] = i[13209];
  assign o[3096] = i[13208];
  assign o[3095] = i[13207];
  assign o[3094] = i[13206];
  assign o[3093] = i[13205];
  assign o[3092] = i[13204];
  assign o[3091] = i[13203];
  assign o[3090] = i[13202];
  assign o[3089] = i[13201];
  assign o[3088] = i[13200];
  assign o[3087] = i[13199];
  assign o[3086] = i[13198];
  assign o[3085] = i[13197];
  assign o[3084] = i[13196];
  assign o[3083] = i[13195];
  assign o[3082] = i[13194];
  assign o[3081] = i[13193];
  assign o[3080] = i[13192];
  assign o[3079] = i[13191];
  assign o[3078] = i[13190];
  assign o[3077] = i[13189];
  assign o[3076] = i[13188];
  assign o[3075] = i[13187];
  assign o[3074] = i[13186];
  assign o[3073] = i[13185];
  assign o[3072] = i[13184];
  assign o[3071] = i[13439];
  assign o[3070] = i[13438];
  assign o[3069] = i[13437];
  assign o[3068] = i[13436];
  assign o[3067] = i[13435];
  assign o[3066] = i[13434];
  assign o[3065] = i[13433];
  assign o[3064] = i[13432];
  assign o[3063] = i[13431];
  assign o[3062] = i[13430];
  assign o[3061] = i[13429];
  assign o[3060] = i[13428];
  assign o[3059] = i[13427];
  assign o[3058] = i[13426];
  assign o[3057] = i[13425];
  assign o[3056] = i[13424];
  assign o[3055] = i[13423];
  assign o[3054] = i[13422];
  assign o[3053] = i[13421];
  assign o[3052] = i[13420];
  assign o[3051] = i[13419];
  assign o[3050] = i[13418];
  assign o[3049] = i[13417];
  assign o[3048] = i[13416];
  assign o[3047] = i[13415];
  assign o[3046] = i[13414];
  assign o[3045] = i[13413];
  assign o[3044] = i[13412];
  assign o[3043] = i[13411];
  assign o[3042] = i[13410];
  assign o[3041] = i[13409];
  assign o[3040] = i[13408];
  assign o[3039] = i[13407];
  assign o[3038] = i[13406];
  assign o[3037] = i[13405];
  assign o[3036] = i[13404];
  assign o[3035] = i[13403];
  assign o[3034] = i[13402];
  assign o[3033] = i[13401];
  assign o[3032] = i[13400];
  assign o[3031] = i[13399];
  assign o[3030] = i[13398];
  assign o[3029] = i[13397];
  assign o[3028] = i[13396];
  assign o[3027] = i[13395];
  assign o[3026] = i[13394];
  assign o[3025] = i[13393];
  assign o[3024] = i[13392];
  assign o[3023] = i[13391];
  assign o[3022] = i[13390];
  assign o[3021] = i[13389];
  assign o[3020] = i[13388];
  assign o[3019] = i[13387];
  assign o[3018] = i[13386];
  assign o[3017] = i[13385];
  assign o[3016] = i[13384];
  assign o[3015] = i[13383];
  assign o[3014] = i[13382];
  assign o[3013] = i[13381];
  assign o[3012] = i[13380];
  assign o[3011] = i[13379];
  assign o[3010] = i[13378];
  assign o[3009] = i[13377];
  assign o[3008] = i[13376];
  assign o[3007] = i[13375];
  assign o[3006] = i[13374];
  assign o[3005] = i[13373];
  assign o[3004] = i[13372];
  assign o[3003] = i[13371];
  assign o[3002] = i[13370];
  assign o[3001] = i[13369];
  assign o[3000] = i[13368];
  assign o[2999] = i[13367];
  assign o[2998] = i[13366];
  assign o[2997] = i[13365];
  assign o[2996] = i[13364];
  assign o[2995] = i[13363];
  assign o[2994] = i[13362];
  assign o[2993] = i[13361];
  assign o[2992] = i[13360];
  assign o[2991] = i[13359];
  assign o[2990] = i[13358];
  assign o[2989] = i[13357];
  assign o[2988] = i[13356];
  assign o[2987] = i[13355];
  assign o[2986] = i[13354];
  assign o[2985] = i[13353];
  assign o[2984] = i[13352];
  assign o[2983] = i[13351];
  assign o[2982] = i[13350];
  assign o[2981] = i[13349];
  assign o[2980] = i[13348];
  assign o[2979] = i[13347];
  assign o[2978] = i[13346];
  assign o[2977] = i[13345];
  assign o[2976] = i[13344];
  assign o[2975] = i[13343];
  assign o[2974] = i[13342];
  assign o[2973] = i[13341];
  assign o[2972] = i[13340];
  assign o[2971] = i[13339];
  assign o[2970] = i[13338];
  assign o[2969] = i[13337];
  assign o[2968] = i[13336];
  assign o[2967] = i[13335];
  assign o[2966] = i[13334];
  assign o[2965] = i[13333];
  assign o[2964] = i[13332];
  assign o[2963] = i[13331];
  assign o[2962] = i[13330];
  assign o[2961] = i[13329];
  assign o[2960] = i[13328];
  assign o[2959] = i[13327];
  assign o[2958] = i[13326];
  assign o[2957] = i[13325];
  assign o[2956] = i[13324];
  assign o[2955] = i[13323];
  assign o[2954] = i[13322];
  assign o[2953] = i[13321];
  assign o[2952] = i[13320];
  assign o[2951] = i[13319];
  assign o[2950] = i[13318];
  assign o[2949] = i[13317];
  assign o[2948] = i[13316];
  assign o[2947] = i[13315];
  assign o[2946] = i[13314];
  assign o[2945] = i[13313];
  assign o[2944] = i[13312];
  assign o[2943] = i[13567];
  assign o[2942] = i[13566];
  assign o[2941] = i[13565];
  assign o[2940] = i[13564];
  assign o[2939] = i[13563];
  assign o[2938] = i[13562];
  assign o[2937] = i[13561];
  assign o[2936] = i[13560];
  assign o[2935] = i[13559];
  assign o[2934] = i[13558];
  assign o[2933] = i[13557];
  assign o[2932] = i[13556];
  assign o[2931] = i[13555];
  assign o[2930] = i[13554];
  assign o[2929] = i[13553];
  assign o[2928] = i[13552];
  assign o[2927] = i[13551];
  assign o[2926] = i[13550];
  assign o[2925] = i[13549];
  assign o[2924] = i[13548];
  assign o[2923] = i[13547];
  assign o[2922] = i[13546];
  assign o[2921] = i[13545];
  assign o[2920] = i[13544];
  assign o[2919] = i[13543];
  assign o[2918] = i[13542];
  assign o[2917] = i[13541];
  assign o[2916] = i[13540];
  assign o[2915] = i[13539];
  assign o[2914] = i[13538];
  assign o[2913] = i[13537];
  assign o[2912] = i[13536];
  assign o[2911] = i[13535];
  assign o[2910] = i[13534];
  assign o[2909] = i[13533];
  assign o[2908] = i[13532];
  assign o[2907] = i[13531];
  assign o[2906] = i[13530];
  assign o[2905] = i[13529];
  assign o[2904] = i[13528];
  assign o[2903] = i[13527];
  assign o[2902] = i[13526];
  assign o[2901] = i[13525];
  assign o[2900] = i[13524];
  assign o[2899] = i[13523];
  assign o[2898] = i[13522];
  assign o[2897] = i[13521];
  assign o[2896] = i[13520];
  assign o[2895] = i[13519];
  assign o[2894] = i[13518];
  assign o[2893] = i[13517];
  assign o[2892] = i[13516];
  assign o[2891] = i[13515];
  assign o[2890] = i[13514];
  assign o[2889] = i[13513];
  assign o[2888] = i[13512];
  assign o[2887] = i[13511];
  assign o[2886] = i[13510];
  assign o[2885] = i[13509];
  assign o[2884] = i[13508];
  assign o[2883] = i[13507];
  assign o[2882] = i[13506];
  assign o[2881] = i[13505];
  assign o[2880] = i[13504];
  assign o[2879] = i[13503];
  assign o[2878] = i[13502];
  assign o[2877] = i[13501];
  assign o[2876] = i[13500];
  assign o[2875] = i[13499];
  assign o[2874] = i[13498];
  assign o[2873] = i[13497];
  assign o[2872] = i[13496];
  assign o[2871] = i[13495];
  assign o[2870] = i[13494];
  assign o[2869] = i[13493];
  assign o[2868] = i[13492];
  assign o[2867] = i[13491];
  assign o[2866] = i[13490];
  assign o[2865] = i[13489];
  assign o[2864] = i[13488];
  assign o[2863] = i[13487];
  assign o[2862] = i[13486];
  assign o[2861] = i[13485];
  assign o[2860] = i[13484];
  assign o[2859] = i[13483];
  assign o[2858] = i[13482];
  assign o[2857] = i[13481];
  assign o[2856] = i[13480];
  assign o[2855] = i[13479];
  assign o[2854] = i[13478];
  assign o[2853] = i[13477];
  assign o[2852] = i[13476];
  assign o[2851] = i[13475];
  assign o[2850] = i[13474];
  assign o[2849] = i[13473];
  assign o[2848] = i[13472];
  assign o[2847] = i[13471];
  assign o[2846] = i[13470];
  assign o[2845] = i[13469];
  assign o[2844] = i[13468];
  assign o[2843] = i[13467];
  assign o[2842] = i[13466];
  assign o[2841] = i[13465];
  assign o[2840] = i[13464];
  assign o[2839] = i[13463];
  assign o[2838] = i[13462];
  assign o[2837] = i[13461];
  assign o[2836] = i[13460];
  assign o[2835] = i[13459];
  assign o[2834] = i[13458];
  assign o[2833] = i[13457];
  assign o[2832] = i[13456];
  assign o[2831] = i[13455];
  assign o[2830] = i[13454];
  assign o[2829] = i[13453];
  assign o[2828] = i[13452];
  assign o[2827] = i[13451];
  assign o[2826] = i[13450];
  assign o[2825] = i[13449];
  assign o[2824] = i[13448];
  assign o[2823] = i[13447];
  assign o[2822] = i[13446];
  assign o[2821] = i[13445];
  assign o[2820] = i[13444];
  assign o[2819] = i[13443];
  assign o[2818] = i[13442];
  assign o[2817] = i[13441];
  assign o[2816] = i[13440];
  assign o[2815] = i[13695];
  assign o[2814] = i[13694];
  assign o[2813] = i[13693];
  assign o[2812] = i[13692];
  assign o[2811] = i[13691];
  assign o[2810] = i[13690];
  assign o[2809] = i[13689];
  assign o[2808] = i[13688];
  assign o[2807] = i[13687];
  assign o[2806] = i[13686];
  assign o[2805] = i[13685];
  assign o[2804] = i[13684];
  assign o[2803] = i[13683];
  assign o[2802] = i[13682];
  assign o[2801] = i[13681];
  assign o[2800] = i[13680];
  assign o[2799] = i[13679];
  assign o[2798] = i[13678];
  assign o[2797] = i[13677];
  assign o[2796] = i[13676];
  assign o[2795] = i[13675];
  assign o[2794] = i[13674];
  assign o[2793] = i[13673];
  assign o[2792] = i[13672];
  assign o[2791] = i[13671];
  assign o[2790] = i[13670];
  assign o[2789] = i[13669];
  assign o[2788] = i[13668];
  assign o[2787] = i[13667];
  assign o[2786] = i[13666];
  assign o[2785] = i[13665];
  assign o[2784] = i[13664];
  assign o[2783] = i[13663];
  assign o[2782] = i[13662];
  assign o[2781] = i[13661];
  assign o[2780] = i[13660];
  assign o[2779] = i[13659];
  assign o[2778] = i[13658];
  assign o[2777] = i[13657];
  assign o[2776] = i[13656];
  assign o[2775] = i[13655];
  assign o[2774] = i[13654];
  assign o[2773] = i[13653];
  assign o[2772] = i[13652];
  assign o[2771] = i[13651];
  assign o[2770] = i[13650];
  assign o[2769] = i[13649];
  assign o[2768] = i[13648];
  assign o[2767] = i[13647];
  assign o[2766] = i[13646];
  assign o[2765] = i[13645];
  assign o[2764] = i[13644];
  assign o[2763] = i[13643];
  assign o[2762] = i[13642];
  assign o[2761] = i[13641];
  assign o[2760] = i[13640];
  assign o[2759] = i[13639];
  assign o[2758] = i[13638];
  assign o[2757] = i[13637];
  assign o[2756] = i[13636];
  assign o[2755] = i[13635];
  assign o[2754] = i[13634];
  assign o[2753] = i[13633];
  assign o[2752] = i[13632];
  assign o[2751] = i[13631];
  assign o[2750] = i[13630];
  assign o[2749] = i[13629];
  assign o[2748] = i[13628];
  assign o[2747] = i[13627];
  assign o[2746] = i[13626];
  assign o[2745] = i[13625];
  assign o[2744] = i[13624];
  assign o[2743] = i[13623];
  assign o[2742] = i[13622];
  assign o[2741] = i[13621];
  assign o[2740] = i[13620];
  assign o[2739] = i[13619];
  assign o[2738] = i[13618];
  assign o[2737] = i[13617];
  assign o[2736] = i[13616];
  assign o[2735] = i[13615];
  assign o[2734] = i[13614];
  assign o[2733] = i[13613];
  assign o[2732] = i[13612];
  assign o[2731] = i[13611];
  assign o[2730] = i[13610];
  assign o[2729] = i[13609];
  assign o[2728] = i[13608];
  assign o[2727] = i[13607];
  assign o[2726] = i[13606];
  assign o[2725] = i[13605];
  assign o[2724] = i[13604];
  assign o[2723] = i[13603];
  assign o[2722] = i[13602];
  assign o[2721] = i[13601];
  assign o[2720] = i[13600];
  assign o[2719] = i[13599];
  assign o[2718] = i[13598];
  assign o[2717] = i[13597];
  assign o[2716] = i[13596];
  assign o[2715] = i[13595];
  assign o[2714] = i[13594];
  assign o[2713] = i[13593];
  assign o[2712] = i[13592];
  assign o[2711] = i[13591];
  assign o[2710] = i[13590];
  assign o[2709] = i[13589];
  assign o[2708] = i[13588];
  assign o[2707] = i[13587];
  assign o[2706] = i[13586];
  assign o[2705] = i[13585];
  assign o[2704] = i[13584];
  assign o[2703] = i[13583];
  assign o[2702] = i[13582];
  assign o[2701] = i[13581];
  assign o[2700] = i[13580];
  assign o[2699] = i[13579];
  assign o[2698] = i[13578];
  assign o[2697] = i[13577];
  assign o[2696] = i[13576];
  assign o[2695] = i[13575];
  assign o[2694] = i[13574];
  assign o[2693] = i[13573];
  assign o[2692] = i[13572];
  assign o[2691] = i[13571];
  assign o[2690] = i[13570];
  assign o[2689] = i[13569];
  assign o[2688] = i[13568];
  assign o[2687] = i[13823];
  assign o[2686] = i[13822];
  assign o[2685] = i[13821];
  assign o[2684] = i[13820];
  assign o[2683] = i[13819];
  assign o[2682] = i[13818];
  assign o[2681] = i[13817];
  assign o[2680] = i[13816];
  assign o[2679] = i[13815];
  assign o[2678] = i[13814];
  assign o[2677] = i[13813];
  assign o[2676] = i[13812];
  assign o[2675] = i[13811];
  assign o[2674] = i[13810];
  assign o[2673] = i[13809];
  assign o[2672] = i[13808];
  assign o[2671] = i[13807];
  assign o[2670] = i[13806];
  assign o[2669] = i[13805];
  assign o[2668] = i[13804];
  assign o[2667] = i[13803];
  assign o[2666] = i[13802];
  assign o[2665] = i[13801];
  assign o[2664] = i[13800];
  assign o[2663] = i[13799];
  assign o[2662] = i[13798];
  assign o[2661] = i[13797];
  assign o[2660] = i[13796];
  assign o[2659] = i[13795];
  assign o[2658] = i[13794];
  assign o[2657] = i[13793];
  assign o[2656] = i[13792];
  assign o[2655] = i[13791];
  assign o[2654] = i[13790];
  assign o[2653] = i[13789];
  assign o[2652] = i[13788];
  assign o[2651] = i[13787];
  assign o[2650] = i[13786];
  assign o[2649] = i[13785];
  assign o[2648] = i[13784];
  assign o[2647] = i[13783];
  assign o[2646] = i[13782];
  assign o[2645] = i[13781];
  assign o[2644] = i[13780];
  assign o[2643] = i[13779];
  assign o[2642] = i[13778];
  assign o[2641] = i[13777];
  assign o[2640] = i[13776];
  assign o[2639] = i[13775];
  assign o[2638] = i[13774];
  assign o[2637] = i[13773];
  assign o[2636] = i[13772];
  assign o[2635] = i[13771];
  assign o[2634] = i[13770];
  assign o[2633] = i[13769];
  assign o[2632] = i[13768];
  assign o[2631] = i[13767];
  assign o[2630] = i[13766];
  assign o[2629] = i[13765];
  assign o[2628] = i[13764];
  assign o[2627] = i[13763];
  assign o[2626] = i[13762];
  assign o[2625] = i[13761];
  assign o[2624] = i[13760];
  assign o[2623] = i[13759];
  assign o[2622] = i[13758];
  assign o[2621] = i[13757];
  assign o[2620] = i[13756];
  assign o[2619] = i[13755];
  assign o[2618] = i[13754];
  assign o[2617] = i[13753];
  assign o[2616] = i[13752];
  assign o[2615] = i[13751];
  assign o[2614] = i[13750];
  assign o[2613] = i[13749];
  assign o[2612] = i[13748];
  assign o[2611] = i[13747];
  assign o[2610] = i[13746];
  assign o[2609] = i[13745];
  assign o[2608] = i[13744];
  assign o[2607] = i[13743];
  assign o[2606] = i[13742];
  assign o[2605] = i[13741];
  assign o[2604] = i[13740];
  assign o[2603] = i[13739];
  assign o[2602] = i[13738];
  assign o[2601] = i[13737];
  assign o[2600] = i[13736];
  assign o[2599] = i[13735];
  assign o[2598] = i[13734];
  assign o[2597] = i[13733];
  assign o[2596] = i[13732];
  assign o[2595] = i[13731];
  assign o[2594] = i[13730];
  assign o[2593] = i[13729];
  assign o[2592] = i[13728];
  assign o[2591] = i[13727];
  assign o[2590] = i[13726];
  assign o[2589] = i[13725];
  assign o[2588] = i[13724];
  assign o[2587] = i[13723];
  assign o[2586] = i[13722];
  assign o[2585] = i[13721];
  assign o[2584] = i[13720];
  assign o[2583] = i[13719];
  assign o[2582] = i[13718];
  assign o[2581] = i[13717];
  assign o[2580] = i[13716];
  assign o[2579] = i[13715];
  assign o[2578] = i[13714];
  assign o[2577] = i[13713];
  assign o[2576] = i[13712];
  assign o[2575] = i[13711];
  assign o[2574] = i[13710];
  assign o[2573] = i[13709];
  assign o[2572] = i[13708];
  assign o[2571] = i[13707];
  assign o[2570] = i[13706];
  assign o[2569] = i[13705];
  assign o[2568] = i[13704];
  assign o[2567] = i[13703];
  assign o[2566] = i[13702];
  assign o[2565] = i[13701];
  assign o[2564] = i[13700];
  assign o[2563] = i[13699];
  assign o[2562] = i[13698];
  assign o[2561] = i[13697];
  assign o[2560] = i[13696];
  assign o[2559] = i[13951];
  assign o[2558] = i[13950];
  assign o[2557] = i[13949];
  assign o[2556] = i[13948];
  assign o[2555] = i[13947];
  assign o[2554] = i[13946];
  assign o[2553] = i[13945];
  assign o[2552] = i[13944];
  assign o[2551] = i[13943];
  assign o[2550] = i[13942];
  assign o[2549] = i[13941];
  assign o[2548] = i[13940];
  assign o[2547] = i[13939];
  assign o[2546] = i[13938];
  assign o[2545] = i[13937];
  assign o[2544] = i[13936];
  assign o[2543] = i[13935];
  assign o[2542] = i[13934];
  assign o[2541] = i[13933];
  assign o[2540] = i[13932];
  assign o[2539] = i[13931];
  assign o[2538] = i[13930];
  assign o[2537] = i[13929];
  assign o[2536] = i[13928];
  assign o[2535] = i[13927];
  assign o[2534] = i[13926];
  assign o[2533] = i[13925];
  assign o[2532] = i[13924];
  assign o[2531] = i[13923];
  assign o[2530] = i[13922];
  assign o[2529] = i[13921];
  assign o[2528] = i[13920];
  assign o[2527] = i[13919];
  assign o[2526] = i[13918];
  assign o[2525] = i[13917];
  assign o[2524] = i[13916];
  assign o[2523] = i[13915];
  assign o[2522] = i[13914];
  assign o[2521] = i[13913];
  assign o[2520] = i[13912];
  assign o[2519] = i[13911];
  assign o[2518] = i[13910];
  assign o[2517] = i[13909];
  assign o[2516] = i[13908];
  assign o[2515] = i[13907];
  assign o[2514] = i[13906];
  assign o[2513] = i[13905];
  assign o[2512] = i[13904];
  assign o[2511] = i[13903];
  assign o[2510] = i[13902];
  assign o[2509] = i[13901];
  assign o[2508] = i[13900];
  assign o[2507] = i[13899];
  assign o[2506] = i[13898];
  assign o[2505] = i[13897];
  assign o[2504] = i[13896];
  assign o[2503] = i[13895];
  assign o[2502] = i[13894];
  assign o[2501] = i[13893];
  assign o[2500] = i[13892];
  assign o[2499] = i[13891];
  assign o[2498] = i[13890];
  assign o[2497] = i[13889];
  assign o[2496] = i[13888];
  assign o[2495] = i[13887];
  assign o[2494] = i[13886];
  assign o[2493] = i[13885];
  assign o[2492] = i[13884];
  assign o[2491] = i[13883];
  assign o[2490] = i[13882];
  assign o[2489] = i[13881];
  assign o[2488] = i[13880];
  assign o[2487] = i[13879];
  assign o[2486] = i[13878];
  assign o[2485] = i[13877];
  assign o[2484] = i[13876];
  assign o[2483] = i[13875];
  assign o[2482] = i[13874];
  assign o[2481] = i[13873];
  assign o[2480] = i[13872];
  assign o[2479] = i[13871];
  assign o[2478] = i[13870];
  assign o[2477] = i[13869];
  assign o[2476] = i[13868];
  assign o[2475] = i[13867];
  assign o[2474] = i[13866];
  assign o[2473] = i[13865];
  assign o[2472] = i[13864];
  assign o[2471] = i[13863];
  assign o[2470] = i[13862];
  assign o[2469] = i[13861];
  assign o[2468] = i[13860];
  assign o[2467] = i[13859];
  assign o[2466] = i[13858];
  assign o[2465] = i[13857];
  assign o[2464] = i[13856];
  assign o[2463] = i[13855];
  assign o[2462] = i[13854];
  assign o[2461] = i[13853];
  assign o[2460] = i[13852];
  assign o[2459] = i[13851];
  assign o[2458] = i[13850];
  assign o[2457] = i[13849];
  assign o[2456] = i[13848];
  assign o[2455] = i[13847];
  assign o[2454] = i[13846];
  assign o[2453] = i[13845];
  assign o[2452] = i[13844];
  assign o[2451] = i[13843];
  assign o[2450] = i[13842];
  assign o[2449] = i[13841];
  assign o[2448] = i[13840];
  assign o[2447] = i[13839];
  assign o[2446] = i[13838];
  assign o[2445] = i[13837];
  assign o[2444] = i[13836];
  assign o[2443] = i[13835];
  assign o[2442] = i[13834];
  assign o[2441] = i[13833];
  assign o[2440] = i[13832];
  assign o[2439] = i[13831];
  assign o[2438] = i[13830];
  assign o[2437] = i[13829];
  assign o[2436] = i[13828];
  assign o[2435] = i[13827];
  assign o[2434] = i[13826];
  assign o[2433] = i[13825];
  assign o[2432] = i[13824];
  assign o[2431] = i[14079];
  assign o[2430] = i[14078];
  assign o[2429] = i[14077];
  assign o[2428] = i[14076];
  assign o[2427] = i[14075];
  assign o[2426] = i[14074];
  assign o[2425] = i[14073];
  assign o[2424] = i[14072];
  assign o[2423] = i[14071];
  assign o[2422] = i[14070];
  assign o[2421] = i[14069];
  assign o[2420] = i[14068];
  assign o[2419] = i[14067];
  assign o[2418] = i[14066];
  assign o[2417] = i[14065];
  assign o[2416] = i[14064];
  assign o[2415] = i[14063];
  assign o[2414] = i[14062];
  assign o[2413] = i[14061];
  assign o[2412] = i[14060];
  assign o[2411] = i[14059];
  assign o[2410] = i[14058];
  assign o[2409] = i[14057];
  assign o[2408] = i[14056];
  assign o[2407] = i[14055];
  assign o[2406] = i[14054];
  assign o[2405] = i[14053];
  assign o[2404] = i[14052];
  assign o[2403] = i[14051];
  assign o[2402] = i[14050];
  assign o[2401] = i[14049];
  assign o[2400] = i[14048];
  assign o[2399] = i[14047];
  assign o[2398] = i[14046];
  assign o[2397] = i[14045];
  assign o[2396] = i[14044];
  assign o[2395] = i[14043];
  assign o[2394] = i[14042];
  assign o[2393] = i[14041];
  assign o[2392] = i[14040];
  assign o[2391] = i[14039];
  assign o[2390] = i[14038];
  assign o[2389] = i[14037];
  assign o[2388] = i[14036];
  assign o[2387] = i[14035];
  assign o[2386] = i[14034];
  assign o[2385] = i[14033];
  assign o[2384] = i[14032];
  assign o[2383] = i[14031];
  assign o[2382] = i[14030];
  assign o[2381] = i[14029];
  assign o[2380] = i[14028];
  assign o[2379] = i[14027];
  assign o[2378] = i[14026];
  assign o[2377] = i[14025];
  assign o[2376] = i[14024];
  assign o[2375] = i[14023];
  assign o[2374] = i[14022];
  assign o[2373] = i[14021];
  assign o[2372] = i[14020];
  assign o[2371] = i[14019];
  assign o[2370] = i[14018];
  assign o[2369] = i[14017];
  assign o[2368] = i[14016];
  assign o[2367] = i[14015];
  assign o[2366] = i[14014];
  assign o[2365] = i[14013];
  assign o[2364] = i[14012];
  assign o[2363] = i[14011];
  assign o[2362] = i[14010];
  assign o[2361] = i[14009];
  assign o[2360] = i[14008];
  assign o[2359] = i[14007];
  assign o[2358] = i[14006];
  assign o[2357] = i[14005];
  assign o[2356] = i[14004];
  assign o[2355] = i[14003];
  assign o[2354] = i[14002];
  assign o[2353] = i[14001];
  assign o[2352] = i[14000];
  assign o[2351] = i[13999];
  assign o[2350] = i[13998];
  assign o[2349] = i[13997];
  assign o[2348] = i[13996];
  assign o[2347] = i[13995];
  assign o[2346] = i[13994];
  assign o[2345] = i[13993];
  assign o[2344] = i[13992];
  assign o[2343] = i[13991];
  assign o[2342] = i[13990];
  assign o[2341] = i[13989];
  assign o[2340] = i[13988];
  assign o[2339] = i[13987];
  assign o[2338] = i[13986];
  assign o[2337] = i[13985];
  assign o[2336] = i[13984];
  assign o[2335] = i[13983];
  assign o[2334] = i[13982];
  assign o[2333] = i[13981];
  assign o[2332] = i[13980];
  assign o[2331] = i[13979];
  assign o[2330] = i[13978];
  assign o[2329] = i[13977];
  assign o[2328] = i[13976];
  assign o[2327] = i[13975];
  assign o[2326] = i[13974];
  assign o[2325] = i[13973];
  assign o[2324] = i[13972];
  assign o[2323] = i[13971];
  assign o[2322] = i[13970];
  assign o[2321] = i[13969];
  assign o[2320] = i[13968];
  assign o[2319] = i[13967];
  assign o[2318] = i[13966];
  assign o[2317] = i[13965];
  assign o[2316] = i[13964];
  assign o[2315] = i[13963];
  assign o[2314] = i[13962];
  assign o[2313] = i[13961];
  assign o[2312] = i[13960];
  assign o[2311] = i[13959];
  assign o[2310] = i[13958];
  assign o[2309] = i[13957];
  assign o[2308] = i[13956];
  assign o[2307] = i[13955];
  assign o[2306] = i[13954];
  assign o[2305] = i[13953];
  assign o[2304] = i[13952];
  assign o[2303] = i[14207];
  assign o[2302] = i[14206];
  assign o[2301] = i[14205];
  assign o[2300] = i[14204];
  assign o[2299] = i[14203];
  assign o[2298] = i[14202];
  assign o[2297] = i[14201];
  assign o[2296] = i[14200];
  assign o[2295] = i[14199];
  assign o[2294] = i[14198];
  assign o[2293] = i[14197];
  assign o[2292] = i[14196];
  assign o[2291] = i[14195];
  assign o[2290] = i[14194];
  assign o[2289] = i[14193];
  assign o[2288] = i[14192];
  assign o[2287] = i[14191];
  assign o[2286] = i[14190];
  assign o[2285] = i[14189];
  assign o[2284] = i[14188];
  assign o[2283] = i[14187];
  assign o[2282] = i[14186];
  assign o[2281] = i[14185];
  assign o[2280] = i[14184];
  assign o[2279] = i[14183];
  assign o[2278] = i[14182];
  assign o[2277] = i[14181];
  assign o[2276] = i[14180];
  assign o[2275] = i[14179];
  assign o[2274] = i[14178];
  assign o[2273] = i[14177];
  assign o[2272] = i[14176];
  assign o[2271] = i[14175];
  assign o[2270] = i[14174];
  assign o[2269] = i[14173];
  assign o[2268] = i[14172];
  assign o[2267] = i[14171];
  assign o[2266] = i[14170];
  assign o[2265] = i[14169];
  assign o[2264] = i[14168];
  assign o[2263] = i[14167];
  assign o[2262] = i[14166];
  assign o[2261] = i[14165];
  assign o[2260] = i[14164];
  assign o[2259] = i[14163];
  assign o[2258] = i[14162];
  assign o[2257] = i[14161];
  assign o[2256] = i[14160];
  assign o[2255] = i[14159];
  assign o[2254] = i[14158];
  assign o[2253] = i[14157];
  assign o[2252] = i[14156];
  assign o[2251] = i[14155];
  assign o[2250] = i[14154];
  assign o[2249] = i[14153];
  assign o[2248] = i[14152];
  assign o[2247] = i[14151];
  assign o[2246] = i[14150];
  assign o[2245] = i[14149];
  assign o[2244] = i[14148];
  assign o[2243] = i[14147];
  assign o[2242] = i[14146];
  assign o[2241] = i[14145];
  assign o[2240] = i[14144];
  assign o[2239] = i[14143];
  assign o[2238] = i[14142];
  assign o[2237] = i[14141];
  assign o[2236] = i[14140];
  assign o[2235] = i[14139];
  assign o[2234] = i[14138];
  assign o[2233] = i[14137];
  assign o[2232] = i[14136];
  assign o[2231] = i[14135];
  assign o[2230] = i[14134];
  assign o[2229] = i[14133];
  assign o[2228] = i[14132];
  assign o[2227] = i[14131];
  assign o[2226] = i[14130];
  assign o[2225] = i[14129];
  assign o[2224] = i[14128];
  assign o[2223] = i[14127];
  assign o[2222] = i[14126];
  assign o[2221] = i[14125];
  assign o[2220] = i[14124];
  assign o[2219] = i[14123];
  assign o[2218] = i[14122];
  assign o[2217] = i[14121];
  assign o[2216] = i[14120];
  assign o[2215] = i[14119];
  assign o[2214] = i[14118];
  assign o[2213] = i[14117];
  assign o[2212] = i[14116];
  assign o[2211] = i[14115];
  assign o[2210] = i[14114];
  assign o[2209] = i[14113];
  assign o[2208] = i[14112];
  assign o[2207] = i[14111];
  assign o[2206] = i[14110];
  assign o[2205] = i[14109];
  assign o[2204] = i[14108];
  assign o[2203] = i[14107];
  assign o[2202] = i[14106];
  assign o[2201] = i[14105];
  assign o[2200] = i[14104];
  assign o[2199] = i[14103];
  assign o[2198] = i[14102];
  assign o[2197] = i[14101];
  assign o[2196] = i[14100];
  assign o[2195] = i[14099];
  assign o[2194] = i[14098];
  assign o[2193] = i[14097];
  assign o[2192] = i[14096];
  assign o[2191] = i[14095];
  assign o[2190] = i[14094];
  assign o[2189] = i[14093];
  assign o[2188] = i[14092];
  assign o[2187] = i[14091];
  assign o[2186] = i[14090];
  assign o[2185] = i[14089];
  assign o[2184] = i[14088];
  assign o[2183] = i[14087];
  assign o[2182] = i[14086];
  assign o[2181] = i[14085];
  assign o[2180] = i[14084];
  assign o[2179] = i[14083];
  assign o[2178] = i[14082];
  assign o[2177] = i[14081];
  assign o[2176] = i[14080];
  assign o[2175] = i[14335];
  assign o[2174] = i[14334];
  assign o[2173] = i[14333];
  assign o[2172] = i[14332];
  assign o[2171] = i[14331];
  assign o[2170] = i[14330];
  assign o[2169] = i[14329];
  assign o[2168] = i[14328];
  assign o[2167] = i[14327];
  assign o[2166] = i[14326];
  assign o[2165] = i[14325];
  assign o[2164] = i[14324];
  assign o[2163] = i[14323];
  assign o[2162] = i[14322];
  assign o[2161] = i[14321];
  assign o[2160] = i[14320];
  assign o[2159] = i[14319];
  assign o[2158] = i[14318];
  assign o[2157] = i[14317];
  assign o[2156] = i[14316];
  assign o[2155] = i[14315];
  assign o[2154] = i[14314];
  assign o[2153] = i[14313];
  assign o[2152] = i[14312];
  assign o[2151] = i[14311];
  assign o[2150] = i[14310];
  assign o[2149] = i[14309];
  assign o[2148] = i[14308];
  assign o[2147] = i[14307];
  assign o[2146] = i[14306];
  assign o[2145] = i[14305];
  assign o[2144] = i[14304];
  assign o[2143] = i[14303];
  assign o[2142] = i[14302];
  assign o[2141] = i[14301];
  assign o[2140] = i[14300];
  assign o[2139] = i[14299];
  assign o[2138] = i[14298];
  assign o[2137] = i[14297];
  assign o[2136] = i[14296];
  assign o[2135] = i[14295];
  assign o[2134] = i[14294];
  assign o[2133] = i[14293];
  assign o[2132] = i[14292];
  assign o[2131] = i[14291];
  assign o[2130] = i[14290];
  assign o[2129] = i[14289];
  assign o[2128] = i[14288];
  assign o[2127] = i[14287];
  assign o[2126] = i[14286];
  assign o[2125] = i[14285];
  assign o[2124] = i[14284];
  assign o[2123] = i[14283];
  assign o[2122] = i[14282];
  assign o[2121] = i[14281];
  assign o[2120] = i[14280];
  assign o[2119] = i[14279];
  assign o[2118] = i[14278];
  assign o[2117] = i[14277];
  assign o[2116] = i[14276];
  assign o[2115] = i[14275];
  assign o[2114] = i[14274];
  assign o[2113] = i[14273];
  assign o[2112] = i[14272];
  assign o[2111] = i[14271];
  assign o[2110] = i[14270];
  assign o[2109] = i[14269];
  assign o[2108] = i[14268];
  assign o[2107] = i[14267];
  assign o[2106] = i[14266];
  assign o[2105] = i[14265];
  assign o[2104] = i[14264];
  assign o[2103] = i[14263];
  assign o[2102] = i[14262];
  assign o[2101] = i[14261];
  assign o[2100] = i[14260];
  assign o[2099] = i[14259];
  assign o[2098] = i[14258];
  assign o[2097] = i[14257];
  assign o[2096] = i[14256];
  assign o[2095] = i[14255];
  assign o[2094] = i[14254];
  assign o[2093] = i[14253];
  assign o[2092] = i[14252];
  assign o[2091] = i[14251];
  assign o[2090] = i[14250];
  assign o[2089] = i[14249];
  assign o[2088] = i[14248];
  assign o[2087] = i[14247];
  assign o[2086] = i[14246];
  assign o[2085] = i[14245];
  assign o[2084] = i[14244];
  assign o[2083] = i[14243];
  assign o[2082] = i[14242];
  assign o[2081] = i[14241];
  assign o[2080] = i[14240];
  assign o[2079] = i[14239];
  assign o[2078] = i[14238];
  assign o[2077] = i[14237];
  assign o[2076] = i[14236];
  assign o[2075] = i[14235];
  assign o[2074] = i[14234];
  assign o[2073] = i[14233];
  assign o[2072] = i[14232];
  assign o[2071] = i[14231];
  assign o[2070] = i[14230];
  assign o[2069] = i[14229];
  assign o[2068] = i[14228];
  assign o[2067] = i[14227];
  assign o[2066] = i[14226];
  assign o[2065] = i[14225];
  assign o[2064] = i[14224];
  assign o[2063] = i[14223];
  assign o[2062] = i[14222];
  assign o[2061] = i[14221];
  assign o[2060] = i[14220];
  assign o[2059] = i[14219];
  assign o[2058] = i[14218];
  assign o[2057] = i[14217];
  assign o[2056] = i[14216];
  assign o[2055] = i[14215];
  assign o[2054] = i[14214];
  assign o[2053] = i[14213];
  assign o[2052] = i[14212];
  assign o[2051] = i[14211];
  assign o[2050] = i[14210];
  assign o[2049] = i[14209];
  assign o[2048] = i[14208];
  assign o[2047] = i[14463];
  assign o[2046] = i[14462];
  assign o[2045] = i[14461];
  assign o[2044] = i[14460];
  assign o[2043] = i[14459];
  assign o[2042] = i[14458];
  assign o[2041] = i[14457];
  assign o[2040] = i[14456];
  assign o[2039] = i[14455];
  assign o[2038] = i[14454];
  assign o[2037] = i[14453];
  assign o[2036] = i[14452];
  assign o[2035] = i[14451];
  assign o[2034] = i[14450];
  assign o[2033] = i[14449];
  assign o[2032] = i[14448];
  assign o[2031] = i[14447];
  assign o[2030] = i[14446];
  assign o[2029] = i[14445];
  assign o[2028] = i[14444];
  assign o[2027] = i[14443];
  assign o[2026] = i[14442];
  assign o[2025] = i[14441];
  assign o[2024] = i[14440];
  assign o[2023] = i[14439];
  assign o[2022] = i[14438];
  assign o[2021] = i[14437];
  assign o[2020] = i[14436];
  assign o[2019] = i[14435];
  assign o[2018] = i[14434];
  assign o[2017] = i[14433];
  assign o[2016] = i[14432];
  assign o[2015] = i[14431];
  assign o[2014] = i[14430];
  assign o[2013] = i[14429];
  assign o[2012] = i[14428];
  assign o[2011] = i[14427];
  assign o[2010] = i[14426];
  assign o[2009] = i[14425];
  assign o[2008] = i[14424];
  assign o[2007] = i[14423];
  assign o[2006] = i[14422];
  assign o[2005] = i[14421];
  assign o[2004] = i[14420];
  assign o[2003] = i[14419];
  assign o[2002] = i[14418];
  assign o[2001] = i[14417];
  assign o[2000] = i[14416];
  assign o[1999] = i[14415];
  assign o[1998] = i[14414];
  assign o[1997] = i[14413];
  assign o[1996] = i[14412];
  assign o[1995] = i[14411];
  assign o[1994] = i[14410];
  assign o[1993] = i[14409];
  assign o[1992] = i[14408];
  assign o[1991] = i[14407];
  assign o[1990] = i[14406];
  assign o[1989] = i[14405];
  assign o[1988] = i[14404];
  assign o[1987] = i[14403];
  assign o[1986] = i[14402];
  assign o[1985] = i[14401];
  assign o[1984] = i[14400];
  assign o[1983] = i[14399];
  assign o[1982] = i[14398];
  assign o[1981] = i[14397];
  assign o[1980] = i[14396];
  assign o[1979] = i[14395];
  assign o[1978] = i[14394];
  assign o[1977] = i[14393];
  assign o[1976] = i[14392];
  assign o[1975] = i[14391];
  assign o[1974] = i[14390];
  assign o[1973] = i[14389];
  assign o[1972] = i[14388];
  assign o[1971] = i[14387];
  assign o[1970] = i[14386];
  assign o[1969] = i[14385];
  assign o[1968] = i[14384];
  assign o[1967] = i[14383];
  assign o[1966] = i[14382];
  assign o[1965] = i[14381];
  assign o[1964] = i[14380];
  assign o[1963] = i[14379];
  assign o[1962] = i[14378];
  assign o[1961] = i[14377];
  assign o[1960] = i[14376];
  assign o[1959] = i[14375];
  assign o[1958] = i[14374];
  assign o[1957] = i[14373];
  assign o[1956] = i[14372];
  assign o[1955] = i[14371];
  assign o[1954] = i[14370];
  assign o[1953] = i[14369];
  assign o[1952] = i[14368];
  assign o[1951] = i[14367];
  assign o[1950] = i[14366];
  assign o[1949] = i[14365];
  assign o[1948] = i[14364];
  assign o[1947] = i[14363];
  assign o[1946] = i[14362];
  assign o[1945] = i[14361];
  assign o[1944] = i[14360];
  assign o[1943] = i[14359];
  assign o[1942] = i[14358];
  assign o[1941] = i[14357];
  assign o[1940] = i[14356];
  assign o[1939] = i[14355];
  assign o[1938] = i[14354];
  assign o[1937] = i[14353];
  assign o[1936] = i[14352];
  assign o[1935] = i[14351];
  assign o[1934] = i[14350];
  assign o[1933] = i[14349];
  assign o[1932] = i[14348];
  assign o[1931] = i[14347];
  assign o[1930] = i[14346];
  assign o[1929] = i[14345];
  assign o[1928] = i[14344];
  assign o[1927] = i[14343];
  assign o[1926] = i[14342];
  assign o[1925] = i[14341];
  assign o[1924] = i[14340];
  assign o[1923] = i[14339];
  assign o[1922] = i[14338];
  assign o[1921] = i[14337];
  assign o[1920] = i[14336];
  assign o[1919] = i[14591];
  assign o[1918] = i[14590];
  assign o[1917] = i[14589];
  assign o[1916] = i[14588];
  assign o[1915] = i[14587];
  assign o[1914] = i[14586];
  assign o[1913] = i[14585];
  assign o[1912] = i[14584];
  assign o[1911] = i[14583];
  assign o[1910] = i[14582];
  assign o[1909] = i[14581];
  assign o[1908] = i[14580];
  assign o[1907] = i[14579];
  assign o[1906] = i[14578];
  assign o[1905] = i[14577];
  assign o[1904] = i[14576];
  assign o[1903] = i[14575];
  assign o[1902] = i[14574];
  assign o[1901] = i[14573];
  assign o[1900] = i[14572];
  assign o[1899] = i[14571];
  assign o[1898] = i[14570];
  assign o[1897] = i[14569];
  assign o[1896] = i[14568];
  assign o[1895] = i[14567];
  assign o[1894] = i[14566];
  assign o[1893] = i[14565];
  assign o[1892] = i[14564];
  assign o[1891] = i[14563];
  assign o[1890] = i[14562];
  assign o[1889] = i[14561];
  assign o[1888] = i[14560];
  assign o[1887] = i[14559];
  assign o[1886] = i[14558];
  assign o[1885] = i[14557];
  assign o[1884] = i[14556];
  assign o[1883] = i[14555];
  assign o[1882] = i[14554];
  assign o[1881] = i[14553];
  assign o[1880] = i[14552];
  assign o[1879] = i[14551];
  assign o[1878] = i[14550];
  assign o[1877] = i[14549];
  assign o[1876] = i[14548];
  assign o[1875] = i[14547];
  assign o[1874] = i[14546];
  assign o[1873] = i[14545];
  assign o[1872] = i[14544];
  assign o[1871] = i[14543];
  assign o[1870] = i[14542];
  assign o[1869] = i[14541];
  assign o[1868] = i[14540];
  assign o[1867] = i[14539];
  assign o[1866] = i[14538];
  assign o[1865] = i[14537];
  assign o[1864] = i[14536];
  assign o[1863] = i[14535];
  assign o[1862] = i[14534];
  assign o[1861] = i[14533];
  assign o[1860] = i[14532];
  assign o[1859] = i[14531];
  assign o[1858] = i[14530];
  assign o[1857] = i[14529];
  assign o[1856] = i[14528];
  assign o[1855] = i[14527];
  assign o[1854] = i[14526];
  assign o[1853] = i[14525];
  assign o[1852] = i[14524];
  assign o[1851] = i[14523];
  assign o[1850] = i[14522];
  assign o[1849] = i[14521];
  assign o[1848] = i[14520];
  assign o[1847] = i[14519];
  assign o[1846] = i[14518];
  assign o[1845] = i[14517];
  assign o[1844] = i[14516];
  assign o[1843] = i[14515];
  assign o[1842] = i[14514];
  assign o[1841] = i[14513];
  assign o[1840] = i[14512];
  assign o[1839] = i[14511];
  assign o[1838] = i[14510];
  assign o[1837] = i[14509];
  assign o[1836] = i[14508];
  assign o[1835] = i[14507];
  assign o[1834] = i[14506];
  assign o[1833] = i[14505];
  assign o[1832] = i[14504];
  assign o[1831] = i[14503];
  assign o[1830] = i[14502];
  assign o[1829] = i[14501];
  assign o[1828] = i[14500];
  assign o[1827] = i[14499];
  assign o[1826] = i[14498];
  assign o[1825] = i[14497];
  assign o[1824] = i[14496];
  assign o[1823] = i[14495];
  assign o[1822] = i[14494];
  assign o[1821] = i[14493];
  assign o[1820] = i[14492];
  assign o[1819] = i[14491];
  assign o[1818] = i[14490];
  assign o[1817] = i[14489];
  assign o[1816] = i[14488];
  assign o[1815] = i[14487];
  assign o[1814] = i[14486];
  assign o[1813] = i[14485];
  assign o[1812] = i[14484];
  assign o[1811] = i[14483];
  assign o[1810] = i[14482];
  assign o[1809] = i[14481];
  assign o[1808] = i[14480];
  assign o[1807] = i[14479];
  assign o[1806] = i[14478];
  assign o[1805] = i[14477];
  assign o[1804] = i[14476];
  assign o[1803] = i[14475];
  assign o[1802] = i[14474];
  assign o[1801] = i[14473];
  assign o[1800] = i[14472];
  assign o[1799] = i[14471];
  assign o[1798] = i[14470];
  assign o[1797] = i[14469];
  assign o[1796] = i[14468];
  assign o[1795] = i[14467];
  assign o[1794] = i[14466];
  assign o[1793] = i[14465];
  assign o[1792] = i[14464];
  assign o[1791] = i[14719];
  assign o[1790] = i[14718];
  assign o[1789] = i[14717];
  assign o[1788] = i[14716];
  assign o[1787] = i[14715];
  assign o[1786] = i[14714];
  assign o[1785] = i[14713];
  assign o[1784] = i[14712];
  assign o[1783] = i[14711];
  assign o[1782] = i[14710];
  assign o[1781] = i[14709];
  assign o[1780] = i[14708];
  assign o[1779] = i[14707];
  assign o[1778] = i[14706];
  assign o[1777] = i[14705];
  assign o[1776] = i[14704];
  assign o[1775] = i[14703];
  assign o[1774] = i[14702];
  assign o[1773] = i[14701];
  assign o[1772] = i[14700];
  assign o[1771] = i[14699];
  assign o[1770] = i[14698];
  assign o[1769] = i[14697];
  assign o[1768] = i[14696];
  assign o[1767] = i[14695];
  assign o[1766] = i[14694];
  assign o[1765] = i[14693];
  assign o[1764] = i[14692];
  assign o[1763] = i[14691];
  assign o[1762] = i[14690];
  assign o[1761] = i[14689];
  assign o[1760] = i[14688];
  assign o[1759] = i[14687];
  assign o[1758] = i[14686];
  assign o[1757] = i[14685];
  assign o[1756] = i[14684];
  assign o[1755] = i[14683];
  assign o[1754] = i[14682];
  assign o[1753] = i[14681];
  assign o[1752] = i[14680];
  assign o[1751] = i[14679];
  assign o[1750] = i[14678];
  assign o[1749] = i[14677];
  assign o[1748] = i[14676];
  assign o[1747] = i[14675];
  assign o[1746] = i[14674];
  assign o[1745] = i[14673];
  assign o[1744] = i[14672];
  assign o[1743] = i[14671];
  assign o[1742] = i[14670];
  assign o[1741] = i[14669];
  assign o[1740] = i[14668];
  assign o[1739] = i[14667];
  assign o[1738] = i[14666];
  assign o[1737] = i[14665];
  assign o[1736] = i[14664];
  assign o[1735] = i[14663];
  assign o[1734] = i[14662];
  assign o[1733] = i[14661];
  assign o[1732] = i[14660];
  assign o[1731] = i[14659];
  assign o[1730] = i[14658];
  assign o[1729] = i[14657];
  assign o[1728] = i[14656];
  assign o[1727] = i[14655];
  assign o[1726] = i[14654];
  assign o[1725] = i[14653];
  assign o[1724] = i[14652];
  assign o[1723] = i[14651];
  assign o[1722] = i[14650];
  assign o[1721] = i[14649];
  assign o[1720] = i[14648];
  assign o[1719] = i[14647];
  assign o[1718] = i[14646];
  assign o[1717] = i[14645];
  assign o[1716] = i[14644];
  assign o[1715] = i[14643];
  assign o[1714] = i[14642];
  assign o[1713] = i[14641];
  assign o[1712] = i[14640];
  assign o[1711] = i[14639];
  assign o[1710] = i[14638];
  assign o[1709] = i[14637];
  assign o[1708] = i[14636];
  assign o[1707] = i[14635];
  assign o[1706] = i[14634];
  assign o[1705] = i[14633];
  assign o[1704] = i[14632];
  assign o[1703] = i[14631];
  assign o[1702] = i[14630];
  assign o[1701] = i[14629];
  assign o[1700] = i[14628];
  assign o[1699] = i[14627];
  assign o[1698] = i[14626];
  assign o[1697] = i[14625];
  assign o[1696] = i[14624];
  assign o[1695] = i[14623];
  assign o[1694] = i[14622];
  assign o[1693] = i[14621];
  assign o[1692] = i[14620];
  assign o[1691] = i[14619];
  assign o[1690] = i[14618];
  assign o[1689] = i[14617];
  assign o[1688] = i[14616];
  assign o[1687] = i[14615];
  assign o[1686] = i[14614];
  assign o[1685] = i[14613];
  assign o[1684] = i[14612];
  assign o[1683] = i[14611];
  assign o[1682] = i[14610];
  assign o[1681] = i[14609];
  assign o[1680] = i[14608];
  assign o[1679] = i[14607];
  assign o[1678] = i[14606];
  assign o[1677] = i[14605];
  assign o[1676] = i[14604];
  assign o[1675] = i[14603];
  assign o[1674] = i[14602];
  assign o[1673] = i[14601];
  assign o[1672] = i[14600];
  assign o[1671] = i[14599];
  assign o[1670] = i[14598];
  assign o[1669] = i[14597];
  assign o[1668] = i[14596];
  assign o[1667] = i[14595];
  assign o[1666] = i[14594];
  assign o[1665] = i[14593];
  assign o[1664] = i[14592];
  assign o[1663] = i[14847];
  assign o[1662] = i[14846];
  assign o[1661] = i[14845];
  assign o[1660] = i[14844];
  assign o[1659] = i[14843];
  assign o[1658] = i[14842];
  assign o[1657] = i[14841];
  assign o[1656] = i[14840];
  assign o[1655] = i[14839];
  assign o[1654] = i[14838];
  assign o[1653] = i[14837];
  assign o[1652] = i[14836];
  assign o[1651] = i[14835];
  assign o[1650] = i[14834];
  assign o[1649] = i[14833];
  assign o[1648] = i[14832];
  assign o[1647] = i[14831];
  assign o[1646] = i[14830];
  assign o[1645] = i[14829];
  assign o[1644] = i[14828];
  assign o[1643] = i[14827];
  assign o[1642] = i[14826];
  assign o[1641] = i[14825];
  assign o[1640] = i[14824];
  assign o[1639] = i[14823];
  assign o[1638] = i[14822];
  assign o[1637] = i[14821];
  assign o[1636] = i[14820];
  assign o[1635] = i[14819];
  assign o[1634] = i[14818];
  assign o[1633] = i[14817];
  assign o[1632] = i[14816];
  assign o[1631] = i[14815];
  assign o[1630] = i[14814];
  assign o[1629] = i[14813];
  assign o[1628] = i[14812];
  assign o[1627] = i[14811];
  assign o[1626] = i[14810];
  assign o[1625] = i[14809];
  assign o[1624] = i[14808];
  assign o[1623] = i[14807];
  assign o[1622] = i[14806];
  assign o[1621] = i[14805];
  assign o[1620] = i[14804];
  assign o[1619] = i[14803];
  assign o[1618] = i[14802];
  assign o[1617] = i[14801];
  assign o[1616] = i[14800];
  assign o[1615] = i[14799];
  assign o[1614] = i[14798];
  assign o[1613] = i[14797];
  assign o[1612] = i[14796];
  assign o[1611] = i[14795];
  assign o[1610] = i[14794];
  assign o[1609] = i[14793];
  assign o[1608] = i[14792];
  assign o[1607] = i[14791];
  assign o[1606] = i[14790];
  assign o[1605] = i[14789];
  assign o[1604] = i[14788];
  assign o[1603] = i[14787];
  assign o[1602] = i[14786];
  assign o[1601] = i[14785];
  assign o[1600] = i[14784];
  assign o[1599] = i[14783];
  assign o[1598] = i[14782];
  assign o[1597] = i[14781];
  assign o[1596] = i[14780];
  assign o[1595] = i[14779];
  assign o[1594] = i[14778];
  assign o[1593] = i[14777];
  assign o[1592] = i[14776];
  assign o[1591] = i[14775];
  assign o[1590] = i[14774];
  assign o[1589] = i[14773];
  assign o[1588] = i[14772];
  assign o[1587] = i[14771];
  assign o[1586] = i[14770];
  assign o[1585] = i[14769];
  assign o[1584] = i[14768];
  assign o[1583] = i[14767];
  assign o[1582] = i[14766];
  assign o[1581] = i[14765];
  assign o[1580] = i[14764];
  assign o[1579] = i[14763];
  assign o[1578] = i[14762];
  assign o[1577] = i[14761];
  assign o[1576] = i[14760];
  assign o[1575] = i[14759];
  assign o[1574] = i[14758];
  assign o[1573] = i[14757];
  assign o[1572] = i[14756];
  assign o[1571] = i[14755];
  assign o[1570] = i[14754];
  assign o[1569] = i[14753];
  assign o[1568] = i[14752];
  assign o[1567] = i[14751];
  assign o[1566] = i[14750];
  assign o[1565] = i[14749];
  assign o[1564] = i[14748];
  assign o[1563] = i[14747];
  assign o[1562] = i[14746];
  assign o[1561] = i[14745];
  assign o[1560] = i[14744];
  assign o[1559] = i[14743];
  assign o[1558] = i[14742];
  assign o[1557] = i[14741];
  assign o[1556] = i[14740];
  assign o[1555] = i[14739];
  assign o[1554] = i[14738];
  assign o[1553] = i[14737];
  assign o[1552] = i[14736];
  assign o[1551] = i[14735];
  assign o[1550] = i[14734];
  assign o[1549] = i[14733];
  assign o[1548] = i[14732];
  assign o[1547] = i[14731];
  assign o[1546] = i[14730];
  assign o[1545] = i[14729];
  assign o[1544] = i[14728];
  assign o[1543] = i[14727];
  assign o[1542] = i[14726];
  assign o[1541] = i[14725];
  assign o[1540] = i[14724];
  assign o[1539] = i[14723];
  assign o[1538] = i[14722];
  assign o[1537] = i[14721];
  assign o[1536] = i[14720];
  assign o[1535] = i[14975];
  assign o[1534] = i[14974];
  assign o[1533] = i[14973];
  assign o[1532] = i[14972];
  assign o[1531] = i[14971];
  assign o[1530] = i[14970];
  assign o[1529] = i[14969];
  assign o[1528] = i[14968];
  assign o[1527] = i[14967];
  assign o[1526] = i[14966];
  assign o[1525] = i[14965];
  assign o[1524] = i[14964];
  assign o[1523] = i[14963];
  assign o[1522] = i[14962];
  assign o[1521] = i[14961];
  assign o[1520] = i[14960];
  assign o[1519] = i[14959];
  assign o[1518] = i[14958];
  assign o[1517] = i[14957];
  assign o[1516] = i[14956];
  assign o[1515] = i[14955];
  assign o[1514] = i[14954];
  assign o[1513] = i[14953];
  assign o[1512] = i[14952];
  assign o[1511] = i[14951];
  assign o[1510] = i[14950];
  assign o[1509] = i[14949];
  assign o[1508] = i[14948];
  assign o[1507] = i[14947];
  assign o[1506] = i[14946];
  assign o[1505] = i[14945];
  assign o[1504] = i[14944];
  assign o[1503] = i[14943];
  assign o[1502] = i[14942];
  assign o[1501] = i[14941];
  assign o[1500] = i[14940];
  assign o[1499] = i[14939];
  assign o[1498] = i[14938];
  assign o[1497] = i[14937];
  assign o[1496] = i[14936];
  assign o[1495] = i[14935];
  assign o[1494] = i[14934];
  assign o[1493] = i[14933];
  assign o[1492] = i[14932];
  assign o[1491] = i[14931];
  assign o[1490] = i[14930];
  assign o[1489] = i[14929];
  assign o[1488] = i[14928];
  assign o[1487] = i[14927];
  assign o[1486] = i[14926];
  assign o[1485] = i[14925];
  assign o[1484] = i[14924];
  assign o[1483] = i[14923];
  assign o[1482] = i[14922];
  assign o[1481] = i[14921];
  assign o[1480] = i[14920];
  assign o[1479] = i[14919];
  assign o[1478] = i[14918];
  assign o[1477] = i[14917];
  assign o[1476] = i[14916];
  assign o[1475] = i[14915];
  assign o[1474] = i[14914];
  assign o[1473] = i[14913];
  assign o[1472] = i[14912];
  assign o[1471] = i[14911];
  assign o[1470] = i[14910];
  assign o[1469] = i[14909];
  assign o[1468] = i[14908];
  assign o[1467] = i[14907];
  assign o[1466] = i[14906];
  assign o[1465] = i[14905];
  assign o[1464] = i[14904];
  assign o[1463] = i[14903];
  assign o[1462] = i[14902];
  assign o[1461] = i[14901];
  assign o[1460] = i[14900];
  assign o[1459] = i[14899];
  assign o[1458] = i[14898];
  assign o[1457] = i[14897];
  assign o[1456] = i[14896];
  assign o[1455] = i[14895];
  assign o[1454] = i[14894];
  assign o[1453] = i[14893];
  assign o[1452] = i[14892];
  assign o[1451] = i[14891];
  assign o[1450] = i[14890];
  assign o[1449] = i[14889];
  assign o[1448] = i[14888];
  assign o[1447] = i[14887];
  assign o[1446] = i[14886];
  assign o[1445] = i[14885];
  assign o[1444] = i[14884];
  assign o[1443] = i[14883];
  assign o[1442] = i[14882];
  assign o[1441] = i[14881];
  assign o[1440] = i[14880];
  assign o[1439] = i[14879];
  assign o[1438] = i[14878];
  assign o[1437] = i[14877];
  assign o[1436] = i[14876];
  assign o[1435] = i[14875];
  assign o[1434] = i[14874];
  assign o[1433] = i[14873];
  assign o[1432] = i[14872];
  assign o[1431] = i[14871];
  assign o[1430] = i[14870];
  assign o[1429] = i[14869];
  assign o[1428] = i[14868];
  assign o[1427] = i[14867];
  assign o[1426] = i[14866];
  assign o[1425] = i[14865];
  assign o[1424] = i[14864];
  assign o[1423] = i[14863];
  assign o[1422] = i[14862];
  assign o[1421] = i[14861];
  assign o[1420] = i[14860];
  assign o[1419] = i[14859];
  assign o[1418] = i[14858];
  assign o[1417] = i[14857];
  assign o[1416] = i[14856];
  assign o[1415] = i[14855];
  assign o[1414] = i[14854];
  assign o[1413] = i[14853];
  assign o[1412] = i[14852];
  assign o[1411] = i[14851];
  assign o[1410] = i[14850];
  assign o[1409] = i[14849];
  assign o[1408] = i[14848];
  assign o[1407] = i[15103];
  assign o[1406] = i[15102];
  assign o[1405] = i[15101];
  assign o[1404] = i[15100];
  assign o[1403] = i[15099];
  assign o[1402] = i[15098];
  assign o[1401] = i[15097];
  assign o[1400] = i[15096];
  assign o[1399] = i[15095];
  assign o[1398] = i[15094];
  assign o[1397] = i[15093];
  assign o[1396] = i[15092];
  assign o[1395] = i[15091];
  assign o[1394] = i[15090];
  assign o[1393] = i[15089];
  assign o[1392] = i[15088];
  assign o[1391] = i[15087];
  assign o[1390] = i[15086];
  assign o[1389] = i[15085];
  assign o[1388] = i[15084];
  assign o[1387] = i[15083];
  assign o[1386] = i[15082];
  assign o[1385] = i[15081];
  assign o[1384] = i[15080];
  assign o[1383] = i[15079];
  assign o[1382] = i[15078];
  assign o[1381] = i[15077];
  assign o[1380] = i[15076];
  assign o[1379] = i[15075];
  assign o[1378] = i[15074];
  assign o[1377] = i[15073];
  assign o[1376] = i[15072];
  assign o[1375] = i[15071];
  assign o[1374] = i[15070];
  assign o[1373] = i[15069];
  assign o[1372] = i[15068];
  assign o[1371] = i[15067];
  assign o[1370] = i[15066];
  assign o[1369] = i[15065];
  assign o[1368] = i[15064];
  assign o[1367] = i[15063];
  assign o[1366] = i[15062];
  assign o[1365] = i[15061];
  assign o[1364] = i[15060];
  assign o[1363] = i[15059];
  assign o[1362] = i[15058];
  assign o[1361] = i[15057];
  assign o[1360] = i[15056];
  assign o[1359] = i[15055];
  assign o[1358] = i[15054];
  assign o[1357] = i[15053];
  assign o[1356] = i[15052];
  assign o[1355] = i[15051];
  assign o[1354] = i[15050];
  assign o[1353] = i[15049];
  assign o[1352] = i[15048];
  assign o[1351] = i[15047];
  assign o[1350] = i[15046];
  assign o[1349] = i[15045];
  assign o[1348] = i[15044];
  assign o[1347] = i[15043];
  assign o[1346] = i[15042];
  assign o[1345] = i[15041];
  assign o[1344] = i[15040];
  assign o[1343] = i[15039];
  assign o[1342] = i[15038];
  assign o[1341] = i[15037];
  assign o[1340] = i[15036];
  assign o[1339] = i[15035];
  assign o[1338] = i[15034];
  assign o[1337] = i[15033];
  assign o[1336] = i[15032];
  assign o[1335] = i[15031];
  assign o[1334] = i[15030];
  assign o[1333] = i[15029];
  assign o[1332] = i[15028];
  assign o[1331] = i[15027];
  assign o[1330] = i[15026];
  assign o[1329] = i[15025];
  assign o[1328] = i[15024];
  assign o[1327] = i[15023];
  assign o[1326] = i[15022];
  assign o[1325] = i[15021];
  assign o[1324] = i[15020];
  assign o[1323] = i[15019];
  assign o[1322] = i[15018];
  assign o[1321] = i[15017];
  assign o[1320] = i[15016];
  assign o[1319] = i[15015];
  assign o[1318] = i[15014];
  assign o[1317] = i[15013];
  assign o[1316] = i[15012];
  assign o[1315] = i[15011];
  assign o[1314] = i[15010];
  assign o[1313] = i[15009];
  assign o[1312] = i[15008];
  assign o[1311] = i[15007];
  assign o[1310] = i[15006];
  assign o[1309] = i[15005];
  assign o[1308] = i[15004];
  assign o[1307] = i[15003];
  assign o[1306] = i[15002];
  assign o[1305] = i[15001];
  assign o[1304] = i[15000];
  assign o[1303] = i[14999];
  assign o[1302] = i[14998];
  assign o[1301] = i[14997];
  assign o[1300] = i[14996];
  assign o[1299] = i[14995];
  assign o[1298] = i[14994];
  assign o[1297] = i[14993];
  assign o[1296] = i[14992];
  assign o[1295] = i[14991];
  assign o[1294] = i[14990];
  assign o[1293] = i[14989];
  assign o[1292] = i[14988];
  assign o[1291] = i[14987];
  assign o[1290] = i[14986];
  assign o[1289] = i[14985];
  assign o[1288] = i[14984];
  assign o[1287] = i[14983];
  assign o[1286] = i[14982];
  assign o[1285] = i[14981];
  assign o[1284] = i[14980];
  assign o[1283] = i[14979];
  assign o[1282] = i[14978];
  assign o[1281] = i[14977];
  assign o[1280] = i[14976];
  assign o[1279] = i[15231];
  assign o[1278] = i[15230];
  assign o[1277] = i[15229];
  assign o[1276] = i[15228];
  assign o[1275] = i[15227];
  assign o[1274] = i[15226];
  assign o[1273] = i[15225];
  assign o[1272] = i[15224];
  assign o[1271] = i[15223];
  assign o[1270] = i[15222];
  assign o[1269] = i[15221];
  assign o[1268] = i[15220];
  assign o[1267] = i[15219];
  assign o[1266] = i[15218];
  assign o[1265] = i[15217];
  assign o[1264] = i[15216];
  assign o[1263] = i[15215];
  assign o[1262] = i[15214];
  assign o[1261] = i[15213];
  assign o[1260] = i[15212];
  assign o[1259] = i[15211];
  assign o[1258] = i[15210];
  assign o[1257] = i[15209];
  assign o[1256] = i[15208];
  assign o[1255] = i[15207];
  assign o[1254] = i[15206];
  assign o[1253] = i[15205];
  assign o[1252] = i[15204];
  assign o[1251] = i[15203];
  assign o[1250] = i[15202];
  assign o[1249] = i[15201];
  assign o[1248] = i[15200];
  assign o[1247] = i[15199];
  assign o[1246] = i[15198];
  assign o[1245] = i[15197];
  assign o[1244] = i[15196];
  assign o[1243] = i[15195];
  assign o[1242] = i[15194];
  assign o[1241] = i[15193];
  assign o[1240] = i[15192];
  assign o[1239] = i[15191];
  assign o[1238] = i[15190];
  assign o[1237] = i[15189];
  assign o[1236] = i[15188];
  assign o[1235] = i[15187];
  assign o[1234] = i[15186];
  assign o[1233] = i[15185];
  assign o[1232] = i[15184];
  assign o[1231] = i[15183];
  assign o[1230] = i[15182];
  assign o[1229] = i[15181];
  assign o[1228] = i[15180];
  assign o[1227] = i[15179];
  assign o[1226] = i[15178];
  assign o[1225] = i[15177];
  assign o[1224] = i[15176];
  assign o[1223] = i[15175];
  assign o[1222] = i[15174];
  assign o[1221] = i[15173];
  assign o[1220] = i[15172];
  assign o[1219] = i[15171];
  assign o[1218] = i[15170];
  assign o[1217] = i[15169];
  assign o[1216] = i[15168];
  assign o[1215] = i[15167];
  assign o[1214] = i[15166];
  assign o[1213] = i[15165];
  assign o[1212] = i[15164];
  assign o[1211] = i[15163];
  assign o[1210] = i[15162];
  assign o[1209] = i[15161];
  assign o[1208] = i[15160];
  assign o[1207] = i[15159];
  assign o[1206] = i[15158];
  assign o[1205] = i[15157];
  assign o[1204] = i[15156];
  assign o[1203] = i[15155];
  assign o[1202] = i[15154];
  assign o[1201] = i[15153];
  assign o[1200] = i[15152];
  assign o[1199] = i[15151];
  assign o[1198] = i[15150];
  assign o[1197] = i[15149];
  assign o[1196] = i[15148];
  assign o[1195] = i[15147];
  assign o[1194] = i[15146];
  assign o[1193] = i[15145];
  assign o[1192] = i[15144];
  assign o[1191] = i[15143];
  assign o[1190] = i[15142];
  assign o[1189] = i[15141];
  assign o[1188] = i[15140];
  assign o[1187] = i[15139];
  assign o[1186] = i[15138];
  assign o[1185] = i[15137];
  assign o[1184] = i[15136];
  assign o[1183] = i[15135];
  assign o[1182] = i[15134];
  assign o[1181] = i[15133];
  assign o[1180] = i[15132];
  assign o[1179] = i[15131];
  assign o[1178] = i[15130];
  assign o[1177] = i[15129];
  assign o[1176] = i[15128];
  assign o[1175] = i[15127];
  assign o[1174] = i[15126];
  assign o[1173] = i[15125];
  assign o[1172] = i[15124];
  assign o[1171] = i[15123];
  assign o[1170] = i[15122];
  assign o[1169] = i[15121];
  assign o[1168] = i[15120];
  assign o[1167] = i[15119];
  assign o[1166] = i[15118];
  assign o[1165] = i[15117];
  assign o[1164] = i[15116];
  assign o[1163] = i[15115];
  assign o[1162] = i[15114];
  assign o[1161] = i[15113];
  assign o[1160] = i[15112];
  assign o[1159] = i[15111];
  assign o[1158] = i[15110];
  assign o[1157] = i[15109];
  assign o[1156] = i[15108];
  assign o[1155] = i[15107];
  assign o[1154] = i[15106];
  assign o[1153] = i[15105];
  assign o[1152] = i[15104];
  assign o[1151] = i[15359];
  assign o[1150] = i[15358];
  assign o[1149] = i[15357];
  assign o[1148] = i[15356];
  assign o[1147] = i[15355];
  assign o[1146] = i[15354];
  assign o[1145] = i[15353];
  assign o[1144] = i[15352];
  assign o[1143] = i[15351];
  assign o[1142] = i[15350];
  assign o[1141] = i[15349];
  assign o[1140] = i[15348];
  assign o[1139] = i[15347];
  assign o[1138] = i[15346];
  assign o[1137] = i[15345];
  assign o[1136] = i[15344];
  assign o[1135] = i[15343];
  assign o[1134] = i[15342];
  assign o[1133] = i[15341];
  assign o[1132] = i[15340];
  assign o[1131] = i[15339];
  assign o[1130] = i[15338];
  assign o[1129] = i[15337];
  assign o[1128] = i[15336];
  assign o[1127] = i[15335];
  assign o[1126] = i[15334];
  assign o[1125] = i[15333];
  assign o[1124] = i[15332];
  assign o[1123] = i[15331];
  assign o[1122] = i[15330];
  assign o[1121] = i[15329];
  assign o[1120] = i[15328];
  assign o[1119] = i[15327];
  assign o[1118] = i[15326];
  assign o[1117] = i[15325];
  assign o[1116] = i[15324];
  assign o[1115] = i[15323];
  assign o[1114] = i[15322];
  assign o[1113] = i[15321];
  assign o[1112] = i[15320];
  assign o[1111] = i[15319];
  assign o[1110] = i[15318];
  assign o[1109] = i[15317];
  assign o[1108] = i[15316];
  assign o[1107] = i[15315];
  assign o[1106] = i[15314];
  assign o[1105] = i[15313];
  assign o[1104] = i[15312];
  assign o[1103] = i[15311];
  assign o[1102] = i[15310];
  assign o[1101] = i[15309];
  assign o[1100] = i[15308];
  assign o[1099] = i[15307];
  assign o[1098] = i[15306];
  assign o[1097] = i[15305];
  assign o[1096] = i[15304];
  assign o[1095] = i[15303];
  assign o[1094] = i[15302];
  assign o[1093] = i[15301];
  assign o[1092] = i[15300];
  assign o[1091] = i[15299];
  assign o[1090] = i[15298];
  assign o[1089] = i[15297];
  assign o[1088] = i[15296];
  assign o[1087] = i[15295];
  assign o[1086] = i[15294];
  assign o[1085] = i[15293];
  assign o[1084] = i[15292];
  assign o[1083] = i[15291];
  assign o[1082] = i[15290];
  assign o[1081] = i[15289];
  assign o[1080] = i[15288];
  assign o[1079] = i[15287];
  assign o[1078] = i[15286];
  assign o[1077] = i[15285];
  assign o[1076] = i[15284];
  assign o[1075] = i[15283];
  assign o[1074] = i[15282];
  assign o[1073] = i[15281];
  assign o[1072] = i[15280];
  assign o[1071] = i[15279];
  assign o[1070] = i[15278];
  assign o[1069] = i[15277];
  assign o[1068] = i[15276];
  assign o[1067] = i[15275];
  assign o[1066] = i[15274];
  assign o[1065] = i[15273];
  assign o[1064] = i[15272];
  assign o[1063] = i[15271];
  assign o[1062] = i[15270];
  assign o[1061] = i[15269];
  assign o[1060] = i[15268];
  assign o[1059] = i[15267];
  assign o[1058] = i[15266];
  assign o[1057] = i[15265];
  assign o[1056] = i[15264];
  assign o[1055] = i[15263];
  assign o[1054] = i[15262];
  assign o[1053] = i[15261];
  assign o[1052] = i[15260];
  assign o[1051] = i[15259];
  assign o[1050] = i[15258];
  assign o[1049] = i[15257];
  assign o[1048] = i[15256];
  assign o[1047] = i[15255];
  assign o[1046] = i[15254];
  assign o[1045] = i[15253];
  assign o[1044] = i[15252];
  assign o[1043] = i[15251];
  assign o[1042] = i[15250];
  assign o[1041] = i[15249];
  assign o[1040] = i[15248];
  assign o[1039] = i[15247];
  assign o[1038] = i[15246];
  assign o[1037] = i[15245];
  assign o[1036] = i[15244];
  assign o[1035] = i[15243];
  assign o[1034] = i[15242];
  assign o[1033] = i[15241];
  assign o[1032] = i[15240];
  assign o[1031] = i[15239];
  assign o[1030] = i[15238];
  assign o[1029] = i[15237];
  assign o[1028] = i[15236];
  assign o[1027] = i[15235];
  assign o[1026] = i[15234];
  assign o[1025] = i[15233];
  assign o[1024] = i[15232];
  assign o[1023] = i[15487];
  assign o[1022] = i[15486];
  assign o[1021] = i[15485];
  assign o[1020] = i[15484];
  assign o[1019] = i[15483];
  assign o[1018] = i[15482];
  assign o[1017] = i[15481];
  assign o[1016] = i[15480];
  assign o[1015] = i[15479];
  assign o[1014] = i[15478];
  assign o[1013] = i[15477];
  assign o[1012] = i[15476];
  assign o[1011] = i[15475];
  assign o[1010] = i[15474];
  assign o[1009] = i[15473];
  assign o[1008] = i[15472];
  assign o[1007] = i[15471];
  assign o[1006] = i[15470];
  assign o[1005] = i[15469];
  assign o[1004] = i[15468];
  assign o[1003] = i[15467];
  assign o[1002] = i[15466];
  assign o[1001] = i[15465];
  assign o[1000] = i[15464];
  assign o[999] = i[15463];
  assign o[998] = i[15462];
  assign o[997] = i[15461];
  assign o[996] = i[15460];
  assign o[995] = i[15459];
  assign o[994] = i[15458];
  assign o[993] = i[15457];
  assign o[992] = i[15456];
  assign o[991] = i[15455];
  assign o[990] = i[15454];
  assign o[989] = i[15453];
  assign o[988] = i[15452];
  assign o[987] = i[15451];
  assign o[986] = i[15450];
  assign o[985] = i[15449];
  assign o[984] = i[15448];
  assign o[983] = i[15447];
  assign o[982] = i[15446];
  assign o[981] = i[15445];
  assign o[980] = i[15444];
  assign o[979] = i[15443];
  assign o[978] = i[15442];
  assign o[977] = i[15441];
  assign o[976] = i[15440];
  assign o[975] = i[15439];
  assign o[974] = i[15438];
  assign o[973] = i[15437];
  assign o[972] = i[15436];
  assign o[971] = i[15435];
  assign o[970] = i[15434];
  assign o[969] = i[15433];
  assign o[968] = i[15432];
  assign o[967] = i[15431];
  assign o[966] = i[15430];
  assign o[965] = i[15429];
  assign o[964] = i[15428];
  assign o[963] = i[15427];
  assign o[962] = i[15426];
  assign o[961] = i[15425];
  assign o[960] = i[15424];
  assign o[959] = i[15423];
  assign o[958] = i[15422];
  assign o[957] = i[15421];
  assign o[956] = i[15420];
  assign o[955] = i[15419];
  assign o[954] = i[15418];
  assign o[953] = i[15417];
  assign o[952] = i[15416];
  assign o[951] = i[15415];
  assign o[950] = i[15414];
  assign o[949] = i[15413];
  assign o[948] = i[15412];
  assign o[947] = i[15411];
  assign o[946] = i[15410];
  assign o[945] = i[15409];
  assign o[944] = i[15408];
  assign o[943] = i[15407];
  assign o[942] = i[15406];
  assign o[941] = i[15405];
  assign o[940] = i[15404];
  assign o[939] = i[15403];
  assign o[938] = i[15402];
  assign o[937] = i[15401];
  assign o[936] = i[15400];
  assign o[935] = i[15399];
  assign o[934] = i[15398];
  assign o[933] = i[15397];
  assign o[932] = i[15396];
  assign o[931] = i[15395];
  assign o[930] = i[15394];
  assign o[929] = i[15393];
  assign o[928] = i[15392];
  assign o[927] = i[15391];
  assign o[926] = i[15390];
  assign o[925] = i[15389];
  assign o[924] = i[15388];
  assign o[923] = i[15387];
  assign o[922] = i[15386];
  assign o[921] = i[15385];
  assign o[920] = i[15384];
  assign o[919] = i[15383];
  assign o[918] = i[15382];
  assign o[917] = i[15381];
  assign o[916] = i[15380];
  assign o[915] = i[15379];
  assign o[914] = i[15378];
  assign o[913] = i[15377];
  assign o[912] = i[15376];
  assign o[911] = i[15375];
  assign o[910] = i[15374];
  assign o[909] = i[15373];
  assign o[908] = i[15372];
  assign o[907] = i[15371];
  assign o[906] = i[15370];
  assign o[905] = i[15369];
  assign o[904] = i[15368];
  assign o[903] = i[15367];
  assign o[902] = i[15366];
  assign o[901] = i[15365];
  assign o[900] = i[15364];
  assign o[899] = i[15363];
  assign o[898] = i[15362];
  assign o[897] = i[15361];
  assign o[896] = i[15360];
  assign o[895] = i[15615];
  assign o[894] = i[15614];
  assign o[893] = i[15613];
  assign o[892] = i[15612];
  assign o[891] = i[15611];
  assign o[890] = i[15610];
  assign o[889] = i[15609];
  assign o[888] = i[15608];
  assign o[887] = i[15607];
  assign o[886] = i[15606];
  assign o[885] = i[15605];
  assign o[884] = i[15604];
  assign o[883] = i[15603];
  assign o[882] = i[15602];
  assign o[881] = i[15601];
  assign o[880] = i[15600];
  assign o[879] = i[15599];
  assign o[878] = i[15598];
  assign o[877] = i[15597];
  assign o[876] = i[15596];
  assign o[875] = i[15595];
  assign o[874] = i[15594];
  assign o[873] = i[15593];
  assign o[872] = i[15592];
  assign o[871] = i[15591];
  assign o[870] = i[15590];
  assign o[869] = i[15589];
  assign o[868] = i[15588];
  assign o[867] = i[15587];
  assign o[866] = i[15586];
  assign o[865] = i[15585];
  assign o[864] = i[15584];
  assign o[863] = i[15583];
  assign o[862] = i[15582];
  assign o[861] = i[15581];
  assign o[860] = i[15580];
  assign o[859] = i[15579];
  assign o[858] = i[15578];
  assign o[857] = i[15577];
  assign o[856] = i[15576];
  assign o[855] = i[15575];
  assign o[854] = i[15574];
  assign o[853] = i[15573];
  assign o[852] = i[15572];
  assign o[851] = i[15571];
  assign o[850] = i[15570];
  assign o[849] = i[15569];
  assign o[848] = i[15568];
  assign o[847] = i[15567];
  assign o[846] = i[15566];
  assign o[845] = i[15565];
  assign o[844] = i[15564];
  assign o[843] = i[15563];
  assign o[842] = i[15562];
  assign o[841] = i[15561];
  assign o[840] = i[15560];
  assign o[839] = i[15559];
  assign o[838] = i[15558];
  assign o[837] = i[15557];
  assign o[836] = i[15556];
  assign o[835] = i[15555];
  assign o[834] = i[15554];
  assign o[833] = i[15553];
  assign o[832] = i[15552];
  assign o[831] = i[15551];
  assign o[830] = i[15550];
  assign o[829] = i[15549];
  assign o[828] = i[15548];
  assign o[827] = i[15547];
  assign o[826] = i[15546];
  assign o[825] = i[15545];
  assign o[824] = i[15544];
  assign o[823] = i[15543];
  assign o[822] = i[15542];
  assign o[821] = i[15541];
  assign o[820] = i[15540];
  assign o[819] = i[15539];
  assign o[818] = i[15538];
  assign o[817] = i[15537];
  assign o[816] = i[15536];
  assign o[815] = i[15535];
  assign o[814] = i[15534];
  assign o[813] = i[15533];
  assign o[812] = i[15532];
  assign o[811] = i[15531];
  assign o[810] = i[15530];
  assign o[809] = i[15529];
  assign o[808] = i[15528];
  assign o[807] = i[15527];
  assign o[806] = i[15526];
  assign o[805] = i[15525];
  assign o[804] = i[15524];
  assign o[803] = i[15523];
  assign o[802] = i[15522];
  assign o[801] = i[15521];
  assign o[800] = i[15520];
  assign o[799] = i[15519];
  assign o[798] = i[15518];
  assign o[797] = i[15517];
  assign o[796] = i[15516];
  assign o[795] = i[15515];
  assign o[794] = i[15514];
  assign o[793] = i[15513];
  assign o[792] = i[15512];
  assign o[791] = i[15511];
  assign o[790] = i[15510];
  assign o[789] = i[15509];
  assign o[788] = i[15508];
  assign o[787] = i[15507];
  assign o[786] = i[15506];
  assign o[785] = i[15505];
  assign o[784] = i[15504];
  assign o[783] = i[15503];
  assign o[782] = i[15502];
  assign o[781] = i[15501];
  assign o[780] = i[15500];
  assign o[779] = i[15499];
  assign o[778] = i[15498];
  assign o[777] = i[15497];
  assign o[776] = i[15496];
  assign o[775] = i[15495];
  assign o[774] = i[15494];
  assign o[773] = i[15493];
  assign o[772] = i[15492];
  assign o[771] = i[15491];
  assign o[770] = i[15490];
  assign o[769] = i[15489];
  assign o[768] = i[15488];
  assign o[767] = i[15743];
  assign o[766] = i[15742];
  assign o[765] = i[15741];
  assign o[764] = i[15740];
  assign o[763] = i[15739];
  assign o[762] = i[15738];
  assign o[761] = i[15737];
  assign o[760] = i[15736];
  assign o[759] = i[15735];
  assign o[758] = i[15734];
  assign o[757] = i[15733];
  assign o[756] = i[15732];
  assign o[755] = i[15731];
  assign o[754] = i[15730];
  assign o[753] = i[15729];
  assign o[752] = i[15728];
  assign o[751] = i[15727];
  assign o[750] = i[15726];
  assign o[749] = i[15725];
  assign o[748] = i[15724];
  assign o[747] = i[15723];
  assign o[746] = i[15722];
  assign o[745] = i[15721];
  assign o[744] = i[15720];
  assign o[743] = i[15719];
  assign o[742] = i[15718];
  assign o[741] = i[15717];
  assign o[740] = i[15716];
  assign o[739] = i[15715];
  assign o[738] = i[15714];
  assign o[737] = i[15713];
  assign o[736] = i[15712];
  assign o[735] = i[15711];
  assign o[734] = i[15710];
  assign o[733] = i[15709];
  assign o[732] = i[15708];
  assign o[731] = i[15707];
  assign o[730] = i[15706];
  assign o[729] = i[15705];
  assign o[728] = i[15704];
  assign o[727] = i[15703];
  assign o[726] = i[15702];
  assign o[725] = i[15701];
  assign o[724] = i[15700];
  assign o[723] = i[15699];
  assign o[722] = i[15698];
  assign o[721] = i[15697];
  assign o[720] = i[15696];
  assign o[719] = i[15695];
  assign o[718] = i[15694];
  assign o[717] = i[15693];
  assign o[716] = i[15692];
  assign o[715] = i[15691];
  assign o[714] = i[15690];
  assign o[713] = i[15689];
  assign o[712] = i[15688];
  assign o[711] = i[15687];
  assign o[710] = i[15686];
  assign o[709] = i[15685];
  assign o[708] = i[15684];
  assign o[707] = i[15683];
  assign o[706] = i[15682];
  assign o[705] = i[15681];
  assign o[704] = i[15680];
  assign o[703] = i[15679];
  assign o[702] = i[15678];
  assign o[701] = i[15677];
  assign o[700] = i[15676];
  assign o[699] = i[15675];
  assign o[698] = i[15674];
  assign o[697] = i[15673];
  assign o[696] = i[15672];
  assign o[695] = i[15671];
  assign o[694] = i[15670];
  assign o[693] = i[15669];
  assign o[692] = i[15668];
  assign o[691] = i[15667];
  assign o[690] = i[15666];
  assign o[689] = i[15665];
  assign o[688] = i[15664];
  assign o[687] = i[15663];
  assign o[686] = i[15662];
  assign o[685] = i[15661];
  assign o[684] = i[15660];
  assign o[683] = i[15659];
  assign o[682] = i[15658];
  assign o[681] = i[15657];
  assign o[680] = i[15656];
  assign o[679] = i[15655];
  assign o[678] = i[15654];
  assign o[677] = i[15653];
  assign o[676] = i[15652];
  assign o[675] = i[15651];
  assign o[674] = i[15650];
  assign o[673] = i[15649];
  assign o[672] = i[15648];
  assign o[671] = i[15647];
  assign o[670] = i[15646];
  assign o[669] = i[15645];
  assign o[668] = i[15644];
  assign o[667] = i[15643];
  assign o[666] = i[15642];
  assign o[665] = i[15641];
  assign o[664] = i[15640];
  assign o[663] = i[15639];
  assign o[662] = i[15638];
  assign o[661] = i[15637];
  assign o[660] = i[15636];
  assign o[659] = i[15635];
  assign o[658] = i[15634];
  assign o[657] = i[15633];
  assign o[656] = i[15632];
  assign o[655] = i[15631];
  assign o[654] = i[15630];
  assign o[653] = i[15629];
  assign o[652] = i[15628];
  assign o[651] = i[15627];
  assign o[650] = i[15626];
  assign o[649] = i[15625];
  assign o[648] = i[15624];
  assign o[647] = i[15623];
  assign o[646] = i[15622];
  assign o[645] = i[15621];
  assign o[644] = i[15620];
  assign o[643] = i[15619];
  assign o[642] = i[15618];
  assign o[641] = i[15617];
  assign o[640] = i[15616];
  assign o[639] = i[15871];
  assign o[638] = i[15870];
  assign o[637] = i[15869];
  assign o[636] = i[15868];
  assign o[635] = i[15867];
  assign o[634] = i[15866];
  assign o[633] = i[15865];
  assign o[632] = i[15864];
  assign o[631] = i[15863];
  assign o[630] = i[15862];
  assign o[629] = i[15861];
  assign o[628] = i[15860];
  assign o[627] = i[15859];
  assign o[626] = i[15858];
  assign o[625] = i[15857];
  assign o[624] = i[15856];
  assign o[623] = i[15855];
  assign o[622] = i[15854];
  assign o[621] = i[15853];
  assign o[620] = i[15852];
  assign o[619] = i[15851];
  assign o[618] = i[15850];
  assign o[617] = i[15849];
  assign o[616] = i[15848];
  assign o[615] = i[15847];
  assign o[614] = i[15846];
  assign o[613] = i[15845];
  assign o[612] = i[15844];
  assign o[611] = i[15843];
  assign o[610] = i[15842];
  assign o[609] = i[15841];
  assign o[608] = i[15840];
  assign o[607] = i[15839];
  assign o[606] = i[15838];
  assign o[605] = i[15837];
  assign o[604] = i[15836];
  assign o[603] = i[15835];
  assign o[602] = i[15834];
  assign o[601] = i[15833];
  assign o[600] = i[15832];
  assign o[599] = i[15831];
  assign o[598] = i[15830];
  assign o[597] = i[15829];
  assign o[596] = i[15828];
  assign o[595] = i[15827];
  assign o[594] = i[15826];
  assign o[593] = i[15825];
  assign o[592] = i[15824];
  assign o[591] = i[15823];
  assign o[590] = i[15822];
  assign o[589] = i[15821];
  assign o[588] = i[15820];
  assign o[587] = i[15819];
  assign o[586] = i[15818];
  assign o[585] = i[15817];
  assign o[584] = i[15816];
  assign o[583] = i[15815];
  assign o[582] = i[15814];
  assign o[581] = i[15813];
  assign o[580] = i[15812];
  assign o[579] = i[15811];
  assign o[578] = i[15810];
  assign o[577] = i[15809];
  assign o[576] = i[15808];
  assign o[575] = i[15807];
  assign o[574] = i[15806];
  assign o[573] = i[15805];
  assign o[572] = i[15804];
  assign o[571] = i[15803];
  assign o[570] = i[15802];
  assign o[569] = i[15801];
  assign o[568] = i[15800];
  assign o[567] = i[15799];
  assign o[566] = i[15798];
  assign o[565] = i[15797];
  assign o[564] = i[15796];
  assign o[563] = i[15795];
  assign o[562] = i[15794];
  assign o[561] = i[15793];
  assign o[560] = i[15792];
  assign o[559] = i[15791];
  assign o[558] = i[15790];
  assign o[557] = i[15789];
  assign o[556] = i[15788];
  assign o[555] = i[15787];
  assign o[554] = i[15786];
  assign o[553] = i[15785];
  assign o[552] = i[15784];
  assign o[551] = i[15783];
  assign o[550] = i[15782];
  assign o[549] = i[15781];
  assign o[548] = i[15780];
  assign o[547] = i[15779];
  assign o[546] = i[15778];
  assign o[545] = i[15777];
  assign o[544] = i[15776];
  assign o[543] = i[15775];
  assign o[542] = i[15774];
  assign o[541] = i[15773];
  assign o[540] = i[15772];
  assign o[539] = i[15771];
  assign o[538] = i[15770];
  assign o[537] = i[15769];
  assign o[536] = i[15768];
  assign o[535] = i[15767];
  assign o[534] = i[15766];
  assign o[533] = i[15765];
  assign o[532] = i[15764];
  assign o[531] = i[15763];
  assign o[530] = i[15762];
  assign o[529] = i[15761];
  assign o[528] = i[15760];
  assign o[527] = i[15759];
  assign o[526] = i[15758];
  assign o[525] = i[15757];
  assign o[524] = i[15756];
  assign o[523] = i[15755];
  assign o[522] = i[15754];
  assign o[521] = i[15753];
  assign o[520] = i[15752];
  assign o[519] = i[15751];
  assign o[518] = i[15750];
  assign o[517] = i[15749];
  assign o[516] = i[15748];
  assign o[515] = i[15747];
  assign o[514] = i[15746];
  assign o[513] = i[15745];
  assign o[512] = i[15744];
  assign o[511] = i[15999];
  assign o[510] = i[15998];
  assign o[509] = i[15997];
  assign o[508] = i[15996];
  assign o[507] = i[15995];
  assign o[506] = i[15994];
  assign o[505] = i[15993];
  assign o[504] = i[15992];
  assign o[503] = i[15991];
  assign o[502] = i[15990];
  assign o[501] = i[15989];
  assign o[500] = i[15988];
  assign o[499] = i[15987];
  assign o[498] = i[15986];
  assign o[497] = i[15985];
  assign o[496] = i[15984];
  assign o[495] = i[15983];
  assign o[494] = i[15982];
  assign o[493] = i[15981];
  assign o[492] = i[15980];
  assign o[491] = i[15979];
  assign o[490] = i[15978];
  assign o[489] = i[15977];
  assign o[488] = i[15976];
  assign o[487] = i[15975];
  assign o[486] = i[15974];
  assign o[485] = i[15973];
  assign o[484] = i[15972];
  assign o[483] = i[15971];
  assign o[482] = i[15970];
  assign o[481] = i[15969];
  assign o[480] = i[15968];
  assign o[479] = i[15967];
  assign o[478] = i[15966];
  assign o[477] = i[15965];
  assign o[476] = i[15964];
  assign o[475] = i[15963];
  assign o[474] = i[15962];
  assign o[473] = i[15961];
  assign o[472] = i[15960];
  assign o[471] = i[15959];
  assign o[470] = i[15958];
  assign o[469] = i[15957];
  assign o[468] = i[15956];
  assign o[467] = i[15955];
  assign o[466] = i[15954];
  assign o[465] = i[15953];
  assign o[464] = i[15952];
  assign o[463] = i[15951];
  assign o[462] = i[15950];
  assign o[461] = i[15949];
  assign o[460] = i[15948];
  assign o[459] = i[15947];
  assign o[458] = i[15946];
  assign o[457] = i[15945];
  assign o[456] = i[15944];
  assign o[455] = i[15943];
  assign o[454] = i[15942];
  assign o[453] = i[15941];
  assign o[452] = i[15940];
  assign o[451] = i[15939];
  assign o[450] = i[15938];
  assign o[449] = i[15937];
  assign o[448] = i[15936];
  assign o[447] = i[15935];
  assign o[446] = i[15934];
  assign o[445] = i[15933];
  assign o[444] = i[15932];
  assign o[443] = i[15931];
  assign o[442] = i[15930];
  assign o[441] = i[15929];
  assign o[440] = i[15928];
  assign o[439] = i[15927];
  assign o[438] = i[15926];
  assign o[437] = i[15925];
  assign o[436] = i[15924];
  assign o[435] = i[15923];
  assign o[434] = i[15922];
  assign o[433] = i[15921];
  assign o[432] = i[15920];
  assign o[431] = i[15919];
  assign o[430] = i[15918];
  assign o[429] = i[15917];
  assign o[428] = i[15916];
  assign o[427] = i[15915];
  assign o[426] = i[15914];
  assign o[425] = i[15913];
  assign o[424] = i[15912];
  assign o[423] = i[15911];
  assign o[422] = i[15910];
  assign o[421] = i[15909];
  assign o[420] = i[15908];
  assign o[419] = i[15907];
  assign o[418] = i[15906];
  assign o[417] = i[15905];
  assign o[416] = i[15904];
  assign o[415] = i[15903];
  assign o[414] = i[15902];
  assign o[413] = i[15901];
  assign o[412] = i[15900];
  assign o[411] = i[15899];
  assign o[410] = i[15898];
  assign o[409] = i[15897];
  assign o[408] = i[15896];
  assign o[407] = i[15895];
  assign o[406] = i[15894];
  assign o[405] = i[15893];
  assign o[404] = i[15892];
  assign o[403] = i[15891];
  assign o[402] = i[15890];
  assign o[401] = i[15889];
  assign o[400] = i[15888];
  assign o[399] = i[15887];
  assign o[398] = i[15886];
  assign o[397] = i[15885];
  assign o[396] = i[15884];
  assign o[395] = i[15883];
  assign o[394] = i[15882];
  assign o[393] = i[15881];
  assign o[392] = i[15880];
  assign o[391] = i[15879];
  assign o[390] = i[15878];
  assign o[389] = i[15877];
  assign o[388] = i[15876];
  assign o[387] = i[15875];
  assign o[386] = i[15874];
  assign o[385] = i[15873];
  assign o[384] = i[15872];
  assign o[383] = i[16127];
  assign o[382] = i[16126];
  assign o[381] = i[16125];
  assign o[380] = i[16124];
  assign o[379] = i[16123];
  assign o[378] = i[16122];
  assign o[377] = i[16121];
  assign o[376] = i[16120];
  assign o[375] = i[16119];
  assign o[374] = i[16118];
  assign o[373] = i[16117];
  assign o[372] = i[16116];
  assign o[371] = i[16115];
  assign o[370] = i[16114];
  assign o[369] = i[16113];
  assign o[368] = i[16112];
  assign o[367] = i[16111];
  assign o[366] = i[16110];
  assign o[365] = i[16109];
  assign o[364] = i[16108];
  assign o[363] = i[16107];
  assign o[362] = i[16106];
  assign o[361] = i[16105];
  assign o[360] = i[16104];
  assign o[359] = i[16103];
  assign o[358] = i[16102];
  assign o[357] = i[16101];
  assign o[356] = i[16100];
  assign o[355] = i[16099];
  assign o[354] = i[16098];
  assign o[353] = i[16097];
  assign o[352] = i[16096];
  assign o[351] = i[16095];
  assign o[350] = i[16094];
  assign o[349] = i[16093];
  assign o[348] = i[16092];
  assign o[347] = i[16091];
  assign o[346] = i[16090];
  assign o[345] = i[16089];
  assign o[344] = i[16088];
  assign o[343] = i[16087];
  assign o[342] = i[16086];
  assign o[341] = i[16085];
  assign o[340] = i[16084];
  assign o[339] = i[16083];
  assign o[338] = i[16082];
  assign o[337] = i[16081];
  assign o[336] = i[16080];
  assign o[335] = i[16079];
  assign o[334] = i[16078];
  assign o[333] = i[16077];
  assign o[332] = i[16076];
  assign o[331] = i[16075];
  assign o[330] = i[16074];
  assign o[329] = i[16073];
  assign o[328] = i[16072];
  assign o[327] = i[16071];
  assign o[326] = i[16070];
  assign o[325] = i[16069];
  assign o[324] = i[16068];
  assign o[323] = i[16067];
  assign o[322] = i[16066];
  assign o[321] = i[16065];
  assign o[320] = i[16064];
  assign o[319] = i[16063];
  assign o[318] = i[16062];
  assign o[317] = i[16061];
  assign o[316] = i[16060];
  assign o[315] = i[16059];
  assign o[314] = i[16058];
  assign o[313] = i[16057];
  assign o[312] = i[16056];
  assign o[311] = i[16055];
  assign o[310] = i[16054];
  assign o[309] = i[16053];
  assign o[308] = i[16052];
  assign o[307] = i[16051];
  assign o[306] = i[16050];
  assign o[305] = i[16049];
  assign o[304] = i[16048];
  assign o[303] = i[16047];
  assign o[302] = i[16046];
  assign o[301] = i[16045];
  assign o[300] = i[16044];
  assign o[299] = i[16043];
  assign o[298] = i[16042];
  assign o[297] = i[16041];
  assign o[296] = i[16040];
  assign o[295] = i[16039];
  assign o[294] = i[16038];
  assign o[293] = i[16037];
  assign o[292] = i[16036];
  assign o[291] = i[16035];
  assign o[290] = i[16034];
  assign o[289] = i[16033];
  assign o[288] = i[16032];
  assign o[287] = i[16031];
  assign o[286] = i[16030];
  assign o[285] = i[16029];
  assign o[284] = i[16028];
  assign o[283] = i[16027];
  assign o[282] = i[16026];
  assign o[281] = i[16025];
  assign o[280] = i[16024];
  assign o[279] = i[16023];
  assign o[278] = i[16022];
  assign o[277] = i[16021];
  assign o[276] = i[16020];
  assign o[275] = i[16019];
  assign o[274] = i[16018];
  assign o[273] = i[16017];
  assign o[272] = i[16016];
  assign o[271] = i[16015];
  assign o[270] = i[16014];
  assign o[269] = i[16013];
  assign o[268] = i[16012];
  assign o[267] = i[16011];
  assign o[266] = i[16010];
  assign o[265] = i[16009];
  assign o[264] = i[16008];
  assign o[263] = i[16007];
  assign o[262] = i[16006];
  assign o[261] = i[16005];
  assign o[260] = i[16004];
  assign o[259] = i[16003];
  assign o[258] = i[16002];
  assign o[257] = i[16001];
  assign o[256] = i[16000];
  assign o[255] = i[16255];
  assign o[254] = i[16254];
  assign o[253] = i[16253];
  assign o[252] = i[16252];
  assign o[251] = i[16251];
  assign o[250] = i[16250];
  assign o[249] = i[16249];
  assign o[248] = i[16248];
  assign o[247] = i[16247];
  assign o[246] = i[16246];
  assign o[245] = i[16245];
  assign o[244] = i[16244];
  assign o[243] = i[16243];
  assign o[242] = i[16242];
  assign o[241] = i[16241];
  assign o[240] = i[16240];
  assign o[239] = i[16239];
  assign o[238] = i[16238];
  assign o[237] = i[16237];
  assign o[236] = i[16236];
  assign o[235] = i[16235];
  assign o[234] = i[16234];
  assign o[233] = i[16233];
  assign o[232] = i[16232];
  assign o[231] = i[16231];
  assign o[230] = i[16230];
  assign o[229] = i[16229];
  assign o[228] = i[16228];
  assign o[227] = i[16227];
  assign o[226] = i[16226];
  assign o[225] = i[16225];
  assign o[224] = i[16224];
  assign o[223] = i[16223];
  assign o[222] = i[16222];
  assign o[221] = i[16221];
  assign o[220] = i[16220];
  assign o[219] = i[16219];
  assign o[218] = i[16218];
  assign o[217] = i[16217];
  assign o[216] = i[16216];
  assign o[215] = i[16215];
  assign o[214] = i[16214];
  assign o[213] = i[16213];
  assign o[212] = i[16212];
  assign o[211] = i[16211];
  assign o[210] = i[16210];
  assign o[209] = i[16209];
  assign o[208] = i[16208];
  assign o[207] = i[16207];
  assign o[206] = i[16206];
  assign o[205] = i[16205];
  assign o[204] = i[16204];
  assign o[203] = i[16203];
  assign o[202] = i[16202];
  assign o[201] = i[16201];
  assign o[200] = i[16200];
  assign o[199] = i[16199];
  assign o[198] = i[16198];
  assign o[197] = i[16197];
  assign o[196] = i[16196];
  assign o[195] = i[16195];
  assign o[194] = i[16194];
  assign o[193] = i[16193];
  assign o[192] = i[16192];
  assign o[191] = i[16191];
  assign o[190] = i[16190];
  assign o[189] = i[16189];
  assign o[188] = i[16188];
  assign o[187] = i[16187];
  assign o[186] = i[16186];
  assign o[185] = i[16185];
  assign o[184] = i[16184];
  assign o[183] = i[16183];
  assign o[182] = i[16182];
  assign o[181] = i[16181];
  assign o[180] = i[16180];
  assign o[179] = i[16179];
  assign o[178] = i[16178];
  assign o[177] = i[16177];
  assign o[176] = i[16176];
  assign o[175] = i[16175];
  assign o[174] = i[16174];
  assign o[173] = i[16173];
  assign o[172] = i[16172];
  assign o[171] = i[16171];
  assign o[170] = i[16170];
  assign o[169] = i[16169];
  assign o[168] = i[16168];
  assign o[167] = i[16167];
  assign o[166] = i[16166];
  assign o[165] = i[16165];
  assign o[164] = i[16164];
  assign o[163] = i[16163];
  assign o[162] = i[16162];
  assign o[161] = i[16161];
  assign o[160] = i[16160];
  assign o[159] = i[16159];
  assign o[158] = i[16158];
  assign o[157] = i[16157];
  assign o[156] = i[16156];
  assign o[155] = i[16155];
  assign o[154] = i[16154];
  assign o[153] = i[16153];
  assign o[152] = i[16152];
  assign o[151] = i[16151];
  assign o[150] = i[16150];
  assign o[149] = i[16149];
  assign o[148] = i[16148];
  assign o[147] = i[16147];
  assign o[146] = i[16146];
  assign o[145] = i[16145];
  assign o[144] = i[16144];
  assign o[143] = i[16143];
  assign o[142] = i[16142];
  assign o[141] = i[16141];
  assign o[140] = i[16140];
  assign o[139] = i[16139];
  assign o[138] = i[16138];
  assign o[137] = i[16137];
  assign o[136] = i[16136];
  assign o[135] = i[16135];
  assign o[134] = i[16134];
  assign o[133] = i[16133];
  assign o[132] = i[16132];
  assign o[131] = i[16131];
  assign o[130] = i[16130];
  assign o[129] = i[16129];
  assign o[128] = i[16128];
  assign o[127] = i[16383];
  assign o[126] = i[16382];
  assign o[125] = i[16381];
  assign o[124] = i[16380];
  assign o[123] = i[16379];
  assign o[122] = i[16378];
  assign o[121] = i[16377];
  assign o[120] = i[16376];
  assign o[119] = i[16375];
  assign o[118] = i[16374];
  assign o[117] = i[16373];
  assign o[116] = i[16372];
  assign o[115] = i[16371];
  assign o[114] = i[16370];
  assign o[113] = i[16369];
  assign o[112] = i[16368];
  assign o[111] = i[16367];
  assign o[110] = i[16366];
  assign o[109] = i[16365];
  assign o[108] = i[16364];
  assign o[107] = i[16363];
  assign o[106] = i[16362];
  assign o[105] = i[16361];
  assign o[104] = i[16360];
  assign o[103] = i[16359];
  assign o[102] = i[16358];
  assign o[101] = i[16357];
  assign o[100] = i[16356];
  assign o[99] = i[16355];
  assign o[98] = i[16354];
  assign o[97] = i[16353];
  assign o[96] = i[16352];
  assign o[95] = i[16351];
  assign o[94] = i[16350];
  assign o[93] = i[16349];
  assign o[92] = i[16348];
  assign o[91] = i[16347];
  assign o[90] = i[16346];
  assign o[89] = i[16345];
  assign o[88] = i[16344];
  assign o[87] = i[16343];
  assign o[86] = i[16342];
  assign o[85] = i[16341];
  assign o[84] = i[16340];
  assign o[83] = i[16339];
  assign o[82] = i[16338];
  assign o[81] = i[16337];
  assign o[80] = i[16336];
  assign o[79] = i[16335];
  assign o[78] = i[16334];
  assign o[77] = i[16333];
  assign o[76] = i[16332];
  assign o[75] = i[16331];
  assign o[74] = i[16330];
  assign o[73] = i[16329];
  assign o[72] = i[16328];
  assign o[71] = i[16327];
  assign o[70] = i[16326];
  assign o[69] = i[16325];
  assign o[68] = i[16324];
  assign o[67] = i[16323];
  assign o[66] = i[16322];
  assign o[65] = i[16321];
  assign o[64] = i[16320];
  assign o[63] = i[16319];
  assign o[62] = i[16318];
  assign o[61] = i[16317];
  assign o[60] = i[16316];
  assign o[59] = i[16315];
  assign o[58] = i[16314];
  assign o[57] = i[16313];
  assign o[56] = i[16312];
  assign o[55] = i[16311];
  assign o[54] = i[16310];
  assign o[53] = i[16309];
  assign o[52] = i[16308];
  assign o[51] = i[16307];
  assign o[50] = i[16306];
  assign o[49] = i[16305];
  assign o[48] = i[16304];
  assign o[47] = i[16303];
  assign o[46] = i[16302];
  assign o[45] = i[16301];
  assign o[44] = i[16300];
  assign o[43] = i[16299];
  assign o[42] = i[16298];
  assign o[41] = i[16297];
  assign o[40] = i[16296];
  assign o[39] = i[16295];
  assign o[38] = i[16294];
  assign o[37] = i[16293];
  assign o[36] = i[16292];
  assign o[35] = i[16291];
  assign o[34] = i[16290];
  assign o[33] = i[16289];
  assign o[32] = i[16288];
  assign o[31] = i[16287];
  assign o[30] = i[16286];
  assign o[29] = i[16285];
  assign o[28] = i[16284];
  assign o[27] = i[16283];
  assign o[26] = i[16282];
  assign o[25] = i[16281];
  assign o[24] = i[16280];
  assign o[23] = i[16279];
  assign o[22] = i[16278];
  assign o[21] = i[16277];
  assign o[20] = i[16276];
  assign o[19] = i[16275];
  assign o[18] = i[16274];
  assign o[17] = i[16273];
  assign o[16] = i[16272];
  assign o[15] = i[16271];
  assign o[14] = i[16270];
  assign o[13] = i[16269];
  assign o[12] = i[16268];
  assign o[11] = i[16267];
  assign o[10] = i[16266];
  assign o[9] = i[16265];
  assign o[8] = i[16264];
  assign o[7] = i[16263];
  assign o[6] = i[16262];
  assign o[5] = i[16261];
  assign o[4] = i[16260];
  assign o[3] = i[16259];
  assign o[2] = i[16258];
  assign o[1] = i[16257];
  assign o[0] = i[16256];

endmodule

