

module top
(
  i,
  sel_oi_one_hot_i,
  o
);

  input [4095:0] i;
  input [4095:0] sel_oi_one_hot_i;
  output [4095:0] o;

  bsg_crossbar_o_by_i
  wrapper
  (
    .i(i),
    .sel_oi_one_hot_i(sel_oi_one_hot_i),
    .o(o)
  );


endmodule



module bsg_mux_one_hot_width_p64_els_p64
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [4095:0] data_i;
  input [63:0] sel_one_hot_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
  N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,
  N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,
  N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,
  N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,
  N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,
  N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,
  N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,
  N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,
  N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,
  N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,
  N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,
  N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,
  N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,
  N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,
  N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,
  N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,
  N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
  N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,
  N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,
  N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,
  N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,
  N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,
  N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,
  N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,
  N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,
  N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,
  N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,
  N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,
  N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,
  N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,
  N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,
  N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,
  N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,
  N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,
  N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,
  N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,
  N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,
  N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,
  N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,
  N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,
  N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,
  N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,
  N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,
  N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,
  N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,
  N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,
  N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,
  N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,
  N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,
  N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,
  N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,
  N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,
  N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,
  N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,
  N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,
  N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,
  N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,
  N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,
  N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,
  N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,
  N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,
  N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,
  N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,
  N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,
  N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,
  N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,
  N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,
  N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,
  N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,
  N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,
  N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,
  N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,
  N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,
  N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,
  N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,
  N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,
  N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,
  N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,
  N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,
  N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,
  N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,
  N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,
  N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144,
  N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,
  N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,N2170,
  N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,N2184,
  N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197,
  N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,N2210,
  N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,N2224,
  N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,
  N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,
  N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,N2264,
  N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,
  N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290,
  N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302,N2303,N2304,
  N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,
  N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,
  N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,
  N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,
  N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2369,N2370,
  N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382,N2383,N2384,
  N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,N2394,N2395,N2396,N2397,
  N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407,N2408,N2409,N2410,
  N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422,N2423,N2424,
  N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,
  N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447,N2448,N2449,N2450,
  N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,N2460,N2461,N2462,N2463,N2464,
  N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,N2474,N2475,N2476,N2477,
  N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,N2488,N2489,N2490,
  N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,N2500,N2501,N2502,N2503,N2504,
  N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,N2514,N2515,N2516,N2517,
  N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528,N2529,N2530,
  N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539,N2540,N2541,N2542,N2543,N2544,
  N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2554,N2555,N2556,N2557,
  N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,N2567,N2568,N2569,N2570,
  N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579,N2580,N2581,N2582,N2583,N2584,
  N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,N2594,N2595,N2596,N2597,
  N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,N2609,N2610,
  N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,N2620,N2621,N2622,N2623,N2624,
  N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2637,
  N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,N2649,N2650,
  N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662,N2663,N2664,
  N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,
  N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,N2687,N2688,N2689,N2690,
  N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2704,
  N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,N2714,N2715,N2716,N2717,
  N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,N2727,N2728,N2729,N2730,
  N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,
  N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,N2754,N2755,N2756,N2757,
  N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,N2767,N2768,N2769,N2770,
  N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2779,N2780,N2781,N2782,N2783,N2784,
  N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793,N2794,N2795,N2796,N2797,
  N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,N2807,N2808,N2809,N2810,
  N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,N2819,N2820,N2821,N2822,N2823,N2824,
  N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,N2834,N2835,N2836,N2837,
  N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,N2847,N2848,N2849,N2850,
  N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,N2859,N2860,N2861,N2862,N2863,N2864,
  N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877,
  N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,N2887,N2888,N2889,N2890,
  N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,N2899,N2900,N2901,N2902,N2903,N2904,
  N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,N2917,
  N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,N2930,
  N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,N2939,N2940,N2941,N2942,N2943,N2944,
  N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952,N2953,N2954,N2955,N2956,N2957,
  N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2965,N2966,N2967,N2968,N2969,N2970,
  N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980,N2981,N2982,N2983,N2984,
  N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,
  N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,N3010,
  N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022,N3023,N3024,
  N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3036,N3037,
  N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,N3050,
  N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3062,N3063,N3064,
  N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,N3076,N3077,
  N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,N3090,
  N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,N3101,N3102,N3103,N3104,
  N3105,N3106,N3107,N3108,N3109,N3110,N3111,N3112,N3113,N3114,N3115,N3116,N3117,
  N3118,N3119,N3120,N3121,N3122,N3123,N3124,N3125,N3126,N3127,N3128,N3129,N3130,
  N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,N3139,N3140,N3141,N3142,N3143,N3144,
  N3145,N3146,N3147,N3148,N3149,N3150,N3151,N3152,N3153,N3154,N3155,N3156,N3157,
  N3158,N3159,N3160,N3161,N3162,N3163,N3164,N3165,N3166,N3167,N3168,N3169,N3170,
  N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,N3179,N3180,N3181,N3182,N3183,N3184,
  N3185,N3186,N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194,N3195,N3196,N3197,
  N3198,N3199,N3200,N3201,N3202,N3203,N3204,N3205,N3206,N3207,N3208,N3209,N3210,
  N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,N3220,N3221,N3222,N3223,N3224,
  N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,
  N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,N3249,N3250,
  N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,N3260,N3261,N3262,N3263,N3264,
  N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,
  N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,N3290,
  N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,N3300,N3301,N3302,N3303,N3304,
  N3305,N3306,N3307,N3308,N3309,N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,
  N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,N3330,
  N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,N3339,N3340,N3341,N3342,N3343,N3344,
  N3345,N3346,N3347,N3348,N3349,N3350,N3351,N3352,N3353,N3354,N3355,N3356,N3357,
  N3358,N3359,N3360,N3361,N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,N3370,
  N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,N3379,N3380,N3381,N3382,N3383,N3384,
  N3385,N3386,N3387,N3388,N3389,N3390,N3391,N3392,N3393,N3394,N3395,N3396,N3397,
  N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3408,N3409,N3410,
  N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,N3419,N3420,N3421,N3422,N3423,N3424,
  N3425,N3426,N3427,N3428,N3429,N3430,N3431,N3432,N3433,N3434,N3435,N3436,N3437,
  N3438,N3439,N3440,N3441,N3442,N3443,N3444,N3445,N3446,N3447,N3448,N3449,N3450,
  N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,N3459,N3460,N3461,N3462,N3463,N3464,
  N3465,N3466,N3467,N3468,N3469,N3470,N3471,N3472,N3473,N3474,N3475,N3476,N3477,
  N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,N3487,N3488,N3489,N3490,
  N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,N3499,N3500,N3501,N3502,N3503,N3504,
  N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,N3513,N3514,N3515,N3516,N3517,
  N3518,N3519,N3520,N3521,N3522,N3523,N3524,N3525,N3526,N3527,N3528,N3529,N3530,
  N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,N3539,N3540,N3541,N3542,N3543,N3544,
  N3545,N3546,N3547,N3548,N3549,N3550,N3551,N3552,N3553,N3554,N3555,N3556,N3557,
  N3558,N3559,N3560,N3561,N3562,N3563,N3564,N3565,N3566,N3567,N3568,N3569,N3570,
  N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,N3579,N3580,N3581,N3582,N3583,N3584,
  N3585,N3586,N3587,N3588,N3589,N3590,N3591,N3592,N3593,N3594,N3595,N3596,N3597,
  N3598,N3599,N3600,N3601,N3602,N3603,N3604,N3605,N3606,N3607,N3608,N3609,N3610,
  N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,N3619,N3620,N3621,N3622,N3623,N3624,
  N3625,N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3636,N3637,
  N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3646,N3647,N3648,N3649,N3650,
  N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,N3659,N3660,N3661,N3662,N3663,N3664,
  N3665,N3666,N3667,N3668,N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3676,N3677,
  N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685,N3686,N3687,N3688,N3689,N3690,
  N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,N3699,N3700,N3701,N3702,N3703,N3704,
  N3705,N3706,N3707,N3708,N3709,N3710,N3711,N3712,N3713,N3714,N3715,N3716,N3717,
  N3718,N3719,N3720,N3721,N3722,N3723,N3724,N3725,N3726,N3727,N3728,N3729,N3730,
  N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,N3739,N3740,N3741,N3742,N3743,N3744,
  N3745,N3746,N3747,N3748,N3749,N3750,N3751,N3752,N3753,N3754,N3755,N3756,N3757,
  N3758,N3759,N3760,N3761,N3762,N3763,N3764,N3765,N3766,N3767,N3768,N3769,N3770,
  N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,N3779,N3780,N3781,N3782,N3783,N3784,
  N3785,N3786,N3787,N3788,N3789,N3790,N3791,N3792,N3793,N3794,N3795,N3796,N3797,
  N3798,N3799,N3800,N3801,N3802,N3803,N3804,N3805,N3806,N3807,N3808,N3809,N3810,
  N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,N3819,N3820,N3821,N3822,N3823,N3824,
  N3825,N3826,N3827,N3828,N3829,N3830,N3831,N3832,N3833,N3834,N3835,N3836,N3837,
  N3838,N3839,N3840,N3841,N3842,N3843,N3844,N3845,N3846,N3847,N3848,N3849,N3850,
  N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,N3859,N3860,N3861,N3862,N3863,N3864,
  N3865,N3866,N3867,N3868,N3869,N3870,N3871,N3872,N3873,N3874,N3875,N3876,N3877,
  N3878,N3879,N3880,N3881,N3882,N3883,N3884,N3885,N3886,N3887,N3888,N3889,N3890,
  N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,N3899,N3900,N3901,N3902,N3903,N3904,
  N3905,N3906,N3907,N3908,N3909,N3910,N3911,N3912,N3913,N3914,N3915,N3916,N3917,
  N3918,N3919,N3920,N3921,N3922,N3923,N3924,N3925,N3926,N3927,N3928,N3929,N3930,
  N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,N3939,N3940,N3941,N3942,N3943,N3944,
  N3945,N3946,N3947,N3948,N3949,N3950,N3951,N3952,N3953,N3954,N3955,N3956,N3957,
  N3958,N3959,N3960,N3961,N3962,N3963,N3964,N3965,N3966,N3967;
  wire [4095:0] data_masked;
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[1];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[1];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[1];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[1];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[1];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[1];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[1];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[1];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[1];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[1];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[1];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[1];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[1];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[1];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[1];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[1];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[1];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[1];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[1];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[1];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[1];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[1];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[1];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[2];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[2];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[2];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[2];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[2];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[2];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[2];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[2];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[2];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[2];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[2];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[2];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[2];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[2];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[2];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[2];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[2];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[2];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[2];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[2];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[2];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[2];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[2];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[2];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[2];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[2];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[2];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[2];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[2];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[2];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[2];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[2];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[2];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[2];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[2];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[2];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[2];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[2];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[2];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[2];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[2];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[2];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[2];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[2];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[2];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[2];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[2];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[2];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[2];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[2];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[2];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[2];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[2];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[2];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[2];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[2];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[2];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[2];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[2];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[2];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[2];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[2];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[2];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[2];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[3];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[3];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[3];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[3];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[3];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[3];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[3];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[3];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[3];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[3];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[3];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[3];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[3];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[3];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[3];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[3];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[3];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[3];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[3];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[3];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[3];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[3];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[3];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[3];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[3];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[3];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[3];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[3];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[3];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[3];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[3];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[3];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[3];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[3];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[3];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[3];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[3];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[3];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[3];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[3];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[3];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[3];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[3];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[3];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[3];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[3];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[3];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[3];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[3];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[3];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[3];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[3];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[3];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[3];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[3];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[3];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[3];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[3];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[3];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[3];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[3];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[3];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[3];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[3];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[4];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[4];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[4];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[4];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[4];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[4];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[4];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[4];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[4];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[4];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[4];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[4];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[4];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[4];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[4];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[4];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[4];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[4];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[4];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[4];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[4];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[4];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[4];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[4];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[4];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[4];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[4];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[4];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[4];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[4];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[4];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[4];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[4];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[4];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[4];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[4];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[4];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[4];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[4];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[4];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[4];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[4];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[4];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[4];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[4];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[4];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[4];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[4];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[4];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[4];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[4];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[4];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[4];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[4];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[4];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[4];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[4];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[4];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[4];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[4];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[4];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[4];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[4];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[4];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[5];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[5];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[5];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[5];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[5];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[5];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[5];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[5];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[5];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[5];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[5];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[5];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[5];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[5];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[5];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[5];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[5];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[5];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[5];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[5];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[5];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[5];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[5];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[5];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[5];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[5];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[5];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[5];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[5];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[5];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[5];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[5];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[5];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[5];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[5];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[5];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[5];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[5];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[5];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[5];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[5];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[5];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[5];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[5];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[5];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[5];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[5];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[5];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[5];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[5];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[5];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[5];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[5];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[5];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[5];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[5];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[5];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[5];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[5];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[5];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[5];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[5];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[5];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[5];
  assign data_masked[447] = data_i[447] & sel_one_hot_i[6];
  assign data_masked[446] = data_i[446] & sel_one_hot_i[6];
  assign data_masked[445] = data_i[445] & sel_one_hot_i[6];
  assign data_masked[444] = data_i[444] & sel_one_hot_i[6];
  assign data_masked[443] = data_i[443] & sel_one_hot_i[6];
  assign data_masked[442] = data_i[442] & sel_one_hot_i[6];
  assign data_masked[441] = data_i[441] & sel_one_hot_i[6];
  assign data_masked[440] = data_i[440] & sel_one_hot_i[6];
  assign data_masked[439] = data_i[439] & sel_one_hot_i[6];
  assign data_masked[438] = data_i[438] & sel_one_hot_i[6];
  assign data_masked[437] = data_i[437] & sel_one_hot_i[6];
  assign data_masked[436] = data_i[436] & sel_one_hot_i[6];
  assign data_masked[435] = data_i[435] & sel_one_hot_i[6];
  assign data_masked[434] = data_i[434] & sel_one_hot_i[6];
  assign data_masked[433] = data_i[433] & sel_one_hot_i[6];
  assign data_masked[432] = data_i[432] & sel_one_hot_i[6];
  assign data_masked[431] = data_i[431] & sel_one_hot_i[6];
  assign data_masked[430] = data_i[430] & sel_one_hot_i[6];
  assign data_masked[429] = data_i[429] & sel_one_hot_i[6];
  assign data_masked[428] = data_i[428] & sel_one_hot_i[6];
  assign data_masked[427] = data_i[427] & sel_one_hot_i[6];
  assign data_masked[426] = data_i[426] & sel_one_hot_i[6];
  assign data_masked[425] = data_i[425] & sel_one_hot_i[6];
  assign data_masked[424] = data_i[424] & sel_one_hot_i[6];
  assign data_masked[423] = data_i[423] & sel_one_hot_i[6];
  assign data_masked[422] = data_i[422] & sel_one_hot_i[6];
  assign data_masked[421] = data_i[421] & sel_one_hot_i[6];
  assign data_masked[420] = data_i[420] & sel_one_hot_i[6];
  assign data_masked[419] = data_i[419] & sel_one_hot_i[6];
  assign data_masked[418] = data_i[418] & sel_one_hot_i[6];
  assign data_masked[417] = data_i[417] & sel_one_hot_i[6];
  assign data_masked[416] = data_i[416] & sel_one_hot_i[6];
  assign data_masked[415] = data_i[415] & sel_one_hot_i[6];
  assign data_masked[414] = data_i[414] & sel_one_hot_i[6];
  assign data_masked[413] = data_i[413] & sel_one_hot_i[6];
  assign data_masked[412] = data_i[412] & sel_one_hot_i[6];
  assign data_masked[411] = data_i[411] & sel_one_hot_i[6];
  assign data_masked[410] = data_i[410] & sel_one_hot_i[6];
  assign data_masked[409] = data_i[409] & sel_one_hot_i[6];
  assign data_masked[408] = data_i[408] & sel_one_hot_i[6];
  assign data_masked[407] = data_i[407] & sel_one_hot_i[6];
  assign data_masked[406] = data_i[406] & sel_one_hot_i[6];
  assign data_masked[405] = data_i[405] & sel_one_hot_i[6];
  assign data_masked[404] = data_i[404] & sel_one_hot_i[6];
  assign data_masked[403] = data_i[403] & sel_one_hot_i[6];
  assign data_masked[402] = data_i[402] & sel_one_hot_i[6];
  assign data_masked[401] = data_i[401] & sel_one_hot_i[6];
  assign data_masked[400] = data_i[400] & sel_one_hot_i[6];
  assign data_masked[399] = data_i[399] & sel_one_hot_i[6];
  assign data_masked[398] = data_i[398] & sel_one_hot_i[6];
  assign data_masked[397] = data_i[397] & sel_one_hot_i[6];
  assign data_masked[396] = data_i[396] & sel_one_hot_i[6];
  assign data_masked[395] = data_i[395] & sel_one_hot_i[6];
  assign data_masked[394] = data_i[394] & sel_one_hot_i[6];
  assign data_masked[393] = data_i[393] & sel_one_hot_i[6];
  assign data_masked[392] = data_i[392] & sel_one_hot_i[6];
  assign data_masked[391] = data_i[391] & sel_one_hot_i[6];
  assign data_masked[390] = data_i[390] & sel_one_hot_i[6];
  assign data_masked[389] = data_i[389] & sel_one_hot_i[6];
  assign data_masked[388] = data_i[388] & sel_one_hot_i[6];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[6];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[6];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[6];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[6];
  assign data_masked[511] = data_i[511] & sel_one_hot_i[7];
  assign data_masked[510] = data_i[510] & sel_one_hot_i[7];
  assign data_masked[509] = data_i[509] & sel_one_hot_i[7];
  assign data_masked[508] = data_i[508] & sel_one_hot_i[7];
  assign data_masked[507] = data_i[507] & sel_one_hot_i[7];
  assign data_masked[506] = data_i[506] & sel_one_hot_i[7];
  assign data_masked[505] = data_i[505] & sel_one_hot_i[7];
  assign data_masked[504] = data_i[504] & sel_one_hot_i[7];
  assign data_masked[503] = data_i[503] & sel_one_hot_i[7];
  assign data_masked[502] = data_i[502] & sel_one_hot_i[7];
  assign data_masked[501] = data_i[501] & sel_one_hot_i[7];
  assign data_masked[500] = data_i[500] & sel_one_hot_i[7];
  assign data_masked[499] = data_i[499] & sel_one_hot_i[7];
  assign data_masked[498] = data_i[498] & sel_one_hot_i[7];
  assign data_masked[497] = data_i[497] & sel_one_hot_i[7];
  assign data_masked[496] = data_i[496] & sel_one_hot_i[7];
  assign data_masked[495] = data_i[495] & sel_one_hot_i[7];
  assign data_masked[494] = data_i[494] & sel_one_hot_i[7];
  assign data_masked[493] = data_i[493] & sel_one_hot_i[7];
  assign data_masked[492] = data_i[492] & sel_one_hot_i[7];
  assign data_masked[491] = data_i[491] & sel_one_hot_i[7];
  assign data_masked[490] = data_i[490] & sel_one_hot_i[7];
  assign data_masked[489] = data_i[489] & sel_one_hot_i[7];
  assign data_masked[488] = data_i[488] & sel_one_hot_i[7];
  assign data_masked[487] = data_i[487] & sel_one_hot_i[7];
  assign data_masked[486] = data_i[486] & sel_one_hot_i[7];
  assign data_masked[485] = data_i[485] & sel_one_hot_i[7];
  assign data_masked[484] = data_i[484] & sel_one_hot_i[7];
  assign data_masked[483] = data_i[483] & sel_one_hot_i[7];
  assign data_masked[482] = data_i[482] & sel_one_hot_i[7];
  assign data_masked[481] = data_i[481] & sel_one_hot_i[7];
  assign data_masked[480] = data_i[480] & sel_one_hot_i[7];
  assign data_masked[479] = data_i[479] & sel_one_hot_i[7];
  assign data_masked[478] = data_i[478] & sel_one_hot_i[7];
  assign data_masked[477] = data_i[477] & sel_one_hot_i[7];
  assign data_masked[476] = data_i[476] & sel_one_hot_i[7];
  assign data_masked[475] = data_i[475] & sel_one_hot_i[7];
  assign data_masked[474] = data_i[474] & sel_one_hot_i[7];
  assign data_masked[473] = data_i[473] & sel_one_hot_i[7];
  assign data_masked[472] = data_i[472] & sel_one_hot_i[7];
  assign data_masked[471] = data_i[471] & sel_one_hot_i[7];
  assign data_masked[470] = data_i[470] & sel_one_hot_i[7];
  assign data_masked[469] = data_i[469] & sel_one_hot_i[7];
  assign data_masked[468] = data_i[468] & sel_one_hot_i[7];
  assign data_masked[467] = data_i[467] & sel_one_hot_i[7];
  assign data_masked[466] = data_i[466] & sel_one_hot_i[7];
  assign data_masked[465] = data_i[465] & sel_one_hot_i[7];
  assign data_masked[464] = data_i[464] & sel_one_hot_i[7];
  assign data_masked[463] = data_i[463] & sel_one_hot_i[7];
  assign data_masked[462] = data_i[462] & sel_one_hot_i[7];
  assign data_masked[461] = data_i[461] & sel_one_hot_i[7];
  assign data_masked[460] = data_i[460] & sel_one_hot_i[7];
  assign data_masked[459] = data_i[459] & sel_one_hot_i[7];
  assign data_masked[458] = data_i[458] & sel_one_hot_i[7];
  assign data_masked[457] = data_i[457] & sel_one_hot_i[7];
  assign data_masked[456] = data_i[456] & sel_one_hot_i[7];
  assign data_masked[455] = data_i[455] & sel_one_hot_i[7];
  assign data_masked[454] = data_i[454] & sel_one_hot_i[7];
  assign data_masked[453] = data_i[453] & sel_one_hot_i[7];
  assign data_masked[452] = data_i[452] & sel_one_hot_i[7];
  assign data_masked[451] = data_i[451] & sel_one_hot_i[7];
  assign data_masked[450] = data_i[450] & sel_one_hot_i[7];
  assign data_masked[449] = data_i[449] & sel_one_hot_i[7];
  assign data_masked[448] = data_i[448] & sel_one_hot_i[7];
  assign data_masked[575] = data_i[575] & sel_one_hot_i[8];
  assign data_masked[574] = data_i[574] & sel_one_hot_i[8];
  assign data_masked[573] = data_i[573] & sel_one_hot_i[8];
  assign data_masked[572] = data_i[572] & sel_one_hot_i[8];
  assign data_masked[571] = data_i[571] & sel_one_hot_i[8];
  assign data_masked[570] = data_i[570] & sel_one_hot_i[8];
  assign data_masked[569] = data_i[569] & sel_one_hot_i[8];
  assign data_masked[568] = data_i[568] & sel_one_hot_i[8];
  assign data_masked[567] = data_i[567] & sel_one_hot_i[8];
  assign data_masked[566] = data_i[566] & sel_one_hot_i[8];
  assign data_masked[565] = data_i[565] & sel_one_hot_i[8];
  assign data_masked[564] = data_i[564] & sel_one_hot_i[8];
  assign data_masked[563] = data_i[563] & sel_one_hot_i[8];
  assign data_masked[562] = data_i[562] & sel_one_hot_i[8];
  assign data_masked[561] = data_i[561] & sel_one_hot_i[8];
  assign data_masked[560] = data_i[560] & sel_one_hot_i[8];
  assign data_masked[559] = data_i[559] & sel_one_hot_i[8];
  assign data_masked[558] = data_i[558] & sel_one_hot_i[8];
  assign data_masked[557] = data_i[557] & sel_one_hot_i[8];
  assign data_masked[556] = data_i[556] & sel_one_hot_i[8];
  assign data_masked[555] = data_i[555] & sel_one_hot_i[8];
  assign data_masked[554] = data_i[554] & sel_one_hot_i[8];
  assign data_masked[553] = data_i[553] & sel_one_hot_i[8];
  assign data_masked[552] = data_i[552] & sel_one_hot_i[8];
  assign data_masked[551] = data_i[551] & sel_one_hot_i[8];
  assign data_masked[550] = data_i[550] & sel_one_hot_i[8];
  assign data_masked[549] = data_i[549] & sel_one_hot_i[8];
  assign data_masked[548] = data_i[548] & sel_one_hot_i[8];
  assign data_masked[547] = data_i[547] & sel_one_hot_i[8];
  assign data_masked[546] = data_i[546] & sel_one_hot_i[8];
  assign data_masked[545] = data_i[545] & sel_one_hot_i[8];
  assign data_masked[544] = data_i[544] & sel_one_hot_i[8];
  assign data_masked[543] = data_i[543] & sel_one_hot_i[8];
  assign data_masked[542] = data_i[542] & sel_one_hot_i[8];
  assign data_masked[541] = data_i[541] & sel_one_hot_i[8];
  assign data_masked[540] = data_i[540] & sel_one_hot_i[8];
  assign data_masked[539] = data_i[539] & sel_one_hot_i[8];
  assign data_masked[538] = data_i[538] & sel_one_hot_i[8];
  assign data_masked[537] = data_i[537] & sel_one_hot_i[8];
  assign data_masked[536] = data_i[536] & sel_one_hot_i[8];
  assign data_masked[535] = data_i[535] & sel_one_hot_i[8];
  assign data_masked[534] = data_i[534] & sel_one_hot_i[8];
  assign data_masked[533] = data_i[533] & sel_one_hot_i[8];
  assign data_masked[532] = data_i[532] & sel_one_hot_i[8];
  assign data_masked[531] = data_i[531] & sel_one_hot_i[8];
  assign data_masked[530] = data_i[530] & sel_one_hot_i[8];
  assign data_masked[529] = data_i[529] & sel_one_hot_i[8];
  assign data_masked[528] = data_i[528] & sel_one_hot_i[8];
  assign data_masked[527] = data_i[527] & sel_one_hot_i[8];
  assign data_masked[526] = data_i[526] & sel_one_hot_i[8];
  assign data_masked[525] = data_i[525] & sel_one_hot_i[8];
  assign data_masked[524] = data_i[524] & sel_one_hot_i[8];
  assign data_masked[523] = data_i[523] & sel_one_hot_i[8];
  assign data_masked[522] = data_i[522] & sel_one_hot_i[8];
  assign data_masked[521] = data_i[521] & sel_one_hot_i[8];
  assign data_masked[520] = data_i[520] & sel_one_hot_i[8];
  assign data_masked[519] = data_i[519] & sel_one_hot_i[8];
  assign data_masked[518] = data_i[518] & sel_one_hot_i[8];
  assign data_masked[517] = data_i[517] & sel_one_hot_i[8];
  assign data_masked[516] = data_i[516] & sel_one_hot_i[8];
  assign data_masked[515] = data_i[515] & sel_one_hot_i[8];
  assign data_masked[514] = data_i[514] & sel_one_hot_i[8];
  assign data_masked[513] = data_i[513] & sel_one_hot_i[8];
  assign data_masked[512] = data_i[512] & sel_one_hot_i[8];
  assign data_masked[639] = data_i[639] & sel_one_hot_i[9];
  assign data_masked[638] = data_i[638] & sel_one_hot_i[9];
  assign data_masked[637] = data_i[637] & sel_one_hot_i[9];
  assign data_masked[636] = data_i[636] & sel_one_hot_i[9];
  assign data_masked[635] = data_i[635] & sel_one_hot_i[9];
  assign data_masked[634] = data_i[634] & sel_one_hot_i[9];
  assign data_masked[633] = data_i[633] & sel_one_hot_i[9];
  assign data_masked[632] = data_i[632] & sel_one_hot_i[9];
  assign data_masked[631] = data_i[631] & sel_one_hot_i[9];
  assign data_masked[630] = data_i[630] & sel_one_hot_i[9];
  assign data_masked[629] = data_i[629] & sel_one_hot_i[9];
  assign data_masked[628] = data_i[628] & sel_one_hot_i[9];
  assign data_masked[627] = data_i[627] & sel_one_hot_i[9];
  assign data_masked[626] = data_i[626] & sel_one_hot_i[9];
  assign data_masked[625] = data_i[625] & sel_one_hot_i[9];
  assign data_masked[624] = data_i[624] & sel_one_hot_i[9];
  assign data_masked[623] = data_i[623] & sel_one_hot_i[9];
  assign data_masked[622] = data_i[622] & sel_one_hot_i[9];
  assign data_masked[621] = data_i[621] & sel_one_hot_i[9];
  assign data_masked[620] = data_i[620] & sel_one_hot_i[9];
  assign data_masked[619] = data_i[619] & sel_one_hot_i[9];
  assign data_masked[618] = data_i[618] & sel_one_hot_i[9];
  assign data_masked[617] = data_i[617] & sel_one_hot_i[9];
  assign data_masked[616] = data_i[616] & sel_one_hot_i[9];
  assign data_masked[615] = data_i[615] & sel_one_hot_i[9];
  assign data_masked[614] = data_i[614] & sel_one_hot_i[9];
  assign data_masked[613] = data_i[613] & sel_one_hot_i[9];
  assign data_masked[612] = data_i[612] & sel_one_hot_i[9];
  assign data_masked[611] = data_i[611] & sel_one_hot_i[9];
  assign data_masked[610] = data_i[610] & sel_one_hot_i[9];
  assign data_masked[609] = data_i[609] & sel_one_hot_i[9];
  assign data_masked[608] = data_i[608] & sel_one_hot_i[9];
  assign data_masked[607] = data_i[607] & sel_one_hot_i[9];
  assign data_masked[606] = data_i[606] & sel_one_hot_i[9];
  assign data_masked[605] = data_i[605] & sel_one_hot_i[9];
  assign data_masked[604] = data_i[604] & sel_one_hot_i[9];
  assign data_masked[603] = data_i[603] & sel_one_hot_i[9];
  assign data_masked[602] = data_i[602] & sel_one_hot_i[9];
  assign data_masked[601] = data_i[601] & sel_one_hot_i[9];
  assign data_masked[600] = data_i[600] & sel_one_hot_i[9];
  assign data_masked[599] = data_i[599] & sel_one_hot_i[9];
  assign data_masked[598] = data_i[598] & sel_one_hot_i[9];
  assign data_masked[597] = data_i[597] & sel_one_hot_i[9];
  assign data_masked[596] = data_i[596] & sel_one_hot_i[9];
  assign data_masked[595] = data_i[595] & sel_one_hot_i[9];
  assign data_masked[594] = data_i[594] & sel_one_hot_i[9];
  assign data_masked[593] = data_i[593] & sel_one_hot_i[9];
  assign data_masked[592] = data_i[592] & sel_one_hot_i[9];
  assign data_masked[591] = data_i[591] & sel_one_hot_i[9];
  assign data_masked[590] = data_i[590] & sel_one_hot_i[9];
  assign data_masked[589] = data_i[589] & sel_one_hot_i[9];
  assign data_masked[588] = data_i[588] & sel_one_hot_i[9];
  assign data_masked[587] = data_i[587] & sel_one_hot_i[9];
  assign data_masked[586] = data_i[586] & sel_one_hot_i[9];
  assign data_masked[585] = data_i[585] & sel_one_hot_i[9];
  assign data_masked[584] = data_i[584] & sel_one_hot_i[9];
  assign data_masked[583] = data_i[583] & sel_one_hot_i[9];
  assign data_masked[582] = data_i[582] & sel_one_hot_i[9];
  assign data_masked[581] = data_i[581] & sel_one_hot_i[9];
  assign data_masked[580] = data_i[580] & sel_one_hot_i[9];
  assign data_masked[579] = data_i[579] & sel_one_hot_i[9];
  assign data_masked[578] = data_i[578] & sel_one_hot_i[9];
  assign data_masked[577] = data_i[577] & sel_one_hot_i[9];
  assign data_masked[576] = data_i[576] & sel_one_hot_i[9];
  assign data_masked[703] = data_i[703] & sel_one_hot_i[10];
  assign data_masked[702] = data_i[702] & sel_one_hot_i[10];
  assign data_masked[701] = data_i[701] & sel_one_hot_i[10];
  assign data_masked[700] = data_i[700] & sel_one_hot_i[10];
  assign data_masked[699] = data_i[699] & sel_one_hot_i[10];
  assign data_masked[698] = data_i[698] & sel_one_hot_i[10];
  assign data_masked[697] = data_i[697] & sel_one_hot_i[10];
  assign data_masked[696] = data_i[696] & sel_one_hot_i[10];
  assign data_masked[695] = data_i[695] & sel_one_hot_i[10];
  assign data_masked[694] = data_i[694] & sel_one_hot_i[10];
  assign data_masked[693] = data_i[693] & sel_one_hot_i[10];
  assign data_masked[692] = data_i[692] & sel_one_hot_i[10];
  assign data_masked[691] = data_i[691] & sel_one_hot_i[10];
  assign data_masked[690] = data_i[690] & sel_one_hot_i[10];
  assign data_masked[689] = data_i[689] & sel_one_hot_i[10];
  assign data_masked[688] = data_i[688] & sel_one_hot_i[10];
  assign data_masked[687] = data_i[687] & sel_one_hot_i[10];
  assign data_masked[686] = data_i[686] & sel_one_hot_i[10];
  assign data_masked[685] = data_i[685] & sel_one_hot_i[10];
  assign data_masked[684] = data_i[684] & sel_one_hot_i[10];
  assign data_masked[683] = data_i[683] & sel_one_hot_i[10];
  assign data_masked[682] = data_i[682] & sel_one_hot_i[10];
  assign data_masked[681] = data_i[681] & sel_one_hot_i[10];
  assign data_masked[680] = data_i[680] & sel_one_hot_i[10];
  assign data_masked[679] = data_i[679] & sel_one_hot_i[10];
  assign data_masked[678] = data_i[678] & sel_one_hot_i[10];
  assign data_masked[677] = data_i[677] & sel_one_hot_i[10];
  assign data_masked[676] = data_i[676] & sel_one_hot_i[10];
  assign data_masked[675] = data_i[675] & sel_one_hot_i[10];
  assign data_masked[674] = data_i[674] & sel_one_hot_i[10];
  assign data_masked[673] = data_i[673] & sel_one_hot_i[10];
  assign data_masked[672] = data_i[672] & sel_one_hot_i[10];
  assign data_masked[671] = data_i[671] & sel_one_hot_i[10];
  assign data_masked[670] = data_i[670] & sel_one_hot_i[10];
  assign data_masked[669] = data_i[669] & sel_one_hot_i[10];
  assign data_masked[668] = data_i[668] & sel_one_hot_i[10];
  assign data_masked[667] = data_i[667] & sel_one_hot_i[10];
  assign data_masked[666] = data_i[666] & sel_one_hot_i[10];
  assign data_masked[665] = data_i[665] & sel_one_hot_i[10];
  assign data_masked[664] = data_i[664] & sel_one_hot_i[10];
  assign data_masked[663] = data_i[663] & sel_one_hot_i[10];
  assign data_masked[662] = data_i[662] & sel_one_hot_i[10];
  assign data_masked[661] = data_i[661] & sel_one_hot_i[10];
  assign data_masked[660] = data_i[660] & sel_one_hot_i[10];
  assign data_masked[659] = data_i[659] & sel_one_hot_i[10];
  assign data_masked[658] = data_i[658] & sel_one_hot_i[10];
  assign data_masked[657] = data_i[657] & sel_one_hot_i[10];
  assign data_masked[656] = data_i[656] & sel_one_hot_i[10];
  assign data_masked[655] = data_i[655] & sel_one_hot_i[10];
  assign data_masked[654] = data_i[654] & sel_one_hot_i[10];
  assign data_masked[653] = data_i[653] & sel_one_hot_i[10];
  assign data_masked[652] = data_i[652] & sel_one_hot_i[10];
  assign data_masked[651] = data_i[651] & sel_one_hot_i[10];
  assign data_masked[650] = data_i[650] & sel_one_hot_i[10];
  assign data_masked[649] = data_i[649] & sel_one_hot_i[10];
  assign data_masked[648] = data_i[648] & sel_one_hot_i[10];
  assign data_masked[647] = data_i[647] & sel_one_hot_i[10];
  assign data_masked[646] = data_i[646] & sel_one_hot_i[10];
  assign data_masked[645] = data_i[645] & sel_one_hot_i[10];
  assign data_masked[644] = data_i[644] & sel_one_hot_i[10];
  assign data_masked[643] = data_i[643] & sel_one_hot_i[10];
  assign data_masked[642] = data_i[642] & sel_one_hot_i[10];
  assign data_masked[641] = data_i[641] & sel_one_hot_i[10];
  assign data_masked[640] = data_i[640] & sel_one_hot_i[10];
  assign data_masked[767] = data_i[767] & sel_one_hot_i[11];
  assign data_masked[766] = data_i[766] & sel_one_hot_i[11];
  assign data_masked[765] = data_i[765] & sel_one_hot_i[11];
  assign data_masked[764] = data_i[764] & sel_one_hot_i[11];
  assign data_masked[763] = data_i[763] & sel_one_hot_i[11];
  assign data_masked[762] = data_i[762] & sel_one_hot_i[11];
  assign data_masked[761] = data_i[761] & sel_one_hot_i[11];
  assign data_masked[760] = data_i[760] & sel_one_hot_i[11];
  assign data_masked[759] = data_i[759] & sel_one_hot_i[11];
  assign data_masked[758] = data_i[758] & sel_one_hot_i[11];
  assign data_masked[757] = data_i[757] & sel_one_hot_i[11];
  assign data_masked[756] = data_i[756] & sel_one_hot_i[11];
  assign data_masked[755] = data_i[755] & sel_one_hot_i[11];
  assign data_masked[754] = data_i[754] & sel_one_hot_i[11];
  assign data_masked[753] = data_i[753] & sel_one_hot_i[11];
  assign data_masked[752] = data_i[752] & sel_one_hot_i[11];
  assign data_masked[751] = data_i[751] & sel_one_hot_i[11];
  assign data_masked[750] = data_i[750] & sel_one_hot_i[11];
  assign data_masked[749] = data_i[749] & sel_one_hot_i[11];
  assign data_masked[748] = data_i[748] & sel_one_hot_i[11];
  assign data_masked[747] = data_i[747] & sel_one_hot_i[11];
  assign data_masked[746] = data_i[746] & sel_one_hot_i[11];
  assign data_masked[745] = data_i[745] & sel_one_hot_i[11];
  assign data_masked[744] = data_i[744] & sel_one_hot_i[11];
  assign data_masked[743] = data_i[743] & sel_one_hot_i[11];
  assign data_masked[742] = data_i[742] & sel_one_hot_i[11];
  assign data_masked[741] = data_i[741] & sel_one_hot_i[11];
  assign data_masked[740] = data_i[740] & sel_one_hot_i[11];
  assign data_masked[739] = data_i[739] & sel_one_hot_i[11];
  assign data_masked[738] = data_i[738] & sel_one_hot_i[11];
  assign data_masked[737] = data_i[737] & sel_one_hot_i[11];
  assign data_masked[736] = data_i[736] & sel_one_hot_i[11];
  assign data_masked[735] = data_i[735] & sel_one_hot_i[11];
  assign data_masked[734] = data_i[734] & sel_one_hot_i[11];
  assign data_masked[733] = data_i[733] & sel_one_hot_i[11];
  assign data_masked[732] = data_i[732] & sel_one_hot_i[11];
  assign data_masked[731] = data_i[731] & sel_one_hot_i[11];
  assign data_masked[730] = data_i[730] & sel_one_hot_i[11];
  assign data_masked[729] = data_i[729] & sel_one_hot_i[11];
  assign data_masked[728] = data_i[728] & sel_one_hot_i[11];
  assign data_masked[727] = data_i[727] & sel_one_hot_i[11];
  assign data_masked[726] = data_i[726] & sel_one_hot_i[11];
  assign data_masked[725] = data_i[725] & sel_one_hot_i[11];
  assign data_masked[724] = data_i[724] & sel_one_hot_i[11];
  assign data_masked[723] = data_i[723] & sel_one_hot_i[11];
  assign data_masked[722] = data_i[722] & sel_one_hot_i[11];
  assign data_masked[721] = data_i[721] & sel_one_hot_i[11];
  assign data_masked[720] = data_i[720] & sel_one_hot_i[11];
  assign data_masked[719] = data_i[719] & sel_one_hot_i[11];
  assign data_masked[718] = data_i[718] & sel_one_hot_i[11];
  assign data_masked[717] = data_i[717] & sel_one_hot_i[11];
  assign data_masked[716] = data_i[716] & sel_one_hot_i[11];
  assign data_masked[715] = data_i[715] & sel_one_hot_i[11];
  assign data_masked[714] = data_i[714] & sel_one_hot_i[11];
  assign data_masked[713] = data_i[713] & sel_one_hot_i[11];
  assign data_masked[712] = data_i[712] & sel_one_hot_i[11];
  assign data_masked[711] = data_i[711] & sel_one_hot_i[11];
  assign data_masked[710] = data_i[710] & sel_one_hot_i[11];
  assign data_masked[709] = data_i[709] & sel_one_hot_i[11];
  assign data_masked[708] = data_i[708] & sel_one_hot_i[11];
  assign data_masked[707] = data_i[707] & sel_one_hot_i[11];
  assign data_masked[706] = data_i[706] & sel_one_hot_i[11];
  assign data_masked[705] = data_i[705] & sel_one_hot_i[11];
  assign data_masked[704] = data_i[704] & sel_one_hot_i[11];
  assign data_masked[831] = data_i[831] & sel_one_hot_i[12];
  assign data_masked[830] = data_i[830] & sel_one_hot_i[12];
  assign data_masked[829] = data_i[829] & sel_one_hot_i[12];
  assign data_masked[828] = data_i[828] & sel_one_hot_i[12];
  assign data_masked[827] = data_i[827] & sel_one_hot_i[12];
  assign data_masked[826] = data_i[826] & sel_one_hot_i[12];
  assign data_masked[825] = data_i[825] & sel_one_hot_i[12];
  assign data_masked[824] = data_i[824] & sel_one_hot_i[12];
  assign data_masked[823] = data_i[823] & sel_one_hot_i[12];
  assign data_masked[822] = data_i[822] & sel_one_hot_i[12];
  assign data_masked[821] = data_i[821] & sel_one_hot_i[12];
  assign data_masked[820] = data_i[820] & sel_one_hot_i[12];
  assign data_masked[819] = data_i[819] & sel_one_hot_i[12];
  assign data_masked[818] = data_i[818] & sel_one_hot_i[12];
  assign data_masked[817] = data_i[817] & sel_one_hot_i[12];
  assign data_masked[816] = data_i[816] & sel_one_hot_i[12];
  assign data_masked[815] = data_i[815] & sel_one_hot_i[12];
  assign data_masked[814] = data_i[814] & sel_one_hot_i[12];
  assign data_masked[813] = data_i[813] & sel_one_hot_i[12];
  assign data_masked[812] = data_i[812] & sel_one_hot_i[12];
  assign data_masked[811] = data_i[811] & sel_one_hot_i[12];
  assign data_masked[810] = data_i[810] & sel_one_hot_i[12];
  assign data_masked[809] = data_i[809] & sel_one_hot_i[12];
  assign data_masked[808] = data_i[808] & sel_one_hot_i[12];
  assign data_masked[807] = data_i[807] & sel_one_hot_i[12];
  assign data_masked[806] = data_i[806] & sel_one_hot_i[12];
  assign data_masked[805] = data_i[805] & sel_one_hot_i[12];
  assign data_masked[804] = data_i[804] & sel_one_hot_i[12];
  assign data_masked[803] = data_i[803] & sel_one_hot_i[12];
  assign data_masked[802] = data_i[802] & sel_one_hot_i[12];
  assign data_masked[801] = data_i[801] & sel_one_hot_i[12];
  assign data_masked[800] = data_i[800] & sel_one_hot_i[12];
  assign data_masked[799] = data_i[799] & sel_one_hot_i[12];
  assign data_masked[798] = data_i[798] & sel_one_hot_i[12];
  assign data_masked[797] = data_i[797] & sel_one_hot_i[12];
  assign data_masked[796] = data_i[796] & sel_one_hot_i[12];
  assign data_masked[795] = data_i[795] & sel_one_hot_i[12];
  assign data_masked[794] = data_i[794] & sel_one_hot_i[12];
  assign data_masked[793] = data_i[793] & sel_one_hot_i[12];
  assign data_masked[792] = data_i[792] & sel_one_hot_i[12];
  assign data_masked[791] = data_i[791] & sel_one_hot_i[12];
  assign data_masked[790] = data_i[790] & sel_one_hot_i[12];
  assign data_masked[789] = data_i[789] & sel_one_hot_i[12];
  assign data_masked[788] = data_i[788] & sel_one_hot_i[12];
  assign data_masked[787] = data_i[787] & sel_one_hot_i[12];
  assign data_masked[786] = data_i[786] & sel_one_hot_i[12];
  assign data_masked[785] = data_i[785] & sel_one_hot_i[12];
  assign data_masked[784] = data_i[784] & sel_one_hot_i[12];
  assign data_masked[783] = data_i[783] & sel_one_hot_i[12];
  assign data_masked[782] = data_i[782] & sel_one_hot_i[12];
  assign data_masked[781] = data_i[781] & sel_one_hot_i[12];
  assign data_masked[780] = data_i[780] & sel_one_hot_i[12];
  assign data_masked[779] = data_i[779] & sel_one_hot_i[12];
  assign data_masked[778] = data_i[778] & sel_one_hot_i[12];
  assign data_masked[777] = data_i[777] & sel_one_hot_i[12];
  assign data_masked[776] = data_i[776] & sel_one_hot_i[12];
  assign data_masked[775] = data_i[775] & sel_one_hot_i[12];
  assign data_masked[774] = data_i[774] & sel_one_hot_i[12];
  assign data_masked[773] = data_i[773] & sel_one_hot_i[12];
  assign data_masked[772] = data_i[772] & sel_one_hot_i[12];
  assign data_masked[771] = data_i[771] & sel_one_hot_i[12];
  assign data_masked[770] = data_i[770] & sel_one_hot_i[12];
  assign data_masked[769] = data_i[769] & sel_one_hot_i[12];
  assign data_masked[768] = data_i[768] & sel_one_hot_i[12];
  assign data_masked[895] = data_i[895] & sel_one_hot_i[13];
  assign data_masked[894] = data_i[894] & sel_one_hot_i[13];
  assign data_masked[893] = data_i[893] & sel_one_hot_i[13];
  assign data_masked[892] = data_i[892] & sel_one_hot_i[13];
  assign data_masked[891] = data_i[891] & sel_one_hot_i[13];
  assign data_masked[890] = data_i[890] & sel_one_hot_i[13];
  assign data_masked[889] = data_i[889] & sel_one_hot_i[13];
  assign data_masked[888] = data_i[888] & sel_one_hot_i[13];
  assign data_masked[887] = data_i[887] & sel_one_hot_i[13];
  assign data_masked[886] = data_i[886] & sel_one_hot_i[13];
  assign data_masked[885] = data_i[885] & sel_one_hot_i[13];
  assign data_masked[884] = data_i[884] & sel_one_hot_i[13];
  assign data_masked[883] = data_i[883] & sel_one_hot_i[13];
  assign data_masked[882] = data_i[882] & sel_one_hot_i[13];
  assign data_masked[881] = data_i[881] & sel_one_hot_i[13];
  assign data_masked[880] = data_i[880] & sel_one_hot_i[13];
  assign data_masked[879] = data_i[879] & sel_one_hot_i[13];
  assign data_masked[878] = data_i[878] & sel_one_hot_i[13];
  assign data_masked[877] = data_i[877] & sel_one_hot_i[13];
  assign data_masked[876] = data_i[876] & sel_one_hot_i[13];
  assign data_masked[875] = data_i[875] & sel_one_hot_i[13];
  assign data_masked[874] = data_i[874] & sel_one_hot_i[13];
  assign data_masked[873] = data_i[873] & sel_one_hot_i[13];
  assign data_masked[872] = data_i[872] & sel_one_hot_i[13];
  assign data_masked[871] = data_i[871] & sel_one_hot_i[13];
  assign data_masked[870] = data_i[870] & sel_one_hot_i[13];
  assign data_masked[869] = data_i[869] & sel_one_hot_i[13];
  assign data_masked[868] = data_i[868] & sel_one_hot_i[13];
  assign data_masked[867] = data_i[867] & sel_one_hot_i[13];
  assign data_masked[866] = data_i[866] & sel_one_hot_i[13];
  assign data_masked[865] = data_i[865] & sel_one_hot_i[13];
  assign data_masked[864] = data_i[864] & sel_one_hot_i[13];
  assign data_masked[863] = data_i[863] & sel_one_hot_i[13];
  assign data_masked[862] = data_i[862] & sel_one_hot_i[13];
  assign data_masked[861] = data_i[861] & sel_one_hot_i[13];
  assign data_masked[860] = data_i[860] & sel_one_hot_i[13];
  assign data_masked[859] = data_i[859] & sel_one_hot_i[13];
  assign data_masked[858] = data_i[858] & sel_one_hot_i[13];
  assign data_masked[857] = data_i[857] & sel_one_hot_i[13];
  assign data_masked[856] = data_i[856] & sel_one_hot_i[13];
  assign data_masked[855] = data_i[855] & sel_one_hot_i[13];
  assign data_masked[854] = data_i[854] & sel_one_hot_i[13];
  assign data_masked[853] = data_i[853] & sel_one_hot_i[13];
  assign data_masked[852] = data_i[852] & sel_one_hot_i[13];
  assign data_masked[851] = data_i[851] & sel_one_hot_i[13];
  assign data_masked[850] = data_i[850] & sel_one_hot_i[13];
  assign data_masked[849] = data_i[849] & sel_one_hot_i[13];
  assign data_masked[848] = data_i[848] & sel_one_hot_i[13];
  assign data_masked[847] = data_i[847] & sel_one_hot_i[13];
  assign data_masked[846] = data_i[846] & sel_one_hot_i[13];
  assign data_masked[845] = data_i[845] & sel_one_hot_i[13];
  assign data_masked[844] = data_i[844] & sel_one_hot_i[13];
  assign data_masked[843] = data_i[843] & sel_one_hot_i[13];
  assign data_masked[842] = data_i[842] & sel_one_hot_i[13];
  assign data_masked[841] = data_i[841] & sel_one_hot_i[13];
  assign data_masked[840] = data_i[840] & sel_one_hot_i[13];
  assign data_masked[839] = data_i[839] & sel_one_hot_i[13];
  assign data_masked[838] = data_i[838] & sel_one_hot_i[13];
  assign data_masked[837] = data_i[837] & sel_one_hot_i[13];
  assign data_masked[836] = data_i[836] & sel_one_hot_i[13];
  assign data_masked[835] = data_i[835] & sel_one_hot_i[13];
  assign data_masked[834] = data_i[834] & sel_one_hot_i[13];
  assign data_masked[833] = data_i[833] & sel_one_hot_i[13];
  assign data_masked[832] = data_i[832] & sel_one_hot_i[13];
  assign data_masked[959] = data_i[959] & sel_one_hot_i[14];
  assign data_masked[958] = data_i[958] & sel_one_hot_i[14];
  assign data_masked[957] = data_i[957] & sel_one_hot_i[14];
  assign data_masked[956] = data_i[956] & sel_one_hot_i[14];
  assign data_masked[955] = data_i[955] & sel_one_hot_i[14];
  assign data_masked[954] = data_i[954] & sel_one_hot_i[14];
  assign data_masked[953] = data_i[953] & sel_one_hot_i[14];
  assign data_masked[952] = data_i[952] & sel_one_hot_i[14];
  assign data_masked[951] = data_i[951] & sel_one_hot_i[14];
  assign data_masked[950] = data_i[950] & sel_one_hot_i[14];
  assign data_masked[949] = data_i[949] & sel_one_hot_i[14];
  assign data_masked[948] = data_i[948] & sel_one_hot_i[14];
  assign data_masked[947] = data_i[947] & sel_one_hot_i[14];
  assign data_masked[946] = data_i[946] & sel_one_hot_i[14];
  assign data_masked[945] = data_i[945] & sel_one_hot_i[14];
  assign data_masked[944] = data_i[944] & sel_one_hot_i[14];
  assign data_masked[943] = data_i[943] & sel_one_hot_i[14];
  assign data_masked[942] = data_i[942] & sel_one_hot_i[14];
  assign data_masked[941] = data_i[941] & sel_one_hot_i[14];
  assign data_masked[940] = data_i[940] & sel_one_hot_i[14];
  assign data_masked[939] = data_i[939] & sel_one_hot_i[14];
  assign data_masked[938] = data_i[938] & sel_one_hot_i[14];
  assign data_masked[937] = data_i[937] & sel_one_hot_i[14];
  assign data_masked[936] = data_i[936] & sel_one_hot_i[14];
  assign data_masked[935] = data_i[935] & sel_one_hot_i[14];
  assign data_masked[934] = data_i[934] & sel_one_hot_i[14];
  assign data_masked[933] = data_i[933] & sel_one_hot_i[14];
  assign data_masked[932] = data_i[932] & sel_one_hot_i[14];
  assign data_masked[931] = data_i[931] & sel_one_hot_i[14];
  assign data_masked[930] = data_i[930] & sel_one_hot_i[14];
  assign data_masked[929] = data_i[929] & sel_one_hot_i[14];
  assign data_masked[928] = data_i[928] & sel_one_hot_i[14];
  assign data_masked[927] = data_i[927] & sel_one_hot_i[14];
  assign data_masked[926] = data_i[926] & sel_one_hot_i[14];
  assign data_masked[925] = data_i[925] & sel_one_hot_i[14];
  assign data_masked[924] = data_i[924] & sel_one_hot_i[14];
  assign data_masked[923] = data_i[923] & sel_one_hot_i[14];
  assign data_masked[922] = data_i[922] & sel_one_hot_i[14];
  assign data_masked[921] = data_i[921] & sel_one_hot_i[14];
  assign data_masked[920] = data_i[920] & sel_one_hot_i[14];
  assign data_masked[919] = data_i[919] & sel_one_hot_i[14];
  assign data_masked[918] = data_i[918] & sel_one_hot_i[14];
  assign data_masked[917] = data_i[917] & sel_one_hot_i[14];
  assign data_masked[916] = data_i[916] & sel_one_hot_i[14];
  assign data_masked[915] = data_i[915] & sel_one_hot_i[14];
  assign data_masked[914] = data_i[914] & sel_one_hot_i[14];
  assign data_masked[913] = data_i[913] & sel_one_hot_i[14];
  assign data_masked[912] = data_i[912] & sel_one_hot_i[14];
  assign data_masked[911] = data_i[911] & sel_one_hot_i[14];
  assign data_masked[910] = data_i[910] & sel_one_hot_i[14];
  assign data_masked[909] = data_i[909] & sel_one_hot_i[14];
  assign data_masked[908] = data_i[908] & sel_one_hot_i[14];
  assign data_masked[907] = data_i[907] & sel_one_hot_i[14];
  assign data_masked[906] = data_i[906] & sel_one_hot_i[14];
  assign data_masked[905] = data_i[905] & sel_one_hot_i[14];
  assign data_masked[904] = data_i[904] & sel_one_hot_i[14];
  assign data_masked[903] = data_i[903] & sel_one_hot_i[14];
  assign data_masked[902] = data_i[902] & sel_one_hot_i[14];
  assign data_masked[901] = data_i[901] & sel_one_hot_i[14];
  assign data_masked[900] = data_i[900] & sel_one_hot_i[14];
  assign data_masked[899] = data_i[899] & sel_one_hot_i[14];
  assign data_masked[898] = data_i[898] & sel_one_hot_i[14];
  assign data_masked[897] = data_i[897] & sel_one_hot_i[14];
  assign data_masked[896] = data_i[896] & sel_one_hot_i[14];
  assign data_masked[1023] = data_i[1023] & sel_one_hot_i[15];
  assign data_masked[1022] = data_i[1022] & sel_one_hot_i[15];
  assign data_masked[1021] = data_i[1021] & sel_one_hot_i[15];
  assign data_masked[1020] = data_i[1020] & sel_one_hot_i[15];
  assign data_masked[1019] = data_i[1019] & sel_one_hot_i[15];
  assign data_masked[1018] = data_i[1018] & sel_one_hot_i[15];
  assign data_masked[1017] = data_i[1017] & sel_one_hot_i[15];
  assign data_masked[1016] = data_i[1016] & sel_one_hot_i[15];
  assign data_masked[1015] = data_i[1015] & sel_one_hot_i[15];
  assign data_masked[1014] = data_i[1014] & sel_one_hot_i[15];
  assign data_masked[1013] = data_i[1013] & sel_one_hot_i[15];
  assign data_masked[1012] = data_i[1012] & sel_one_hot_i[15];
  assign data_masked[1011] = data_i[1011] & sel_one_hot_i[15];
  assign data_masked[1010] = data_i[1010] & sel_one_hot_i[15];
  assign data_masked[1009] = data_i[1009] & sel_one_hot_i[15];
  assign data_masked[1008] = data_i[1008] & sel_one_hot_i[15];
  assign data_masked[1007] = data_i[1007] & sel_one_hot_i[15];
  assign data_masked[1006] = data_i[1006] & sel_one_hot_i[15];
  assign data_masked[1005] = data_i[1005] & sel_one_hot_i[15];
  assign data_masked[1004] = data_i[1004] & sel_one_hot_i[15];
  assign data_masked[1003] = data_i[1003] & sel_one_hot_i[15];
  assign data_masked[1002] = data_i[1002] & sel_one_hot_i[15];
  assign data_masked[1001] = data_i[1001] & sel_one_hot_i[15];
  assign data_masked[1000] = data_i[1000] & sel_one_hot_i[15];
  assign data_masked[999] = data_i[999] & sel_one_hot_i[15];
  assign data_masked[998] = data_i[998] & sel_one_hot_i[15];
  assign data_masked[997] = data_i[997] & sel_one_hot_i[15];
  assign data_masked[996] = data_i[996] & sel_one_hot_i[15];
  assign data_masked[995] = data_i[995] & sel_one_hot_i[15];
  assign data_masked[994] = data_i[994] & sel_one_hot_i[15];
  assign data_masked[993] = data_i[993] & sel_one_hot_i[15];
  assign data_masked[992] = data_i[992] & sel_one_hot_i[15];
  assign data_masked[991] = data_i[991] & sel_one_hot_i[15];
  assign data_masked[990] = data_i[990] & sel_one_hot_i[15];
  assign data_masked[989] = data_i[989] & sel_one_hot_i[15];
  assign data_masked[988] = data_i[988] & sel_one_hot_i[15];
  assign data_masked[987] = data_i[987] & sel_one_hot_i[15];
  assign data_masked[986] = data_i[986] & sel_one_hot_i[15];
  assign data_masked[985] = data_i[985] & sel_one_hot_i[15];
  assign data_masked[984] = data_i[984] & sel_one_hot_i[15];
  assign data_masked[983] = data_i[983] & sel_one_hot_i[15];
  assign data_masked[982] = data_i[982] & sel_one_hot_i[15];
  assign data_masked[981] = data_i[981] & sel_one_hot_i[15];
  assign data_masked[980] = data_i[980] & sel_one_hot_i[15];
  assign data_masked[979] = data_i[979] & sel_one_hot_i[15];
  assign data_masked[978] = data_i[978] & sel_one_hot_i[15];
  assign data_masked[977] = data_i[977] & sel_one_hot_i[15];
  assign data_masked[976] = data_i[976] & sel_one_hot_i[15];
  assign data_masked[975] = data_i[975] & sel_one_hot_i[15];
  assign data_masked[974] = data_i[974] & sel_one_hot_i[15];
  assign data_masked[973] = data_i[973] & sel_one_hot_i[15];
  assign data_masked[972] = data_i[972] & sel_one_hot_i[15];
  assign data_masked[971] = data_i[971] & sel_one_hot_i[15];
  assign data_masked[970] = data_i[970] & sel_one_hot_i[15];
  assign data_masked[969] = data_i[969] & sel_one_hot_i[15];
  assign data_masked[968] = data_i[968] & sel_one_hot_i[15];
  assign data_masked[967] = data_i[967] & sel_one_hot_i[15];
  assign data_masked[966] = data_i[966] & sel_one_hot_i[15];
  assign data_masked[965] = data_i[965] & sel_one_hot_i[15];
  assign data_masked[964] = data_i[964] & sel_one_hot_i[15];
  assign data_masked[963] = data_i[963] & sel_one_hot_i[15];
  assign data_masked[962] = data_i[962] & sel_one_hot_i[15];
  assign data_masked[961] = data_i[961] & sel_one_hot_i[15];
  assign data_masked[960] = data_i[960] & sel_one_hot_i[15];
  assign data_masked[1087] = data_i[1087] & sel_one_hot_i[16];
  assign data_masked[1086] = data_i[1086] & sel_one_hot_i[16];
  assign data_masked[1085] = data_i[1085] & sel_one_hot_i[16];
  assign data_masked[1084] = data_i[1084] & sel_one_hot_i[16];
  assign data_masked[1083] = data_i[1083] & sel_one_hot_i[16];
  assign data_masked[1082] = data_i[1082] & sel_one_hot_i[16];
  assign data_masked[1081] = data_i[1081] & sel_one_hot_i[16];
  assign data_masked[1080] = data_i[1080] & sel_one_hot_i[16];
  assign data_masked[1079] = data_i[1079] & sel_one_hot_i[16];
  assign data_masked[1078] = data_i[1078] & sel_one_hot_i[16];
  assign data_masked[1077] = data_i[1077] & sel_one_hot_i[16];
  assign data_masked[1076] = data_i[1076] & sel_one_hot_i[16];
  assign data_masked[1075] = data_i[1075] & sel_one_hot_i[16];
  assign data_masked[1074] = data_i[1074] & sel_one_hot_i[16];
  assign data_masked[1073] = data_i[1073] & sel_one_hot_i[16];
  assign data_masked[1072] = data_i[1072] & sel_one_hot_i[16];
  assign data_masked[1071] = data_i[1071] & sel_one_hot_i[16];
  assign data_masked[1070] = data_i[1070] & sel_one_hot_i[16];
  assign data_masked[1069] = data_i[1069] & sel_one_hot_i[16];
  assign data_masked[1068] = data_i[1068] & sel_one_hot_i[16];
  assign data_masked[1067] = data_i[1067] & sel_one_hot_i[16];
  assign data_masked[1066] = data_i[1066] & sel_one_hot_i[16];
  assign data_masked[1065] = data_i[1065] & sel_one_hot_i[16];
  assign data_masked[1064] = data_i[1064] & sel_one_hot_i[16];
  assign data_masked[1063] = data_i[1063] & sel_one_hot_i[16];
  assign data_masked[1062] = data_i[1062] & sel_one_hot_i[16];
  assign data_masked[1061] = data_i[1061] & sel_one_hot_i[16];
  assign data_masked[1060] = data_i[1060] & sel_one_hot_i[16];
  assign data_masked[1059] = data_i[1059] & sel_one_hot_i[16];
  assign data_masked[1058] = data_i[1058] & sel_one_hot_i[16];
  assign data_masked[1057] = data_i[1057] & sel_one_hot_i[16];
  assign data_masked[1056] = data_i[1056] & sel_one_hot_i[16];
  assign data_masked[1055] = data_i[1055] & sel_one_hot_i[16];
  assign data_masked[1054] = data_i[1054] & sel_one_hot_i[16];
  assign data_masked[1053] = data_i[1053] & sel_one_hot_i[16];
  assign data_masked[1052] = data_i[1052] & sel_one_hot_i[16];
  assign data_masked[1051] = data_i[1051] & sel_one_hot_i[16];
  assign data_masked[1050] = data_i[1050] & sel_one_hot_i[16];
  assign data_masked[1049] = data_i[1049] & sel_one_hot_i[16];
  assign data_masked[1048] = data_i[1048] & sel_one_hot_i[16];
  assign data_masked[1047] = data_i[1047] & sel_one_hot_i[16];
  assign data_masked[1046] = data_i[1046] & sel_one_hot_i[16];
  assign data_masked[1045] = data_i[1045] & sel_one_hot_i[16];
  assign data_masked[1044] = data_i[1044] & sel_one_hot_i[16];
  assign data_masked[1043] = data_i[1043] & sel_one_hot_i[16];
  assign data_masked[1042] = data_i[1042] & sel_one_hot_i[16];
  assign data_masked[1041] = data_i[1041] & sel_one_hot_i[16];
  assign data_masked[1040] = data_i[1040] & sel_one_hot_i[16];
  assign data_masked[1039] = data_i[1039] & sel_one_hot_i[16];
  assign data_masked[1038] = data_i[1038] & sel_one_hot_i[16];
  assign data_masked[1037] = data_i[1037] & sel_one_hot_i[16];
  assign data_masked[1036] = data_i[1036] & sel_one_hot_i[16];
  assign data_masked[1035] = data_i[1035] & sel_one_hot_i[16];
  assign data_masked[1034] = data_i[1034] & sel_one_hot_i[16];
  assign data_masked[1033] = data_i[1033] & sel_one_hot_i[16];
  assign data_masked[1032] = data_i[1032] & sel_one_hot_i[16];
  assign data_masked[1031] = data_i[1031] & sel_one_hot_i[16];
  assign data_masked[1030] = data_i[1030] & sel_one_hot_i[16];
  assign data_masked[1029] = data_i[1029] & sel_one_hot_i[16];
  assign data_masked[1028] = data_i[1028] & sel_one_hot_i[16];
  assign data_masked[1027] = data_i[1027] & sel_one_hot_i[16];
  assign data_masked[1026] = data_i[1026] & sel_one_hot_i[16];
  assign data_masked[1025] = data_i[1025] & sel_one_hot_i[16];
  assign data_masked[1024] = data_i[1024] & sel_one_hot_i[16];
  assign data_masked[1151] = data_i[1151] & sel_one_hot_i[17];
  assign data_masked[1150] = data_i[1150] & sel_one_hot_i[17];
  assign data_masked[1149] = data_i[1149] & sel_one_hot_i[17];
  assign data_masked[1148] = data_i[1148] & sel_one_hot_i[17];
  assign data_masked[1147] = data_i[1147] & sel_one_hot_i[17];
  assign data_masked[1146] = data_i[1146] & sel_one_hot_i[17];
  assign data_masked[1145] = data_i[1145] & sel_one_hot_i[17];
  assign data_masked[1144] = data_i[1144] & sel_one_hot_i[17];
  assign data_masked[1143] = data_i[1143] & sel_one_hot_i[17];
  assign data_masked[1142] = data_i[1142] & sel_one_hot_i[17];
  assign data_masked[1141] = data_i[1141] & sel_one_hot_i[17];
  assign data_masked[1140] = data_i[1140] & sel_one_hot_i[17];
  assign data_masked[1139] = data_i[1139] & sel_one_hot_i[17];
  assign data_masked[1138] = data_i[1138] & sel_one_hot_i[17];
  assign data_masked[1137] = data_i[1137] & sel_one_hot_i[17];
  assign data_masked[1136] = data_i[1136] & sel_one_hot_i[17];
  assign data_masked[1135] = data_i[1135] & sel_one_hot_i[17];
  assign data_masked[1134] = data_i[1134] & sel_one_hot_i[17];
  assign data_masked[1133] = data_i[1133] & sel_one_hot_i[17];
  assign data_masked[1132] = data_i[1132] & sel_one_hot_i[17];
  assign data_masked[1131] = data_i[1131] & sel_one_hot_i[17];
  assign data_masked[1130] = data_i[1130] & sel_one_hot_i[17];
  assign data_masked[1129] = data_i[1129] & sel_one_hot_i[17];
  assign data_masked[1128] = data_i[1128] & sel_one_hot_i[17];
  assign data_masked[1127] = data_i[1127] & sel_one_hot_i[17];
  assign data_masked[1126] = data_i[1126] & sel_one_hot_i[17];
  assign data_masked[1125] = data_i[1125] & sel_one_hot_i[17];
  assign data_masked[1124] = data_i[1124] & sel_one_hot_i[17];
  assign data_masked[1123] = data_i[1123] & sel_one_hot_i[17];
  assign data_masked[1122] = data_i[1122] & sel_one_hot_i[17];
  assign data_masked[1121] = data_i[1121] & sel_one_hot_i[17];
  assign data_masked[1120] = data_i[1120] & sel_one_hot_i[17];
  assign data_masked[1119] = data_i[1119] & sel_one_hot_i[17];
  assign data_masked[1118] = data_i[1118] & sel_one_hot_i[17];
  assign data_masked[1117] = data_i[1117] & sel_one_hot_i[17];
  assign data_masked[1116] = data_i[1116] & sel_one_hot_i[17];
  assign data_masked[1115] = data_i[1115] & sel_one_hot_i[17];
  assign data_masked[1114] = data_i[1114] & sel_one_hot_i[17];
  assign data_masked[1113] = data_i[1113] & sel_one_hot_i[17];
  assign data_masked[1112] = data_i[1112] & sel_one_hot_i[17];
  assign data_masked[1111] = data_i[1111] & sel_one_hot_i[17];
  assign data_masked[1110] = data_i[1110] & sel_one_hot_i[17];
  assign data_masked[1109] = data_i[1109] & sel_one_hot_i[17];
  assign data_masked[1108] = data_i[1108] & sel_one_hot_i[17];
  assign data_masked[1107] = data_i[1107] & sel_one_hot_i[17];
  assign data_masked[1106] = data_i[1106] & sel_one_hot_i[17];
  assign data_masked[1105] = data_i[1105] & sel_one_hot_i[17];
  assign data_masked[1104] = data_i[1104] & sel_one_hot_i[17];
  assign data_masked[1103] = data_i[1103] & sel_one_hot_i[17];
  assign data_masked[1102] = data_i[1102] & sel_one_hot_i[17];
  assign data_masked[1101] = data_i[1101] & sel_one_hot_i[17];
  assign data_masked[1100] = data_i[1100] & sel_one_hot_i[17];
  assign data_masked[1099] = data_i[1099] & sel_one_hot_i[17];
  assign data_masked[1098] = data_i[1098] & sel_one_hot_i[17];
  assign data_masked[1097] = data_i[1097] & sel_one_hot_i[17];
  assign data_masked[1096] = data_i[1096] & sel_one_hot_i[17];
  assign data_masked[1095] = data_i[1095] & sel_one_hot_i[17];
  assign data_masked[1094] = data_i[1094] & sel_one_hot_i[17];
  assign data_masked[1093] = data_i[1093] & sel_one_hot_i[17];
  assign data_masked[1092] = data_i[1092] & sel_one_hot_i[17];
  assign data_masked[1091] = data_i[1091] & sel_one_hot_i[17];
  assign data_masked[1090] = data_i[1090] & sel_one_hot_i[17];
  assign data_masked[1089] = data_i[1089] & sel_one_hot_i[17];
  assign data_masked[1088] = data_i[1088] & sel_one_hot_i[17];
  assign data_masked[1215] = data_i[1215] & sel_one_hot_i[18];
  assign data_masked[1214] = data_i[1214] & sel_one_hot_i[18];
  assign data_masked[1213] = data_i[1213] & sel_one_hot_i[18];
  assign data_masked[1212] = data_i[1212] & sel_one_hot_i[18];
  assign data_masked[1211] = data_i[1211] & sel_one_hot_i[18];
  assign data_masked[1210] = data_i[1210] & sel_one_hot_i[18];
  assign data_masked[1209] = data_i[1209] & sel_one_hot_i[18];
  assign data_masked[1208] = data_i[1208] & sel_one_hot_i[18];
  assign data_masked[1207] = data_i[1207] & sel_one_hot_i[18];
  assign data_masked[1206] = data_i[1206] & sel_one_hot_i[18];
  assign data_masked[1205] = data_i[1205] & sel_one_hot_i[18];
  assign data_masked[1204] = data_i[1204] & sel_one_hot_i[18];
  assign data_masked[1203] = data_i[1203] & sel_one_hot_i[18];
  assign data_masked[1202] = data_i[1202] & sel_one_hot_i[18];
  assign data_masked[1201] = data_i[1201] & sel_one_hot_i[18];
  assign data_masked[1200] = data_i[1200] & sel_one_hot_i[18];
  assign data_masked[1199] = data_i[1199] & sel_one_hot_i[18];
  assign data_masked[1198] = data_i[1198] & sel_one_hot_i[18];
  assign data_masked[1197] = data_i[1197] & sel_one_hot_i[18];
  assign data_masked[1196] = data_i[1196] & sel_one_hot_i[18];
  assign data_masked[1195] = data_i[1195] & sel_one_hot_i[18];
  assign data_masked[1194] = data_i[1194] & sel_one_hot_i[18];
  assign data_masked[1193] = data_i[1193] & sel_one_hot_i[18];
  assign data_masked[1192] = data_i[1192] & sel_one_hot_i[18];
  assign data_masked[1191] = data_i[1191] & sel_one_hot_i[18];
  assign data_masked[1190] = data_i[1190] & sel_one_hot_i[18];
  assign data_masked[1189] = data_i[1189] & sel_one_hot_i[18];
  assign data_masked[1188] = data_i[1188] & sel_one_hot_i[18];
  assign data_masked[1187] = data_i[1187] & sel_one_hot_i[18];
  assign data_masked[1186] = data_i[1186] & sel_one_hot_i[18];
  assign data_masked[1185] = data_i[1185] & sel_one_hot_i[18];
  assign data_masked[1184] = data_i[1184] & sel_one_hot_i[18];
  assign data_masked[1183] = data_i[1183] & sel_one_hot_i[18];
  assign data_masked[1182] = data_i[1182] & sel_one_hot_i[18];
  assign data_masked[1181] = data_i[1181] & sel_one_hot_i[18];
  assign data_masked[1180] = data_i[1180] & sel_one_hot_i[18];
  assign data_masked[1179] = data_i[1179] & sel_one_hot_i[18];
  assign data_masked[1178] = data_i[1178] & sel_one_hot_i[18];
  assign data_masked[1177] = data_i[1177] & sel_one_hot_i[18];
  assign data_masked[1176] = data_i[1176] & sel_one_hot_i[18];
  assign data_masked[1175] = data_i[1175] & sel_one_hot_i[18];
  assign data_masked[1174] = data_i[1174] & sel_one_hot_i[18];
  assign data_masked[1173] = data_i[1173] & sel_one_hot_i[18];
  assign data_masked[1172] = data_i[1172] & sel_one_hot_i[18];
  assign data_masked[1171] = data_i[1171] & sel_one_hot_i[18];
  assign data_masked[1170] = data_i[1170] & sel_one_hot_i[18];
  assign data_masked[1169] = data_i[1169] & sel_one_hot_i[18];
  assign data_masked[1168] = data_i[1168] & sel_one_hot_i[18];
  assign data_masked[1167] = data_i[1167] & sel_one_hot_i[18];
  assign data_masked[1166] = data_i[1166] & sel_one_hot_i[18];
  assign data_masked[1165] = data_i[1165] & sel_one_hot_i[18];
  assign data_masked[1164] = data_i[1164] & sel_one_hot_i[18];
  assign data_masked[1163] = data_i[1163] & sel_one_hot_i[18];
  assign data_masked[1162] = data_i[1162] & sel_one_hot_i[18];
  assign data_masked[1161] = data_i[1161] & sel_one_hot_i[18];
  assign data_masked[1160] = data_i[1160] & sel_one_hot_i[18];
  assign data_masked[1159] = data_i[1159] & sel_one_hot_i[18];
  assign data_masked[1158] = data_i[1158] & sel_one_hot_i[18];
  assign data_masked[1157] = data_i[1157] & sel_one_hot_i[18];
  assign data_masked[1156] = data_i[1156] & sel_one_hot_i[18];
  assign data_masked[1155] = data_i[1155] & sel_one_hot_i[18];
  assign data_masked[1154] = data_i[1154] & sel_one_hot_i[18];
  assign data_masked[1153] = data_i[1153] & sel_one_hot_i[18];
  assign data_masked[1152] = data_i[1152] & sel_one_hot_i[18];
  assign data_masked[1279] = data_i[1279] & sel_one_hot_i[19];
  assign data_masked[1278] = data_i[1278] & sel_one_hot_i[19];
  assign data_masked[1277] = data_i[1277] & sel_one_hot_i[19];
  assign data_masked[1276] = data_i[1276] & sel_one_hot_i[19];
  assign data_masked[1275] = data_i[1275] & sel_one_hot_i[19];
  assign data_masked[1274] = data_i[1274] & sel_one_hot_i[19];
  assign data_masked[1273] = data_i[1273] & sel_one_hot_i[19];
  assign data_masked[1272] = data_i[1272] & sel_one_hot_i[19];
  assign data_masked[1271] = data_i[1271] & sel_one_hot_i[19];
  assign data_masked[1270] = data_i[1270] & sel_one_hot_i[19];
  assign data_masked[1269] = data_i[1269] & sel_one_hot_i[19];
  assign data_masked[1268] = data_i[1268] & sel_one_hot_i[19];
  assign data_masked[1267] = data_i[1267] & sel_one_hot_i[19];
  assign data_masked[1266] = data_i[1266] & sel_one_hot_i[19];
  assign data_masked[1265] = data_i[1265] & sel_one_hot_i[19];
  assign data_masked[1264] = data_i[1264] & sel_one_hot_i[19];
  assign data_masked[1263] = data_i[1263] & sel_one_hot_i[19];
  assign data_masked[1262] = data_i[1262] & sel_one_hot_i[19];
  assign data_masked[1261] = data_i[1261] & sel_one_hot_i[19];
  assign data_masked[1260] = data_i[1260] & sel_one_hot_i[19];
  assign data_masked[1259] = data_i[1259] & sel_one_hot_i[19];
  assign data_masked[1258] = data_i[1258] & sel_one_hot_i[19];
  assign data_masked[1257] = data_i[1257] & sel_one_hot_i[19];
  assign data_masked[1256] = data_i[1256] & sel_one_hot_i[19];
  assign data_masked[1255] = data_i[1255] & sel_one_hot_i[19];
  assign data_masked[1254] = data_i[1254] & sel_one_hot_i[19];
  assign data_masked[1253] = data_i[1253] & sel_one_hot_i[19];
  assign data_masked[1252] = data_i[1252] & sel_one_hot_i[19];
  assign data_masked[1251] = data_i[1251] & sel_one_hot_i[19];
  assign data_masked[1250] = data_i[1250] & sel_one_hot_i[19];
  assign data_masked[1249] = data_i[1249] & sel_one_hot_i[19];
  assign data_masked[1248] = data_i[1248] & sel_one_hot_i[19];
  assign data_masked[1247] = data_i[1247] & sel_one_hot_i[19];
  assign data_masked[1246] = data_i[1246] & sel_one_hot_i[19];
  assign data_masked[1245] = data_i[1245] & sel_one_hot_i[19];
  assign data_masked[1244] = data_i[1244] & sel_one_hot_i[19];
  assign data_masked[1243] = data_i[1243] & sel_one_hot_i[19];
  assign data_masked[1242] = data_i[1242] & sel_one_hot_i[19];
  assign data_masked[1241] = data_i[1241] & sel_one_hot_i[19];
  assign data_masked[1240] = data_i[1240] & sel_one_hot_i[19];
  assign data_masked[1239] = data_i[1239] & sel_one_hot_i[19];
  assign data_masked[1238] = data_i[1238] & sel_one_hot_i[19];
  assign data_masked[1237] = data_i[1237] & sel_one_hot_i[19];
  assign data_masked[1236] = data_i[1236] & sel_one_hot_i[19];
  assign data_masked[1235] = data_i[1235] & sel_one_hot_i[19];
  assign data_masked[1234] = data_i[1234] & sel_one_hot_i[19];
  assign data_masked[1233] = data_i[1233] & sel_one_hot_i[19];
  assign data_masked[1232] = data_i[1232] & sel_one_hot_i[19];
  assign data_masked[1231] = data_i[1231] & sel_one_hot_i[19];
  assign data_masked[1230] = data_i[1230] & sel_one_hot_i[19];
  assign data_masked[1229] = data_i[1229] & sel_one_hot_i[19];
  assign data_masked[1228] = data_i[1228] & sel_one_hot_i[19];
  assign data_masked[1227] = data_i[1227] & sel_one_hot_i[19];
  assign data_masked[1226] = data_i[1226] & sel_one_hot_i[19];
  assign data_masked[1225] = data_i[1225] & sel_one_hot_i[19];
  assign data_masked[1224] = data_i[1224] & sel_one_hot_i[19];
  assign data_masked[1223] = data_i[1223] & sel_one_hot_i[19];
  assign data_masked[1222] = data_i[1222] & sel_one_hot_i[19];
  assign data_masked[1221] = data_i[1221] & sel_one_hot_i[19];
  assign data_masked[1220] = data_i[1220] & sel_one_hot_i[19];
  assign data_masked[1219] = data_i[1219] & sel_one_hot_i[19];
  assign data_masked[1218] = data_i[1218] & sel_one_hot_i[19];
  assign data_masked[1217] = data_i[1217] & sel_one_hot_i[19];
  assign data_masked[1216] = data_i[1216] & sel_one_hot_i[19];
  assign data_masked[1343] = data_i[1343] & sel_one_hot_i[20];
  assign data_masked[1342] = data_i[1342] & sel_one_hot_i[20];
  assign data_masked[1341] = data_i[1341] & sel_one_hot_i[20];
  assign data_masked[1340] = data_i[1340] & sel_one_hot_i[20];
  assign data_masked[1339] = data_i[1339] & sel_one_hot_i[20];
  assign data_masked[1338] = data_i[1338] & sel_one_hot_i[20];
  assign data_masked[1337] = data_i[1337] & sel_one_hot_i[20];
  assign data_masked[1336] = data_i[1336] & sel_one_hot_i[20];
  assign data_masked[1335] = data_i[1335] & sel_one_hot_i[20];
  assign data_masked[1334] = data_i[1334] & sel_one_hot_i[20];
  assign data_masked[1333] = data_i[1333] & sel_one_hot_i[20];
  assign data_masked[1332] = data_i[1332] & sel_one_hot_i[20];
  assign data_masked[1331] = data_i[1331] & sel_one_hot_i[20];
  assign data_masked[1330] = data_i[1330] & sel_one_hot_i[20];
  assign data_masked[1329] = data_i[1329] & sel_one_hot_i[20];
  assign data_masked[1328] = data_i[1328] & sel_one_hot_i[20];
  assign data_masked[1327] = data_i[1327] & sel_one_hot_i[20];
  assign data_masked[1326] = data_i[1326] & sel_one_hot_i[20];
  assign data_masked[1325] = data_i[1325] & sel_one_hot_i[20];
  assign data_masked[1324] = data_i[1324] & sel_one_hot_i[20];
  assign data_masked[1323] = data_i[1323] & sel_one_hot_i[20];
  assign data_masked[1322] = data_i[1322] & sel_one_hot_i[20];
  assign data_masked[1321] = data_i[1321] & sel_one_hot_i[20];
  assign data_masked[1320] = data_i[1320] & sel_one_hot_i[20];
  assign data_masked[1319] = data_i[1319] & sel_one_hot_i[20];
  assign data_masked[1318] = data_i[1318] & sel_one_hot_i[20];
  assign data_masked[1317] = data_i[1317] & sel_one_hot_i[20];
  assign data_masked[1316] = data_i[1316] & sel_one_hot_i[20];
  assign data_masked[1315] = data_i[1315] & sel_one_hot_i[20];
  assign data_masked[1314] = data_i[1314] & sel_one_hot_i[20];
  assign data_masked[1313] = data_i[1313] & sel_one_hot_i[20];
  assign data_masked[1312] = data_i[1312] & sel_one_hot_i[20];
  assign data_masked[1311] = data_i[1311] & sel_one_hot_i[20];
  assign data_masked[1310] = data_i[1310] & sel_one_hot_i[20];
  assign data_masked[1309] = data_i[1309] & sel_one_hot_i[20];
  assign data_masked[1308] = data_i[1308] & sel_one_hot_i[20];
  assign data_masked[1307] = data_i[1307] & sel_one_hot_i[20];
  assign data_masked[1306] = data_i[1306] & sel_one_hot_i[20];
  assign data_masked[1305] = data_i[1305] & sel_one_hot_i[20];
  assign data_masked[1304] = data_i[1304] & sel_one_hot_i[20];
  assign data_masked[1303] = data_i[1303] & sel_one_hot_i[20];
  assign data_masked[1302] = data_i[1302] & sel_one_hot_i[20];
  assign data_masked[1301] = data_i[1301] & sel_one_hot_i[20];
  assign data_masked[1300] = data_i[1300] & sel_one_hot_i[20];
  assign data_masked[1299] = data_i[1299] & sel_one_hot_i[20];
  assign data_masked[1298] = data_i[1298] & sel_one_hot_i[20];
  assign data_masked[1297] = data_i[1297] & sel_one_hot_i[20];
  assign data_masked[1296] = data_i[1296] & sel_one_hot_i[20];
  assign data_masked[1295] = data_i[1295] & sel_one_hot_i[20];
  assign data_masked[1294] = data_i[1294] & sel_one_hot_i[20];
  assign data_masked[1293] = data_i[1293] & sel_one_hot_i[20];
  assign data_masked[1292] = data_i[1292] & sel_one_hot_i[20];
  assign data_masked[1291] = data_i[1291] & sel_one_hot_i[20];
  assign data_masked[1290] = data_i[1290] & sel_one_hot_i[20];
  assign data_masked[1289] = data_i[1289] & sel_one_hot_i[20];
  assign data_masked[1288] = data_i[1288] & sel_one_hot_i[20];
  assign data_masked[1287] = data_i[1287] & sel_one_hot_i[20];
  assign data_masked[1286] = data_i[1286] & sel_one_hot_i[20];
  assign data_masked[1285] = data_i[1285] & sel_one_hot_i[20];
  assign data_masked[1284] = data_i[1284] & sel_one_hot_i[20];
  assign data_masked[1283] = data_i[1283] & sel_one_hot_i[20];
  assign data_masked[1282] = data_i[1282] & sel_one_hot_i[20];
  assign data_masked[1281] = data_i[1281] & sel_one_hot_i[20];
  assign data_masked[1280] = data_i[1280] & sel_one_hot_i[20];
  assign data_masked[1407] = data_i[1407] & sel_one_hot_i[21];
  assign data_masked[1406] = data_i[1406] & sel_one_hot_i[21];
  assign data_masked[1405] = data_i[1405] & sel_one_hot_i[21];
  assign data_masked[1404] = data_i[1404] & sel_one_hot_i[21];
  assign data_masked[1403] = data_i[1403] & sel_one_hot_i[21];
  assign data_masked[1402] = data_i[1402] & sel_one_hot_i[21];
  assign data_masked[1401] = data_i[1401] & sel_one_hot_i[21];
  assign data_masked[1400] = data_i[1400] & sel_one_hot_i[21];
  assign data_masked[1399] = data_i[1399] & sel_one_hot_i[21];
  assign data_masked[1398] = data_i[1398] & sel_one_hot_i[21];
  assign data_masked[1397] = data_i[1397] & sel_one_hot_i[21];
  assign data_masked[1396] = data_i[1396] & sel_one_hot_i[21];
  assign data_masked[1395] = data_i[1395] & sel_one_hot_i[21];
  assign data_masked[1394] = data_i[1394] & sel_one_hot_i[21];
  assign data_masked[1393] = data_i[1393] & sel_one_hot_i[21];
  assign data_masked[1392] = data_i[1392] & sel_one_hot_i[21];
  assign data_masked[1391] = data_i[1391] & sel_one_hot_i[21];
  assign data_masked[1390] = data_i[1390] & sel_one_hot_i[21];
  assign data_masked[1389] = data_i[1389] & sel_one_hot_i[21];
  assign data_masked[1388] = data_i[1388] & sel_one_hot_i[21];
  assign data_masked[1387] = data_i[1387] & sel_one_hot_i[21];
  assign data_masked[1386] = data_i[1386] & sel_one_hot_i[21];
  assign data_masked[1385] = data_i[1385] & sel_one_hot_i[21];
  assign data_masked[1384] = data_i[1384] & sel_one_hot_i[21];
  assign data_masked[1383] = data_i[1383] & sel_one_hot_i[21];
  assign data_masked[1382] = data_i[1382] & sel_one_hot_i[21];
  assign data_masked[1381] = data_i[1381] & sel_one_hot_i[21];
  assign data_masked[1380] = data_i[1380] & sel_one_hot_i[21];
  assign data_masked[1379] = data_i[1379] & sel_one_hot_i[21];
  assign data_masked[1378] = data_i[1378] & sel_one_hot_i[21];
  assign data_masked[1377] = data_i[1377] & sel_one_hot_i[21];
  assign data_masked[1376] = data_i[1376] & sel_one_hot_i[21];
  assign data_masked[1375] = data_i[1375] & sel_one_hot_i[21];
  assign data_masked[1374] = data_i[1374] & sel_one_hot_i[21];
  assign data_masked[1373] = data_i[1373] & sel_one_hot_i[21];
  assign data_masked[1372] = data_i[1372] & sel_one_hot_i[21];
  assign data_masked[1371] = data_i[1371] & sel_one_hot_i[21];
  assign data_masked[1370] = data_i[1370] & sel_one_hot_i[21];
  assign data_masked[1369] = data_i[1369] & sel_one_hot_i[21];
  assign data_masked[1368] = data_i[1368] & sel_one_hot_i[21];
  assign data_masked[1367] = data_i[1367] & sel_one_hot_i[21];
  assign data_masked[1366] = data_i[1366] & sel_one_hot_i[21];
  assign data_masked[1365] = data_i[1365] & sel_one_hot_i[21];
  assign data_masked[1364] = data_i[1364] & sel_one_hot_i[21];
  assign data_masked[1363] = data_i[1363] & sel_one_hot_i[21];
  assign data_masked[1362] = data_i[1362] & sel_one_hot_i[21];
  assign data_masked[1361] = data_i[1361] & sel_one_hot_i[21];
  assign data_masked[1360] = data_i[1360] & sel_one_hot_i[21];
  assign data_masked[1359] = data_i[1359] & sel_one_hot_i[21];
  assign data_masked[1358] = data_i[1358] & sel_one_hot_i[21];
  assign data_masked[1357] = data_i[1357] & sel_one_hot_i[21];
  assign data_masked[1356] = data_i[1356] & sel_one_hot_i[21];
  assign data_masked[1355] = data_i[1355] & sel_one_hot_i[21];
  assign data_masked[1354] = data_i[1354] & sel_one_hot_i[21];
  assign data_masked[1353] = data_i[1353] & sel_one_hot_i[21];
  assign data_masked[1352] = data_i[1352] & sel_one_hot_i[21];
  assign data_masked[1351] = data_i[1351] & sel_one_hot_i[21];
  assign data_masked[1350] = data_i[1350] & sel_one_hot_i[21];
  assign data_masked[1349] = data_i[1349] & sel_one_hot_i[21];
  assign data_masked[1348] = data_i[1348] & sel_one_hot_i[21];
  assign data_masked[1347] = data_i[1347] & sel_one_hot_i[21];
  assign data_masked[1346] = data_i[1346] & sel_one_hot_i[21];
  assign data_masked[1345] = data_i[1345] & sel_one_hot_i[21];
  assign data_masked[1344] = data_i[1344] & sel_one_hot_i[21];
  assign data_masked[1471] = data_i[1471] & sel_one_hot_i[22];
  assign data_masked[1470] = data_i[1470] & sel_one_hot_i[22];
  assign data_masked[1469] = data_i[1469] & sel_one_hot_i[22];
  assign data_masked[1468] = data_i[1468] & sel_one_hot_i[22];
  assign data_masked[1467] = data_i[1467] & sel_one_hot_i[22];
  assign data_masked[1466] = data_i[1466] & sel_one_hot_i[22];
  assign data_masked[1465] = data_i[1465] & sel_one_hot_i[22];
  assign data_masked[1464] = data_i[1464] & sel_one_hot_i[22];
  assign data_masked[1463] = data_i[1463] & sel_one_hot_i[22];
  assign data_masked[1462] = data_i[1462] & sel_one_hot_i[22];
  assign data_masked[1461] = data_i[1461] & sel_one_hot_i[22];
  assign data_masked[1460] = data_i[1460] & sel_one_hot_i[22];
  assign data_masked[1459] = data_i[1459] & sel_one_hot_i[22];
  assign data_masked[1458] = data_i[1458] & sel_one_hot_i[22];
  assign data_masked[1457] = data_i[1457] & sel_one_hot_i[22];
  assign data_masked[1456] = data_i[1456] & sel_one_hot_i[22];
  assign data_masked[1455] = data_i[1455] & sel_one_hot_i[22];
  assign data_masked[1454] = data_i[1454] & sel_one_hot_i[22];
  assign data_masked[1453] = data_i[1453] & sel_one_hot_i[22];
  assign data_masked[1452] = data_i[1452] & sel_one_hot_i[22];
  assign data_masked[1451] = data_i[1451] & sel_one_hot_i[22];
  assign data_masked[1450] = data_i[1450] & sel_one_hot_i[22];
  assign data_masked[1449] = data_i[1449] & sel_one_hot_i[22];
  assign data_masked[1448] = data_i[1448] & sel_one_hot_i[22];
  assign data_masked[1447] = data_i[1447] & sel_one_hot_i[22];
  assign data_masked[1446] = data_i[1446] & sel_one_hot_i[22];
  assign data_masked[1445] = data_i[1445] & sel_one_hot_i[22];
  assign data_masked[1444] = data_i[1444] & sel_one_hot_i[22];
  assign data_masked[1443] = data_i[1443] & sel_one_hot_i[22];
  assign data_masked[1442] = data_i[1442] & sel_one_hot_i[22];
  assign data_masked[1441] = data_i[1441] & sel_one_hot_i[22];
  assign data_masked[1440] = data_i[1440] & sel_one_hot_i[22];
  assign data_masked[1439] = data_i[1439] & sel_one_hot_i[22];
  assign data_masked[1438] = data_i[1438] & sel_one_hot_i[22];
  assign data_masked[1437] = data_i[1437] & sel_one_hot_i[22];
  assign data_masked[1436] = data_i[1436] & sel_one_hot_i[22];
  assign data_masked[1435] = data_i[1435] & sel_one_hot_i[22];
  assign data_masked[1434] = data_i[1434] & sel_one_hot_i[22];
  assign data_masked[1433] = data_i[1433] & sel_one_hot_i[22];
  assign data_masked[1432] = data_i[1432] & sel_one_hot_i[22];
  assign data_masked[1431] = data_i[1431] & sel_one_hot_i[22];
  assign data_masked[1430] = data_i[1430] & sel_one_hot_i[22];
  assign data_masked[1429] = data_i[1429] & sel_one_hot_i[22];
  assign data_masked[1428] = data_i[1428] & sel_one_hot_i[22];
  assign data_masked[1427] = data_i[1427] & sel_one_hot_i[22];
  assign data_masked[1426] = data_i[1426] & sel_one_hot_i[22];
  assign data_masked[1425] = data_i[1425] & sel_one_hot_i[22];
  assign data_masked[1424] = data_i[1424] & sel_one_hot_i[22];
  assign data_masked[1423] = data_i[1423] & sel_one_hot_i[22];
  assign data_masked[1422] = data_i[1422] & sel_one_hot_i[22];
  assign data_masked[1421] = data_i[1421] & sel_one_hot_i[22];
  assign data_masked[1420] = data_i[1420] & sel_one_hot_i[22];
  assign data_masked[1419] = data_i[1419] & sel_one_hot_i[22];
  assign data_masked[1418] = data_i[1418] & sel_one_hot_i[22];
  assign data_masked[1417] = data_i[1417] & sel_one_hot_i[22];
  assign data_masked[1416] = data_i[1416] & sel_one_hot_i[22];
  assign data_masked[1415] = data_i[1415] & sel_one_hot_i[22];
  assign data_masked[1414] = data_i[1414] & sel_one_hot_i[22];
  assign data_masked[1413] = data_i[1413] & sel_one_hot_i[22];
  assign data_masked[1412] = data_i[1412] & sel_one_hot_i[22];
  assign data_masked[1411] = data_i[1411] & sel_one_hot_i[22];
  assign data_masked[1410] = data_i[1410] & sel_one_hot_i[22];
  assign data_masked[1409] = data_i[1409] & sel_one_hot_i[22];
  assign data_masked[1408] = data_i[1408] & sel_one_hot_i[22];
  assign data_masked[1535] = data_i[1535] & sel_one_hot_i[23];
  assign data_masked[1534] = data_i[1534] & sel_one_hot_i[23];
  assign data_masked[1533] = data_i[1533] & sel_one_hot_i[23];
  assign data_masked[1532] = data_i[1532] & sel_one_hot_i[23];
  assign data_masked[1531] = data_i[1531] & sel_one_hot_i[23];
  assign data_masked[1530] = data_i[1530] & sel_one_hot_i[23];
  assign data_masked[1529] = data_i[1529] & sel_one_hot_i[23];
  assign data_masked[1528] = data_i[1528] & sel_one_hot_i[23];
  assign data_masked[1527] = data_i[1527] & sel_one_hot_i[23];
  assign data_masked[1526] = data_i[1526] & sel_one_hot_i[23];
  assign data_masked[1525] = data_i[1525] & sel_one_hot_i[23];
  assign data_masked[1524] = data_i[1524] & sel_one_hot_i[23];
  assign data_masked[1523] = data_i[1523] & sel_one_hot_i[23];
  assign data_masked[1522] = data_i[1522] & sel_one_hot_i[23];
  assign data_masked[1521] = data_i[1521] & sel_one_hot_i[23];
  assign data_masked[1520] = data_i[1520] & sel_one_hot_i[23];
  assign data_masked[1519] = data_i[1519] & sel_one_hot_i[23];
  assign data_masked[1518] = data_i[1518] & sel_one_hot_i[23];
  assign data_masked[1517] = data_i[1517] & sel_one_hot_i[23];
  assign data_masked[1516] = data_i[1516] & sel_one_hot_i[23];
  assign data_masked[1515] = data_i[1515] & sel_one_hot_i[23];
  assign data_masked[1514] = data_i[1514] & sel_one_hot_i[23];
  assign data_masked[1513] = data_i[1513] & sel_one_hot_i[23];
  assign data_masked[1512] = data_i[1512] & sel_one_hot_i[23];
  assign data_masked[1511] = data_i[1511] & sel_one_hot_i[23];
  assign data_masked[1510] = data_i[1510] & sel_one_hot_i[23];
  assign data_masked[1509] = data_i[1509] & sel_one_hot_i[23];
  assign data_masked[1508] = data_i[1508] & sel_one_hot_i[23];
  assign data_masked[1507] = data_i[1507] & sel_one_hot_i[23];
  assign data_masked[1506] = data_i[1506] & sel_one_hot_i[23];
  assign data_masked[1505] = data_i[1505] & sel_one_hot_i[23];
  assign data_masked[1504] = data_i[1504] & sel_one_hot_i[23];
  assign data_masked[1503] = data_i[1503] & sel_one_hot_i[23];
  assign data_masked[1502] = data_i[1502] & sel_one_hot_i[23];
  assign data_masked[1501] = data_i[1501] & sel_one_hot_i[23];
  assign data_masked[1500] = data_i[1500] & sel_one_hot_i[23];
  assign data_masked[1499] = data_i[1499] & sel_one_hot_i[23];
  assign data_masked[1498] = data_i[1498] & sel_one_hot_i[23];
  assign data_masked[1497] = data_i[1497] & sel_one_hot_i[23];
  assign data_masked[1496] = data_i[1496] & sel_one_hot_i[23];
  assign data_masked[1495] = data_i[1495] & sel_one_hot_i[23];
  assign data_masked[1494] = data_i[1494] & sel_one_hot_i[23];
  assign data_masked[1493] = data_i[1493] & sel_one_hot_i[23];
  assign data_masked[1492] = data_i[1492] & sel_one_hot_i[23];
  assign data_masked[1491] = data_i[1491] & sel_one_hot_i[23];
  assign data_masked[1490] = data_i[1490] & sel_one_hot_i[23];
  assign data_masked[1489] = data_i[1489] & sel_one_hot_i[23];
  assign data_masked[1488] = data_i[1488] & sel_one_hot_i[23];
  assign data_masked[1487] = data_i[1487] & sel_one_hot_i[23];
  assign data_masked[1486] = data_i[1486] & sel_one_hot_i[23];
  assign data_masked[1485] = data_i[1485] & sel_one_hot_i[23];
  assign data_masked[1484] = data_i[1484] & sel_one_hot_i[23];
  assign data_masked[1483] = data_i[1483] & sel_one_hot_i[23];
  assign data_masked[1482] = data_i[1482] & sel_one_hot_i[23];
  assign data_masked[1481] = data_i[1481] & sel_one_hot_i[23];
  assign data_masked[1480] = data_i[1480] & sel_one_hot_i[23];
  assign data_masked[1479] = data_i[1479] & sel_one_hot_i[23];
  assign data_masked[1478] = data_i[1478] & sel_one_hot_i[23];
  assign data_masked[1477] = data_i[1477] & sel_one_hot_i[23];
  assign data_masked[1476] = data_i[1476] & sel_one_hot_i[23];
  assign data_masked[1475] = data_i[1475] & sel_one_hot_i[23];
  assign data_masked[1474] = data_i[1474] & sel_one_hot_i[23];
  assign data_masked[1473] = data_i[1473] & sel_one_hot_i[23];
  assign data_masked[1472] = data_i[1472] & sel_one_hot_i[23];
  assign data_masked[1599] = data_i[1599] & sel_one_hot_i[24];
  assign data_masked[1598] = data_i[1598] & sel_one_hot_i[24];
  assign data_masked[1597] = data_i[1597] & sel_one_hot_i[24];
  assign data_masked[1596] = data_i[1596] & sel_one_hot_i[24];
  assign data_masked[1595] = data_i[1595] & sel_one_hot_i[24];
  assign data_masked[1594] = data_i[1594] & sel_one_hot_i[24];
  assign data_masked[1593] = data_i[1593] & sel_one_hot_i[24];
  assign data_masked[1592] = data_i[1592] & sel_one_hot_i[24];
  assign data_masked[1591] = data_i[1591] & sel_one_hot_i[24];
  assign data_masked[1590] = data_i[1590] & sel_one_hot_i[24];
  assign data_masked[1589] = data_i[1589] & sel_one_hot_i[24];
  assign data_masked[1588] = data_i[1588] & sel_one_hot_i[24];
  assign data_masked[1587] = data_i[1587] & sel_one_hot_i[24];
  assign data_masked[1586] = data_i[1586] & sel_one_hot_i[24];
  assign data_masked[1585] = data_i[1585] & sel_one_hot_i[24];
  assign data_masked[1584] = data_i[1584] & sel_one_hot_i[24];
  assign data_masked[1583] = data_i[1583] & sel_one_hot_i[24];
  assign data_masked[1582] = data_i[1582] & sel_one_hot_i[24];
  assign data_masked[1581] = data_i[1581] & sel_one_hot_i[24];
  assign data_masked[1580] = data_i[1580] & sel_one_hot_i[24];
  assign data_masked[1579] = data_i[1579] & sel_one_hot_i[24];
  assign data_masked[1578] = data_i[1578] & sel_one_hot_i[24];
  assign data_masked[1577] = data_i[1577] & sel_one_hot_i[24];
  assign data_masked[1576] = data_i[1576] & sel_one_hot_i[24];
  assign data_masked[1575] = data_i[1575] & sel_one_hot_i[24];
  assign data_masked[1574] = data_i[1574] & sel_one_hot_i[24];
  assign data_masked[1573] = data_i[1573] & sel_one_hot_i[24];
  assign data_masked[1572] = data_i[1572] & sel_one_hot_i[24];
  assign data_masked[1571] = data_i[1571] & sel_one_hot_i[24];
  assign data_masked[1570] = data_i[1570] & sel_one_hot_i[24];
  assign data_masked[1569] = data_i[1569] & sel_one_hot_i[24];
  assign data_masked[1568] = data_i[1568] & sel_one_hot_i[24];
  assign data_masked[1567] = data_i[1567] & sel_one_hot_i[24];
  assign data_masked[1566] = data_i[1566] & sel_one_hot_i[24];
  assign data_masked[1565] = data_i[1565] & sel_one_hot_i[24];
  assign data_masked[1564] = data_i[1564] & sel_one_hot_i[24];
  assign data_masked[1563] = data_i[1563] & sel_one_hot_i[24];
  assign data_masked[1562] = data_i[1562] & sel_one_hot_i[24];
  assign data_masked[1561] = data_i[1561] & sel_one_hot_i[24];
  assign data_masked[1560] = data_i[1560] & sel_one_hot_i[24];
  assign data_masked[1559] = data_i[1559] & sel_one_hot_i[24];
  assign data_masked[1558] = data_i[1558] & sel_one_hot_i[24];
  assign data_masked[1557] = data_i[1557] & sel_one_hot_i[24];
  assign data_masked[1556] = data_i[1556] & sel_one_hot_i[24];
  assign data_masked[1555] = data_i[1555] & sel_one_hot_i[24];
  assign data_masked[1554] = data_i[1554] & sel_one_hot_i[24];
  assign data_masked[1553] = data_i[1553] & sel_one_hot_i[24];
  assign data_masked[1552] = data_i[1552] & sel_one_hot_i[24];
  assign data_masked[1551] = data_i[1551] & sel_one_hot_i[24];
  assign data_masked[1550] = data_i[1550] & sel_one_hot_i[24];
  assign data_masked[1549] = data_i[1549] & sel_one_hot_i[24];
  assign data_masked[1548] = data_i[1548] & sel_one_hot_i[24];
  assign data_masked[1547] = data_i[1547] & sel_one_hot_i[24];
  assign data_masked[1546] = data_i[1546] & sel_one_hot_i[24];
  assign data_masked[1545] = data_i[1545] & sel_one_hot_i[24];
  assign data_masked[1544] = data_i[1544] & sel_one_hot_i[24];
  assign data_masked[1543] = data_i[1543] & sel_one_hot_i[24];
  assign data_masked[1542] = data_i[1542] & sel_one_hot_i[24];
  assign data_masked[1541] = data_i[1541] & sel_one_hot_i[24];
  assign data_masked[1540] = data_i[1540] & sel_one_hot_i[24];
  assign data_masked[1539] = data_i[1539] & sel_one_hot_i[24];
  assign data_masked[1538] = data_i[1538] & sel_one_hot_i[24];
  assign data_masked[1537] = data_i[1537] & sel_one_hot_i[24];
  assign data_masked[1536] = data_i[1536] & sel_one_hot_i[24];
  assign data_masked[1663] = data_i[1663] & sel_one_hot_i[25];
  assign data_masked[1662] = data_i[1662] & sel_one_hot_i[25];
  assign data_masked[1661] = data_i[1661] & sel_one_hot_i[25];
  assign data_masked[1660] = data_i[1660] & sel_one_hot_i[25];
  assign data_masked[1659] = data_i[1659] & sel_one_hot_i[25];
  assign data_masked[1658] = data_i[1658] & sel_one_hot_i[25];
  assign data_masked[1657] = data_i[1657] & sel_one_hot_i[25];
  assign data_masked[1656] = data_i[1656] & sel_one_hot_i[25];
  assign data_masked[1655] = data_i[1655] & sel_one_hot_i[25];
  assign data_masked[1654] = data_i[1654] & sel_one_hot_i[25];
  assign data_masked[1653] = data_i[1653] & sel_one_hot_i[25];
  assign data_masked[1652] = data_i[1652] & sel_one_hot_i[25];
  assign data_masked[1651] = data_i[1651] & sel_one_hot_i[25];
  assign data_masked[1650] = data_i[1650] & sel_one_hot_i[25];
  assign data_masked[1649] = data_i[1649] & sel_one_hot_i[25];
  assign data_masked[1648] = data_i[1648] & sel_one_hot_i[25];
  assign data_masked[1647] = data_i[1647] & sel_one_hot_i[25];
  assign data_masked[1646] = data_i[1646] & sel_one_hot_i[25];
  assign data_masked[1645] = data_i[1645] & sel_one_hot_i[25];
  assign data_masked[1644] = data_i[1644] & sel_one_hot_i[25];
  assign data_masked[1643] = data_i[1643] & sel_one_hot_i[25];
  assign data_masked[1642] = data_i[1642] & sel_one_hot_i[25];
  assign data_masked[1641] = data_i[1641] & sel_one_hot_i[25];
  assign data_masked[1640] = data_i[1640] & sel_one_hot_i[25];
  assign data_masked[1639] = data_i[1639] & sel_one_hot_i[25];
  assign data_masked[1638] = data_i[1638] & sel_one_hot_i[25];
  assign data_masked[1637] = data_i[1637] & sel_one_hot_i[25];
  assign data_masked[1636] = data_i[1636] & sel_one_hot_i[25];
  assign data_masked[1635] = data_i[1635] & sel_one_hot_i[25];
  assign data_masked[1634] = data_i[1634] & sel_one_hot_i[25];
  assign data_masked[1633] = data_i[1633] & sel_one_hot_i[25];
  assign data_masked[1632] = data_i[1632] & sel_one_hot_i[25];
  assign data_masked[1631] = data_i[1631] & sel_one_hot_i[25];
  assign data_masked[1630] = data_i[1630] & sel_one_hot_i[25];
  assign data_masked[1629] = data_i[1629] & sel_one_hot_i[25];
  assign data_masked[1628] = data_i[1628] & sel_one_hot_i[25];
  assign data_masked[1627] = data_i[1627] & sel_one_hot_i[25];
  assign data_masked[1626] = data_i[1626] & sel_one_hot_i[25];
  assign data_masked[1625] = data_i[1625] & sel_one_hot_i[25];
  assign data_masked[1624] = data_i[1624] & sel_one_hot_i[25];
  assign data_masked[1623] = data_i[1623] & sel_one_hot_i[25];
  assign data_masked[1622] = data_i[1622] & sel_one_hot_i[25];
  assign data_masked[1621] = data_i[1621] & sel_one_hot_i[25];
  assign data_masked[1620] = data_i[1620] & sel_one_hot_i[25];
  assign data_masked[1619] = data_i[1619] & sel_one_hot_i[25];
  assign data_masked[1618] = data_i[1618] & sel_one_hot_i[25];
  assign data_masked[1617] = data_i[1617] & sel_one_hot_i[25];
  assign data_masked[1616] = data_i[1616] & sel_one_hot_i[25];
  assign data_masked[1615] = data_i[1615] & sel_one_hot_i[25];
  assign data_masked[1614] = data_i[1614] & sel_one_hot_i[25];
  assign data_masked[1613] = data_i[1613] & sel_one_hot_i[25];
  assign data_masked[1612] = data_i[1612] & sel_one_hot_i[25];
  assign data_masked[1611] = data_i[1611] & sel_one_hot_i[25];
  assign data_masked[1610] = data_i[1610] & sel_one_hot_i[25];
  assign data_masked[1609] = data_i[1609] & sel_one_hot_i[25];
  assign data_masked[1608] = data_i[1608] & sel_one_hot_i[25];
  assign data_masked[1607] = data_i[1607] & sel_one_hot_i[25];
  assign data_masked[1606] = data_i[1606] & sel_one_hot_i[25];
  assign data_masked[1605] = data_i[1605] & sel_one_hot_i[25];
  assign data_masked[1604] = data_i[1604] & sel_one_hot_i[25];
  assign data_masked[1603] = data_i[1603] & sel_one_hot_i[25];
  assign data_masked[1602] = data_i[1602] & sel_one_hot_i[25];
  assign data_masked[1601] = data_i[1601] & sel_one_hot_i[25];
  assign data_masked[1600] = data_i[1600] & sel_one_hot_i[25];
  assign data_masked[1727] = data_i[1727] & sel_one_hot_i[26];
  assign data_masked[1726] = data_i[1726] & sel_one_hot_i[26];
  assign data_masked[1725] = data_i[1725] & sel_one_hot_i[26];
  assign data_masked[1724] = data_i[1724] & sel_one_hot_i[26];
  assign data_masked[1723] = data_i[1723] & sel_one_hot_i[26];
  assign data_masked[1722] = data_i[1722] & sel_one_hot_i[26];
  assign data_masked[1721] = data_i[1721] & sel_one_hot_i[26];
  assign data_masked[1720] = data_i[1720] & sel_one_hot_i[26];
  assign data_masked[1719] = data_i[1719] & sel_one_hot_i[26];
  assign data_masked[1718] = data_i[1718] & sel_one_hot_i[26];
  assign data_masked[1717] = data_i[1717] & sel_one_hot_i[26];
  assign data_masked[1716] = data_i[1716] & sel_one_hot_i[26];
  assign data_masked[1715] = data_i[1715] & sel_one_hot_i[26];
  assign data_masked[1714] = data_i[1714] & sel_one_hot_i[26];
  assign data_masked[1713] = data_i[1713] & sel_one_hot_i[26];
  assign data_masked[1712] = data_i[1712] & sel_one_hot_i[26];
  assign data_masked[1711] = data_i[1711] & sel_one_hot_i[26];
  assign data_masked[1710] = data_i[1710] & sel_one_hot_i[26];
  assign data_masked[1709] = data_i[1709] & sel_one_hot_i[26];
  assign data_masked[1708] = data_i[1708] & sel_one_hot_i[26];
  assign data_masked[1707] = data_i[1707] & sel_one_hot_i[26];
  assign data_masked[1706] = data_i[1706] & sel_one_hot_i[26];
  assign data_masked[1705] = data_i[1705] & sel_one_hot_i[26];
  assign data_masked[1704] = data_i[1704] & sel_one_hot_i[26];
  assign data_masked[1703] = data_i[1703] & sel_one_hot_i[26];
  assign data_masked[1702] = data_i[1702] & sel_one_hot_i[26];
  assign data_masked[1701] = data_i[1701] & sel_one_hot_i[26];
  assign data_masked[1700] = data_i[1700] & sel_one_hot_i[26];
  assign data_masked[1699] = data_i[1699] & sel_one_hot_i[26];
  assign data_masked[1698] = data_i[1698] & sel_one_hot_i[26];
  assign data_masked[1697] = data_i[1697] & sel_one_hot_i[26];
  assign data_masked[1696] = data_i[1696] & sel_one_hot_i[26];
  assign data_masked[1695] = data_i[1695] & sel_one_hot_i[26];
  assign data_masked[1694] = data_i[1694] & sel_one_hot_i[26];
  assign data_masked[1693] = data_i[1693] & sel_one_hot_i[26];
  assign data_masked[1692] = data_i[1692] & sel_one_hot_i[26];
  assign data_masked[1691] = data_i[1691] & sel_one_hot_i[26];
  assign data_masked[1690] = data_i[1690] & sel_one_hot_i[26];
  assign data_masked[1689] = data_i[1689] & sel_one_hot_i[26];
  assign data_masked[1688] = data_i[1688] & sel_one_hot_i[26];
  assign data_masked[1687] = data_i[1687] & sel_one_hot_i[26];
  assign data_masked[1686] = data_i[1686] & sel_one_hot_i[26];
  assign data_masked[1685] = data_i[1685] & sel_one_hot_i[26];
  assign data_masked[1684] = data_i[1684] & sel_one_hot_i[26];
  assign data_masked[1683] = data_i[1683] & sel_one_hot_i[26];
  assign data_masked[1682] = data_i[1682] & sel_one_hot_i[26];
  assign data_masked[1681] = data_i[1681] & sel_one_hot_i[26];
  assign data_masked[1680] = data_i[1680] & sel_one_hot_i[26];
  assign data_masked[1679] = data_i[1679] & sel_one_hot_i[26];
  assign data_masked[1678] = data_i[1678] & sel_one_hot_i[26];
  assign data_masked[1677] = data_i[1677] & sel_one_hot_i[26];
  assign data_masked[1676] = data_i[1676] & sel_one_hot_i[26];
  assign data_masked[1675] = data_i[1675] & sel_one_hot_i[26];
  assign data_masked[1674] = data_i[1674] & sel_one_hot_i[26];
  assign data_masked[1673] = data_i[1673] & sel_one_hot_i[26];
  assign data_masked[1672] = data_i[1672] & sel_one_hot_i[26];
  assign data_masked[1671] = data_i[1671] & sel_one_hot_i[26];
  assign data_masked[1670] = data_i[1670] & sel_one_hot_i[26];
  assign data_masked[1669] = data_i[1669] & sel_one_hot_i[26];
  assign data_masked[1668] = data_i[1668] & sel_one_hot_i[26];
  assign data_masked[1667] = data_i[1667] & sel_one_hot_i[26];
  assign data_masked[1666] = data_i[1666] & sel_one_hot_i[26];
  assign data_masked[1665] = data_i[1665] & sel_one_hot_i[26];
  assign data_masked[1664] = data_i[1664] & sel_one_hot_i[26];
  assign data_masked[1791] = data_i[1791] & sel_one_hot_i[27];
  assign data_masked[1790] = data_i[1790] & sel_one_hot_i[27];
  assign data_masked[1789] = data_i[1789] & sel_one_hot_i[27];
  assign data_masked[1788] = data_i[1788] & sel_one_hot_i[27];
  assign data_masked[1787] = data_i[1787] & sel_one_hot_i[27];
  assign data_masked[1786] = data_i[1786] & sel_one_hot_i[27];
  assign data_masked[1785] = data_i[1785] & sel_one_hot_i[27];
  assign data_masked[1784] = data_i[1784] & sel_one_hot_i[27];
  assign data_masked[1783] = data_i[1783] & sel_one_hot_i[27];
  assign data_masked[1782] = data_i[1782] & sel_one_hot_i[27];
  assign data_masked[1781] = data_i[1781] & sel_one_hot_i[27];
  assign data_masked[1780] = data_i[1780] & sel_one_hot_i[27];
  assign data_masked[1779] = data_i[1779] & sel_one_hot_i[27];
  assign data_masked[1778] = data_i[1778] & sel_one_hot_i[27];
  assign data_masked[1777] = data_i[1777] & sel_one_hot_i[27];
  assign data_masked[1776] = data_i[1776] & sel_one_hot_i[27];
  assign data_masked[1775] = data_i[1775] & sel_one_hot_i[27];
  assign data_masked[1774] = data_i[1774] & sel_one_hot_i[27];
  assign data_masked[1773] = data_i[1773] & sel_one_hot_i[27];
  assign data_masked[1772] = data_i[1772] & sel_one_hot_i[27];
  assign data_masked[1771] = data_i[1771] & sel_one_hot_i[27];
  assign data_masked[1770] = data_i[1770] & sel_one_hot_i[27];
  assign data_masked[1769] = data_i[1769] & sel_one_hot_i[27];
  assign data_masked[1768] = data_i[1768] & sel_one_hot_i[27];
  assign data_masked[1767] = data_i[1767] & sel_one_hot_i[27];
  assign data_masked[1766] = data_i[1766] & sel_one_hot_i[27];
  assign data_masked[1765] = data_i[1765] & sel_one_hot_i[27];
  assign data_masked[1764] = data_i[1764] & sel_one_hot_i[27];
  assign data_masked[1763] = data_i[1763] & sel_one_hot_i[27];
  assign data_masked[1762] = data_i[1762] & sel_one_hot_i[27];
  assign data_masked[1761] = data_i[1761] & sel_one_hot_i[27];
  assign data_masked[1760] = data_i[1760] & sel_one_hot_i[27];
  assign data_masked[1759] = data_i[1759] & sel_one_hot_i[27];
  assign data_masked[1758] = data_i[1758] & sel_one_hot_i[27];
  assign data_masked[1757] = data_i[1757] & sel_one_hot_i[27];
  assign data_masked[1756] = data_i[1756] & sel_one_hot_i[27];
  assign data_masked[1755] = data_i[1755] & sel_one_hot_i[27];
  assign data_masked[1754] = data_i[1754] & sel_one_hot_i[27];
  assign data_masked[1753] = data_i[1753] & sel_one_hot_i[27];
  assign data_masked[1752] = data_i[1752] & sel_one_hot_i[27];
  assign data_masked[1751] = data_i[1751] & sel_one_hot_i[27];
  assign data_masked[1750] = data_i[1750] & sel_one_hot_i[27];
  assign data_masked[1749] = data_i[1749] & sel_one_hot_i[27];
  assign data_masked[1748] = data_i[1748] & sel_one_hot_i[27];
  assign data_masked[1747] = data_i[1747] & sel_one_hot_i[27];
  assign data_masked[1746] = data_i[1746] & sel_one_hot_i[27];
  assign data_masked[1745] = data_i[1745] & sel_one_hot_i[27];
  assign data_masked[1744] = data_i[1744] & sel_one_hot_i[27];
  assign data_masked[1743] = data_i[1743] & sel_one_hot_i[27];
  assign data_masked[1742] = data_i[1742] & sel_one_hot_i[27];
  assign data_masked[1741] = data_i[1741] & sel_one_hot_i[27];
  assign data_masked[1740] = data_i[1740] & sel_one_hot_i[27];
  assign data_masked[1739] = data_i[1739] & sel_one_hot_i[27];
  assign data_masked[1738] = data_i[1738] & sel_one_hot_i[27];
  assign data_masked[1737] = data_i[1737] & sel_one_hot_i[27];
  assign data_masked[1736] = data_i[1736] & sel_one_hot_i[27];
  assign data_masked[1735] = data_i[1735] & sel_one_hot_i[27];
  assign data_masked[1734] = data_i[1734] & sel_one_hot_i[27];
  assign data_masked[1733] = data_i[1733] & sel_one_hot_i[27];
  assign data_masked[1732] = data_i[1732] & sel_one_hot_i[27];
  assign data_masked[1731] = data_i[1731] & sel_one_hot_i[27];
  assign data_masked[1730] = data_i[1730] & sel_one_hot_i[27];
  assign data_masked[1729] = data_i[1729] & sel_one_hot_i[27];
  assign data_masked[1728] = data_i[1728] & sel_one_hot_i[27];
  assign data_masked[1855] = data_i[1855] & sel_one_hot_i[28];
  assign data_masked[1854] = data_i[1854] & sel_one_hot_i[28];
  assign data_masked[1853] = data_i[1853] & sel_one_hot_i[28];
  assign data_masked[1852] = data_i[1852] & sel_one_hot_i[28];
  assign data_masked[1851] = data_i[1851] & sel_one_hot_i[28];
  assign data_masked[1850] = data_i[1850] & sel_one_hot_i[28];
  assign data_masked[1849] = data_i[1849] & sel_one_hot_i[28];
  assign data_masked[1848] = data_i[1848] & sel_one_hot_i[28];
  assign data_masked[1847] = data_i[1847] & sel_one_hot_i[28];
  assign data_masked[1846] = data_i[1846] & sel_one_hot_i[28];
  assign data_masked[1845] = data_i[1845] & sel_one_hot_i[28];
  assign data_masked[1844] = data_i[1844] & sel_one_hot_i[28];
  assign data_masked[1843] = data_i[1843] & sel_one_hot_i[28];
  assign data_masked[1842] = data_i[1842] & sel_one_hot_i[28];
  assign data_masked[1841] = data_i[1841] & sel_one_hot_i[28];
  assign data_masked[1840] = data_i[1840] & sel_one_hot_i[28];
  assign data_masked[1839] = data_i[1839] & sel_one_hot_i[28];
  assign data_masked[1838] = data_i[1838] & sel_one_hot_i[28];
  assign data_masked[1837] = data_i[1837] & sel_one_hot_i[28];
  assign data_masked[1836] = data_i[1836] & sel_one_hot_i[28];
  assign data_masked[1835] = data_i[1835] & sel_one_hot_i[28];
  assign data_masked[1834] = data_i[1834] & sel_one_hot_i[28];
  assign data_masked[1833] = data_i[1833] & sel_one_hot_i[28];
  assign data_masked[1832] = data_i[1832] & sel_one_hot_i[28];
  assign data_masked[1831] = data_i[1831] & sel_one_hot_i[28];
  assign data_masked[1830] = data_i[1830] & sel_one_hot_i[28];
  assign data_masked[1829] = data_i[1829] & sel_one_hot_i[28];
  assign data_masked[1828] = data_i[1828] & sel_one_hot_i[28];
  assign data_masked[1827] = data_i[1827] & sel_one_hot_i[28];
  assign data_masked[1826] = data_i[1826] & sel_one_hot_i[28];
  assign data_masked[1825] = data_i[1825] & sel_one_hot_i[28];
  assign data_masked[1824] = data_i[1824] & sel_one_hot_i[28];
  assign data_masked[1823] = data_i[1823] & sel_one_hot_i[28];
  assign data_masked[1822] = data_i[1822] & sel_one_hot_i[28];
  assign data_masked[1821] = data_i[1821] & sel_one_hot_i[28];
  assign data_masked[1820] = data_i[1820] & sel_one_hot_i[28];
  assign data_masked[1819] = data_i[1819] & sel_one_hot_i[28];
  assign data_masked[1818] = data_i[1818] & sel_one_hot_i[28];
  assign data_masked[1817] = data_i[1817] & sel_one_hot_i[28];
  assign data_masked[1816] = data_i[1816] & sel_one_hot_i[28];
  assign data_masked[1815] = data_i[1815] & sel_one_hot_i[28];
  assign data_masked[1814] = data_i[1814] & sel_one_hot_i[28];
  assign data_masked[1813] = data_i[1813] & sel_one_hot_i[28];
  assign data_masked[1812] = data_i[1812] & sel_one_hot_i[28];
  assign data_masked[1811] = data_i[1811] & sel_one_hot_i[28];
  assign data_masked[1810] = data_i[1810] & sel_one_hot_i[28];
  assign data_masked[1809] = data_i[1809] & sel_one_hot_i[28];
  assign data_masked[1808] = data_i[1808] & sel_one_hot_i[28];
  assign data_masked[1807] = data_i[1807] & sel_one_hot_i[28];
  assign data_masked[1806] = data_i[1806] & sel_one_hot_i[28];
  assign data_masked[1805] = data_i[1805] & sel_one_hot_i[28];
  assign data_masked[1804] = data_i[1804] & sel_one_hot_i[28];
  assign data_masked[1803] = data_i[1803] & sel_one_hot_i[28];
  assign data_masked[1802] = data_i[1802] & sel_one_hot_i[28];
  assign data_masked[1801] = data_i[1801] & sel_one_hot_i[28];
  assign data_masked[1800] = data_i[1800] & sel_one_hot_i[28];
  assign data_masked[1799] = data_i[1799] & sel_one_hot_i[28];
  assign data_masked[1798] = data_i[1798] & sel_one_hot_i[28];
  assign data_masked[1797] = data_i[1797] & sel_one_hot_i[28];
  assign data_masked[1796] = data_i[1796] & sel_one_hot_i[28];
  assign data_masked[1795] = data_i[1795] & sel_one_hot_i[28];
  assign data_masked[1794] = data_i[1794] & sel_one_hot_i[28];
  assign data_masked[1793] = data_i[1793] & sel_one_hot_i[28];
  assign data_masked[1792] = data_i[1792] & sel_one_hot_i[28];
  assign data_masked[1919] = data_i[1919] & sel_one_hot_i[29];
  assign data_masked[1918] = data_i[1918] & sel_one_hot_i[29];
  assign data_masked[1917] = data_i[1917] & sel_one_hot_i[29];
  assign data_masked[1916] = data_i[1916] & sel_one_hot_i[29];
  assign data_masked[1915] = data_i[1915] & sel_one_hot_i[29];
  assign data_masked[1914] = data_i[1914] & sel_one_hot_i[29];
  assign data_masked[1913] = data_i[1913] & sel_one_hot_i[29];
  assign data_masked[1912] = data_i[1912] & sel_one_hot_i[29];
  assign data_masked[1911] = data_i[1911] & sel_one_hot_i[29];
  assign data_masked[1910] = data_i[1910] & sel_one_hot_i[29];
  assign data_masked[1909] = data_i[1909] & sel_one_hot_i[29];
  assign data_masked[1908] = data_i[1908] & sel_one_hot_i[29];
  assign data_masked[1907] = data_i[1907] & sel_one_hot_i[29];
  assign data_masked[1906] = data_i[1906] & sel_one_hot_i[29];
  assign data_masked[1905] = data_i[1905] & sel_one_hot_i[29];
  assign data_masked[1904] = data_i[1904] & sel_one_hot_i[29];
  assign data_masked[1903] = data_i[1903] & sel_one_hot_i[29];
  assign data_masked[1902] = data_i[1902] & sel_one_hot_i[29];
  assign data_masked[1901] = data_i[1901] & sel_one_hot_i[29];
  assign data_masked[1900] = data_i[1900] & sel_one_hot_i[29];
  assign data_masked[1899] = data_i[1899] & sel_one_hot_i[29];
  assign data_masked[1898] = data_i[1898] & sel_one_hot_i[29];
  assign data_masked[1897] = data_i[1897] & sel_one_hot_i[29];
  assign data_masked[1896] = data_i[1896] & sel_one_hot_i[29];
  assign data_masked[1895] = data_i[1895] & sel_one_hot_i[29];
  assign data_masked[1894] = data_i[1894] & sel_one_hot_i[29];
  assign data_masked[1893] = data_i[1893] & sel_one_hot_i[29];
  assign data_masked[1892] = data_i[1892] & sel_one_hot_i[29];
  assign data_masked[1891] = data_i[1891] & sel_one_hot_i[29];
  assign data_masked[1890] = data_i[1890] & sel_one_hot_i[29];
  assign data_masked[1889] = data_i[1889] & sel_one_hot_i[29];
  assign data_masked[1888] = data_i[1888] & sel_one_hot_i[29];
  assign data_masked[1887] = data_i[1887] & sel_one_hot_i[29];
  assign data_masked[1886] = data_i[1886] & sel_one_hot_i[29];
  assign data_masked[1885] = data_i[1885] & sel_one_hot_i[29];
  assign data_masked[1884] = data_i[1884] & sel_one_hot_i[29];
  assign data_masked[1883] = data_i[1883] & sel_one_hot_i[29];
  assign data_masked[1882] = data_i[1882] & sel_one_hot_i[29];
  assign data_masked[1881] = data_i[1881] & sel_one_hot_i[29];
  assign data_masked[1880] = data_i[1880] & sel_one_hot_i[29];
  assign data_masked[1879] = data_i[1879] & sel_one_hot_i[29];
  assign data_masked[1878] = data_i[1878] & sel_one_hot_i[29];
  assign data_masked[1877] = data_i[1877] & sel_one_hot_i[29];
  assign data_masked[1876] = data_i[1876] & sel_one_hot_i[29];
  assign data_masked[1875] = data_i[1875] & sel_one_hot_i[29];
  assign data_masked[1874] = data_i[1874] & sel_one_hot_i[29];
  assign data_masked[1873] = data_i[1873] & sel_one_hot_i[29];
  assign data_masked[1872] = data_i[1872] & sel_one_hot_i[29];
  assign data_masked[1871] = data_i[1871] & sel_one_hot_i[29];
  assign data_masked[1870] = data_i[1870] & sel_one_hot_i[29];
  assign data_masked[1869] = data_i[1869] & sel_one_hot_i[29];
  assign data_masked[1868] = data_i[1868] & sel_one_hot_i[29];
  assign data_masked[1867] = data_i[1867] & sel_one_hot_i[29];
  assign data_masked[1866] = data_i[1866] & sel_one_hot_i[29];
  assign data_masked[1865] = data_i[1865] & sel_one_hot_i[29];
  assign data_masked[1864] = data_i[1864] & sel_one_hot_i[29];
  assign data_masked[1863] = data_i[1863] & sel_one_hot_i[29];
  assign data_masked[1862] = data_i[1862] & sel_one_hot_i[29];
  assign data_masked[1861] = data_i[1861] & sel_one_hot_i[29];
  assign data_masked[1860] = data_i[1860] & sel_one_hot_i[29];
  assign data_masked[1859] = data_i[1859] & sel_one_hot_i[29];
  assign data_masked[1858] = data_i[1858] & sel_one_hot_i[29];
  assign data_masked[1857] = data_i[1857] & sel_one_hot_i[29];
  assign data_masked[1856] = data_i[1856] & sel_one_hot_i[29];
  assign data_masked[1983] = data_i[1983] & sel_one_hot_i[30];
  assign data_masked[1982] = data_i[1982] & sel_one_hot_i[30];
  assign data_masked[1981] = data_i[1981] & sel_one_hot_i[30];
  assign data_masked[1980] = data_i[1980] & sel_one_hot_i[30];
  assign data_masked[1979] = data_i[1979] & sel_one_hot_i[30];
  assign data_masked[1978] = data_i[1978] & sel_one_hot_i[30];
  assign data_masked[1977] = data_i[1977] & sel_one_hot_i[30];
  assign data_masked[1976] = data_i[1976] & sel_one_hot_i[30];
  assign data_masked[1975] = data_i[1975] & sel_one_hot_i[30];
  assign data_masked[1974] = data_i[1974] & sel_one_hot_i[30];
  assign data_masked[1973] = data_i[1973] & sel_one_hot_i[30];
  assign data_masked[1972] = data_i[1972] & sel_one_hot_i[30];
  assign data_masked[1971] = data_i[1971] & sel_one_hot_i[30];
  assign data_masked[1970] = data_i[1970] & sel_one_hot_i[30];
  assign data_masked[1969] = data_i[1969] & sel_one_hot_i[30];
  assign data_masked[1968] = data_i[1968] & sel_one_hot_i[30];
  assign data_masked[1967] = data_i[1967] & sel_one_hot_i[30];
  assign data_masked[1966] = data_i[1966] & sel_one_hot_i[30];
  assign data_masked[1965] = data_i[1965] & sel_one_hot_i[30];
  assign data_masked[1964] = data_i[1964] & sel_one_hot_i[30];
  assign data_masked[1963] = data_i[1963] & sel_one_hot_i[30];
  assign data_masked[1962] = data_i[1962] & sel_one_hot_i[30];
  assign data_masked[1961] = data_i[1961] & sel_one_hot_i[30];
  assign data_masked[1960] = data_i[1960] & sel_one_hot_i[30];
  assign data_masked[1959] = data_i[1959] & sel_one_hot_i[30];
  assign data_masked[1958] = data_i[1958] & sel_one_hot_i[30];
  assign data_masked[1957] = data_i[1957] & sel_one_hot_i[30];
  assign data_masked[1956] = data_i[1956] & sel_one_hot_i[30];
  assign data_masked[1955] = data_i[1955] & sel_one_hot_i[30];
  assign data_masked[1954] = data_i[1954] & sel_one_hot_i[30];
  assign data_masked[1953] = data_i[1953] & sel_one_hot_i[30];
  assign data_masked[1952] = data_i[1952] & sel_one_hot_i[30];
  assign data_masked[1951] = data_i[1951] & sel_one_hot_i[30];
  assign data_masked[1950] = data_i[1950] & sel_one_hot_i[30];
  assign data_masked[1949] = data_i[1949] & sel_one_hot_i[30];
  assign data_masked[1948] = data_i[1948] & sel_one_hot_i[30];
  assign data_masked[1947] = data_i[1947] & sel_one_hot_i[30];
  assign data_masked[1946] = data_i[1946] & sel_one_hot_i[30];
  assign data_masked[1945] = data_i[1945] & sel_one_hot_i[30];
  assign data_masked[1944] = data_i[1944] & sel_one_hot_i[30];
  assign data_masked[1943] = data_i[1943] & sel_one_hot_i[30];
  assign data_masked[1942] = data_i[1942] & sel_one_hot_i[30];
  assign data_masked[1941] = data_i[1941] & sel_one_hot_i[30];
  assign data_masked[1940] = data_i[1940] & sel_one_hot_i[30];
  assign data_masked[1939] = data_i[1939] & sel_one_hot_i[30];
  assign data_masked[1938] = data_i[1938] & sel_one_hot_i[30];
  assign data_masked[1937] = data_i[1937] & sel_one_hot_i[30];
  assign data_masked[1936] = data_i[1936] & sel_one_hot_i[30];
  assign data_masked[1935] = data_i[1935] & sel_one_hot_i[30];
  assign data_masked[1934] = data_i[1934] & sel_one_hot_i[30];
  assign data_masked[1933] = data_i[1933] & sel_one_hot_i[30];
  assign data_masked[1932] = data_i[1932] & sel_one_hot_i[30];
  assign data_masked[1931] = data_i[1931] & sel_one_hot_i[30];
  assign data_masked[1930] = data_i[1930] & sel_one_hot_i[30];
  assign data_masked[1929] = data_i[1929] & sel_one_hot_i[30];
  assign data_masked[1928] = data_i[1928] & sel_one_hot_i[30];
  assign data_masked[1927] = data_i[1927] & sel_one_hot_i[30];
  assign data_masked[1926] = data_i[1926] & sel_one_hot_i[30];
  assign data_masked[1925] = data_i[1925] & sel_one_hot_i[30];
  assign data_masked[1924] = data_i[1924] & sel_one_hot_i[30];
  assign data_masked[1923] = data_i[1923] & sel_one_hot_i[30];
  assign data_masked[1922] = data_i[1922] & sel_one_hot_i[30];
  assign data_masked[1921] = data_i[1921] & sel_one_hot_i[30];
  assign data_masked[1920] = data_i[1920] & sel_one_hot_i[30];
  assign data_masked[2047] = data_i[2047] & sel_one_hot_i[31];
  assign data_masked[2046] = data_i[2046] & sel_one_hot_i[31];
  assign data_masked[2045] = data_i[2045] & sel_one_hot_i[31];
  assign data_masked[2044] = data_i[2044] & sel_one_hot_i[31];
  assign data_masked[2043] = data_i[2043] & sel_one_hot_i[31];
  assign data_masked[2042] = data_i[2042] & sel_one_hot_i[31];
  assign data_masked[2041] = data_i[2041] & sel_one_hot_i[31];
  assign data_masked[2040] = data_i[2040] & sel_one_hot_i[31];
  assign data_masked[2039] = data_i[2039] & sel_one_hot_i[31];
  assign data_masked[2038] = data_i[2038] & sel_one_hot_i[31];
  assign data_masked[2037] = data_i[2037] & sel_one_hot_i[31];
  assign data_masked[2036] = data_i[2036] & sel_one_hot_i[31];
  assign data_masked[2035] = data_i[2035] & sel_one_hot_i[31];
  assign data_masked[2034] = data_i[2034] & sel_one_hot_i[31];
  assign data_masked[2033] = data_i[2033] & sel_one_hot_i[31];
  assign data_masked[2032] = data_i[2032] & sel_one_hot_i[31];
  assign data_masked[2031] = data_i[2031] & sel_one_hot_i[31];
  assign data_masked[2030] = data_i[2030] & sel_one_hot_i[31];
  assign data_masked[2029] = data_i[2029] & sel_one_hot_i[31];
  assign data_masked[2028] = data_i[2028] & sel_one_hot_i[31];
  assign data_masked[2027] = data_i[2027] & sel_one_hot_i[31];
  assign data_masked[2026] = data_i[2026] & sel_one_hot_i[31];
  assign data_masked[2025] = data_i[2025] & sel_one_hot_i[31];
  assign data_masked[2024] = data_i[2024] & sel_one_hot_i[31];
  assign data_masked[2023] = data_i[2023] & sel_one_hot_i[31];
  assign data_masked[2022] = data_i[2022] & sel_one_hot_i[31];
  assign data_masked[2021] = data_i[2021] & sel_one_hot_i[31];
  assign data_masked[2020] = data_i[2020] & sel_one_hot_i[31];
  assign data_masked[2019] = data_i[2019] & sel_one_hot_i[31];
  assign data_masked[2018] = data_i[2018] & sel_one_hot_i[31];
  assign data_masked[2017] = data_i[2017] & sel_one_hot_i[31];
  assign data_masked[2016] = data_i[2016] & sel_one_hot_i[31];
  assign data_masked[2015] = data_i[2015] & sel_one_hot_i[31];
  assign data_masked[2014] = data_i[2014] & sel_one_hot_i[31];
  assign data_masked[2013] = data_i[2013] & sel_one_hot_i[31];
  assign data_masked[2012] = data_i[2012] & sel_one_hot_i[31];
  assign data_masked[2011] = data_i[2011] & sel_one_hot_i[31];
  assign data_masked[2010] = data_i[2010] & sel_one_hot_i[31];
  assign data_masked[2009] = data_i[2009] & sel_one_hot_i[31];
  assign data_masked[2008] = data_i[2008] & sel_one_hot_i[31];
  assign data_masked[2007] = data_i[2007] & sel_one_hot_i[31];
  assign data_masked[2006] = data_i[2006] & sel_one_hot_i[31];
  assign data_masked[2005] = data_i[2005] & sel_one_hot_i[31];
  assign data_masked[2004] = data_i[2004] & sel_one_hot_i[31];
  assign data_masked[2003] = data_i[2003] & sel_one_hot_i[31];
  assign data_masked[2002] = data_i[2002] & sel_one_hot_i[31];
  assign data_masked[2001] = data_i[2001] & sel_one_hot_i[31];
  assign data_masked[2000] = data_i[2000] & sel_one_hot_i[31];
  assign data_masked[1999] = data_i[1999] & sel_one_hot_i[31];
  assign data_masked[1998] = data_i[1998] & sel_one_hot_i[31];
  assign data_masked[1997] = data_i[1997] & sel_one_hot_i[31];
  assign data_masked[1996] = data_i[1996] & sel_one_hot_i[31];
  assign data_masked[1995] = data_i[1995] & sel_one_hot_i[31];
  assign data_masked[1994] = data_i[1994] & sel_one_hot_i[31];
  assign data_masked[1993] = data_i[1993] & sel_one_hot_i[31];
  assign data_masked[1992] = data_i[1992] & sel_one_hot_i[31];
  assign data_masked[1991] = data_i[1991] & sel_one_hot_i[31];
  assign data_masked[1990] = data_i[1990] & sel_one_hot_i[31];
  assign data_masked[1989] = data_i[1989] & sel_one_hot_i[31];
  assign data_masked[1988] = data_i[1988] & sel_one_hot_i[31];
  assign data_masked[1987] = data_i[1987] & sel_one_hot_i[31];
  assign data_masked[1986] = data_i[1986] & sel_one_hot_i[31];
  assign data_masked[1985] = data_i[1985] & sel_one_hot_i[31];
  assign data_masked[1984] = data_i[1984] & sel_one_hot_i[31];
  assign data_masked[2111] = data_i[2111] & sel_one_hot_i[32];
  assign data_masked[2110] = data_i[2110] & sel_one_hot_i[32];
  assign data_masked[2109] = data_i[2109] & sel_one_hot_i[32];
  assign data_masked[2108] = data_i[2108] & sel_one_hot_i[32];
  assign data_masked[2107] = data_i[2107] & sel_one_hot_i[32];
  assign data_masked[2106] = data_i[2106] & sel_one_hot_i[32];
  assign data_masked[2105] = data_i[2105] & sel_one_hot_i[32];
  assign data_masked[2104] = data_i[2104] & sel_one_hot_i[32];
  assign data_masked[2103] = data_i[2103] & sel_one_hot_i[32];
  assign data_masked[2102] = data_i[2102] & sel_one_hot_i[32];
  assign data_masked[2101] = data_i[2101] & sel_one_hot_i[32];
  assign data_masked[2100] = data_i[2100] & sel_one_hot_i[32];
  assign data_masked[2099] = data_i[2099] & sel_one_hot_i[32];
  assign data_masked[2098] = data_i[2098] & sel_one_hot_i[32];
  assign data_masked[2097] = data_i[2097] & sel_one_hot_i[32];
  assign data_masked[2096] = data_i[2096] & sel_one_hot_i[32];
  assign data_masked[2095] = data_i[2095] & sel_one_hot_i[32];
  assign data_masked[2094] = data_i[2094] & sel_one_hot_i[32];
  assign data_masked[2093] = data_i[2093] & sel_one_hot_i[32];
  assign data_masked[2092] = data_i[2092] & sel_one_hot_i[32];
  assign data_masked[2091] = data_i[2091] & sel_one_hot_i[32];
  assign data_masked[2090] = data_i[2090] & sel_one_hot_i[32];
  assign data_masked[2089] = data_i[2089] & sel_one_hot_i[32];
  assign data_masked[2088] = data_i[2088] & sel_one_hot_i[32];
  assign data_masked[2087] = data_i[2087] & sel_one_hot_i[32];
  assign data_masked[2086] = data_i[2086] & sel_one_hot_i[32];
  assign data_masked[2085] = data_i[2085] & sel_one_hot_i[32];
  assign data_masked[2084] = data_i[2084] & sel_one_hot_i[32];
  assign data_masked[2083] = data_i[2083] & sel_one_hot_i[32];
  assign data_masked[2082] = data_i[2082] & sel_one_hot_i[32];
  assign data_masked[2081] = data_i[2081] & sel_one_hot_i[32];
  assign data_masked[2080] = data_i[2080] & sel_one_hot_i[32];
  assign data_masked[2079] = data_i[2079] & sel_one_hot_i[32];
  assign data_masked[2078] = data_i[2078] & sel_one_hot_i[32];
  assign data_masked[2077] = data_i[2077] & sel_one_hot_i[32];
  assign data_masked[2076] = data_i[2076] & sel_one_hot_i[32];
  assign data_masked[2075] = data_i[2075] & sel_one_hot_i[32];
  assign data_masked[2074] = data_i[2074] & sel_one_hot_i[32];
  assign data_masked[2073] = data_i[2073] & sel_one_hot_i[32];
  assign data_masked[2072] = data_i[2072] & sel_one_hot_i[32];
  assign data_masked[2071] = data_i[2071] & sel_one_hot_i[32];
  assign data_masked[2070] = data_i[2070] & sel_one_hot_i[32];
  assign data_masked[2069] = data_i[2069] & sel_one_hot_i[32];
  assign data_masked[2068] = data_i[2068] & sel_one_hot_i[32];
  assign data_masked[2067] = data_i[2067] & sel_one_hot_i[32];
  assign data_masked[2066] = data_i[2066] & sel_one_hot_i[32];
  assign data_masked[2065] = data_i[2065] & sel_one_hot_i[32];
  assign data_masked[2064] = data_i[2064] & sel_one_hot_i[32];
  assign data_masked[2063] = data_i[2063] & sel_one_hot_i[32];
  assign data_masked[2062] = data_i[2062] & sel_one_hot_i[32];
  assign data_masked[2061] = data_i[2061] & sel_one_hot_i[32];
  assign data_masked[2060] = data_i[2060] & sel_one_hot_i[32];
  assign data_masked[2059] = data_i[2059] & sel_one_hot_i[32];
  assign data_masked[2058] = data_i[2058] & sel_one_hot_i[32];
  assign data_masked[2057] = data_i[2057] & sel_one_hot_i[32];
  assign data_masked[2056] = data_i[2056] & sel_one_hot_i[32];
  assign data_masked[2055] = data_i[2055] & sel_one_hot_i[32];
  assign data_masked[2054] = data_i[2054] & sel_one_hot_i[32];
  assign data_masked[2053] = data_i[2053] & sel_one_hot_i[32];
  assign data_masked[2052] = data_i[2052] & sel_one_hot_i[32];
  assign data_masked[2051] = data_i[2051] & sel_one_hot_i[32];
  assign data_masked[2050] = data_i[2050] & sel_one_hot_i[32];
  assign data_masked[2049] = data_i[2049] & sel_one_hot_i[32];
  assign data_masked[2048] = data_i[2048] & sel_one_hot_i[32];
  assign data_masked[2175] = data_i[2175] & sel_one_hot_i[33];
  assign data_masked[2174] = data_i[2174] & sel_one_hot_i[33];
  assign data_masked[2173] = data_i[2173] & sel_one_hot_i[33];
  assign data_masked[2172] = data_i[2172] & sel_one_hot_i[33];
  assign data_masked[2171] = data_i[2171] & sel_one_hot_i[33];
  assign data_masked[2170] = data_i[2170] & sel_one_hot_i[33];
  assign data_masked[2169] = data_i[2169] & sel_one_hot_i[33];
  assign data_masked[2168] = data_i[2168] & sel_one_hot_i[33];
  assign data_masked[2167] = data_i[2167] & sel_one_hot_i[33];
  assign data_masked[2166] = data_i[2166] & sel_one_hot_i[33];
  assign data_masked[2165] = data_i[2165] & sel_one_hot_i[33];
  assign data_masked[2164] = data_i[2164] & sel_one_hot_i[33];
  assign data_masked[2163] = data_i[2163] & sel_one_hot_i[33];
  assign data_masked[2162] = data_i[2162] & sel_one_hot_i[33];
  assign data_masked[2161] = data_i[2161] & sel_one_hot_i[33];
  assign data_masked[2160] = data_i[2160] & sel_one_hot_i[33];
  assign data_masked[2159] = data_i[2159] & sel_one_hot_i[33];
  assign data_masked[2158] = data_i[2158] & sel_one_hot_i[33];
  assign data_masked[2157] = data_i[2157] & sel_one_hot_i[33];
  assign data_masked[2156] = data_i[2156] & sel_one_hot_i[33];
  assign data_masked[2155] = data_i[2155] & sel_one_hot_i[33];
  assign data_masked[2154] = data_i[2154] & sel_one_hot_i[33];
  assign data_masked[2153] = data_i[2153] & sel_one_hot_i[33];
  assign data_masked[2152] = data_i[2152] & sel_one_hot_i[33];
  assign data_masked[2151] = data_i[2151] & sel_one_hot_i[33];
  assign data_masked[2150] = data_i[2150] & sel_one_hot_i[33];
  assign data_masked[2149] = data_i[2149] & sel_one_hot_i[33];
  assign data_masked[2148] = data_i[2148] & sel_one_hot_i[33];
  assign data_masked[2147] = data_i[2147] & sel_one_hot_i[33];
  assign data_masked[2146] = data_i[2146] & sel_one_hot_i[33];
  assign data_masked[2145] = data_i[2145] & sel_one_hot_i[33];
  assign data_masked[2144] = data_i[2144] & sel_one_hot_i[33];
  assign data_masked[2143] = data_i[2143] & sel_one_hot_i[33];
  assign data_masked[2142] = data_i[2142] & sel_one_hot_i[33];
  assign data_masked[2141] = data_i[2141] & sel_one_hot_i[33];
  assign data_masked[2140] = data_i[2140] & sel_one_hot_i[33];
  assign data_masked[2139] = data_i[2139] & sel_one_hot_i[33];
  assign data_masked[2138] = data_i[2138] & sel_one_hot_i[33];
  assign data_masked[2137] = data_i[2137] & sel_one_hot_i[33];
  assign data_masked[2136] = data_i[2136] & sel_one_hot_i[33];
  assign data_masked[2135] = data_i[2135] & sel_one_hot_i[33];
  assign data_masked[2134] = data_i[2134] & sel_one_hot_i[33];
  assign data_masked[2133] = data_i[2133] & sel_one_hot_i[33];
  assign data_masked[2132] = data_i[2132] & sel_one_hot_i[33];
  assign data_masked[2131] = data_i[2131] & sel_one_hot_i[33];
  assign data_masked[2130] = data_i[2130] & sel_one_hot_i[33];
  assign data_masked[2129] = data_i[2129] & sel_one_hot_i[33];
  assign data_masked[2128] = data_i[2128] & sel_one_hot_i[33];
  assign data_masked[2127] = data_i[2127] & sel_one_hot_i[33];
  assign data_masked[2126] = data_i[2126] & sel_one_hot_i[33];
  assign data_masked[2125] = data_i[2125] & sel_one_hot_i[33];
  assign data_masked[2124] = data_i[2124] & sel_one_hot_i[33];
  assign data_masked[2123] = data_i[2123] & sel_one_hot_i[33];
  assign data_masked[2122] = data_i[2122] & sel_one_hot_i[33];
  assign data_masked[2121] = data_i[2121] & sel_one_hot_i[33];
  assign data_masked[2120] = data_i[2120] & sel_one_hot_i[33];
  assign data_masked[2119] = data_i[2119] & sel_one_hot_i[33];
  assign data_masked[2118] = data_i[2118] & sel_one_hot_i[33];
  assign data_masked[2117] = data_i[2117] & sel_one_hot_i[33];
  assign data_masked[2116] = data_i[2116] & sel_one_hot_i[33];
  assign data_masked[2115] = data_i[2115] & sel_one_hot_i[33];
  assign data_masked[2114] = data_i[2114] & sel_one_hot_i[33];
  assign data_masked[2113] = data_i[2113] & sel_one_hot_i[33];
  assign data_masked[2112] = data_i[2112] & sel_one_hot_i[33];
  assign data_masked[2239] = data_i[2239] & sel_one_hot_i[34];
  assign data_masked[2238] = data_i[2238] & sel_one_hot_i[34];
  assign data_masked[2237] = data_i[2237] & sel_one_hot_i[34];
  assign data_masked[2236] = data_i[2236] & sel_one_hot_i[34];
  assign data_masked[2235] = data_i[2235] & sel_one_hot_i[34];
  assign data_masked[2234] = data_i[2234] & sel_one_hot_i[34];
  assign data_masked[2233] = data_i[2233] & sel_one_hot_i[34];
  assign data_masked[2232] = data_i[2232] & sel_one_hot_i[34];
  assign data_masked[2231] = data_i[2231] & sel_one_hot_i[34];
  assign data_masked[2230] = data_i[2230] & sel_one_hot_i[34];
  assign data_masked[2229] = data_i[2229] & sel_one_hot_i[34];
  assign data_masked[2228] = data_i[2228] & sel_one_hot_i[34];
  assign data_masked[2227] = data_i[2227] & sel_one_hot_i[34];
  assign data_masked[2226] = data_i[2226] & sel_one_hot_i[34];
  assign data_masked[2225] = data_i[2225] & sel_one_hot_i[34];
  assign data_masked[2224] = data_i[2224] & sel_one_hot_i[34];
  assign data_masked[2223] = data_i[2223] & sel_one_hot_i[34];
  assign data_masked[2222] = data_i[2222] & sel_one_hot_i[34];
  assign data_masked[2221] = data_i[2221] & sel_one_hot_i[34];
  assign data_masked[2220] = data_i[2220] & sel_one_hot_i[34];
  assign data_masked[2219] = data_i[2219] & sel_one_hot_i[34];
  assign data_masked[2218] = data_i[2218] & sel_one_hot_i[34];
  assign data_masked[2217] = data_i[2217] & sel_one_hot_i[34];
  assign data_masked[2216] = data_i[2216] & sel_one_hot_i[34];
  assign data_masked[2215] = data_i[2215] & sel_one_hot_i[34];
  assign data_masked[2214] = data_i[2214] & sel_one_hot_i[34];
  assign data_masked[2213] = data_i[2213] & sel_one_hot_i[34];
  assign data_masked[2212] = data_i[2212] & sel_one_hot_i[34];
  assign data_masked[2211] = data_i[2211] & sel_one_hot_i[34];
  assign data_masked[2210] = data_i[2210] & sel_one_hot_i[34];
  assign data_masked[2209] = data_i[2209] & sel_one_hot_i[34];
  assign data_masked[2208] = data_i[2208] & sel_one_hot_i[34];
  assign data_masked[2207] = data_i[2207] & sel_one_hot_i[34];
  assign data_masked[2206] = data_i[2206] & sel_one_hot_i[34];
  assign data_masked[2205] = data_i[2205] & sel_one_hot_i[34];
  assign data_masked[2204] = data_i[2204] & sel_one_hot_i[34];
  assign data_masked[2203] = data_i[2203] & sel_one_hot_i[34];
  assign data_masked[2202] = data_i[2202] & sel_one_hot_i[34];
  assign data_masked[2201] = data_i[2201] & sel_one_hot_i[34];
  assign data_masked[2200] = data_i[2200] & sel_one_hot_i[34];
  assign data_masked[2199] = data_i[2199] & sel_one_hot_i[34];
  assign data_masked[2198] = data_i[2198] & sel_one_hot_i[34];
  assign data_masked[2197] = data_i[2197] & sel_one_hot_i[34];
  assign data_masked[2196] = data_i[2196] & sel_one_hot_i[34];
  assign data_masked[2195] = data_i[2195] & sel_one_hot_i[34];
  assign data_masked[2194] = data_i[2194] & sel_one_hot_i[34];
  assign data_masked[2193] = data_i[2193] & sel_one_hot_i[34];
  assign data_masked[2192] = data_i[2192] & sel_one_hot_i[34];
  assign data_masked[2191] = data_i[2191] & sel_one_hot_i[34];
  assign data_masked[2190] = data_i[2190] & sel_one_hot_i[34];
  assign data_masked[2189] = data_i[2189] & sel_one_hot_i[34];
  assign data_masked[2188] = data_i[2188] & sel_one_hot_i[34];
  assign data_masked[2187] = data_i[2187] & sel_one_hot_i[34];
  assign data_masked[2186] = data_i[2186] & sel_one_hot_i[34];
  assign data_masked[2185] = data_i[2185] & sel_one_hot_i[34];
  assign data_masked[2184] = data_i[2184] & sel_one_hot_i[34];
  assign data_masked[2183] = data_i[2183] & sel_one_hot_i[34];
  assign data_masked[2182] = data_i[2182] & sel_one_hot_i[34];
  assign data_masked[2181] = data_i[2181] & sel_one_hot_i[34];
  assign data_masked[2180] = data_i[2180] & sel_one_hot_i[34];
  assign data_masked[2179] = data_i[2179] & sel_one_hot_i[34];
  assign data_masked[2178] = data_i[2178] & sel_one_hot_i[34];
  assign data_masked[2177] = data_i[2177] & sel_one_hot_i[34];
  assign data_masked[2176] = data_i[2176] & sel_one_hot_i[34];
  assign data_masked[2303] = data_i[2303] & sel_one_hot_i[35];
  assign data_masked[2302] = data_i[2302] & sel_one_hot_i[35];
  assign data_masked[2301] = data_i[2301] & sel_one_hot_i[35];
  assign data_masked[2300] = data_i[2300] & sel_one_hot_i[35];
  assign data_masked[2299] = data_i[2299] & sel_one_hot_i[35];
  assign data_masked[2298] = data_i[2298] & sel_one_hot_i[35];
  assign data_masked[2297] = data_i[2297] & sel_one_hot_i[35];
  assign data_masked[2296] = data_i[2296] & sel_one_hot_i[35];
  assign data_masked[2295] = data_i[2295] & sel_one_hot_i[35];
  assign data_masked[2294] = data_i[2294] & sel_one_hot_i[35];
  assign data_masked[2293] = data_i[2293] & sel_one_hot_i[35];
  assign data_masked[2292] = data_i[2292] & sel_one_hot_i[35];
  assign data_masked[2291] = data_i[2291] & sel_one_hot_i[35];
  assign data_masked[2290] = data_i[2290] & sel_one_hot_i[35];
  assign data_masked[2289] = data_i[2289] & sel_one_hot_i[35];
  assign data_masked[2288] = data_i[2288] & sel_one_hot_i[35];
  assign data_masked[2287] = data_i[2287] & sel_one_hot_i[35];
  assign data_masked[2286] = data_i[2286] & sel_one_hot_i[35];
  assign data_masked[2285] = data_i[2285] & sel_one_hot_i[35];
  assign data_masked[2284] = data_i[2284] & sel_one_hot_i[35];
  assign data_masked[2283] = data_i[2283] & sel_one_hot_i[35];
  assign data_masked[2282] = data_i[2282] & sel_one_hot_i[35];
  assign data_masked[2281] = data_i[2281] & sel_one_hot_i[35];
  assign data_masked[2280] = data_i[2280] & sel_one_hot_i[35];
  assign data_masked[2279] = data_i[2279] & sel_one_hot_i[35];
  assign data_masked[2278] = data_i[2278] & sel_one_hot_i[35];
  assign data_masked[2277] = data_i[2277] & sel_one_hot_i[35];
  assign data_masked[2276] = data_i[2276] & sel_one_hot_i[35];
  assign data_masked[2275] = data_i[2275] & sel_one_hot_i[35];
  assign data_masked[2274] = data_i[2274] & sel_one_hot_i[35];
  assign data_masked[2273] = data_i[2273] & sel_one_hot_i[35];
  assign data_masked[2272] = data_i[2272] & sel_one_hot_i[35];
  assign data_masked[2271] = data_i[2271] & sel_one_hot_i[35];
  assign data_masked[2270] = data_i[2270] & sel_one_hot_i[35];
  assign data_masked[2269] = data_i[2269] & sel_one_hot_i[35];
  assign data_masked[2268] = data_i[2268] & sel_one_hot_i[35];
  assign data_masked[2267] = data_i[2267] & sel_one_hot_i[35];
  assign data_masked[2266] = data_i[2266] & sel_one_hot_i[35];
  assign data_masked[2265] = data_i[2265] & sel_one_hot_i[35];
  assign data_masked[2264] = data_i[2264] & sel_one_hot_i[35];
  assign data_masked[2263] = data_i[2263] & sel_one_hot_i[35];
  assign data_masked[2262] = data_i[2262] & sel_one_hot_i[35];
  assign data_masked[2261] = data_i[2261] & sel_one_hot_i[35];
  assign data_masked[2260] = data_i[2260] & sel_one_hot_i[35];
  assign data_masked[2259] = data_i[2259] & sel_one_hot_i[35];
  assign data_masked[2258] = data_i[2258] & sel_one_hot_i[35];
  assign data_masked[2257] = data_i[2257] & sel_one_hot_i[35];
  assign data_masked[2256] = data_i[2256] & sel_one_hot_i[35];
  assign data_masked[2255] = data_i[2255] & sel_one_hot_i[35];
  assign data_masked[2254] = data_i[2254] & sel_one_hot_i[35];
  assign data_masked[2253] = data_i[2253] & sel_one_hot_i[35];
  assign data_masked[2252] = data_i[2252] & sel_one_hot_i[35];
  assign data_masked[2251] = data_i[2251] & sel_one_hot_i[35];
  assign data_masked[2250] = data_i[2250] & sel_one_hot_i[35];
  assign data_masked[2249] = data_i[2249] & sel_one_hot_i[35];
  assign data_masked[2248] = data_i[2248] & sel_one_hot_i[35];
  assign data_masked[2247] = data_i[2247] & sel_one_hot_i[35];
  assign data_masked[2246] = data_i[2246] & sel_one_hot_i[35];
  assign data_masked[2245] = data_i[2245] & sel_one_hot_i[35];
  assign data_masked[2244] = data_i[2244] & sel_one_hot_i[35];
  assign data_masked[2243] = data_i[2243] & sel_one_hot_i[35];
  assign data_masked[2242] = data_i[2242] & sel_one_hot_i[35];
  assign data_masked[2241] = data_i[2241] & sel_one_hot_i[35];
  assign data_masked[2240] = data_i[2240] & sel_one_hot_i[35];
  assign data_masked[2367] = data_i[2367] & sel_one_hot_i[36];
  assign data_masked[2366] = data_i[2366] & sel_one_hot_i[36];
  assign data_masked[2365] = data_i[2365] & sel_one_hot_i[36];
  assign data_masked[2364] = data_i[2364] & sel_one_hot_i[36];
  assign data_masked[2363] = data_i[2363] & sel_one_hot_i[36];
  assign data_masked[2362] = data_i[2362] & sel_one_hot_i[36];
  assign data_masked[2361] = data_i[2361] & sel_one_hot_i[36];
  assign data_masked[2360] = data_i[2360] & sel_one_hot_i[36];
  assign data_masked[2359] = data_i[2359] & sel_one_hot_i[36];
  assign data_masked[2358] = data_i[2358] & sel_one_hot_i[36];
  assign data_masked[2357] = data_i[2357] & sel_one_hot_i[36];
  assign data_masked[2356] = data_i[2356] & sel_one_hot_i[36];
  assign data_masked[2355] = data_i[2355] & sel_one_hot_i[36];
  assign data_masked[2354] = data_i[2354] & sel_one_hot_i[36];
  assign data_masked[2353] = data_i[2353] & sel_one_hot_i[36];
  assign data_masked[2352] = data_i[2352] & sel_one_hot_i[36];
  assign data_masked[2351] = data_i[2351] & sel_one_hot_i[36];
  assign data_masked[2350] = data_i[2350] & sel_one_hot_i[36];
  assign data_masked[2349] = data_i[2349] & sel_one_hot_i[36];
  assign data_masked[2348] = data_i[2348] & sel_one_hot_i[36];
  assign data_masked[2347] = data_i[2347] & sel_one_hot_i[36];
  assign data_masked[2346] = data_i[2346] & sel_one_hot_i[36];
  assign data_masked[2345] = data_i[2345] & sel_one_hot_i[36];
  assign data_masked[2344] = data_i[2344] & sel_one_hot_i[36];
  assign data_masked[2343] = data_i[2343] & sel_one_hot_i[36];
  assign data_masked[2342] = data_i[2342] & sel_one_hot_i[36];
  assign data_masked[2341] = data_i[2341] & sel_one_hot_i[36];
  assign data_masked[2340] = data_i[2340] & sel_one_hot_i[36];
  assign data_masked[2339] = data_i[2339] & sel_one_hot_i[36];
  assign data_masked[2338] = data_i[2338] & sel_one_hot_i[36];
  assign data_masked[2337] = data_i[2337] & sel_one_hot_i[36];
  assign data_masked[2336] = data_i[2336] & sel_one_hot_i[36];
  assign data_masked[2335] = data_i[2335] & sel_one_hot_i[36];
  assign data_masked[2334] = data_i[2334] & sel_one_hot_i[36];
  assign data_masked[2333] = data_i[2333] & sel_one_hot_i[36];
  assign data_masked[2332] = data_i[2332] & sel_one_hot_i[36];
  assign data_masked[2331] = data_i[2331] & sel_one_hot_i[36];
  assign data_masked[2330] = data_i[2330] & sel_one_hot_i[36];
  assign data_masked[2329] = data_i[2329] & sel_one_hot_i[36];
  assign data_masked[2328] = data_i[2328] & sel_one_hot_i[36];
  assign data_masked[2327] = data_i[2327] & sel_one_hot_i[36];
  assign data_masked[2326] = data_i[2326] & sel_one_hot_i[36];
  assign data_masked[2325] = data_i[2325] & sel_one_hot_i[36];
  assign data_masked[2324] = data_i[2324] & sel_one_hot_i[36];
  assign data_masked[2323] = data_i[2323] & sel_one_hot_i[36];
  assign data_masked[2322] = data_i[2322] & sel_one_hot_i[36];
  assign data_masked[2321] = data_i[2321] & sel_one_hot_i[36];
  assign data_masked[2320] = data_i[2320] & sel_one_hot_i[36];
  assign data_masked[2319] = data_i[2319] & sel_one_hot_i[36];
  assign data_masked[2318] = data_i[2318] & sel_one_hot_i[36];
  assign data_masked[2317] = data_i[2317] & sel_one_hot_i[36];
  assign data_masked[2316] = data_i[2316] & sel_one_hot_i[36];
  assign data_masked[2315] = data_i[2315] & sel_one_hot_i[36];
  assign data_masked[2314] = data_i[2314] & sel_one_hot_i[36];
  assign data_masked[2313] = data_i[2313] & sel_one_hot_i[36];
  assign data_masked[2312] = data_i[2312] & sel_one_hot_i[36];
  assign data_masked[2311] = data_i[2311] & sel_one_hot_i[36];
  assign data_masked[2310] = data_i[2310] & sel_one_hot_i[36];
  assign data_masked[2309] = data_i[2309] & sel_one_hot_i[36];
  assign data_masked[2308] = data_i[2308] & sel_one_hot_i[36];
  assign data_masked[2307] = data_i[2307] & sel_one_hot_i[36];
  assign data_masked[2306] = data_i[2306] & sel_one_hot_i[36];
  assign data_masked[2305] = data_i[2305] & sel_one_hot_i[36];
  assign data_masked[2304] = data_i[2304] & sel_one_hot_i[36];
  assign data_masked[2431] = data_i[2431] & sel_one_hot_i[37];
  assign data_masked[2430] = data_i[2430] & sel_one_hot_i[37];
  assign data_masked[2429] = data_i[2429] & sel_one_hot_i[37];
  assign data_masked[2428] = data_i[2428] & sel_one_hot_i[37];
  assign data_masked[2427] = data_i[2427] & sel_one_hot_i[37];
  assign data_masked[2426] = data_i[2426] & sel_one_hot_i[37];
  assign data_masked[2425] = data_i[2425] & sel_one_hot_i[37];
  assign data_masked[2424] = data_i[2424] & sel_one_hot_i[37];
  assign data_masked[2423] = data_i[2423] & sel_one_hot_i[37];
  assign data_masked[2422] = data_i[2422] & sel_one_hot_i[37];
  assign data_masked[2421] = data_i[2421] & sel_one_hot_i[37];
  assign data_masked[2420] = data_i[2420] & sel_one_hot_i[37];
  assign data_masked[2419] = data_i[2419] & sel_one_hot_i[37];
  assign data_masked[2418] = data_i[2418] & sel_one_hot_i[37];
  assign data_masked[2417] = data_i[2417] & sel_one_hot_i[37];
  assign data_masked[2416] = data_i[2416] & sel_one_hot_i[37];
  assign data_masked[2415] = data_i[2415] & sel_one_hot_i[37];
  assign data_masked[2414] = data_i[2414] & sel_one_hot_i[37];
  assign data_masked[2413] = data_i[2413] & sel_one_hot_i[37];
  assign data_masked[2412] = data_i[2412] & sel_one_hot_i[37];
  assign data_masked[2411] = data_i[2411] & sel_one_hot_i[37];
  assign data_masked[2410] = data_i[2410] & sel_one_hot_i[37];
  assign data_masked[2409] = data_i[2409] & sel_one_hot_i[37];
  assign data_masked[2408] = data_i[2408] & sel_one_hot_i[37];
  assign data_masked[2407] = data_i[2407] & sel_one_hot_i[37];
  assign data_masked[2406] = data_i[2406] & sel_one_hot_i[37];
  assign data_masked[2405] = data_i[2405] & sel_one_hot_i[37];
  assign data_masked[2404] = data_i[2404] & sel_one_hot_i[37];
  assign data_masked[2403] = data_i[2403] & sel_one_hot_i[37];
  assign data_masked[2402] = data_i[2402] & sel_one_hot_i[37];
  assign data_masked[2401] = data_i[2401] & sel_one_hot_i[37];
  assign data_masked[2400] = data_i[2400] & sel_one_hot_i[37];
  assign data_masked[2399] = data_i[2399] & sel_one_hot_i[37];
  assign data_masked[2398] = data_i[2398] & sel_one_hot_i[37];
  assign data_masked[2397] = data_i[2397] & sel_one_hot_i[37];
  assign data_masked[2396] = data_i[2396] & sel_one_hot_i[37];
  assign data_masked[2395] = data_i[2395] & sel_one_hot_i[37];
  assign data_masked[2394] = data_i[2394] & sel_one_hot_i[37];
  assign data_masked[2393] = data_i[2393] & sel_one_hot_i[37];
  assign data_masked[2392] = data_i[2392] & sel_one_hot_i[37];
  assign data_masked[2391] = data_i[2391] & sel_one_hot_i[37];
  assign data_masked[2390] = data_i[2390] & sel_one_hot_i[37];
  assign data_masked[2389] = data_i[2389] & sel_one_hot_i[37];
  assign data_masked[2388] = data_i[2388] & sel_one_hot_i[37];
  assign data_masked[2387] = data_i[2387] & sel_one_hot_i[37];
  assign data_masked[2386] = data_i[2386] & sel_one_hot_i[37];
  assign data_masked[2385] = data_i[2385] & sel_one_hot_i[37];
  assign data_masked[2384] = data_i[2384] & sel_one_hot_i[37];
  assign data_masked[2383] = data_i[2383] & sel_one_hot_i[37];
  assign data_masked[2382] = data_i[2382] & sel_one_hot_i[37];
  assign data_masked[2381] = data_i[2381] & sel_one_hot_i[37];
  assign data_masked[2380] = data_i[2380] & sel_one_hot_i[37];
  assign data_masked[2379] = data_i[2379] & sel_one_hot_i[37];
  assign data_masked[2378] = data_i[2378] & sel_one_hot_i[37];
  assign data_masked[2377] = data_i[2377] & sel_one_hot_i[37];
  assign data_masked[2376] = data_i[2376] & sel_one_hot_i[37];
  assign data_masked[2375] = data_i[2375] & sel_one_hot_i[37];
  assign data_masked[2374] = data_i[2374] & sel_one_hot_i[37];
  assign data_masked[2373] = data_i[2373] & sel_one_hot_i[37];
  assign data_masked[2372] = data_i[2372] & sel_one_hot_i[37];
  assign data_masked[2371] = data_i[2371] & sel_one_hot_i[37];
  assign data_masked[2370] = data_i[2370] & sel_one_hot_i[37];
  assign data_masked[2369] = data_i[2369] & sel_one_hot_i[37];
  assign data_masked[2368] = data_i[2368] & sel_one_hot_i[37];
  assign data_masked[2495] = data_i[2495] & sel_one_hot_i[38];
  assign data_masked[2494] = data_i[2494] & sel_one_hot_i[38];
  assign data_masked[2493] = data_i[2493] & sel_one_hot_i[38];
  assign data_masked[2492] = data_i[2492] & sel_one_hot_i[38];
  assign data_masked[2491] = data_i[2491] & sel_one_hot_i[38];
  assign data_masked[2490] = data_i[2490] & sel_one_hot_i[38];
  assign data_masked[2489] = data_i[2489] & sel_one_hot_i[38];
  assign data_masked[2488] = data_i[2488] & sel_one_hot_i[38];
  assign data_masked[2487] = data_i[2487] & sel_one_hot_i[38];
  assign data_masked[2486] = data_i[2486] & sel_one_hot_i[38];
  assign data_masked[2485] = data_i[2485] & sel_one_hot_i[38];
  assign data_masked[2484] = data_i[2484] & sel_one_hot_i[38];
  assign data_masked[2483] = data_i[2483] & sel_one_hot_i[38];
  assign data_masked[2482] = data_i[2482] & sel_one_hot_i[38];
  assign data_masked[2481] = data_i[2481] & sel_one_hot_i[38];
  assign data_masked[2480] = data_i[2480] & sel_one_hot_i[38];
  assign data_masked[2479] = data_i[2479] & sel_one_hot_i[38];
  assign data_masked[2478] = data_i[2478] & sel_one_hot_i[38];
  assign data_masked[2477] = data_i[2477] & sel_one_hot_i[38];
  assign data_masked[2476] = data_i[2476] & sel_one_hot_i[38];
  assign data_masked[2475] = data_i[2475] & sel_one_hot_i[38];
  assign data_masked[2474] = data_i[2474] & sel_one_hot_i[38];
  assign data_masked[2473] = data_i[2473] & sel_one_hot_i[38];
  assign data_masked[2472] = data_i[2472] & sel_one_hot_i[38];
  assign data_masked[2471] = data_i[2471] & sel_one_hot_i[38];
  assign data_masked[2470] = data_i[2470] & sel_one_hot_i[38];
  assign data_masked[2469] = data_i[2469] & sel_one_hot_i[38];
  assign data_masked[2468] = data_i[2468] & sel_one_hot_i[38];
  assign data_masked[2467] = data_i[2467] & sel_one_hot_i[38];
  assign data_masked[2466] = data_i[2466] & sel_one_hot_i[38];
  assign data_masked[2465] = data_i[2465] & sel_one_hot_i[38];
  assign data_masked[2464] = data_i[2464] & sel_one_hot_i[38];
  assign data_masked[2463] = data_i[2463] & sel_one_hot_i[38];
  assign data_masked[2462] = data_i[2462] & sel_one_hot_i[38];
  assign data_masked[2461] = data_i[2461] & sel_one_hot_i[38];
  assign data_masked[2460] = data_i[2460] & sel_one_hot_i[38];
  assign data_masked[2459] = data_i[2459] & sel_one_hot_i[38];
  assign data_masked[2458] = data_i[2458] & sel_one_hot_i[38];
  assign data_masked[2457] = data_i[2457] & sel_one_hot_i[38];
  assign data_masked[2456] = data_i[2456] & sel_one_hot_i[38];
  assign data_masked[2455] = data_i[2455] & sel_one_hot_i[38];
  assign data_masked[2454] = data_i[2454] & sel_one_hot_i[38];
  assign data_masked[2453] = data_i[2453] & sel_one_hot_i[38];
  assign data_masked[2452] = data_i[2452] & sel_one_hot_i[38];
  assign data_masked[2451] = data_i[2451] & sel_one_hot_i[38];
  assign data_masked[2450] = data_i[2450] & sel_one_hot_i[38];
  assign data_masked[2449] = data_i[2449] & sel_one_hot_i[38];
  assign data_masked[2448] = data_i[2448] & sel_one_hot_i[38];
  assign data_masked[2447] = data_i[2447] & sel_one_hot_i[38];
  assign data_masked[2446] = data_i[2446] & sel_one_hot_i[38];
  assign data_masked[2445] = data_i[2445] & sel_one_hot_i[38];
  assign data_masked[2444] = data_i[2444] & sel_one_hot_i[38];
  assign data_masked[2443] = data_i[2443] & sel_one_hot_i[38];
  assign data_masked[2442] = data_i[2442] & sel_one_hot_i[38];
  assign data_masked[2441] = data_i[2441] & sel_one_hot_i[38];
  assign data_masked[2440] = data_i[2440] & sel_one_hot_i[38];
  assign data_masked[2439] = data_i[2439] & sel_one_hot_i[38];
  assign data_masked[2438] = data_i[2438] & sel_one_hot_i[38];
  assign data_masked[2437] = data_i[2437] & sel_one_hot_i[38];
  assign data_masked[2436] = data_i[2436] & sel_one_hot_i[38];
  assign data_masked[2435] = data_i[2435] & sel_one_hot_i[38];
  assign data_masked[2434] = data_i[2434] & sel_one_hot_i[38];
  assign data_masked[2433] = data_i[2433] & sel_one_hot_i[38];
  assign data_masked[2432] = data_i[2432] & sel_one_hot_i[38];
  assign data_masked[2559] = data_i[2559] & sel_one_hot_i[39];
  assign data_masked[2558] = data_i[2558] & sel_one_hot_i[39];
  assign data_masked[2557] = data_i[2557] & sel_one_hot_i[39];
  assign data_masked[2556] = data_i[2556] & sel_one_hot_i[39];
  assign data_masked[2555] = data_i[2555] & sel_one_hot_i[39];
  assign data_masked[2554] = data_i[2554] & sel_one_hot_i[39];
  assign data_masked[2553] = data_i[2553] & sel_one_hot_i[39];
  assign data_masked[2552] = data_i[2552] & sel_one_hot_i[39];
  assign data_masked[2551] = data_i[2551] & sel_one_hot_i[39];
  assign data_masked[2550] = data_i[2550] & sel_one_hot_i[39];
  assign data_masked[2549] = data_i[2549] & sel_one_hot_i[39];
  assign data_masked[2548] = data_i[2548] & sel_one_hot_i[39];
  assign data_masked[2547] = data_i[2547] & sel_one_hot_i[39];
  assign data_masked[2546] = data_i[2546] & sel_one_hot_i[39];
  assign data_masked[2545] = data_i[2545] & sel_one_hot_i[39];
  assign data_masked[2544] = data_i[2544] & sel_one_hot_i[39];
  assign data_masked[2543] = data_i[2543] & sel_one_hot_i[39];
  assign data_masked[2542] = data_i[2542] & sel_one_hot_i[39];
  assign data_masked[2541] = data_i[2541] & sel_one_hot_i[39];
  assign data_masked[2540] = data_i[2540] & sel_one_hot_i[39];
  assign data_masked[2539] = data_i[2539] & sel_one_hot_i[39];
  assign data_masked[2538] = data_i[2538] & sel_one_hot_i[39];
  assign data_masked[2537] = data_i[2537] & sel_one_hot_i[39];
  assign data_masked[2536] = data_i[2536] & sel_one_hot_i[39];
  assign data_masked[2535] = data_i[2535] & sel_one_hot_i[39];
  assign data_masked[2534] = data_i[2534] & sel_one_hot_i[39];
  assign data_masked[2533] = data_i[2533] & sel_one_hot_i[39];
  assign data_masked[2532] = data_i[2532] & sel_one_hot_i[39];
  assign data_masked[2531] = data_i[2531] & sel_one_hot_i[39];
  assign data_masked[2530] = data_i[2530] & sel_one_hot_i[39];
  assign data_masked[2529] = data_i[2529] & sel_one_hot_i[39];
  assign data_masked[2528] = data_i[2528] & sel_one_hot_i[39];
  assign data_masked[2527] = data_i[2527] & sel_one_hot_i[39];
  assign data_masked[2526] = data_i[2526] & sel_one_hot_i[39];
  assign data_masked[2525] = data_i[2525] & sel_one_hot_i[39];
  assign data_masked[2524] = data_i[2524] & sel_one_hot_i[39];
  assign data_masked[2523] = data_i[2523] & sel_one_hot_i[39];
  assign data_masked[2522] = data_i[2522] & sel_one_hot_i[39];
  assign data_masked[2521] = data_i[2521] & sel_one_hot_i[39];
  assign data_masked[2520] = data_i[2520] & sel_one_hot_i[39];
  assign data_masked[2519] = data_i[2519] & sel_one_hot_i[39];
  assign data_masked[2518] = data_i[2518] & sel_one_hot_i[39];
  assign data_masked[2517] = data_i[2517] & sel_one_hot_i[39];
  assign data_masked[2516] = data_i[2516] & sel_one_hot_i[39];
  assign data_masked[2515] = data_i[2515] & sel_one_hot_i[39];
  assign data_masked[2514] = data_i[2514] & sel_one_hot_i[39];
  assign data_masked[2513] = data_i[2513] & sel_one_hot_i[39];
  assign data_masked[2512] = data_i[2512] & sel_one_hot_i[39];
  assign data_masked[2511] = data_i[2511] & sel_one_hot_i[39];
  assign data_masked[2510] = data_i[2510] & sel_one_hot_i[39];
  assign data_masked[2509] = data_i[2509] & sel_one_hot_i[39];
  assign data_masked[2508] = data_i[2508] & sel_one_hot_i[39];
  assign data_masked[2507] = data_i[2507] & sel_one_hot_i[39];
  assign data_masked[2506] = data_i[2506] & sel_one_hot_i[39];
  assign data_masked[2505] = data_i[2505] & sel_one_hot_i[39];
  assign data_masked[2504] = data_i[2504] & sel_one_hot_i[39];
  assign data_masked[2503] = data_i[2503] & sel_one_hot_i[39];
  assign data_masked[2502] = data_i[2502] & sel_one_hot_i[39];
  assign data_masked[2501] = data_i[2501] & sel_one_hot_i[39];
  assign data_masked[2500] = data_i[2500] & sel_one_hot_i[39];
  assign data_masked[2499] = data_i[2499] & sel_one_hot_i[39];
  assign data_masked[2498] = data_i[2498] & sel_one_hot_i[39];
  assign data_masked[2497] = data_i[2497] & sel_one_hot_i[39];
  assign data_masked[2496] = data_i[2496] & sel_one_hot_i[39];
  assign data_masked[2623] = data_i[2623] & sel_one_hot_i[40];
  assign data_masked[2622] = data_i[2622] & sel_one_hot_i[40];
  assign data_masked[2621] = data_i[2621] & sel_one_hot_i[40];
  assign data_masked[2620] = data_i[2620] & sel_one_hot_i[40];
  assign data_masked[2619] = data_i[2619] & sel_one_hot_i[40];
  assign data_masked[2618] = data_i[2618] & sel_one_hot_i[40];
  assign data_masked[2617] = data_i[2617] & sel_one_hot_i[40];
  assign data_masked[2616] = data_i[2616] & sel_one_hot_i[40];
  assign data_masked[2615] = data_i[2615] & sel_one_hot_i[40];
  assign data_masked[2614] = data_i[2614] & sel_one_hot_i[40];
  assign data_masked[2613] = data_i[2613] & sel_one_hot_i[40];
  assign data_masked[2612] = data_i[2612] & sel_one_hot_i[40];
  assign data_masked[2611] = data_i[2611] & sel_one_hot_i[40];
  assign data_masked[2610] = data_i[2610] & sel_one_hot_i[40];
  assign data_masked[2609] = data_i[2609] & sel_one_hot_i[40];
  assign data_masked[2608] = data_i[2608] & sel_one_hot_i[40];
  assign data_masked[2607] = data_i[2607] & sel_one_hot_i[40];
  assign data_masked[2606] = data_i[2606] & sel_one_hot_i[40];
  assign data_masked[2605] = data_i[2605] & sel_one_hot_i[40];
  assign data_masked[2604] = data_i[2604] & sel_one_hot_i[40];
  assign data_masked[2603] = data_i[2603] & sel_one_hot_i[40];
  assign data_masked[2602] = data_i[2602] & sel_one_hot_i[40];
  assign data_masked[2601] = data_i[2601] & sel_one_hot_i[40];
  assign data_masked[2600] = data_i[2600] & sel_one_hot_i[40];
  assign data_masked[2599] = data_i[2599] & sel_one_hot_i[40];
  assign data_masked[2598] = data_i[2598] & sel_one_hot_i[40];
  assign data_masked[2597] = data_i[2597] & sel_one_hot_i[40];
  assign data_masked[2596] = data_i[2596] & sel_one_hot_i[40];
  assign data_masked[2595] = data_i[2595] & sel_one_hot_i[40];
  assign data_masked[2594] = data_i[2594] & sel_one_hot_i[40];
  assign data_masked[2593] = data_i[2593] & sel_one_hot_i[40];
  assign data_masked[2592] = data_i[2592] & sel_one_hot_i[40];
  assign data_masked[2591] = data_i[2591] & sel_one_hot_i[40];
  assign data_masked[2590] = data_i[2590] & sel_one_hot_i[40];
  assign data_masked[2589] = data_i[2589] & sel_one_hot_i[40];
  assign data_masked[2588] = data_i[2588] & sel_one_hot_i[40];
  assign data_masked[2587] = data_i[2587] & sel_one_hot_i[40];
  assign data_masked[2586] = data_i[2586] & sel_one_hot_i[40];
  assign data_masked[2585] = data_i[2585] & sel_one_hot_i[40];
  assign data_masked[2584] = data_i[2584] & sel_one_hot_i[40];
  assign data_masked[2583] = data_i[2583] & sel_one_hot_i[40];
  assign data_masked[2582] = data_i[2582] & sel_one_hot_i[40];
  assign data_masked[2581] = data_i[2581] & sel_one_hot_i[40];
  assign data_masked[2580] = data_i[2580] & sel_one_hot_i[40];
  assign data_masked[2579] = data_i[2579] & sel_one_hot_i[40];
  assign data_masked[2578] = data_i[2578] & sel_one_hot_i[40];
  assign data_masked[2577] = data_i[2577] & sel_one_hot_i[40];
  assign data_masked[2576] = data_i[2576] & sel_one_hot_i[40];
  assign data_masked[2575] = data_i[2575] & sel_one_hot_i[40];
  assign data_masked[2574] = data_i[2574] & sel_one_hot_i[40];
  assign data_masked[2573] = data_i[2573] & sel_one_hot_i[40];
  assign data_masked[2572] = data_i[2572] & sel_one_hot_i[40];
  assign data_masked[2571] = data_i[2571] & sel_one_hot_i[40];
  assign data_masked[2570] = data_i[2570] & sel_one_hot_i[40];
  assign data_masked[2569] = data_i[2569] & sel_one_hot_i[40];
  assign data_masked[2568] = data_i[2568] & sel_one_hot_i[40];
  assign data_masked[2567] = data_i[2567] & sel_one_hot_i[40];
  assign data_masked[2566] = data_i[2566] & sel_one_hot_i[40];
  assign data_masked[2565] = data_i[2565] & sel_one_hot_i[40];
  assign data_masked[2564] = data_i[2564] & sel_one_hot_i[40];
  assign data_masked[2563] = data_i[2563] & sel_one_hot_i[40];
  assign data_masked[2562] = data_i[2562] & sel_one_hot_i[40];
  assign data_masked[2561] = data_i[2561] & sel_one_hot_i[40];
  assign data_masked[2560] = data_i[2560] & sel_one_hot_i[40];
  assign data_masked[2687] = data_i[2687] & sel_one_hot_i[41];
  assign data_masked[2686] = data_i[2686] & sel_one_hot_i[41];
  assign data_masked[2685] = data_i[2685] & sel_one_hot_i[41];
  assign data_masked[2684] = data_i[2684] & sel_one_hot_i[41];
  assign data_masked[2683] = data_i[2683] & sel_one_hot_i[41];
  assign data_masked[2682] = data_i[2682] & sel_one_hot_i[41];
  assign data_masked[2681] = data_i[2681] & sel_one_hot_i[41];
  assign data_masked[2680] = data_i[2680] & sel_one_hot_i[41];
  assign data_masked[2679] = data_i[2679] & sel_one_hot_i[41];
  assign data_masked[2678] = data_i[2678] & sel_one_hot_i[41];
  assign data_masked[2677] = data_i[2677] & sel_one_hot_i[41];
  assign data_masked[2676] = data_i[2676] & sel_one_hot_i[41];
  assign data_masked[2675] = data_i[2675] & sel_one_hot_i[41];
  assign data_masked[2674] = data_i[2674] & sel_one_hot_i[41];
  assign data_masked[2673] = data_i[2673] & sel_one_hot_i[41];
  assign data_masked[2672] = data_i[2672] & sel_one_hot_i[41];
  assign data_masked[2671] = data_i[2671] & sel_one_hot_i[41];
  assign data_masked[2670] = data_i[2670] & sel_one_hot_i[41];
  assign data_masked[2669] = data_i[2669] & sel_one_hot_i[41];
  assign data_masked[2668] = data_i[2668] & sel_one_hot_i[41];
  assign data_masked[2667] = data_i[2667] & sel_one_hot_i[41];
  assign data_masked[2666] = data_i[2666] & sel_one_hot_i[41];
  assign data_masked[2665] = data_i[2665] & sel_one_hot_i[41];
  assign data_masked[2664] = data_i[2664] & sel_one_hot_i[41];
  assign data_masked[2663] = data_i[2663] & sel_one_hot_i[41];
  assign data_masked[2662] = data_i[2662] & sel_one_hot_i[41];
  assign data_masked[2661] = data_i[2661] & sel_one_hot_i[41];
  assign data_masked[2660] = data_i[2660] & sel_one_hot_i[41];
  assign data_masked[2659] = data_i[2659] & sel_one_hot_i[41];
  assign data_masked[2658] = data_i[2658] & sel_one_hot_i[41];
  assign data_masked[2657] = data_i[2657] & sel_one_hot_i[41];
  assign data_masked[2656] = data_i[2656] & sel_one_hot_i[41];
  assign data_masked[2655] = data_i[2655] & sel_one_hot_i[41];
  assign data_masked[2654] = data_i[2654] & sel_one_hot_i[41];
  assign data_masked[2653] = data_i[2653] & sel_one_hot_i[41];
  assign data_masked[2652] = data_i[2652] & sel_one_hot_i[41];
  assign data_masked[2651] = data_i[2651] & sel_one_hot_i[41];
  assign data_masked[2650] = data_i[2650] & sel_one_hot_i[41];
  assign data_masked[2649] = data_i[2649] & sel_one_hot_i[41];
  assign data_masked[2648] = data_i[2648] & sel_one_hot_i[41];
  assign data_masked[2647] = data_i[2647] & sel_one_hot_i[41];
  assign data_masked[2646] = data_i[2646] & sel_one_hot_i[41];
  assign data_masked[2645] = data_i[2645] & sel_one_hot_i[41];
  assign data_masked[2644] = data_i[2644] & sel_one_hot_i[41];
  assign data_masked[2643] = data_i[2643] & sel_one_hot_i[41];
  assign data_masked[2642] = data_i[2642] & sel_one_hot_i[41];
  assign data_masked[2641] = data_i[2641] & sel_one_hot_i[41];
  assign data_masked[2640] = data_i[2640] & sel_one_hot_i[41];
  assign data_masked[2639] = data_i[2639] & sel_one_hot_i[41];
  assign data_masked[2638] = data_i[2638] & sel_one_hot_i[41];
  assign data_masked[2637] = data_i[2637] & sel_one_hot_i[41];
  assign data_masked[2636] = data_i[2636] & sel_one_hot_i[41];
  assign data_masked[2635] = data_i[2635] & sel_one_hot_i[41];
  assign data_masked[2634] = data_i[2634] & sel_one_hot_i[41];
  assign data_masked[2633] = data_i[2633] & sel_one_hot_i[41];
  assign data_masked[2632] = data_i[2632] & sel_one_hot_i[41];
  assign data_masked[2631] = data_i[2631] & sel_one_hot_i[41];
  assign data_masked[2630] = data_i[2630] & sel_one_hot_i[41];
  assign data_masked[2629] = data_i[2629] & sel_one_hot_i[41];
  assign data_masked[2628] = data_i[2628] & sel_one_hot_i[41];
  assign data_masked[2627] = data_i[2627] & sel_one_hot_i[41];
  assign data_masked[2626] = data_i[2626] & sel_one_hot_i[41];
  assign data_masked[2625] = data_i[2625] & sel_one_hot_i[41];
  assign data_masked[2624] = data_i[2624] & sel_one_hot_i[41];
  assign data_masked[2751] = data_i[2751] & sel_one_hot_i[42];
  assign data_masked[2750] = data_i[2750] & sel_one_hot_i[42];
  assign data_masked[2749] = data_i[2749] & sel_one_hot_i[42];
  assign data_masked[2748] = data_i[2748] & sel_one_hot_i[42];
  assign data_masked[2747] = data_i[2747] & sel_one_hot_i[42];
  assign data_masked[2746] = data_i[2746] & sel_one_hot_i[42];
  assign data_masked[2745] = data_i[2745] & sel_one_hot_i[42];
  assign data_masked[2744] = data_i[2744] & sel_one_hot_i[42];
  assign data_masked[2743] = data_i[2743] & sel_one_hot_i[42];
  assign data_masked[2742] = data_i[2742] & sel_one_hot_i[42];
  assign data_masked[2741] = data_i[2741] & sel_one_hot_i[42];
  assign data_masked[2740] = data_i[2740] & sel_one_hot_i[42];
  assign data_masked[2739] = data_i[2739] & sel_one_hot_i[42];
  assign data_masked[2738] = data_i[2738] & sel_one_hot_i[42];
  assign data_masked[2737] = data_i[2737] & sel_one_hot_i[42];
  assign data_masked[2736] = data_i[2736] & sel_one_hot_i[42];
  assign data_masked[2735] = data_i[2735] & sel_one_hot_i[42];
  assign data_masked[2734] = data_i[2734] & sel_one_hot_i[42];
  assign data_masked[2733] = data_i[2733] & sel_one_hot_i[42];
  assign data_masked[2732] = data_i[2732] & sel_one_hot_i[42];
  assign data_masked[2731] = data_i[2731] & sel_one_hot_i[42];
  assign data_masked[2730] = data_i[2730] & sel_one_hot_i[42];
  assign data_masked[2729] = data_i[2729] & sel_one_hot_i[42];
  assign data_masked[2728] = data_i[2728] & sel_one_hot_i[42];
  assign data_masked[2727] = data_i[2727] & sel_one_hot_i[42];
  assign data_masked[2726] = data_i[2726] & sel_one_hot_i[42];
  assign data_masked[2725] = data_i[2725] & sel_one_hot_i[42];
  assign data_masked[2724] = data_i[2724] & sel_one_hot_i[42];
  assign data_masked[2723] = data_i[2723] & sel_one_hot_i[42];
  assign data_masked[2722] = data_i[2722] & sel_one_hot_i[42];
  assign data_masked[2721] = data_i[2721] & sel_one_hot_i[42];
  assign data_masked[2720] = data_i[2720] & sel_one_hot_i[42];
  assign data_masked[2719] = data_i[2719] & sel_one_hot_i[42];
  assign data_masked[2718] = data_i[2718] & sel_one_hot_i[42];
  assign data_masked[2717] = data_i[2717] & sel_one_hot_i[42];
  assign data_masked[2716] = data_i[2716] & sel_one_hot_i[42];
  assign data_masked[2715] = data_i[2715] & sel_one_hot_i[42];
  assign data_masked[2714] = data_i[2714] & sel_one_hot_i[42];
  assign data_masked[2713] = data_i[2713] & sel_one_hot_i[42];
  assign data_masked[2712] = data_i[2712] & sel_one_hot_i[42];
  assign data_masked[2711] = data_i[2711] & sel_one_hot_i[42];
  assign data_masked[2710] = data_i[2710] & sel_one_hot_i[42];
  assign data_masked[2709] = data_i[2709] & sel_one_hot_i[42];
  assign data_masked[2708] = data_i[2708] & sel_one_hot_i[42];
  assign data_masked[2707] = data_i[2707] & sel_one_hot_i[42];
  assign data_masked[2706] = data_i[2706] & sel_one_hot_i[42];
  assign data_masked[2705] = data_i[2705] & sel_one_hot_i[42];
  assign data_masked[2704] = data_i[2704] & sel_one_hot_i[42];
  assign data_masked[2703] = data_i[2703] & sel_one_hot_i[42];
  assign data_masked[2702] = data_i[2702] & sel_one_hot_i[42];
  assign data_masked[2701] = data_i[2701] & sel_one_hot_i[42];
  assign data_masked[2700] = data_i[2700] & sel_one_hot_i[42];
  assign data_masked[2699] = data_i[2699] & sel_one_hot_i[42];
  assign data_masked[2698] = data_i[2698] & sel_one_hot_i[42];
  assign data_masked[2697] = data_i[2697] & sel_one_hot_i[42];
  assign data_masked[2696] = data_i[2696] & sel_one_hot_i[42];
  assign data_masked[2695] = data_i[2695] & sel_one_hot_i[42];
  assign data_masked[2694] = data_i[2694] & sel_one_hot_i[42];
  assign data_masked[2693] = data_i[2693] & sel_one_hot_i[42];
  assign data_masked[2692] = data_i[2692] & sel_one_hot_i[42];
  assign data_masked[2691] = data_i[2691] & sel_one_hot_i[42];
  assign data_masked[2690] = data_i[2690] & sel_one_hot_i[42];
  assign data_masked[2689] = data_i[2689] & sel_one_hot_i[42];
  assign data_masked[2688] = data_i[2688] & sel_one_hot_i[42];
  assign data_masked[2815] = data_i[2815] & sel_one_hot_i[43];
  assign data_masked[2814] = data_i[2814] & sel_one_hot_i[43];
  assign data_masked[2813] = data_i[2813] & sel_one_hot_i[43];
  assign data_masked[2812] = data_i[2812] & sel_one_hot_i[43];
  assign data_masked[2811] = data_i[2811] & sel_one_hot_i[43];
  assign data_masked[2810] = data_i[2810] & sel_one_hot_i[43];
  assign data_masked[2809] = data_i[2809] & sel_one_hot_i[43];
  assign data_masked[2808] = data_i[2808] & sel_one_hot_i[43];
  assign data_masked[2807] = data_i[2807] & sel_one_hot_i[43];
  assign data_masked[2806] = data_i[2806] & sel_one_hot_i[43];
  assign data_masked[2805] = data_i[2805] & sel_one_hot_i[43];
  assign data_masked[2804] = data_i[2804] & sel_one_hot_i[43];
  assign data_masked[2803] = data_i[2803] & sel_one_hot_i[43];
  assign data_masked[2802] = data_i[2802] & sel_one_hot_i[43];
  assign data_masked[2801] = data_i[2801] & sel_one_hot_i[43];
  assign data_masked[2800] = data_i[2800] & sel_one_hot_i[43];
  assign data_masked[2799] = data_i[2799] & sel_one_hot_i[43];
  assign data_masked[2798] = data_i[2798] & sel_one_hot_i[43];
  assign data_masked[2797] = data_i[2797] & sel_one_hot_i[43];
  assign data_masked[2796] = data_i[2796] & sel_one_hot_i[43];
  assign data_masked[2795] = data_i[2795] & sel_one_hot_i[43];
  assign data_masked[2794] = data_i[2794] & sel_one_hot_i[43];
  assign data_masked[2793] = data_i[2793] & sel_one_hot_i[43];
  assign data_masked[2792] = data_i[2792] & sel_one_hot_i[43];
  assign data_masked[2791] = data_i[2791] & sel_one_hot_i[43];
  assign data_masked[2790] = data_i[2790] & sel_one_hot_i[43];
  assign data_masked[2789] = data_i[2789] & sel_one_hot_i[43];
  assign data_masked[2788] = data_i[2788] & sel_one_hot_i[43];
  assign data_masked[2787] = data_i[2787] & sel_one_hot_i[43];
  assign data_masked[2786] = data_i[2786] & sel_one_hot_i[43];
  assign data_masked[2785] = data_i[2785] & sel_one_hot_i[43];
  assign data_masked[2784] = data_i[2784] & sel_one_hot_i[43];
  assign data_masked[2783] = data_i[2783] & sel_one_hot_i[43];
  assign data_masked[2782] = data_i[2782] & sel_one_hot_i[43];
  assign data_masked[2781] = data_i[2781] & sel_one_hot_i[43];
  assign data_masked[2780] = data_i[2780] & sel_one_hot_i[43];
  assign data_masked[2779] = data_i[2779] & sel_one_hot_i[43];
  assign data_masked[2778] = data_i[2778] & sel_one_hot_i[43];
  assign data_masked[2777] = data_i[2777] & sel_one_hot_i[43];
  assign data_masked[2776] = data_i[2776] & sel_one_hot_i[43];
  assign data_masked[2775] = data_i[2775] & sel_one_hot_i[43];
  assign data_masked[2774] = data_i[2774] & sel_one_hot_i[43];
  assign data_masked[2773] = data_i[2773] & sel_one_hot_i[43];
  assign data_masked[2772] = data_i[2772] & sel_one_hot_i[43];
  assign data_masked[2771] = data_i[2771] & sel_one_hot_i[43];
  assign data_masked[2770] = data_i[2770] & sel_one_hot_i[43];
  assign data_masked[2769] = data_i[2769] & sel_one_hot_i[43];
  assign data_masked[2768] = data_i[2768] & sel_one_hot_i[43];
  assign data_masked[2767] = data_i[2767] & sel_one_hot_i[43];
  assign data_masked[2766] = data_i[2766] & sel_one_hot_i[43];
  assign data_masked[2765] = data_i[2765] & sel_one_hot_i[43];
  assign data_masked[2764] = data_i[2764] & sel_one_hot_i[43];
  assign data_masked[2763] = data_i[2763] & sel_one_hot_i[43];
  assign data_masked[2762] = data_i[2762] & sel_one_hot_i[43];
  assign data_masked[2761] = data_i[2761] & sel_one_hot_i[43];
  assign data_masked[2760] = data_i[2760] & sel_one_hot_i[43];
  assign data_masked[2759] = data_i[2759] & sel_one_hot_i[43];
  assign data_masked[2758] = data_i[2758] & sel_one_hot_i[43];
  assign data_masked[2757] = data_i[2757] & sel_one_hot_i[43];
  assign data_masked[2756] = data_i[2756] & sel_one_hot_i[43];
  assign data_masked[2755] = data_i[2755] & sel_one_hot_i[43];
  assign data_masked[2754] = data_i[2754] & sel_one_hot_i[43];
  assign data_masked[2753] = data_i[2753] & sel_one_hot_i[43];
  assign data_masked[2752] = data_i[2752] & sel_one_hot_i[43];
  assign data_masked[2879] = data_i[2879] & sel_one_hot_i[44];
  assign data_masked[2878] = data_i[2878] & sel_one_hot_i[44];
  assign data_masked[2877] = data_i[2877] & sel_one_hot_i[44];
  assign data_masked[2876] = data_i[2876] & sel_one_hot_i[44];
  assign data_masked[2875] = data_i[2875] & sel_one_hot_i[44];
  assign data_masked[2874] = data_i[2874] & sel_one_hot_i[44];
  assign data_masked[2873] = data_i[2873] & sel_one_hot_i[44];
  assign data_masked[2872] = data_i[2872] & sel_one_hot_i[44];
  assign data_masked[2871] = data_i[2871] & sel_one_hot_i[44];
  assign data_masked[2870] = data_i[2870] & sel_one_hot_i[44];
  assign data_masked[2869] = data_i[2869] & sel_one_hot_i[44];
  assign data_masked[2868] = data_i[2868] & sel_one_hot_i[44];
  assign data_masked[2867] = data_i[2867] & sel_one_hot_i[44];
  assign data_masked[2866] = data_i[2866] & sel_one_hot_i[44];
  assign data_masked[2865] = data_i[2865] & sel_one_hot_i[44];
  assign data_masked[2864] = data_i[2864] & sel_one_hot_i[44];
  assign data_masked[2863] = data_i[2863] & sel_one_hot_i[44];
  assign data_masked[2862] = data_i[2862] & sel_one_hot_i[44];
  assign data_masked[2861] = data_i[2861] & sel_one_hot_i[44];
  assign data_masked[2860] = data_i[2860] & sel_one_hot_i[44];
  assign data_masked[2859] = data_i[2859] & sel_one_hot_i[44];
  assign data_masked[2858] = data_i[2858] & sel_one_hot_i[44];
  assign data_masked[2857] = data_i[2857] & sel_one_hot_i[44];
  assign data_masked[2856] = data_i[2856] & sel_one_hot_i[44];
  assign data_masked[2855] = data_i[2855] & sel_one_hot_i[44];
  assign data_masked[2854] = data_i[2854] & sel_one_hot_i[44];
  assign data_masked[2853] = data_i[2853] & sel_one_hot_i[44];
  assign data_masked[2852] = data_i[2852] & sel_one_hot_i[44];
  assign data_masked[2851] = data_i[2851] & sel_one_hot_i[44];
  assign data_masked[2850] = data_i[2850] & sel_one_hot_i[44];
  assign data_masked[2849] = data_i[2849] & sel_one_hot_i[44];
  assign data_masked[2848] = data_i[2848] & sel_one_hot_i[44];
  assign data_masked[2847] = data_i[2847] & sel_one_hot_i[44];
  assign data_masked[2846] = data_i[2846] & sel_one_hot_i[44];
  assign data_masked[2845] = data_i[2845] & sel_one_hot_i[44];
  assign data_masked[2844] = data_i[2844] & sel_one_hot_i[44];
  assign data_masked[2843] = data_i[2843] & sel_one_hot_i[44];
  assign data_masked[2842] = data_i[2842] & sel_one_hot_i[44];
  assign data_masked[2841] = data_i[2841] & sel_one_hot_i[44];
  assign data_masked[2840] = data_i[2840] & sel_one_hot_i[44];
  assign data_masked[2839] = data_i[2839] & sel_one_hot_i[44];
  assign data_masked[2838] = data_i[2838] & sel_one_hot_i[44];
  assign data_masked[2837] = data_i[2837] & sel_one_hot_i[44];
  assign data_masked[2836] = data_i[2836] & sel_one_hot_i[44];
  assign data_masked[2835] = data_i[2835] & sel_one_hot_i[44];
  assign data_masked[2834] = data_i[2834] & sel_one_hot_i[44];
  assign data_masked[2833] = data_i[2833] & sel_one_hot_i[44];
  assign data_masked[2832] = data_i[2832] & sel_one_hot_i[44];
  assign data_masked[2831] = data_i[2831] & sel_one_hot_i[44];
  assign data_masked[2830] = data_i[2830] & sel_one_hot_i[44];
  assign data_masked[2829] = data_i[2829] & sel_one_hot_i[44];
  assign data_masked[2828] = data_i[2828] & sel_one_hot_i[44];
  assign data_masked[2827] = data_i[2827] & sel_one_hot_i[44];
  assign data_masked[2826] = data_i[2826] & sel_one_hot_i[44];
  assign data_masked[2825] = data_i[2825] & sel_one_hot_i[44];
  assign data_masked[2824] = data_i[2824] & sel_one_hot_i[44];
  assign data_masked[2823] = data_i[2823] & sel_one_hot_i[44];
  assign data_masked[2822] = data_i[2822] & sel_one_hot_i[44];
  assign data_masked[2821] = data_i[2821] & sel_one_hot_i[44];
  assign data_masked[2820] = data_i[2820] & sel_one_hot_i[44];
  assign data_masked[2819] = data_i[2819] & sel_one_hot_i[44];
  assign data_masked[2818] = data_i[2818] & sel_one_hot_i[44];
  assign data_masked[2817] = data_i[2817] & sel_one_hot_i[44];
  assign data_masked[2816] = data_i[2816] & sel_one_hot_i[44];
  assign data_masked[2943] = data_i[2943] & sel_one_hot_i[45];
  assign data_masked[2942] = data_i[2942] & sel_one_hot_i[45];
  assign data_masked[2941] = data_i[2941] & sel_one_hot_i[45];
  assign data_masked[2940] = data_i[2940] & sel_one_hot_i[45];
  assign data_masked[2939] = data_i[2939] & sel_one_hot_i[45];
  assign data_masked[2938] = data_i[2938] & sel_one_hot_i[45];
  assign data_masked[2937] = data_i[2937] & sel_one_hot_i[45];
  assign data_masked[2936] = data_i[2936] & sel_one_hot_i[45];
  assign data_masked[2935] = data_i[2935] & sel_one_hot_i[45];
  assign data_masked[2934] = data_i[2934] & sel_one_hot_i[45];
  assign data_masked[2933] = data_i[2933] & sel_one_hot_i[45];
  assign data_masked[2932] = data_i[2932] & sel_one_hot_i[45];
  assign data_masked[2931] = data_i[2931] & sel_one_hot_i[45];
  assign data_masked[2930] = data_i[2930] & sel_one_hot_i[45];
  assign data_masked[2929] = data_i[2929] & sel_one_hot_i[45];
  assign data_masked[2928] = data_i[2928] & sel_one_hot_i[45];
  assign data_masked[2927] = data_i[2927] & sel_one_hot_i[45];
  assign data_masked[2926] = data_i[2926] & sel_one_hot_i[45];
  assign data_masked[2925] = data_i[2925] & sel_one_hot_i[45];
  assign data_masked[2924] = data_i[2924] & sel_one_hot_i[45];
  assign data_masked[2923] = data_i[2923] & sel_one_hot_i[45];
  assign data_masked[2922] = data_i[2922] & sel_one_hot_i[45];
  assign data_masked[2921] = data_i[2921] & sel_one_hot_i[45];
  assign data_masked[2920] = data_i[2920] & sel_one_hot_i[45];
  assign data_masked[2919] = data_i[2919] & sel_one_hot_i[45];
  assign data_masked[2918] = data_i[2918] & sel_one_hot_i[45];
  assign data_masked[2917] = data_i[2917] & sel_one_hot_i[45];
  assign data_masked[2916] = data_i[2916] & sel_one_hot_i[45];
  assign data_masked[2915] = data_i[2915] & sel_one_hot_i[45];
  assign data_masked[2914] = data_i[2914] & sel_one_hot_i[45];
  assign data_masked[2913] = data_i[2913] & sel_one_hot_i[45];
  assign data_masked[2912] = data_i[2912] & sel_one_hot_i[45];
  assign data_masked[2911] = data_i[2911] & sel_one_hot_i[45];
  assign data_masked[2910] = data_i[2910] & sel_one_hot_i[45];
  assign data_masked[2909] = data_i[2909] & sel_one_hot_i[45];
  assign data_masked[2908] = data_i[2908] & sel_one_hot_i[45];
  assign data_masked[2907] = data_i[2907] & sel_one_hot_i[45];
  assign data_masked[2906] = data_i[2906] & sel_one_hot_i[45];
  assign data_masked[2905] = data_i[2905] & sel_one_hot_i[45];
  assign data_masked[2904] = data_i[2904] & sel_one_hot_i[45];
  assign data_masked[2903] = data_i[2903] & sel_one_hot_i[45];
  assign data_masked[2902] = data_i[2902] & sel_one_hot_i[45];
  assign data_masked[2901] = data_i[2901] & sel_one_hot_i[45];
  assign data_masked[2900] = data_i[2900] & sel_one_hot_i[45];
  assign data_masked[2899] = data_i[2899] & sel_one_hot_i[45];
  assign data_masked[2898] = data_i[2898] & sel_one_hot_i[45];
  assign data_masked[2897] = data_i[2897] & sel_one_hot_i[45];
  assign data_masked[2896] = data_i[2896] & sel_one_hot_i[45];
  assign data_masked[2895] = data_i[2895] & sel_one_hot_i[45];
  assign data_masked[2894] = data_i[2894] & sel_one_hot_i[45];
  assign data_masked[2893] = data_i[2893] & sel_one_hot_i[45];
  assign data_masked[2892] = data_i[2892] & sel_one_hot_i[45];
  assign data_masked[2891] = data_i[2891] & sel_one_hot_i[45];
  assign data_masked[2890] = data_i[2890] & sel_one_hot_i[45];
  assign data_masked[2889] = data_i[2889] & sel_one_hot_i[45];
  assign data_masked[2888] = data_i[2888] & sel_one_hot_i[45];
  assign data_masked[2887] = data_i[2887] & sel_one_hot_i[45];
  assign data_masked[2886] = data_i[2886] & sel_one_hot_i[45];
  assign data_masked[2885] = data_i[2885] & sel_one_hot_i[45];
  assign data_masked[2884] = data_i[2884] & sel_one_hot_i[45];
  assign data_masked[2883] = data_i[2883] & sel_one_hot_i[45];
  assign data_masked[2882] = data_i[2882] & sel_one_hot_i[45];
  assign data_masked[2881] = data_i[2881] & sel_one_hot_i[45];
  assign data_masked[2880] = data_i[2880] & sel_one_hot_i[45];
  assign data_masked[3007] = data_i[3007] & sel_one_hot_i[46];
  assign data_masked[3006] = data_i[3006] & sel_one_hot_i[46];
  assign data_masked[3005] = data_i[3005] & sel_one_hot_i[46];
  assign data_masked[3004] = data_i[3004] & sel_one_hot_i[46];
  assign data_masked[3003] = data_i[3003] & sel_one_hot_i[46];
  assign data_masked[3002] = data_i[3002] & sel_one_hot_i[46];
  assign data_masked[3001] = data_i[3001] & sel_one_hot_i[46];
  assign data_masked[3000] = data_i[3000] & sel_one_hot_i[46];
  assign data_masked[2999] = data_i[2999] & sel_one_hot_i[46];
  assign data_masked[2998] = data_i[2998] & sel_one_hot_i[46];
  assign data_masked[2997] = data_i[2997] & sel_one_hot_i[46];
  assign data_masked[2996] = data_i[2996] & sel_one_hot_i[46];
  assign data_masked[2995] = data_i[2995] & sel_one_hot_i[46];
  assign data_masked[2994] = data_i[2994] & sel_one_hot_i[46];
  assign data_masked[2993] = data_i[2993] & sel_one_hot_i[46];
  assign data_masked[2992] = data_i[2992] & sel_one_hot_i[46];
  assign data_masked[2991] = data_i[2991] & sel_one_hot_i[46];
  assign data_masked[2990] = data_i[2990] & sel_one_hot_i[46];
  assign data_masked[2989] = data_i[2989] & sel_one_hot_i[46];
  assign data_masked[2988] = data_i[2988] & sel_one_hot_i[46];
  assign data_masked[2987] = data_i[2987] & sel_one_hot_i[46];
  assign data_masked[2986] = data_i[2986] & sel_one_hot_i[46];
  assign data_masked[2985] = data_i[2985] & sel_one_hot_i[46];
  assign data_masked[2984] = data_i[2984] & sel_one_hot_i[46];
  assign data_masked[2983] = data_i[2983] & sel_one_hot_i[46];
  assign data_masked[2982] = data_i[2982] & sel_one_hot_i[46];
  assign data_masked[2981] = data_i[2981] & sel_one_hot_i[46];
  assign data_masked[2980] = data_i[2980] & sel_one_hot_i[46];
  assign data_masked[2979] = data_i[2979] & sel_one_hot_i[46];
  assign data_masked[2978] = data_i[2978] & sel_one_hot_i[46];
  assign data_masked[2977] = data_i[2977] & sel_one_hot_i[46];
  assign data_masked[2976] = data_i[2976] & sel_one_hot_i[46];
  assign data_masked[2975] = data_i[2975] & sel_one_hot_i[46];
  assign data_masked[2974] = data_i[2974] & sel_one_hot_i[46];
  assign data_masked[2973] = data_i[2973] & sel_one_hot_i[46];
  assign data_masked[2972] = data_i[2972] & sel_one_hot_i[46];
  assign data_masked[2971] = data_i[2971] & sel_one_hot_i[46];
  assign data_masked[2970] = data_i[2970] & sel_one_hot_i[46];
  assign data_masked[2969] = data_i[2969] & sel_one_hot_i[46];
  assign data_masked[2968] = data_i[2968] & sel_one_hot_i[46];
  assign data_masked[2967] = data_i[2967] & sel_one_hot_i[46];
  assign data_masked[2966] = data_i[2966] & sel_one_hot_i[46];
  assign data_masked[2965] = data_i[2965] & sel_one_hot_i[46];
  assign data_masked[2964] = data_i[2964] & sel_one_hot_i[46];
  assign data_masked[2963] = data_i[2963] & sel_one_hot_i[46];
  assign data_masked[2962] = data_i[2962] & sel_one_hot_i[46];
  assign data_masked[2961] = data_i[2961] & sel_one_hot_i[46];
  assign data_masked[2960] = data_i[2960] & sel_one_hot_i[46];
  assign data_masked[2959] = data_i[2959] & sel_one_hot_i[46];
  assign data_masked[2958] = data_i[2958] & sel_one_hot_i[46];
  assign data_masked[2957] = data_i[2957] & sel_one_hot_i[46];
  assign data_masked[2956] = data_i[2956] & sel_one_hot_i[46];
  assign data_masked[2955] = data_i[2955] & sel_one_hot_i[46];
  assign data_masked[2954] = data_i[2954] & sel_one_hot_i[46];
  assign data_masked[2953] = data_i[2953] & sel_one_hot_i[46];
  assign data_masked[2952] = data_i[2952] & sel_one_hot_i[46];
  assign data_masked[2951] = data_i[2951] & sel_one_hot_i[46];
  assign data_masked[2950] = data_i[2950] & sel_one_hot_i[46];
  assign data_masked[2949] = data_i[2949] & sel_one_hot_i[46];
  assign data_masked[2948] = data_i[2948] & sel_one_hot_i[46];
  assign data_masked[2947] = data_i[2947] & sel_one_hot_i[46];
  assign data_masked[2946] = data_i[2946] & sel_one_hot_i[46];
  assign data_masked[2945] = data_i[2945] & sel_one_hot_i[46];
  assign data_masked[2944] = data_i[2944] & sel_one_hot_i[46];
  assign data_masked[3071] = data_i[3071] & sel_one_hot_i[47];
  assign data_masked[3070] = data_i[3070] & sel_one_hot_i[47];
  assign data_masked[3069] = data_i[3069] & sel_one_hot_i[47];
  assign data_masked[3068] = data_i[3068] & sel_one_hot_i[47];
  assign data_masked[3067] = data_i[3067] & sel_one_hot_i[47];
  assign data_masked[3066] = data_i[3066] & sel_one_hot_i[47];
  assign data_masked[3065] = data_i[3065] & sel_one_hot_i[47];
  assign data_masked[3064] = data_i[3064] & sel_one_hot_i[47];
  assign data_masked[3063] = data_i[3063] & sel_one_hot_i[47];
  assign data_masked[3062] = data_i[3062] & sel_one_hot_i[47];
  assign data_masked[3061] = data_i[3061] & sel_one_hot_i[47];
  assign data_masked[3060] = data_i[3060] & sel_one_hot_i[47];
  assign data_masked[3059] = data_i[3059] & sel_one_hot_i[47];
  assign data_masked[3058] = data_i[3058] & sel_one_hot_i[47];
  assign data_masked[3057] = data_i[3057] & sel_one_hot_i[47];
  assign data_masked[3056] = data_i[3056] & sel_one_hot_i[47];
  assign data_masked[3055] = data_i[3055] & sel_one_hot_i[47];
  assign data_masked[3054] = data_i[3054] & sel_one_hot_i[47];
  assign data_masked[3053] = data_i[3053] & sel_one_hot_i[47];
  assign data_masked[3052] = data_i[3052] & sel_one_hot_i[47];
  assign data_masked[3051] = data_i[3051] & sel_one_hot_i[47];
  assign data_masked[3050] = data_i[3050] & sel_one_hot_i[47];
  assign data_masked[3049] = data_i[3049] & sel_one_hot_i[47];
  assign data_masked[3048] = data_i[3048] & sel_one_hot_i[47];
  assign data_masked[3047] = data_i[3047] & sel_one_hot_i[47];
  assign data_masked[3046] = data_i[3046] & sel_one_hot_i[47];
  assign data_masked[3045] = data_i[3045] & sel_one_hot_i[47];
  assign data_masked[3044] = data_i[3044] & sel_one_hot_i[47];
  assign data_masked[3043] = data_i[3043] & sel_one_hot_i[47];
  assign data_masked[3042] = data_i[3042] & sel_one_hot_i[47];
  assign data_masked[3041] = data_i[3041] & sel_one_hot_i[47];
  assign data_masked[3040] = data_i[3040] & sel_one_hot_i[47];
  assign data_masked[3039] = data_i[3039] & sel_one_hot_i[47];
  assign data_masked[3038] = data_i[3038] & sel_one_hot_i[47];
  assign data_masked[3037] = data_i[3037] & sel_one_hot_i[47];
  assign data_masked[3036] = data_i[3036] & sel_one_hot_i[47];
  assign data_masked[3035] = data_i[3035] & sel_one_hot_i[47];
  assign data_masked[3034] = data_i[3034] & sel_one_hot_i[47];
  assign data_masked[3033] = data_i[3033] & sel_one_hot_i[47];
  assign data_masked[3032] = data_i[3032] & sel_one_hot_i[47];
  assign data_masked[3031] = data_i[3031] & sel_one_hot_i[47];
  assign data_masked[3030] = data_i[3030] & sel_one_hot_i[47];
  assign data_masked[3029] = data_i[3029] & sel_one_hot_i[47];
  assign data_masked[3028] = data_i[3028] & sel_one_hot_i[47];
  assign data_masked[3027] = data_i[3027] & sel_one_hot_i[47];
  assign data_masked[3026] = data_i[3026] & sel_one_hot_i[47];
  assign data_masked[3025] = data_i[3025] & sel_one_hot_i[47];
  assign data_masked[3024] = data_i[3024] & sel_one_hot_i[47];
  assign data_masked[3023] = data_i[3023] & sel_one_hot_i[47];
  assign data_masked[3022] = data_i[3022] & sel_one_hot_i[47];
  assign data_masked[3021] = data_i[3021] & sel_one_hot_i[47];
  assign data_masked[3020] = data_i[3020] & sel_one_hot_i[47];
  assign data_masked[3019] = data_i[3019] & sel_one_hot_i[47];
  assign data_masked[3018] = data_i[3018] & sel_one_hot_i[47];
  assign data_masked[3017] = data_i[3017] & sel_one_hot_i[47];
  assign data_masked[3016] = data_i[3016] & sel_one_hot_i[47];
  assign data_masked[3015] = data_i[3015] & sel_one_hot_i[47];
  assign data_masked[3014] = data_i[3014] & sel_one_hot_i[47];
  assign data_masked[3013] = data_i[3013] & sel_one_hot_i[47];
  assign data_masked[3012] = data_i[3012] & sel_one_hot_i[47];
  assign data_masked[3011] = data_i[3011] & sel_one_hot_i[47];
  assign data_masked[3010] = data_i[3010] & sel_one_hot_i[47];
  assign data_masked[3009] = data_i[3009] & sel_one_hot_i[47];
  assign data_masked[3008] = data_i[3008] & sel_one_hot_i[47];
  assign data_masked[3135] = data_i[3135] & sel_one_hot_i[48];
  assign data_masked[3134] = data_i[3134] & sel_one_hot_i[48];
  assign data_masked[3133] = data_i[3133] & sel_one_hot_i[48];
  assign data_masked[3132] = data_i[3132] & sel_one_hot_i[48];
  assign data_masked[3131] = data_i[3131] & sel_one_hot_i[48];
  assign data_masked[3130] = data_i[3130] & sel_one_hot_i[48];
  assign data_masked[3129] = data_i[3129] & sel_one_hot_i[48];
  assign data_masked[3128] = data_i[3128] & sel_one_hot_i[48];
  assign data_masked[3127] = data_i[3127] & sel_one_hot_i[48];
  assign data_masked[3126] = data_i[3126] & sel_one_hot_i[48];
  assign data_masked[3125] = data_i[3125] & sel_one_hot_i[48];
  assign data_masked[3124] = data_i[3124] & sel_one_hot_i[48];
  assign data_masked[3123] = data_i[3123] & sel_one_hot_i[48];
  assign data_masked[3122] = data_i[3122] & sel_one_hot_i[48];
  assign data_masked[3121] = data_i[3121] & sel_one_hot_i[48];
  assign data_masked[3120] = data_i[3120] & sel_one_hot_i[48];
  assign data_masked[3119] = data_i[3119] & sel_one_hot_i[48];
  assign data_masked[3118] = data_i[3118] & sel_one_hot_i[48];
  assign data_masked[3117] = data_i[3117] & sel_one_hot_i[48];
  assign data_masked[3116] = data_i[3116] & sel_one_hot_i[48];
  assign data_masked[3115] = data_i[3115] & sel_one_hot_i[48];
  assign data_masked[3114] = data_i[3114] & sel_one_hot_i[48];
  assign data_masked[3113] = data_i[3113] & sel_one_hot_i[48];
  assign data_masked[3112] = data_i[3112] & sel_one_hot_i[48];
  assign data_masked[3111] = data_i[3111] & sel_one_hot_i[48];
  assign data_masked[3110] = data_i[3110] & sel_one_hot_i[48];
  assign data_masked[3109] = data_i[3109] & sel_one_hot_i[48];
  assign data_masked[3108] = data_i[3108] & sel_one_hot_i[48];
  assign data_masked[3107] = data_i[3107] & sel_one_hot_i[48];
  assign data_masked[3106] = data_i[3106] & sel_one_hot_i[48];
  assign data_masked[3105] = data_i[3105] & sel_one_hot_i[48];
  assign data_masked[3104] = data_i[3104] & sel_one_hot_i[48];
  assign data_masked[3103] = data_i[3103] & sel_one_hot_i[48];
  assign data_masked[3102] = data_i[3102] & sel_one_hot_i[48];
  assign data_masked[3101] = data_i[3101] & sel_one_hot_i[48];
  assign data_masked[3100] = data_i[3100] & sel_one_hot_i[48];
  assign data_masked[3099] = data_i[3099] & sel_one_hot_i[48];
  assign data_masked[3098] = data_i[3098] & sel_one_hot_i[48];
  assign data_masked[3097] = data_i[3097] & sel_one_hot_i[48];
  assign data_masked[3096] = data_i[3096] & sel_one_hot_i[48];
  assign data_masked[3095] = data_i[3095] & sel_one_hot_i[48];
  assign data_masked[3094] = data_i[3094] & sel_one_hot_i[48];
  assign data_masked[3093] = data_i[3093] & sel_one_hot_i[48];
  assign data_masked[3092] = data_i[3092] & sel_one_hot_i[48];
  assign data_masked[3091] = data_i[3091] & sel_one_hot_i[48];
  assign data_masked[3090] = data_i[3090] & sel_one_hot_i[48];
  assign data_masked[3089] = data_i[3089] & sel_one_hot_i[48];
  assign data_masked[3088] = data_i[3088] & sel_one_hot_i[48];
  assign data_masked[3087] = data_i[3087] & sel_one_hot_i[48];
  assign data_masked[3086] = data_i[3086] & sel_one_hot_i[48];
  assign data_masked[3085] = data_i[3085] & sel_one_hot_i[48];
  assign data_masked[3084] = data_i[3084] & sel_one_hot_i[48];
  assign data_masked[3083] = data_i[3083] & sel_one_hot_i[48];
  assign data_masked[3082] = data_i[3082] & sel_one_hot_i[48];
  assign data_masked[3081] = data_i[3081] & sel_one_hot_i[48];
  assign data_masked[3080] = data_i[3080] & sel_one_hot_i[48];
  assign data_masked[3079] = data_i[3079] & sel_one_hot_i[48];
  assign data_masked[3078] = data_i[3078] & sel_one_hot_i[48];
  assign data_masked[3077] = data_i[3077] & sel_one_hot_i[48];
  assign data_masked[3076] = data_i[3076] & sel_one_hot_i[48];
  assign data_masked[3075] = data_i[3075] & sel_one_hot_i[48];
  assign data_masked[3074] = data_i[3074] & sel_one_hot_i[48];
  assign data_masked[3073] = data_i[3073] & sel_one_hot_i[48];
  assign data_masked[3072] = data_i[3072] & sel_one_hot_i[48];
  assign data_masked[3199] = data_i[3199] & sel_one_hot_i[49];
  assign data_masked[3198] = data_i[3198] & sel_one_hot_i[49];
  assign data_masked[3197] = data_i[3197] & sel_one_hot_i[49];
  assign data_masked[3196] = data_i[3196] & sel_one_hot_i[49];
  assign data_masked[3195] = data_i[3195] & sel_one_hot_i[49];
  assign data_masked[3194] = data_i[3194] & sel_one_hot_i[49];
  assign data_masked[3193] = data_i[3193] & sel_one_hot_i[49];
  assign data_masked[3192] = data_i[3192] & sel_one_hot_i[49];
  assign data_masked[3191] = data_i[3191] & sel_one_hot_i[49];
  assign data_masked[3190] = data_i[3190] & sel_one_hot_i[49];
  assign data_masked[3189] = data_i[3189] & sel_one_hot_i[49];
  assign data_masked[3188] = data_i[3188] & sel_one_hot_i[49];
  assign data_masked[3187] = data_i[3187] & sel_one_hot_i[49];
  assign data_masked[3186] = data_i[3186] & sel_one_hot_i[49];
  assign data_masked[3185] = data_i[3185] & sel_one_hot_i[49];
  assign data_masked[3184] = data_i[3184] & sel_one_hot_i[49];
  assign data_masked[3183] = data_i[3183] & sel_one_hot_i[49];
  assign data_masked[3182] = data_i[3182] & sel_one_hot_i[49];
  assign data_masked[3181] = data_i[3181] & sel_one_hot_i[49];
  assign data_masked[3180] = data_i[3180] & sel_one_hot_i[49];
  assign data_masked[3179] = data_i[3179] & sel_one_hot_i[49];
  assign data_masked[3178] = data_i[3178] & sel_one_hot_i[49];
  assign data_masked[3177] = data_i[3177] & sel_one_hot_i[49];
  assign data_masked[3176] = data_i[3176] & sel_one_hot_i[49];
  assign data_masked[3175] = data_i[3175] & sel_one_hot_i[49];
  assign data_masked[3174] = data_i[3174] & sel_one_hot_i[49];
  assign data_masked[3173] = data_i[3173] & sel_one_hot_i[49];
  assign data_masked[3172] = data_i[3172] & sel_one_hot_i[49];
  assign data_masked[3171] = data_i[3171] & sel_one_hot_i[49];
  assign data_masked[3170] = data_i[3170] & sel_one_hot_i[49];
  assign data_masked[3169] = data_i[3169] & sel_one_hot_i[49];
  assign data_masked[3168] = data_i[3168] & sel_one_hot_i[49];
  assign data_masked[3167] = data_i[3167] & sel_one_hot_i[49];
  assign data_masked[3166] = data_i[3166] & sel_one_hot_i[49];
  assign data_masked[3165] = data_i[3165] & sel_one_hot_i[49];
  assign data_masked[3164] = data_i[3164] & sel_one_hot_i[49];
  assign data_masked[3163] = data_i[3163] & sel_one_hot_i[49];
  assign data_masked[3162] = data_i[3162] & sel_one_hot_i[49];
  assign data_masked[3161] = data_i[3161] & sel_one_hot_i[49];
  assign data_masked[3160] = data_i[3160] & sel_one_hot_i[49];
  assign data_masked[3159] = data_i[3159] & sel_one_hot_i[49];
  assign data_masked[3158] = data_i[3158] & sel_one_hot_i[49];
  assign data_masked[3157] = data_i[3157] & sel_one_hot_i[49];
  assign data_masked[3156] = data_i[3156] & sel_one_hot_i[49];
  assign data_masked[3155] = data_i[3155] & sel_one_hot_i[49];
  assign data_masked[3154] = data_i[3154] & sel_one_hot_i[49];
  assign data_masked[3153] = data_i[3153] & sel_one_hot_i[49];
  assign data_masked[3152] = data_i[3152] & sel_one_hot_i[49];
  assign data_masked[3151] = data_i[3151] & sel_one_hot_i[49];
  assign data_masked[3150] = data_i[3150] & sel_one_hot_i[49];
  assign data_masked[3149] = data_i[3149] & sel_one_hot_i[49];
  assign data_masked[3148] = data_i[3148] & sel_one_hot_i[49];
  assign data_masked[3147] = data_i[3147] & sel_one_hot_i[49];
  assign data_masked[3146] = data_i[3146] & sel_one_hot_i[49];
  assign data_masked[3145] = data_i[3145] & sel_one_hot_i[49];
  assign data_masked[3144] = data_i[3144] & sel_one_hot_i[49];
  assign data_masked[3143] = data_i[3143] & sel_one_hot_i[49];
  assign data_masked[3142] = data_i[3142] & sel_one_hot_i[49];
  assign data_masked[3141] = data_i[3141] & sel_one_hot_i[49];
  assign data_masked[3140] = data_i[3140] & sel_one_hot_i[49];
  assign data_masked[3139] = data_i[3139] & sel_one_hot_i[49];
  assign data_masked[3138] = data_i[3138] & sel_one_hot_i[49];
  assign data_masked[3137] = data_i[3137] & sel_one_hot_i[49];
  assign data_masked[3136] = data_i[3136] & sel_one_hot_i[49];
  assign data_masked[3263] = data_i[3263] & sel_one_hot_i[50];
  assign data_masked[3262] = data_i[3262] & sel_one_hot_i[50];
  assign data_masked[3261] = data_i[3261] & sel_one_hot_i[50];
  assign data_masked[3260] = data_i[3260] & sel_one_hot_i[50];
  assign data_masked[3259] = data_i[3259] & sel_one_hot_i[50];
  assign data_masked[3258] = data_i[3258] & sel_one_hot_i[50];
  assign data_masked[3257] = data_i[3257] & sel_one_hot_i[50];
  assign data_masked[3256] = data_i[3256] & sel_one_hot_i[50];
  assign data_masked[3255] = data_i[3255] & sel_one_hot_i[50];
  assign data_masked[3254] = data_i[3254] & sel_one_hot_i[50];
  assign data_masked[3253] = data_i[3253] & sel_one_hot_i[50];
  assign data_masked[3252] = data_i[3252] & sel_one_hot_i[50];
  assign data_masked[3251] = data_i[3251] & sel_one_hot_i[50];
  assign data_masked[3250] = data_i[3250] & sel_one_hot_i[50];
  assign data_masked[3249] = data_i[3249] & sel_one_hot_i[50];
  assign data_masked[3248] = data_i[3248] & sel_one_hot_i[50];
  assign data_masked[3247] = data_i[3247] & sel_one_hot_i[50];
  assign data_masked[3246] = data_i[3246] & sel_one_hot_i[50];
  assign data_masked[3245] = data_i[3245] & sel_one_hot_i[50];
  assign data_masked[3244] = data_i[3244] & sel_one_hot_i[50];
  assign data_masked[3243] = data_i[3243] & sel_one_hot_i[50];
  assign data_masked[3242] = data_i[3242] & sel_one_hot_i[50];
  assign data_masked[3241] = data_i[3241] & sel_one_hot_i[50];
  assign data_masked[3240] = data_i[3240] & sel_one_hot_i[50];
  assign data_masked[3239] = data_i[3239] & sel_one_hot_i[50];
  assign data_masked[3238] = data_i[3238] & sel_one_hot_i[50];
  assign data_masked[3237] = data_i[3237] & sel_one_hot_i[50];
  assign data_masked[3236] = data_i[3236] & sel_one_hot_i[50];
  assign data_masked[3235] = data_i[3235] & sel_one_hot_i[50];
  assign data_masked[3234] = data_i[3234] & sel_one_hot_i[50];
  assign data_masked[3233] = data_i[3233] & sel_one_hot_i[50];
  assign data_masked[3232] = data_i[3232] & sel_one_hot_i[50];
  assign data_masked[3231] = data_i[3231] & sel_one_hot_i[50];
  assign data_masked[3230] = data_i[3230] & sel_one_hot_i[50];
  assign data_masked[3229] = data_i[3229] & sel_one_hot_i[50];
  assign data_masked[3228] = data_i[3228] & sel_one_hot_i[50];
  assign data_masked[3227] = data_i[3227] & sel_one_hot_i[50];
  assign data_masked[3226] = data_i[3226] & sel_one_hot_i[50];
  assign data_masked[3225] = data_i[3225] & sel_one_hot_i[50];
  assign data_masked[3224] = data_i[3224] & sel_one_hot_i[50];
  assign data_masked[3223] = data_i[3223] & sel_one_hot_i[50];
  assign data_masked[3222] = data_i[3222] & sel_one_hot_i[50];
  assign data_masked[3221] = data_i[3221] & sel_one_hot_i[50];
  assign data_masked[3220] = data_i[3220] & sel_one_hot_i[50];
  assign data_masked[3219] = data_i[3219] & sel_one_hot_i[50];
  assign data_masked[3218] = data_i[3218] & sel_one_hot_i[50];
  assign data_masked[3217] = data_i[3217] & sel_one_hot_i[50];
  assign data_masked[3216] = data_i[3216] & sel_one_hot_i[50];
  assign data_masked[3215] = data_i[3215] & sel_one_hot_i[50];
  assign data_masked[3214] = data_i[3214] & sel_one_hot_i[50];
  assign data_masked[3213] = data_i[3213] & sel_one_hot_i[50];
  assign data_masked[3212] = data_i[3212] & sel_one_hot_i[50];
  assign data_masked[3211] = data_i[3211] & sel_one_hot_i[50];
  assign data_masked[3210] = data_i[3210] & sel_one_hot_i[50];
  assign data_masked[3209] = data_i[3209] & sel_one_hot_i[50];
  assign data_masked[3208] = data_i[3208] & sel_one_hot_i[50];
  assign data_masked[3207] = data_i[3207] & sel_one_hot_i[50];
  assign data_masked[3206] = data_i[3206] & sel_one_hot_i[50];
  assign data_masked[3205] = data_i[3205] & sel_one_hot_i[50];
  assign data_masked[3204] = data_i[3204] & sel_one_hot_i[50];
  assign data_masked[3203] = data_i[3203] & sel_one_hot_i[50];
  assign data_masked[3202] = data_i[3202] & sel_one_hot_i[50];
  assign data_masked[3201] = data_i[3201] & sel_one_hot_i[50];
  assign data_masked[3200] = data_i[3200] & sel_one_hot_i[50];
  assign data_masked[3327] = data_i[3327] & sel_one_hot_i[51];
  assign data_masked[3326] = data_i[3326] & sel_one_hot_i[51];
  assign data_masked[3325] = data_i[3325] & sel_one_hot_i[51];
  assign data_masked[3324] = data_i[3324] & sel_one_hot_i[51];
  assign data_masked[3323] = data_i[3323] & sel_one_hot_i[51];
  assign data_masked[3322] = data_i[3322] & sel_one_hot_i[51];
  assign data_masked[3321] = data_i[3321] & sel_one_hot_i[51];
  assign data_masked[3320] = data_i[3320] & sel_one_hot_i[51];
  assign data_masked[3319] = data_i[3319] & sel_one_hot_i[51];
  assign data_masked[3318] = data_i[3318] & sel_one_hot_i[51];
  assign data_masked[3317] = data_i[3317] & sel_one_hot_i[51];
  assign data_masked[3316] = data_i[3316] & sel_one_hot_i[51];
  assign data_masked[3315] = data_i[3315] & sel_one_hot_i[51];
  assign data_masked[3314] = data_i[3314] & sel_one_hot_i[51];
  assign data_masked[3313] = data_i[3313] & sel_one_hot_i[51];
  assign data_masked[3312] = data_i[3312] & sel_one_hot_i[51];
  assign data_masked[3311] = data_i[3311] & sel_one_hot_i[51];
  assign data_masked[3310] = data_i[3310] & sel_one_hot_i[51];
  assign data_masked[3309] = data_i[3309] & sel_one_hot_i[51];
  assign data_masked[3308] = data_i[3308] & sel_one_hot_i[51];
  assign data_masked[3307] = data_i[3307] & sel_one_hot_i[51];
  assign data_masked[3306] = data_i[3306] & sel_one_hot_i[51];
  assign data_masked[3305] = data_i[3305] & sel_one_hot_i[51];
  assign data_masked[3304] = data_i[3304] & sel_one_hot_i[51];
  assign data_masked[3303] = data_i[3303] & sel_one_hot_i[51];
  assign data_masked[3302] = data_i[3302] & sel_one_hot_i[51];
  assign data_masked[3301] = data_i[3301] & sel_one_hot_i[51];
  assign data_masked[3300] = data_i[3300] & sel_one_hot_i[51];
  assign data_masked[3299] = data_i[3299] & sel_one_hot_i[51];
  assign data_masked[3298] = data_i[3298] & sel_one_hot_i[51];
  assign data_masked[3297] = data_i[3297] & sel_one_hot_i[51];
  assign data_masked[3296] = data_i[3296] & sel_one_hot_i[51];
  assign data_masked[3295] = data_i[3295] & sel_one_hot_i[51];
  assign data_masked[3294] = data_i[3294] & sel_one_hot_i[51];
  assign data_masked[3293] = data_i[3293] & sel_one_hot_i[51];
  assign data_masked[3292] = data_i[3292] & sel_one_hot_i[51];
  assign data_masked[3291] = data_i[3291] & sel_one_hot_i[51];
  assign data_masked[3290] = data_i[3290] & sel_one_hot_i[51];
  assign data_masked[3289] = data_i[3289] & sel_one_hot_i[51];
  assign data_masked[3288] = data_i[3288] & sel_one_hot_i[51];
  assign data_masked[3287] = data_i[3287] & sel_one_hot_i[51];
  assign data_masked[3286] = data_i[3286] & sel_one_hot_i[51];
  assign data_masked[3285] = data_i[3285] & sel_one_hot_i[51];
  assign data_masked[3284] = data_i[3284] & sel_one_hot_i[51];
  assign data_masked[3283] = data_i[3283] & sel_one_hot_i[51];
  assign data_masked[3282] = data_i[3282] & sel_one_hot_i[51];
  assign data_masked[3281] = data_i[3281] & sel_one_hot_i[51];
  assign data_masked[3280] = data_i[3280] & sel_one_hot_i[51];
  assign data_masked[3279] = data_i[3279] & sel_one_hot_i[51];
  assign data_masked[3278] = data_i[3278] & sel_one_hot_i[51];
  assign data_masked[3277] = data_i[3277] & sel_one_hot_i[51];
  assign data_masked[3276] = data_i[3276] & sel_one_hot_i[51];
  assign data_masked[3275] = data_i[3275] & sel_one_hot_i[51];
  assign data_masked[3274] = data_i[3274] & sel_one_hot_i[51];
  assign data_masked[3273] = data_i[3273] & sel_one_hot_i[51];
  assign data_masked[3272] = data_i[3272] & sel_one_hot_i[51];
  assign data_masked[3271] = data_i[3271] & sel_one_hot_i[51];
  assign data_masked[3270] = data_i[3270] & sel_one_hot_i[51];
  assign data_masked[3269] = data_i[3269] & sel_one_hot_i[51];
  assign data_masked[3268] = data_i[3268] & sel_one_hot_i[51];
  assign data_masked[3267] = data_i[3267] & sel_one_hot_i[51];
  assign data_masked[3266] = data_i[3266] & sel_one_hot_i[51];
  assign data_masked[3265] = data_i[3265] & sel_one_hot_i[51];
  assign data_masked[3264] = data_i[3264] & sel_one_hot_i[51];
  assign data_masked[3391] = data_i[3391] & sel_one_hot_i[52];
  assign data_masked[3390] = data_i[3390] & sel_one_hot_i[52];
  assign data_masked[3389] = data_i[3389] & sel_one_hot_i[52];
  assign data_masked[3388] = data_i[3388] & sel_one_hot_i[52];
  assign data_masked[3387] = data_i[3387] & sel_one_hot_i[52];
  assign data_masked[3386] = data_i[3386] & sel_one_hot_i[52];
  assign data_masked[3385] = data_i[3385] & sel_one_hot_i[52];
  assign data_masked[3384] = data_i[3384] & sel_one_hot_i[52];
  assign data_masked[3383] = data_i[3383] & sel_one_hot_i[52];
  assign data_masked[3382] = data_i[3382] & sel_one_hot_i[52];
  assign data_masked[3381] = data_i[3381] & sel_one_hot_i[52];
  assign data_masked[3380] = data_i[3380] & sel_one_hot_i[52];
  assign data_masked[3379] = data_i[3379] & sel_one_hot_i[52];
  assign data_masked[3378] = data_i[3378] & sel_one_hot_i[52];
  assign data_masked[3377] = data_i[3377] & sel_one_hot_i[52];
  assign data_masked[3376] = data_i[3376] & sel_one_hot_i[52];
  assign data_masked[3375] = data_i[3375] & sel_one_hot_i[52];
  assign data_masked[3374] = data_i[3374] & sel_one_hot_i[52];
  assign data_masked[3373] = data_i[3373] & sel_one_hot_i[52];
  assign data_masked[3372] = data_i[3372] & sel_one_hot_i[52];
  assign data_masked[3371] = data_i[3371] & sel_one_hot_i[52];
  assign data_masked[3370] = data_i[3370] & sel_one_hot_i[52];
  assign data_masked[3369] = data_i[3369] & sel_one_hot_i[52];
  assign data_masked[3368] = data_i[3368] & sel_one_hot_i[52];
  assign data_masked[3367] = data_i[3367] & sel_one_hot_i[52];
  assign data_masked[3366] = data_i[3366] & sel_one_hot_i[52];
  assign data_masked[3365] = data_i[3365] & sel_one_hot_i[52];
  assign data_masked[3364] = data_i[3364] & sel_one_hot_i[52];
  assign data_masked[3363] = data_i[3363] & sel_one_hot_i[52];
  assign data_masked[3362] = data_i[3362] & sel_one_hot_i[52];
  assign data_masked[3361] = data_i[3361] & sel_one_hot_i[52];
  assign data_masked[3360] = data_i[3360] & sel_one_hot_i[52];
  assign data_masked[3359] = data_i[3359] & sel_one_hot_i[52];
  assign data_masked[3358] = data_i[3358] & sel_one_hot_i[52];
  assign data_masked[3357] = data_i[3357] & sel_one_hot_i[52];
  assign data_masked[3356] = data_i[3356] & sel_one_hot_i[52];
  assign data_masked[3355] = data_i[3355] & sel_one_hot_i[52];
  assign data_masked[3354] = data_i[3354] & sel_one_hot_i[52];
  assign data_masked[3353] = data_i[3353] & sel_one_hot_i[52];
  assign data_masked[3352] = data_i[3352] & sel_one_hot_i[52];
  assign data_masked[3351] = data_i[3351] & sel_one_hot_i[52];
  assign data_masked[3350] = data_i[3350] & sel_one_hot_i[52];
  assign data_masked[3349] = data_i[3349] & sel_one_hot_i[52];
  assign data_masked[3348] = data_i[3348] & sel_one_hot_i[52];
  assign data_masked[3347] = data_i[3347] & sel_one_hot_i[52];
  assign data_masked[3346] = data_i[3346] & sel_one_hot_i[52];
  assign data_masked[3345] = data_i[3345] & sel_one_hot_i[52];
  assign data_masked[3344] = data_i[3344] & sel_one_hot_i[52];
  assign data_masked[3343] = data_i[3343] & sel_one_hot_i[52];
  assign data_masked[3342] = data_i[3342] & sel_one_hot_i[52];
  assign data_masked[3341] = data_i[3341] & sel_one_hot_i[52];
  assign data_masked[3340] = data_i[3340] & sel_one_hot_i[52];
  assign data_masked[3339] = data_i[3339] & sel_one_hot_i[52];
  assign data_masked[3338] = data_i[3338] & sel_one_hot_i[52];
  assign data_masked[3337] = data_i[3337] & sel_one_hot_i[52];
  assign data_masked[3336] = data_i[3336] & sel_one_hot_i[52];
  assign data_masked[3335] = data_i[3335] & sel_one_hot_i[52];
  assign data_masked[3334] = data_i[3334] & sel_one_hot_i[52];
  assign data_masked[3333] = data_i[3333] & sel_one_hot_i[52];
  assign data_masked[3332] = data_i[3332] & sel_one_hot_i[52];
  assign data_masked[3331] = data_i[3331] & sel_one_hot_i[52];
  assign data_masked[3330] = data_i[3330] & sel_one_hot_i[52];
  assign data_masked[3329] = data_i[3329] & sel_one_hot_i[52];
  assign data_masked[3328] = data_i[3328] & sel_one_hot_i[52];
  assign data_masked[3455] = data_i[3455] & sel_one_hot_i[53];
  assign data_masked[3454] = data_i[3454] & sel_one_hot_i[53];
  assign data_masked[3453] = data_i[3453] & sel_one_hot_i[53];
  assign data_masked[3452] = data_i[3452] & sel_one_hot_i[53];
  assign data_masked[3451] = data_i[3451] & sel_one_hot_i[53];
  assign data_masked[3450] = data_i[3450] & sel_one_hot_i[53];
  assign data_masked[3449] = data_i[3449] & sel_one_hot_i[53];
  assign data_masked[3448] = data_i[3448] & sel_one_hot_i[53];
  assign data_masked[3447] = data_i[3447] & sel_one_hot_i[53];
  assign data_masked[3446] = data_i[3446] & sel_one_hot_i[53];
  assign data_masked[3445] = data_i[3445] & sel_one_hot_i[53];
  assign data_masked[3444] = data_i[3444] & sel_one_hot_i[53];
  assign data_masked[3443] = data_i[3443] & sel_one_hot_i[53];
  assign data_masked[3442] = data_i[3442] & sel_one_hot_i[53];
  assign data_masked[3441] = data_i[3441] & sel_one_hot_i[53];
  assign data_masked[3440] = data_i[3440] & sel_one_hot_i[53];
  assign data_masked[3439] = data_i[3439] & sel_one_hot_i[53];
  assign data_masked[3438] = data_i[3438] & sel_one_hot_i[53];
  assign data_masked[3437] = data_i[3437] & sel_one_hot_i[53];
  assign data_masked[3436] = data_i[3436] & sel_one_hot_i[53];
  assign data_masked[3435] = data_i[3435] & sel_one_hot_i[53];
  assign data_masked[3434] = data_i[3434] & sel_one_hot_i[53];
  assign data_masked[3433] = data_i[3433] & sel_one_hot_i[53];
  assign data_masked[3432] = data_i[3432] & sel_one_hot_i[53];
  assign data_masked[3431] = data_i[3431] & sel_one_hot_i[53];
  assign data_masked[3430] = data_i[3430] & sel_one_hot_i[53];
  assign data_masked[3429] = data_i[3429] & sel_one_hot_i[53];
  assign data_masked[3428] = data_i[3428] & sel_one_hot_i[53];
  assign data_masked[3427] = data_i[3427] & sel_one_hot_i[53];
  assign data_masked[3426] = data_i[3426] & sel_one_hot_i[53];
  assign data_masked[3425] = data_i[3425] & sel_one_hot_i[53];
  assign data_masked[3424] = data_i[3424] & sel_one_hot_i[53];
  assign data_masked[3423] = data_i[3423] & sel_one_hot_i[53];
  assign data_masked[3422] = data_i[3422] & sel_one_hot_i[53];
  assign data_masked[3421] = data_i[3421] & sel_one_hot_i[53];
  assign data_masked[3420] = data_i[3420] & sel_one_hot_i[53];
  assign data_masked[3419] = data_i[3419] & sel_one_hot_i[53];
  assign data_masked[3418] = data_i[3418] & sel_one_hot_i[53];
  assign data_masked[3417] = data_i[3417] & sel_one_hot_i[53];
  assign data_masked[3416] = data_i[3416] & sel_one_hot_i[53];
  assign data_masked[3415] = data_i[3415] & sel_one_hot_i[53];
  assign data_masked[3414] = data_i[3414] & sel_one_hot_i[53];
  assign data_masked[3413] = data_i[3413] & sel_one_hot_i[53];
  assign data_masked[3412] = data_i[3412] & sel_one_hot_i[53];
  assign data_masked[3411] = data_i[3411] & sel_one_hot_i[53];
  assign data_masked[3410] = data_i[3410] & sel_one_hot_i[53];
  assign data_masked[3409] = data_i[3409] & sel_one_hot_i[53];
  assign data_masked[3408] = data_i[3408] & sel_one_hot_i[53];
  assign data_masked[3407] = data_i[3407] & sel_one_hot_i[53];
  assign data_masked[3406] = data_i[3406] & sel_one_hot_i[53];
  assign data_masked[3405] = data_i[3405] & sel_one_hot_i[53];
  assign data_masked[3404] = data_i[3404] & sel_one_hot_i[53];
  assign data_masked[3403] = data_i[3403] & sel_one_hot_i[53];
  assign data_masked[3402] = data_i[3402] & sel_one_hot_i[53];
  assign data_masked[3401] = data_i[3401] & sel_one_hot_i[53];
  assign data_masked[3400] = data_i[3400] & sel_one_hot_i[53];
  assign data_masked[3399] = data_i[3399] & sel_one_hot_i[53];
  assign data_masked[3398] = data_i[3398] & sel_one_hot_i[53];
  assign data_masked[3397] = data_i[3397] & sel_one_hot_i[53];
  assign data_masked[3396] = data_i[3396] & sel_one_hot_i[53];
  assign data_masked[3395] = data_i[3395] & sel_one_hot_i[53];
  assign data_masked[3394] = data_i[3394] & sel_one_hot_i[53];
  assign data_masked[3393] = data_i[3393] & sel_one_hot_i[53];
  assign data_masked[3392] = data_i[3392] & sel_one_hot_i[53];
  assign data_masked[3519] = data_i[3519] & sel_one_hot_i[54];
  assign data_masked[3518] = data_i[3518] & sel_one_hot_i[54];
  assign data_masked[3517] = data_i[3517] & sel_one_hot_i[54];
  assign data_masked[3516] = data_i[3516] & sel_one_hot_i[54];
  assign data_masked[3515] = data_i[3515] & sel_one_hot_i[54];
  assign data_masked[3514] = data_i[3514] & sel_one_hot_i[54];
  assign data_masked[3513] = data_i[3513] & sel_one_hot_i[54];
  assign data_masked[3512] = data_i[3512] & sel_one_hot_i[54];
  assign data_masked[3511] = data_i[3511] & sel_one_hot_i[54];
  assign data_masked[3510] = data_i[3510] & sel_one_hot_i[54];
  assign data_masked[3509] = data_i[3509] & sel_one_hot_i[54];
  assign data_masked[3508] = data_i[3508] & sel_one_hot_i[54];
  assign data_masked[3507] = data_i[3507] & sel_one_hot_i[54];
  assign data_masked[3506] = data_i[3506] & sel_one_hot_i[54];
  assign data_masked[3505] = data_i[3505] & sel_one_hot_i[54];
  assign data_masked[3504] = data_i[3504] & sel_one_hot_i[54];
  assign data_masked[3503] = data_i[3503] & sel_one_hot_i[54];
  assign data_masked[3502] = data_i[3502] & sel_one_hot_i[54];
  assign data_masked[3501] = data_i[3501] & sel_one_hot_i[54];
  assign data_masked[3500] = data_i[3500] & sel_one_hot_i[54];
  assign data_masked[3499] = data_i[3499] & sel_one_hot_i[54];
  assign data_masked[3498] = data_i[3498] & sel_one_hot_i[54];
  assign data_masked[3497] = data_i[3497] & sel_one_hot_i[54];
  assign data_masked[3496] = data_i[3496] & sel_one_hot_i[54];
  assign data_masked[3495] = data_i[3495] & sel_one_hot_i[54];
  assign data_masked[3494] = data_i[3494] & sel_one_hot_i[54];
  assign data_masked[3493] = data_i[3493] & sel_one_hot_i[54];
  assign data_masked[3492] = data_i[3492] & sel_one_hot_i[54];
  assign data_masked[3491] = data_i[3491] & sel_one_hot_i[54];
  assign data_masked[3490] = data_i[3490] & sel_one_hot_i[54];
  assign data_masked[3489] = data_i[3489] & sel_one_hot_i[54];
  assign data_masked[3488] = data_i[3488] & sel_one_hot_i[54];
  assign data_masked[3487] = data_i[3487] & sel_one_hot_i[54];
  assign data_masked[3486] = data_i[3486] & sel_one_hot_i[54];
  assign data_masked[3485] = data_i[3485] & sel_one_hot_i[54];
  assign data_masked[3484] = data_i[3484] & sel_one_hot_i[54];
  assign data_masked[3483] = data_i[3483] & sel_one_hot_i[54];
  assign data_masked[3482] = data_i[3482] & sel_one_hot_i[54];
  assign data_masked[3481] = data_i[3481] & sel_one_hot_i[54];
  assign data_masked[3480] = data_i[3480] & sel_one_hot_i[54];
  assign data_masked[3479] = data_i[3479] & sel_one_hot_i[54];
  assign data_masked[3478] = data_i[3478] & sel_one_hot_i[54];
  assign data_masked[3477] = data_i[3477] & sel_one_hot_i[54];
  assign data_masked[3476] = data_i[3476] & sel_one_hot_i[54];
  assign data_masked[3475] = data_i[3475] & sel_one_hot_i[54];
  assign data_masked[3474] = data_i[3474] & sel_one_hot_i[54];
  assign data_masked[3473] = data_i[3473] & sel_one_hot_i[54];
  assign data_masked[3472] = data_i[3472] & sel_one_hot_i[54];
  assign data_masked[3471] = data_i[3471] & sel_one_hot_i[54];
  assign data_masked[3470] = data_i[3470] & sel_one_hot_i[54];
  assign data_masked[3469] = data_i[3469] & sel_one_hot_i[54];
  assign data_masked[3468] = data_i[3468] & sel_one_hot_i[54];
  assign data_masked[3467] = data_i[3467] & sel_one_hot_i[54];
  assign data_masked[3466] = data_i[3466] & sel_one_hot_i[54];
  assign data_masked[3465] = data_i[3465] & sel_one_hot_i[54];
  assign data_masked[3464] = data_i[3464] & sel_one_hot_i[54];
  assign data_masked[3463] = data_i[3463] & sel_one_hot_i[54];
  assign data_masked[3462] = data_i[3462] & sel_one_hot_i[54];
  assign data_masked[3461] = data_i[3461] & sel_one_hot_i[54];
  assign data_masked[3460] = data_i[3460] & sel_one_hot_i[54];
  assign data_masked[3459] = data_i[3459] & sel_one_hot_i[54];
  assign data_masked[3458] = data_i[3458] & sel_one_hot_i[54];
  assign data_masked[3457] = data_i[3457] & sel_one_hot_i[54];
  assign data_masked[3456] = data_i[3456] & sel_one_hot_i[54];
  assign data_masked[3583] = data_i[3583] & sel_one_hot_i[55];
  assign data_masked[3582] = data_i[3582] & sel_one_hot_i[55];
  assign data_masked[3581] = data_i[3581] & sel_one_hot_i[55];
  assign data_masked[3580] = data_i[3580] & sel_one_hot_i[55];
  assign data_masked[3579] = data_i[3579] & sel_one_hot_i[55];
  assign data_masked[3578] = data_i[3578] & sel_one_hot_i[55];
  assign data_masked[3577] = data_i[3577] & sel_one_hot_i[55];
  assign data_masked[3576] = data_i[3576] & sel_one_hot_i[55];
  assign data_masked[3575] = data_i[3575] & sel_one_hot_i[55];
  assign data_masked[3574] = data_i[3574] & sel_one_hot_i[55];
  assign data_masked[3573] = data_i[3573] & sel_one_hot_i[55];
  assign data_masked[3572] = data_i[3572] & sel_one_hot_i[55];
  assign data_masked[3571] = data_i[3571] & sel_one_hot_i[55];
  assign data_masked[3570] = data_i[3570] & sel_one_hot_i[55];
  assign data_masked[3569] = data_i[3569] & sel_one_hot_i[55];
  assign data_masked[3568] = data_i[3568] & sel_one_hot_i[55];
  assign data_masked[3567] = data_i[3567] & sel_one_hot_i[55];
  assign data_masked[3566] = data_i[3566] & sel_one_hot_i[55];
  assign data_masked[3565] = data_i[3565] & sel_one_hot_i[55];
  assign data_masked[3564] = data_i[3564] & sel_one_hot_i[55];
  assign data_masked[3563] = data_i[3563] & sel_one_hot_i[55];
  assign data_masked[3562] = data_i[3562] & sel_one_hot_i[55];
  assign data_masked[3561] = data_i[3561] & sel_one_hot_i[55];
  assign data_masked[3560] = data_i[3560] & sel_one_hot_i[55];
  assign data_masked[3559] = data_i[3559] & sel_one_hot_i[55];
  assign data_masked[3558] = data_i[3558] & sel_one_hot_i[55];
  assign data_masked[3557] = data_i[3557] & sel_one_hot_i[55];
  assign data_masked[3556] = data_i[3556] & sel_one_hot_i[55];
  assign data_masked[3555] = data_i[3555] & sel_one_hot_i[55];
  assign data_masked[3554] = data_i[3554] & sel_one_hot_i[55];
  assign data_masked[3553] = data_i[3553] & sel_one_hot_i[55];
  assign data_masked[3552] = data_i[3552] & sel_one_hot_i[55];
  assign data_masked[3551] = data_i[3551] & sel_one_hot_i[55];
  assign data_masked[3550] = data_i[3550] & sel_one_hot_i[55];
  assign data_masked[3549] = data_i[3549] & sel_one_hot_i[55];
  assign data_masked[3548] = data_i[3548] & sel_one_hot_i[55];
  assign data_masked[3547] = data_i[3547] & sel_one_hot_i[55];
  assign data_masked[3546] = data_i[3546] & sel_one_hot_i[55];
  assign data_masked[3545] = data_i[3545] & sel_one_hot_i[55];
  assign data_masked[3544] = data_i[3544] & sel_one_hot_i[55];
  assign data_masked[3543] = data_i[3543] & sel_one_hot_i[55];
  assign data_masked[3542] = data_i[3542] & sel_one_hot_i[55];
  assign data_masked[3541] = data_i[3541] & sel_one_hot_i[55];
  assign data_masked[3540] = data_i[3540] & sel_one_hot_i[55];
  assign data_masked[3539] = data_i[3539] & sel_one_hot_i[55];
  assign data_masked[3538] = data_i[3538] & sel_one_hot_i[55];
  assign data_masked[3537] = data_i[3537] & sel_one_hot_i[55];
  assign data_masked[3536] = data_i[3536] & sel_one_hot_i[55];
  assign data_masked[3535] = data_i[3535] & sel_one_hot_i[55];
  assign data_masked[3534] = data_i[3534] & sel_one_hot_i[55];
  assign data_masked[3533] = data_i[3533] & sel_one_hot_i[55];
  assign data_masked[3532] = data_i[3532] & sel_one_hot_i[55];
  assign data_masked[3531] = data_i[3531] & sel_one_hot_i[55];
  assign data_masked[3530] = data_i[3530] & sel_one_hot_i[55];
  assign data_masked[3529] = data_i[3529] & sel_one_hot_i[55];
  assign data_masked[3528] = data_i[3528] & sel_one_hot_i[55];
  assign data_masked[3527] = data_i[3527] & sel_one_hot_i[55];
  assign data_masked[3526] = data_i[3526] & sel_one_hot_i[55];
  assign data_masked[3525] = data_i[3525] & sel_one_hot_i[55];
  assign data_masked[3524] = data_i[3524] & sel_one_hot_i[55];
  assign data_masked[3523] = data_i[3523] & sel_one_hot_i[55];
  assign data_masked[3522] = data_i[3522] & sel_one_hot_i[55];
  assign data_masked[3521] = data_i[3521] & sel_one_hot_i[55];
  assign data_masked[3520] = data_i[3520] & sel_one_hot_i[55];
  assign data_masked[3647] = data_i[3647] & sel_one_hot_i[56];
  assign data_masked[3646] = data_i[3646] & sel_one_hot_i[56];
  assign data_masked[3645] = data_i[3645] & sel_one_hot_i[56];
  assign data_masked[3644] = data_i[3644] & sel_one_hot_i[56];
  assign data_masked[3643] = data_i[3643] & sel_one_hot_i[56];
  assign data_masked[3642] = data_i[3642] & sel_one_hot_i[56];
  assign data_masked[3641] = data_i[3641] & sel_one_hot_i[56];
  assign data_masked[3640] = data_i[3640] & sel_one_hot_i[56];
  assign data_masked[3639] = data_i[3639] & sel_one_hot_i[56];
  assign data_masked[3638] = data_i[3638] & sel_one_hot_i[56];
  assign data_masked[3637] = data_i[3637] & sel_one_hot_i[56];
  assign data_masked[3636] = data_i[3636] & sel_one_hot_i[56];
  assign data_masked[3635] = data_i[3635] & sel_one_hot_i[56];
  assign data_masked[3634] = data_i[3634] & sel_one_hot_i[56];
  assign data_masked[3633] = data_i[3633] & sel_one_hot_i[56];
  assign data_masked[3632] = data_i[3632] & sel_one_hot_i[56];
  assign data_masked[3631] = data_i[3631] & sel_one_hot_i[56];
  assign data_masked[3630] = data_i[3630] & sel_one_hot_i[56];
  assign data_masked[3629] = data_i[3629] & sel_one_hot_i[56];
  assign data_masked[3628] = data_i[3628] & sel_one_hot_i[56];
  assign data_masked[3627] = data_i[3627] & sel_one_hot_i[56];
  assign data_masked[3626] = data_i[3626] & sel_one_hot_i[56];
  assign data_masked[3625] = data_i[3625] & sel_one_hot_i[56];
  assign data_masked[3624] = data_i[3624] & sel_one_hot_i[56];
  assign data_masked[3623] = data_i[3623] & sel_one_hot_i[56];
  assign data_masked[3622] = data_i[3622] & sel_one_hot_i[56];
  assign data_masked[3621] = data_i[3621] & sel_one_hot_i[56];
  assign data_masked[3620] = data_i[3620] & sel_one_hot_i[56];
  assign data_masked[3619] = data_i[3619] & sel_one_hot_i[56];
  assign data_masked[3618] = data_i[3618] & sel_one_hot_i[56];
  assign data_masked[3617] = data_i[3617] & sel_one_hot_i[56];
  assign data_masked[3616] = data_i[3616] & sel_one_hot_i[56];
  assign data_masked[3615] = data_i[3615] & sel_one_hot_i[56];
  assign data_masked[3614] = data_i[3614] & sel_one_hot_i[56];
  assign data_masked[3613] = data_i[3613] & sel_one_hot_i[56];
  assign data_masked[3612] = data_i[3612] & sel_one_hot_i[56];
  assign data_masked[3611] = data_i[3611] & sel_one_hot_i[56];
  assign data_masked[3610] = data_i[3610] & sel_one_hot_i[56];
  assign data_masked[3609] = data_i[3609] & sel_one_hot_i[56];
  assign data_masked[3608] = data_i[3608] & sel_one_hot_i[56];
  assign data_masked[3607] = data_i[3607] & sel_one_hot_i[56];
  assign data_masked[3606] = data_i[3606] & sel_one_hot_i[56];
  assign data_masked[3605] = data_i[3605] & sel_one_hot_i[56];
  assign data_masked[3604] = data_i[3604] & sel_one_hot_i[56];
  assign data_masked[3603] = data_i[3603] & sel_one_hot_i[56];
  assign data_masked[3602] = data_i[3602] & sel_one_hot_i[56];
  assign data_masked[3601] = data_i[3601] & sel_one_hot_i[56];
  assign data_masked[3600] = data_i[3600] & sel_one_hot_i[56];
  assign data_masked[3599] = data_i[3599] & sel_one_hot_i[56];
  assign data_masked[3598] = data_i[3598] & sel_one_hot_i[56];
  assign data_masked[3597] = data_i[3597] & sel_one_hot_i[56];
  assign data_masked[3596] = data_i[3596] & sel_one_hot_i[56];
  assign data_masked[3595] = data_i[3595] & sel_one_hot_i[56];
  assign data_masked[3594] = data_i[3594] & sel_one_hot_i[56];
  assign data_masked[3593] = data_i[3593] & sel_one_hot_i[56];
  assign data_masked[3592] = data_i[3592] & sel_one_hot_i[56];
  assign data_masked[3591] = data_i[3591] & sel_one_hot_i[56];
  assign data_masked[3590] = data_i[3590] & sel_one_hot_i[56];
  assign data_masked[3589] = data_i[3589] & sel_one_hot_i[56];
  assign data_masked[3588] = data_i[3588] & sel_one_hot_i[56];
  assign data_masked[3587] = data_i[3587] & sel_one_hot_i[56];
  assign data_masked[3586] = data_i[3586] & sel_one_hot_i[56];
  assign data_masked[3585] = data_i[3585] & sel_one_hot_i[56];
  assign data_masked[3584] = data_i[3584] & sel_one_hot_i[56];
  assign data_masked[3711] = data_i[3711] & sel_one_hot_i[57];
  assign data_masked[3710] = data_i[3710] & sel_one_hot_i[57];
  assign data_masked[3709] = data_i[3709] & sel_one_hot_i[57];
  assign data_masked[3708] = data_i[3708] & sel_one_hot_i[57];
  assign data_masked[3707] = data_i[3707] & sel_one_hot_i[57];
  assign data_masked[3706] = data_i[3706] & sel_one_hot_i[57];
  assign data_masked[3705] = data_i[3705] & sel_one_hot_i[57];
  assign data_masked[3704] = data_i[3704] & sel_one_hot_i[57];
  assign data_masked[3703] = data_i[3703] & sel_one_hot_i[57];
  assign data_masked[3702] = data_i[3702] & sel_one_hot_i[57];
  assign data_masked[3701] = data_i[3701] & sel_one_hot_i[57];
  assign data_masked[3700] = data_i[3700] & sel_one_hot_i[57];
  assign data_masked[3699] = data_i[3699] & sel_one_hot_i[57];
  assign data_masked[3698] = data_i[3698] & sel_one_hot_i[57];
  assign data_masked[3697] = data_i[3697] & sel_one_hot_i[57];
  assign data_masked[3696] = data_i[3696] & sel_one_hot_i[57];
  assign data_masked[3695] = data_i[3695] & sel_one_hot_i[57];
  assign data_masked[3694] = data_i[3694] & sel_one_hot_i[57];
  assign data_masked[3693] = data_i[3693] & sel_one_hot_i[57];
  assign data_masked[3692] = data_i[3692] & sel_one_hot_i[57];
  assign data_masked[3691] = data_i[3691] & sel_one_hot_i[57];
  assign data_masked[3690] = data_i[3690] & sel_one_hot_i[57];
  assign data_masked[3689] = data_i[3689] & sel_one_hot_i[57];
  assign data_masked[3688] = data_i[3688] & sel_one_hot_i[57];
  assign data_masked[3687] = data_i[3687] & sel_one_hot_i[57];
  assign data_masked[3686] = data_i[3686] & sel_one_hot_i[57];
  assign data_masked[3685] = data_i[3685] & sel_one_hot_i[57];
  assign data_masked[3684] = data_i[3684] & sel_one_hot_i[57];
  assign data_masked[3683] = data_i[3683] & sel_one_hot_i[57];
  assign data_masked[3682] = data_i[3682] & sel_one_hot_i[57];
  assign data_masked[3681] = data_i[3681] & sel_one_hot_i[57];
  assign data_masked[3680] = data_i[3680] & sel_one_hot_i[57];
  assign data_masked[3679] = data_i[3679] & sel_one_hot_i[57];
  assign data_masked[3678] = data_i[3678] & sel_one_hot_i[57];
  assign data_masked[3677] = data_i[3677] & sel_one_hot_i[57];
  assign data_masked[3676] = data_i[3676] & sel_one_hot_i[57];
  assign data_masked[3675] = data_i[3675] & sel_one_hot_i[57];
  assign data_masked[3674] = data_i[3674] & sel_one_hot_i[57];
  assign data_masked[3673] = data_i[3673] & sel_one_hot_i[57];
  assign data_masked[3672] = data_i[3672] & sel_one_hot_i[57];
  assign data_masked[3671] = data_i[3671] & sel_one_hot_i[57];
  assign data_masked[3670] = data_i[3670] & sel_one_hot_i[57];
  assign data_masked[3669] = data_i[3669] & sel_one_hot_i[57];
  assign data_masked[3668] = data_i[3668] & sel_one_hot_i[57];
  assign data_masked[3667] = data_i[3667] & sel_one_hot_i[57];
  assign data_masked[3666] = data_i[3666] & sel_one_hot_i[57];
  assign data_masked[3665] = data_i[3665] & sel_one_hot_i[57];
  assign data_masked[3664] = data_i[3664] & sel_one_hot_i[57];
  assign data_masked[3663] = data_i[3663] & sel_one_hot_i[57];
  assign data_masked[3662] = data_i[3662] & sel_one_hot_i[57];
  assign data_masked[3661] = data_i[3661] & sel_one_hot_i[57];
  assign data_masked[3660] = data_i[3660] & sel_one_hot_i[57];
  assign data_masked[3659] = data_i[3659] & sel_one_hot_i[57];
  assign data_masked[3658] = data_i[3658] & sel_one_hot_i[57];
  assign data_masked[3657] = data_i[3657] & sel_one_hot_i[57];
  assign data_masked[3656] = data_i[3656] & sel_one_hot_i[57];
  assign data_masked[3655] = data_i[3655] & sel_one_hot_i[57];
  assign data_masked[3654] = data_i[3654] & sel_one_hot_i[57];
  assign data_masked[3653] = data_i[3653] & sel_one_hot_i[57];
  assign data_masked[3652] = data_i[3652] & sel_one_hot_i[57];
  assign data_masked[3651] = data_i[3651] & sel_one_hot_i[57];
  assign data_masked[3650] = data_i[3650] & sel_one_hot_i[57];
  assign data_masked[3649] = data_i[3649] & sel_one_hot_i[57];
  assign data_masked[3648] = data_i[3648] & sel_one_hot_i[57];
  assign data_masked[3775] = data_i[3775] & sel_one_hot_i[58];
  assign data_masked[3774] = data_i[3774] & sel_one_hot_i[58];
  assign data_masked[3773] = data_i[3773] & sel_one_hot_i[58];
  assign data_masked[3772] = data_i[3772] & sel_one_hot_i[58];
  assign data_masked[3771] = data_i[3771] & sel_one_hot_i[58];
  assign data_masked[3770] = data_i[3770] & sel_one_hot_i[58];
  assign data_masked[3769] = data_i[3769] & sel_one_hot_i[58];
  assign data_masked[3768] = data_i[3768] & sel_one_hot_i[58];
  assign data_masked[3767] = data_i[3767] & sel_one_hot_i[58];
  assign data_masked[3766] = data_i[3766] & sel_one_hot_i[58];
  assign data_masked[3765] = data_i[3765] & sel_one_hot_i[58];
  assign data_masked[3764] = data_i[3764] & sel_one_hot_i[58];
  assign data_masked[3763] = data_i[3763] & sel_one_hot_i[58];
  assign data_masked[3762] = data_i[3762] & sel_one_hot_i[58];
  assign data_masked[3761] = data_i[3761] & sel_one_hot_i[58];
  assign data_masked[3760] = data_i[3760] & sel_one_hot_i[58];
  assign data_masked[3759] = data_i[3759] & sel_one_hot_i[58];
  assign data_masked[3758] = data_i[3758] & sel_one_hot_i[58];
  assign data_masked[3757] = data_i[3757] & sel_one_hot_i[58];
  assign data_masked[3756] = data_i[3756] & sel_one_hot_i[58];
  assign data_masked[3755] = data_i[3755] & sel_one_hot_i[58];
  assign data_masked[3754] = data_i[3754] & sel_one_hot_i[58];
  assign data_masked[3753] = data_i[3753] & sel_one_hot_i[58];
  assign data_masked[3752] = data_i[3752] & sel_one_hot_i[58];
  assign data_masked[3751] = data_i[3751] & sel_one_hot_i[58];
  assign data_masked[3750] = data_i[3750] & sel_one_hot_i[58];
  assign data_masked[3749] = data_i[3749] & sel_one_hot_i[58];
  assign data_masked[3748] = data_i[3748] & sel_one_hot_i[58];
  assign data_masked[3747] = data_i[3747] & sel_one_hot_i[58];
  assign data_masked[3746] = data_i[3746] & sel_one_hot_i[58];
  assign data_masked[3745] = data_i[3745] & sel_one_hot_i[58];
  assign data_masked[3744] = data_i[3744] & sel_one_hot_i[58];
  assign data_masked[3743] = data_i[3743] & sel_one_hot_i[58];
  assign data_masked[3742] = data_i[3742] & sel_one_hot_i[58];
  assign data_masked[3741] = data_i[3741] & sel_one_hot_i[58];
  assign data_masked[3740] = data_i[3740] & sel_one_hot_i[58];
  assign data_masked[3739] = data_i[3739] & sel_one_hot_i[58];
  assign data_masked[3738] = data_i[3738] & sel_one_hot_i[58];
  assign data_masked[3737] = data_i[3737] & sel_one_hot_i[58];
  assign data_masked[3736] = data_i[3736] & sel_one_hot_i[58];
  assign data_masked[3735] = data_i[3735] & sel_one_hot_i[58];
  assign data_masked[3734] = data_i[3734] & sel_one_hot_i[58];
  assign data_masked[3733] = data_i[3733] & sel_one_hot_i[58];
  assign data_masked[3732] = data_i[3732] & sel_one_hot_i[58];
  assign data_masked[3731] = data_i[3731] & sel_one_hot_i[58];
  assign data_masked[3730] = data_i[3730] & sel_one_hot_i[58];
  assign data_masked[3729] = data_i[3729] & sel_one_hot_i[58];
  assign data_masked[3728] = data_i[3728] & sel_one_hot_i[58];
  assign data_masked[3727] = data_i[3727] & sel_one_hot_i[58];
  assign data_masked[3726] = data_i[3726] & sel_one_hot_i[58];
  assign data_masked[3725] = data_i[3725] & sel_one_hot_i[58];
  assign data_masked[3724] = data_i[3724] & sel_one_hot_i[58];
  assign data_masked[3723] = data_i[3723] & sel_one_hot_i[58];
  assign data_masked[3722] = data_i[3722] & sel_one_hot_i[58];
  assign data_masked[3721] = data_i[3721] & sel_one_hot_i[58];
  assign data_masked[3720] = data_i[3720] & sel_one_hot_i[58];
  assign data_masked[3719] = data_i[3719] & sel_one_hot_i[58];
  assign data_masked[3718] = data_i[3718] & sel_one_hot_i[58];
  assign data_masked[3717] = data_i[3717] & sel_one_hot_i[58];
  assign data_masked[3716] = data_i[3716] & sel_one_hot_i[58];
  assign data_masked[3715] = data_i[3715] & sel_one_hot_i[58];
  assign data_masked[3714] = data_i[3714] & sel_one_hot_i[58];
  assign data_masked[3713] = data_i[3713] & sel_one_hot_i[58];
  assign data_masked[3712] = data_i[3712] & sel_one_hot_i[58];
  assign data_masked[3839] = data_i[3839] & sel_one_hot_i[59];
  assign data_masked[3838] = data_i[3838] & sel_one_hot_i[59];
  assign data_masked[3837] = data_i[3837] & sel_one_hot_i[59];
  assign data_masked[3836] = data_i[3836] & sel_one_hot_i[59];
  assign data_masked[3835] = data_i[3835] & sel_one_hot_i[59];
  assign data_masked[3834] = data_i[3834] & sel_one_hot_i[59];
  assign data_masked[3833] = data_i[3833] & sel_one_hot_i[59];
  assign data_masked[3832] = data_i[3832] & sel_one_hot_i[59];
  assign data_masked[3831] = data_i[3831] & sel_one_hot_i[59];
  assign data_masked[3830] = data_i[3830] & sel_one_hot_i[59];
  assign data_masked[3829] = data_i[3829] & sel_one_hot_i[59];
  assign data_masked[3828] = data_i[3828] & sel_one_hot_i[59];
  assign data_masked[3827] = data_i[3827] & sel_one_hot_i[59];
  assign data_masked[3826] = data_i[3826] & sel_one_hot_i[59];
  assign data_masked[3825] = data_i[3825] & sel_one_hot_i[59];
  assign data_masked[3824] = data_i[3824] & sel_one_hot_i[59];
  assign data_masked[3823] = data_i[3823] & sel_one_hot_i[59];
  assign data_masked[3822] = data_i[3822] & sel_one_hot_i[59];
  assign data_masked[3821] = data_i[3821] & sel_one_hot_i[59];
  assign data_masked[3820] = data_i[3820] & sel_one_hot_i[59];
  assign data_masked[3819] = data_i[3819] & sel_one_hot_i[59];
  assign data_masked[3818] = data_i[3818] & sel_one_hot_i[59];
  assign data_masked[3817] = data_i[3817] & sel_one_hot_i[59];
  assign data_masked[3816] = data_i[3816] & sel_one_hot_i[59];
  assign data_masked[3815] = data_i[3815] & sel_one_hot_i[59];
  assign data_masked[3814] = data_i[3814] & sel_one_hot_i[59];
  assign data_masked[3813] = data_i[3813] & sel_one_hot_i[59];
  assign data_masked[3812] = data_i[3812] & sel_one_hot_i[59];
  assign data_masked[3811] = data_i[3811] & sel_one_hot_i[59];
  assign data_masked[3810] = data_i[3810] & sel_one_hot_i[59];
  assign data_masked[3809] = data_i[3809] & sel_one_hot_i[59];
  assign data_masked[3808] = data_i[3808] & sel_one_hot_i[59];
  assign data_masked[3807] = data_i[3807] & sel_one_hot_i[59];
  assign data_masked[3806] = data_i[3806] & sel_one_hot_i[59];
  assign data_masked[3805] = data_i[3805] & sel_one_hot_i[59];
  assign data_masked[3804] = data_i[3804] & sel_one_hot_i[59];
  assign data_masked[3803] = data_i[3803] & sel_one_hot_i[59];
  assign data_masked[3802] = data_i[3802] & sel_one_hot_i[59];
  assign data_masked[3801] = data_i[3801] & sel_one_hot_i[59];
  assign data_masked[3800] = data_i[3800] & sel_one_hot_i[59];
  assign data_masked[3799] = data_i[3799] & sel_one_hot_i[59];
  assign data_masked[3798] = data_i[3798] & sel_one_hot_i[59];
  assign data_masked[3797] = data_i[3797] & sel_one_hot_i[59];
  assign data_masked[3796] = data_i[3796] & sel_one_hot_i[59];
  assign data_masked[3795] = data_i[3795] & sel_one_hot_i[59];
  assign data_masked[3794] = data_i[3794] & sel_one_hot_i[59];
  assign data_masked[3793] = data_i[3793] & sel_one_hot_i[59];
  assign data_masked[3792] = data_i[3792] & sel_one_hot_i[59];
  assign data_masked[3791] = data_i[3791] & sel_one_hot_i[59];
  assign data_masked[3790] = data_i[3790] & sel_one_hot_i[59];
  assign data_masked[3789] = data_i[3789] & sel_one_hot_i[59];
  assign data_masked[3788] = data_i[3788] & sel_one_hot_i[59];
  assign data_masked[3787] = data_i[3787] & sel_one_hot_i[59];
  assign data_masked[3786] = data_i[3786] & sel_one_hot_i[59];
  assign data_masked[3785] = data_i[3785] & sel_one_hot_i[59];
  assign data_masked[3784] = data_i[3784] & sel_one_hot_i[59];
  assign data_masked[3783] = data_i[3783] & sel_one_hot_i[59];
  assign data_masked[3782] = data_i[3782] & sel_one_hot_i[59];
  assign data_masked[3781] = data_i[3781] & sel_one_hot_i[59];
  assign data_masked[3780] = data_i[3780] & sel_one_hot_i[59];
  assign data_masked[3779] = data_i[3779] & sel_one_hot_i[59];
  assign data_masked[3778] = data_i[3778] & sel_one_hot_i[59];
  assign data_masked[3777] = data_i[3777] & sel_one_hot_i[59];
  assign data_masked[3776] = data_i[3776] & sel_one_hot_i[59];
  assign data_masked[3903] = data_i[3903] & sel_one_hot_i[60];
  assign data_masked[3902] = data_i[3902] & sel_one_hot_i[60];
  assign data_masked[3901] = data_i[3901] & sel_one_hot_i[60];
  assign data_masked[3900] = data_i[3900] & sel_one_hot_i[60];
  assign data_masked[3899] = data_i[3899] & sel_one_hot_i[60];
  assign data_masked[3898] = data_i[3898] & sel_one_hot_i[60];
  assign data_masked[3897] = data_i[3897] & sel_one_hot_i[60];
  assign data_masked[3896] = data_i[3896] & sel_one_hot_i[60];
  assign data_masked[3895] = data_i[3895] & sel_one_hot_i[60];
  assign data_masked[3894] = data_i[3894] & sel_one_hot_i[60];
  assign data_masked[3893] = data_i[3893] & sel_one_hot_i[60];
  assign data_masked[3892] = data_i[3892] & sel_one_hot_i[60];
  assign data_masked[3891] = data_i[3891] & sel_one_hot_i[60];
  assign data_masked[3890] = data_i[3890] & sel_one_hot_i[60];
  assign data_masked[3889] = data_i[3889] & sel_one_hot_i[60];
  assign data_masked[3888] = data_i[3888] & sel_one_hot_i[60];
  assign data_masked[3887] = data_i[3887] & sel_one_hot_i[60];
  assign data_masked[3886] = data_i[3886] & sel_one_hot_i[60];
  assign data_masked[3885] = data_i[3885] & sel_one_hot_i[60];
  assign data_masked[3884] = data_i[3884] & sel_one_hot_i[60];
  assign data_masked[3883] = data_i[3883] & sel_one_hot_i[60];
  assign data_masked[3882] = data_i[3882] & sel_one_hot_i[60];
  assign data_masked[3881] = data_i[3881] & sel_one_hot_i[60];
  assign data_masked[3880] = data_i[3880] & sel_one_hot_i[60];
  assign data_masked[3879] = data_i[3879] & sel_one_hot_i[60];
  assign data_masked[3878] = data_i[3878] & sel_one_hot_i[60];
  assign data_masked[3877] = data_i[3877] & sel_one_hot_i[60];
  assign data_masked[3876] = data_i[3876] & sel_one_hot_i[60];
  assign data_masked[3875] = data_i[3875] & sel_one_hot_i[60];
  assign data_masked[3874] = data_i[3874] & sel_one_hot_i[60];
  assign data_masked[3873] = data_i[3873] & sel_one_hot_i[60];
  assign data_masked[3872] = data_i[3872] & sel_one_hot_i[60];
  assign data_masked[3871] = data_i[3871] & sel_one_hot_i[60];
  assign data_masked[3870] = data_i[3870] & sel_one_hot_i[60];
  assign data_masked[3869] = data_i[3869] & sel_one_hot_i[60];
  assign data_masked[3868] = data_i[3868] & sel_one_hot_i[60];
  assign data_masked[3867] = data_i[3867] & sel_one_hot_i[60];
  assign data_masked[3866] = data_i[3866] & sel_one_hot_i[60];
  assign data_masked[3865] = data_i[3865] & sel_one_hot_i[60];
  assign data_masked[3864] = data_i[3864] & sel_one_hot_i[60];
  assign data_masked[3863] = data_i[3863] & sel_one_hot_i[60];
  assign data_masked[3862] = data_i[3862] & sel_one_hot_i[60];
  assign data_masked[3861] = data_i[3861] & sel_one_hot_i[60];
  assign data_masked[3860] = data_i[3860] & sel_one_hot_i[60];
  assign data_masked[3859] = data_i[3859] & sel_one_hot_i[60];
  assign data_masked[3858] = data_i[3858] & sel_one_hot_i[60];
  assign data_masked[3857] = data_i[3857] & sel_one_hot_i[60];
  assign data_masked[3856] = data_i[3856] & sel_one_hot_i[60];
  assign data_masked[3855] = data_i[3855] & sel_one_hot_i[60];
  assign data_masked[3854] = data_i[3854] & sel_one_hot_i[60];
  assign data_masked[3853] = data_i[3853] & sel_one_hot_i[60];
  assign data_masked[3852] = data_i[3852] & sel_one_hot_i[60];
  assign data_masked[3851] = data_i[3851] & sel_one_hot_i[60];
  assign data_masked[3850] = data_i[3850] & sel_one_hot_i[60];
  assign data_masked[3849] = data_i[3849] & sel_one_hot_i[60];
  assign data_masked[3848] = data_i[3848] & sel_one_hot_i[60];
  assign data_masked[3847] = data_i[3847] & sel_one_hot_i[60];
  assign data_masked[3846] = data_i[3846] & sel_one_hot_i[60];
  assign data_masked[3845] = data_i[3845] & sel_one_hot_i[60];
  assign data_masked[3844] = data_i[3844] & sel_one_hot_i[60];
  assign data_masked[3843] = data_i[3843] & sel_one_hot_i[60];
  assign data_masked[3842] = data_i[3842] & sel_one_hot_i[60];
  assign data_masked[3841] = data_i[3841] & sel_one_hot_i[60];
  assign data_masked[3840] = data_i[3840] & sel_one_hot_i[60];
  assign data_masked[3967] = data_i[3967] & sel_one_hot_i[61];
  assign data_masked[3966] = data_i[3966] & sel_one_hot_i[61];
  assign data_masked[3965] = data_i[3965] & sel_one_hot_i[61];
  assign data_masked[3964] = data_i[3964] & sel_one_hot_i[61];
  assign data_masked[3963] = data_i[3963] & sel_one_hot_i[61];
  assign data_masked[3962] = data_i[3962] & sel_one_hot_i[61];
  assign data_masked[3961] = data_i[3961] & sel_one_hot_i[61];
  assign data_masked[3960] = data_i[3960] & sel_one_hot_i[61];
  assign data_masked[3959] = data_i[3959] & sel_one_hot_i[61];
  assign data_masked[3958] = data_i[3958] & sel_one_hot_i[61];
  assign data_masked[3957] = data_i[3957] & sel_one_hot_i[61];
  assign data_masked[3956] = data_i[3956] & sel_one_hot_i[61];
  assign data_masked[3955] = data_i[3955] & sel_one_hot_i[61];
  assign data_masked[3954] = data_i[3954] & sel_one_hot_i[61];
  assign data_masked[3953] = data_i[3953] & sel_one_hot_i[61];
  assign data_masked[3952] = data_i[3952] & sel_one_hot_i[61];
  assign data_masked[3951] = data_i[3951] & sel_one_hot_i[61];
  assign data_masked[3950] = data_i[3950] & sel_one_hot_i[61];
  assign data_masked[3949] = data_i[3949] & sel_one_hot_i[61];
  assign data_masked[3948] = data_i[3948] & sel_one_hot_i[61];
  assign data_masked[3947] = data_i[3947] & sel_one_hot_i[61];
  assign data_masked[3946] = data_i[3946] & sel_one_hot_i[61];
  assign data_masked[3945] = data_i[3945] & sel_one_hot_i[61];
  assign data_masked[3944] = data_i[3944] & sel_one_hot_i[61];
  assign data_masked[3943] = data_i[3943] & sel_one_hot_i[61];
  assign data_masked[3942] = data_i[3942] & sel_one_hot_i[61];
  assign data_masked[3941] = data_i[3941] & sel_one_hot_i[61];
  assign data_masked[3940] = data_i[3940] & sel_one_hot_i[61];
  assign data_masked[3939] = data_i[3939] & sel_one_hot_i[61];
  assign data_masked[3938] = data_i[3938] & sel_one_hot_i[61];
  assign data_masked[3937] = data_i[3937] & sel_one_hot_i[61];
  assign data_masked[3936] = data_i[3936] & sel_one_hot_i[61];
  assign data_masked[3935] = data_i[3935] & sel_one_hot_i[61];
  assign data_masked[3934] = data_i[3934] & sel_one_hot_i[61];
  assign data_masked[3933] = data_i[3933] & sel_one_hot_i[61];
  assign data_masked[3932] = data_i[3932] & sel_one_hot_i[61];
  assign data_masked[3931] = data_i[3931] & sel_one_hot_i[61];
  assign data_masked[3930] = data_i[3930] & sel_one_hot_i[61];
  assign data_masked[3929] = data_i[3929] & sel_one_hot_i[61];
  assign data_masked[3928] = data_i[3928] & sel_one_hot_i[61];
  assign data_masked[3927] = data_i[3927] & sel_one_hot_i[61];
  assign data_masked[3926] = data_i[3926] & sel_one_hot_i[61];
  assign data_masked[3925] = data_i[3925] & sel_one_hot_i[61];
  assign data_masked[3924] = data_i[3924] & sel_one_hot_i[61];
  assign data_masked[3923] = data_i[3923] & sel_one_hot_i[61];
  assign data_masked[3922] = data_i[3922] & sel_one_hot_i[61];
  assign data_masked[3921] = data_i[3921] & sel_one_hot_i[61];
  assign data_masked[3920] = data_i[3920] & sel_one_hot_i[61];
  assign data_masked[3919] = data_i[3919] & sel_one_hot_i[61];
  assign data_masked[3918] = data_i[3918] & sel_one_hot_i[61];
  assign data_masked[3917] = data_i[3917] & sel_one_hot_i[61];
  assign data_masked[3916] = data_i[3916] & sel_one_hot_i[61];
  assign data_masked[3915] = data_i[3915] & sel_one_hot_i[61];
  assign data_masked[3914] = data_i[3914] & sel_one_hot_i[61];
  assign data_masked[3913] = data_i[3913] & sel_one_hot_i[61];
  assign data_masked[3912] = data_i[3912] & sel_one_hot_i[61];
  assign data_masked[3911] = data_i[3911] & sel_one_hot_i[61];
  assign data_masked[3910] = data_i[3910] & sel_one_hot_i[61];
  assign data_masked[3909] = data_i[3909] & sel_one_hot_i[61];
  assign data_masked[3908] = data_i[3908] & sel_one_hot_i[61];
  assign data_masked[3907] = data_i[3907] & sel_one_hot_i[61];
  assign data_masked[3906] = data_i[3906] & sel_one_hot_i[61];
  assign data_masked[3905] = data_i[3905] & sel_one_hot_i[61];
  assign data_masked[3904] = data_i[3904] & sel_one_hot_i[61];
  assign data_masked[4031] = data_i[4031] & sel_one_hot_i[62];
  assign data_masked[4030] = data_i[4030] & sel_one_hot_i[62];
  assign data_masked[4029] = data_i[4029] & sel_one_hot_i[62];
  assign data_masked[4028] = data_i[4028] & sel_one_hot_i[62];
  assign data_masked[4027] = data_i[4027] & sel_one_hot_i[62];
  assign data_masked[4026] = data_i[4026] & sel_one_hot_i[62];
  assign data_masked[4025] = data_i[4025] & sel_one_hot_i[62];
  assign data_masked[4024] = data_i[4024] & sel_one_hot_i[62];
  assign data_masked[4023] = data_i[4023] & sel_one_hot_i[62];
  assign data_masked[4022] = data_i[4022] & sel_one_hot_i[62];
  assign data_masked[4021] = data_i[4021] & sel_one_hot_i[62];
  assign data_masked[4020] = data_i[4020] & sel_one_hot_i[62];
  assign data_masked[4019] = data_i[4019] & sel_one_hot_i[62];
  assign data_masked[4018] = data_i[4018] & sel_one_hot_i[62];
  assign data_masked[4017] = data_i[4017] & sel_one_hot_i[62];
  assign data_masked[4016] = data_i[4016] & sel_one_hot_i[62];
  assign data_masked[4015] = data_i[4015] & sel_one_hot_i[62];
  assign data_masked[4014] = data_i[4014] & sel_one_hot_i[62];
  assign data_masked[4013] = data_i[4013] & sel_one_hot_i[62];
  assign data_masked[4012] = data_i[4012] & sel_one_hot_i[62];
  assign data_masked[4011] = data_i[4011] & sel_one_hot_i[62];
  assign data_masked[4010] = data_i[4010] & sel_one_hot_i[62];
  assign data_masked[4009] = data_i[4009] & sel_one_hot_i[62];
  assign data_masked[4008] = data_i[4008] & sel_one_hot_i[62];
  assign data_masked[4007] = data_i[4007] & sel_one_hot_i[62];
  assign data_masked[4006] = data_i[4006] & sel_one_hot_i[62];
  assign data_masked[4005] = data_i[4005] & sel_one_hot_i[62];
  assign data_masked[4004] = data_i[4004] & sel_one_hot_i[62];
  assign data_masked[4003] = data_i[4003] & sel_one_hot_i[62];
  assign data_masked[4002] = data_i[4002] & sel_one_hot_i[62];
  assign data_masked[4001] = data_i[4001] & sel_one_hot_i[62];
  assign data_masked[4000] = data_i[4000] & sel_one_hot_i[62];
  assign data_masked[3999] = data_i[3999] & sel_one_hot_i[62];
  assign data_masked[3998] = data_i[3998] & sel_one_hot_i[62];
  assign data_masked[3997] = data_i[3997] & sel_one_hot_i[62];
  assign data_masked[3996] = data_i[3996] & sel_one_hot_i[62];
  assign data_masked[3995] = data_i[3995] & sel_one_hot_i[62];
  assign data_masked[3994] = data_i[3994] & sel_one_hot_i[62];
  assign data_masked[3993] = data_i[3993] & sel_one_hot_i[62];
  assign data_masked[3992] = data_i[3992] & sel_one_hot_i[62];
  assign data_masked[3991] = data_i[3991] & sel_one_hot_i[62];
  assign data_masked[3990] = data_i[3990] & sel_one_hot_i[62];
  assign data_masked[3989] = data_i[3989] & sel_one_hot_i[62];
  assign data_masked[3988] = data_i[3988] & sel_one_hot_i[62];
  assign data_masked[3987] = data_i[3987] & sel_one_hot_i[62];
  assign data_masked[3986] = data_i[3986] & sel_one_hot_i[62];
  assign data_masked[3985] = data_i[3985] & sel_one_hot_i[62];
  assign data_masked[3984] = data_i[3984] & sel_one_hot_i[62];
  assign data_masked[3983] = data_i[3983] & sel_one_hot_i[62];
  assign data_masked[3982] = data_i[3982] & sel_one_hot_i[62];
  assign data_masked[3981] = data_i[3981] & sel_one_hot_i[62];
  assign data_masked[3980] = data_i[3980] & sel_one_hot_i[62];
  assign data_masked[3979] = data_i[3979] & sel_one_hot_i[62];
  assign data_masked[3978] = data_i[3978] & sel_one_hot_i[62];
  assign data_masked[3977] = data_i[3977] & sel_one_hot_i[62];
  assign data_masked[3976] = data_i[3976] & sel_one_hot_i[62];
  assign data_masked[3975] = data_i[3975] & sel_one_hot_i[62];
  assign data_masked[3974] = data_i[3974] & sel_one_hot_i[62];
  assign data_masked[3973] = data_i[3973] & sel_one_hot_i[62];
  assign data_masked[3972] = data_i[3972] & sel_one_hot_i[62];
  assign data_masked[3971] = data_i[3971] & sel_one_hot_i[62];
  assign data_masked[3970] = data_i[3970] & sel_one_hot_i[62];
  assign data_masked[3969] = data_i[3969] & sel_one_hot_i[62];
  assign data_masked[3968] = data_i[3968] & sel_one_hot_i[62];
  assign data_masked[4095] = data_i[4095] & sel_one_hot_i[63];
  assign data_masked[4094] = data_i[4094] & sel_one_hot_i[63];
  assign data_masked[4093] = data_i[4093] & sel_one_hot_i[63];
  assign data_masked[4092] = data_i[4092] & sel_one_hot_i[63];
  assign data_masked[4091] = data_i[4091] & sel_one_hot_i[63];
  assign data_masked[4090] = data_i[4090] & sel_one_hot_i[63];
  assign data_masked[4089] = data_i[4089] & sel_one_hot_i[63];
  assign data_masked[4088] = data_i[4088] & sel_one_hot_i[63];
  assign data_masked[4087] = data_i[4087] & sel_one_hot_i[63];
  assign data_masked[4086] = data_i[4086] & sel_one_hot_i[63];
  assign data_masked[4085] = data_i[4085] & sel_one_hot_i[63];
  assign data_masked[4084] = data_i[4084] & sel_one_hot_i[63];
  assign data_masked[4083] = data_i[4083] & sel_one_hot_i[63];
  assign data_masked[4082] = data_i[4082] & sel_one_hot_i[63];
  assign data_masked[4081] = data_i[4081] & sel_one_hot_i[63];
  assign data_masked[4080] = data_i[4080] & sel_one_hot_i[63];
  assign data_masked[4079] = data_i[4079] & sel_one_hot_i[63];
  assign data_masked[4078] = data_i[4078] & sel_one_hot_i[63];
  assign data_masked[4077] = data_i[4077] & sel_one_hot_i[63];
  assign data_masked[4076] = data_i[4076] & sel_one_hot_i[63];
  assign data_masked[4075] = data_i[4075] & sel_one_hot_i[63];
  assign data_masked[4074] = data_i[4074] & sel_one_hot_i[63];
  assign data_masked[4073] = data_i[4073] & sel_one_hot_i[63];
  assign data_masked[4072] = data_i[4072] & sel_one_hot_i[63];
  assign data_masked[4071] = data_i[4071] & sel_one_hot_i[63];
  assign data_masked[4070] = data_i[4070] & sel_one_hot_i[63];
  assign data_masked[4069] = data_i[4069] & sel_one_hot_i[63];
  assign data_masked[4068] = data_i[4068] & sel_one_hot_i[63];
  assign data_masked[4067] = data_i[4067] & sel_one_hot_i[63];
  assign data_masked[4066] = data_i[4066] & sel_one_hot_i[63];
  assign data_masked[4065] = data_i[4065] & sel_one_hot_i[63];
  assign data_masked[4064] = data_i[4064] & sel_one_hot_i[63];
  assign data_masked[4063] = data_i[4063] & sel_one_hot_i[63];
  assign data_masked[4062] = data_i[4062] & sel_one_hot_i[63];
  assign data_masked[4061] = data_i[4061] & sel_one_hot_i[63];
  assign data_masked[4060] = data_i[4060] & sel_one_hot_i[63];
  assign data_masked[4059] = data_i[4059] & sel_one_hot_i[63];
  assign data_masked[4058] = data_i[4058] & sel_one_hot_i[63];
  assign data_masked[4057] = data_i[4057] & sel_one_hot_i[63];
  assign data_masked[4056] = data_i[4056] & sel_one_hot_i[63];
  assign data_masked[4055] = data_i[4055] & sel_one_hot_i[63];
  assign data_masked[4054] = data_i[4054] & sel_one_hot_i[63];
  assign data_masked[4053] = data_i[4053] & sel_one_hot_i[63];
  assign data_masked[4052] = data_i[4052] & sel_one_hot_i[63];
  assign data_masked[4051] = data_i[4051] & sel_one_hot_i[63];
  assign data_masked[4050] = data_i[4050] & sel_one_hot_i[63];
  assign data_masked[4049] = data_i[4049] & sel_one_hot_i[63];
  assign data_masked[4048] = data_i[4048] & sel_one_hot_i[63];
  assign data_masked[4047] = data_i[4047] & sel_one_hot_i[63];
  assign data_masked[4046] = data_i[4046] & sel_one_hot_i[63];
  assign data_masked[4045] = data_i[4045] & sel_one_hot_i[63];
  assign data_masked[4044] = data_i[4044] & sel_one_hot_i[63];
  assign data_masked[4043] = data_i[4043] & sel_one_hot_i[63];
  assign data_masked[4042] = data_i[4042] & sel_one_hot_i[63];
  assign data_masked[4041] = data_i[4041] & sel_one_hot_i[63];
  assign data_masked[4040] = data_i[4040] & sel_one_hot_i[63];
  assign data_masked[4039] = data_i[4039] & sel_one_hot_i[63];
  assign data_masked[4038] = data_i[4038] & sel_one_hot_i[63];
  assign data_masked[4037] = data_i[4037] & sel_one_hot_i[63];
  assign data_masked[4036] = data_i[4036] & sel_one_hot_i[63];
  assign data_masked[4035] = data_i[4035] & sel_one_hot_i[63];
  assign data_masked[4034] = data_i[4034] & sel_one_hot_i[63];
  assign data_masked[4033] = data_i[4033] & sel_one_hot_i[63];
  assign data_masked[4032] = data_i[4032] & sel_one_hot_i[63];
  assign data_o[0] = N61 | data_masked[0];
  assign N61 = N60 | data_masked[64];
  assign N60 = N59 | data_masked[128];
  assign N59 = N58 | data_masked[192];
  assign N58 = N57 | data_masked[256];
  assign N57 = N56 | data_masked[320];
  assign N56 = N55 | data_masked[384];
  assign N55 = N54 | data_masked[448];
  assign N54 = N53 | data_masked[512];
  assign N53 = N52 | data_masked[576];
  assign N52 = N51 | data_masked[640];
  assign N51 = N50 | data_masked[704];
  assign N50 = N49 | data_masked[768];
  assign N49 = N48 | data_masked[832];
  assign N48 = N47 | data_masked[896];
  assign N47 = N46 | data_masked[960];
  assign N46 = N45 | data_masked[1024];
  assign N45 = N44 | data_masked[1088];
  assign N44 = N43 | data_masked[1152];
  assign N43 = N42 | data_masked[1216];
  assign N42 = N41 | data_masked[1280];
  assign N41 = N40 | data_masked[1344];
  assign N40 = N39 | data_masked[1408];
  assign N39 = N38 | data_masked[1472];
  assign N38 = N37 | data_masked[1536];
  assign N37 = N36 | data_masked[1600];
  assign N36 = N35 | data_masked[1664];
  assign N35 = N34 | data_masked[1728];
  assign N34 = N33 | data_masked[1792];
  assign N33 = N32 | data_masked[1856];
  assign N32 = N31 | data_masked[1920];
  assign N31 = N30 | data_masked[1984];
  assign N30 = N29 | data_masked[2048];
  assign N29 = N28 | data_masked[2112];
  assign N28 = N27 | data_masked[2176];
  assign N27 = N26 | data_masked[2240];
  assign N26 = N25 | data_masked[2304];
  assign N25 = N24 | data_masked[2368];
  assign N24 = N23 | data_masked[2432];
  assign N23 = N22 | data_masked[2496];
  assign N22 = N21 | data_masked[2560];
  assign N21 = N20 | data_masked[2624];
  assign N20 = N19 | data_masked[2688];
  assign N19 = N18 | data_masked[2752];
  assign N18 = N17 | data_masked[2816];
  assign N17 = N16 | data_masked[2880];
  assign N16 = N15 | data_masked[2944];
  assign N15 = N14 | data_masked[3008];
  assign N14 = N13 | data_masked[3072];
  assign N13 = N12 | data_masked[3136];
  assign N12 = N11 | data_masked[3200];
  assign N11 = N10 | data_masked[3264];
  assign N10 = N9 | data_masked[3328];
  assign N9 = N8 | data_masked[3392];
  assign N8 = N7 | data_masked[3456];
  assign N7 = N6 | data_masked[3520];
  assign N6 = N5 | data_masked[3584];
  assign N5 = N4 | data_masked[3648];
  assign N4 = N3 | data_masked[3712];
  assign N3 = N2 | data_masked[3776];
  assign N2 = N1 | data_masked[3840];
  assign N1 = N0 | data_masked[3904];
  assign N0 = data_masked[4032] | data_masked[3968];
  assign data_o[1] = N123 | data_masked[1];
  assign N123 = N122 | data_masked[65];
  assign N122 = N121 | data_masked[129];
  assign N121 = N120 | data_masked[193];
  assign N120 = N119 | data_masked[257];
  assign N119 = N118 | data_masked[321];
  assign N118 = N117 | data_masked[385];
  assign N117 = N116 | data_masked[449];
  assign N116 = N115 | data_masked[513];
  assign N115 = N114 | data_masked[577];
  assign N114 = N113 | data_masked[641];
  assign N113 = N112 | data_masked[705];
  assign N112 = N111 | data_masked[769];
  assign N111 = N110 | data_masked[833];
  assign N110 = N109 | data_masked[897];
  assign N109 = N108 | data_masked[961];
  assign N108 = N107 | data_masked[1025];
  assign N107 = N106 | data_masked[1089];
  assign N106 = N105 | data_masked[1153];
  assign N105 = N104 | data_masked[1217];
  assign N104 = N103 | data_masked[1281];
  assign N103 = N102 | data_masked[1345];
  assign N102 = N101 | data_masked[1409];
  assign N101 = N100 | data_masked[1473];
  assign N100 = N99 | data_masked[1537];
  assign N99 = N98 | data_masked[1601];
  assign N98 = N97 | data_masked[1665];
  assign N97 = N96 | data_masked[1729];
  assign N96 = N95 | data_masked[1793];
  assign N95 = N94 | data_masked[1857];
  assign N94 = N93 | data_masked[1921];
  assign N93 = N92 | data_masked[1985];
  assign N92 = N91 | data_masked[2049];
  assign N91 = N90 | data_masked[2113];
  assign N90 = N89 | data_masked[2177];
  assign N89 = N88 | data_masked[2241];
  assign N88 = N87 | data_masked[2305];
  assign N87 = N86 | data_masked[2369];
  assign N86 = N85 | data_masked[2433];
  assign N85 = N84 | data_masked[2497];
  assign N84 = N83 | data_masked[2561];
  assign N83 = N82 | data_masked[2625];
  assign N82 = N81 | data_masked[2689];
  assign N81 = N80 | data_masked[2753];
  assign N80 = N79 | data_masked[2817];
  assign N79 = N78 | data_masked[2881];
  assign N78 = N77 | data_masked[2945];
  assign N77 = N76 | data_masked[3009];
  assign N76 = N75 | data_masked[3073];
  assign N75 = N74 | data_masked[3137];
  assign N74 = N73 | data_masked[3201];
  assign N73 = N72 | data_masked[3265];
  assign N72 = N71 | data_masked[3329];
  assign N71 = N70 | data_masked[3393];
  assign N70 = N69 | data_masked[3457];
  assign N69 = N68 | data_masked[3521];
  assign N68 = N67 | data_masked[3585];
  assign N67 = N66 | data_masked[3649];
  assign N66 = N65 | data_masked[3713];
  assign N65 = N64 | data_masked[3777];
  assign N64 = N63 | data_masked[3841];
  assign N63 = N62 | data_masked[3905];
  assign N62 = data_masked[4033] | data_masked[3969];
  assign data_o[2] = N185 | data_masked[2];
  assign N185 = N184 | data_masked[66];
  assign N184 = N183 | data_masked[130];
  assign N183 = N182 | data_masked[194];
  assign N182 = N181 | data_masked[258];
  assign N181 = N180 | data_masked[322];
  assign N180 = N179 | data_masked[386];
  assign N179 = N178 | data_masked[450];
  assign N178 = N177 | data_masked[514];
  assign N177 = N176 | data_masked[578];
  assign N176 = N175 | data_masked[642];
  assign N175 = N174 | data_masked[706];
  assign N174 = N173 | data_masked[770];
  assign N173 = N172 | data_masked[834];
  assign N172 = N171 | data_masked[898];
  assign N171 = N170 | data_masked[962];
  assign N170 = N169 | data_masked[1026];
  assign N169 = N168 | data_masked[1090];
  assign N168 = N167 | data_masked[1154];
  assign N167 = N166 | data_masked[1218];
  assign N166 = N165 | data_masked[1282];
  assign N165 = N164 | data_masked[1346];
  assign N164 = N163 | data_masked[1410];
  assign N163 = N162 | data_masked[1474];
  assign N162 = N161 | data_masked[1538];
  assign N161 = N160 | data_masked[1602];
  assign N160 = N159 | data_masked[1666];
  assign N159 = N158 | data_masked[1730];
  assign N158 = N157 | data_masked[1794];
  assign N157 = N156 | data_masked[1858];
  assign N156 = N155 | data_masked[1922];
  assign N155 = N154 | data_masked[1986];
  assign N154 = N153 | data_masked[2050];
  assign N153 = N152 | data_masked[2114];
  assign N152 = N151 | data_masked[2178];
  assign N151 = N150 | data_masked[2242];
  assign N150 = N149 | data_masked[2306];
  assign N149 = N148 | data_masked[2370];
  assign N148 = N147 | data_masked[2434];
  assign N147 = N146 | data_masked[2498];
  assign N146 = N145 | data_masked[2562];
  assign N145 = N144 | data_masked[2626];
  assign N144 = N143 | data_masked[2690];
  assign N143 = N142 | data_masked[2754];
  assign N142 = N141 | data_masked[2818];
  assign N141 = N140 | data_masked[2882];
  assign N140 = N139 | data_masked[2946];
  assign N139 = N138 | data_masked[3010];
  assign N138 = N137 | data_masked[3074];
  assign N137 = N136 | data_masked[3138];
  assign N136 = N135 | data_masked[3202];
  assign N135 = N134 | data_masked[3266];
  assign N134 = N133 | data_masked[3330];
  assign N133 = N132 | data_masked[3394];
  assign N132 = N131 | data_masked[3458];
  assign N131 = N130 | data_masked[3522];
  assign N130 = N129 | data_masked[3586];
  assign N129 = N128 | data_masked[3650];
  assign N128 = N127 | data_masked[3714];
  assign N127 = N126 | data_masked[3778];
  assign N126 = N125 | data_masked[3842];
  assign N125 = N124 | data_masked[3906];
  assign N124 = data_masked[4034] | data_masked[3970];
  assign data_o[3] = N247 | data_masked[3];
  assign N247 = N246 | data_masked[67];
  assign N246 = N245 | data_masked[131];
  assign N245 = N244 | data_masked[195];
  assign N244 = N243 | data_masked[259];
  assign N243 = N242 | data_masked[323];
  assign N242 = N241 | data_masked[387];
  assign N241 = N240 | data_masked[451];
  assign N240 = N239 | data_masked[515];
  assign N239 = N238 | data_masked[579];
  assign N238 = N237 | data_masked[643];
  assign N237 = N236 | data_masked[707];
  assign N236 = N235 | data_masked[771];
  assign N235 = N234 | data_masked[835];
  assign N234 = N233 | data_masked[899];
  assign N233 = N232 | data_masked[963];
  assign N232 = N231 | data_masked[1027];
  assign N231 = N230 | data_masked[1091];
  assign N230 = N229 | data_masked[1155];
  assign N229 = N228 | data_masked[1219];
  assign N228 = N227 | data_masked[1283];
  assign N227 = N226 | data_masked[1347];
  assign N226 = N225 | data_masked[1411];
  assign N225 = N224 | data_masked[1475];
  assign N224 = N223 | data_masked[1539];
  assign N223 = N222 | data_masked[1603];
  assign N222 = N221 | data_masked[1667];
  assign N221 = N220 | data_masked[1731];
  assign N220 = N219 | data_masked[1795];
  assign N219 = N218 | data_masked[1859];
  assign N218 = N217 | data_masked[1923];
  assign N217 = N216 | data_masked[1987];
  assign N216 = N215 | data_masked[2051];
  assign N215 = N214 | data_masked[2115];
  assign N214 = N213 | data_masked[2179];
  assign N213 = N212 | data_masked[2243];
  assign N212 = N211 | data_masked[2307];
  assign N211 = N210 | data_masked[2371];
  assign N210 = N209 | data_masked[2435];
  assign N209 = N208 | data_masked[2499];
  assign N208 = N207 | data_masked[2563];
  assign N207 = N206 | data_masked[2627];
  assign N206 = N205 | data_masked[2691];
  assign N205 = N204 | data_masked[2755];
  assign N204 = N203 | data_masked[2819];
  assign N203 = N202 | data_masked[2883];
  assign N202 = N201 | data_masked[2947];
  assign N201 = N200 | data_masked[3011];
  assign N200 = N199 | data_masked[3075];
  assign N199 = N198 | data_masked[3139];
  assign N198 = N197 | data_masked[3203];
  assign N197 = N196 | data_masked[3267];
  assign N196 = N195 | data_masked[3331];
  assign N195 = N194 | data_masked[3395];
  assign N194 = N193 | data_masked[3459];
  assign N193 = N192 | data_masked[3523];
  assign N192 = N191 | data_masked[3587];
  assign N191 = N190 | data_masked[3651];
  assign N190 = N189 | data_masked[3715];
  assign N189 = N188 | data_masked[3779];
  assign N188 = N187 | data_masked[3843];
  assign N187 = N186 | data_masked[3907];
  assign N186 = data_masked[4035] | data_masked[3971];
  assign data_o[4] = N309 | data_masked[4];
  assign N309 = N308 | data_masked[68];
  assign N308 = N307 | data_masked[132];
  assign N307 = N306 | data_masked[196];
  assign N306 = N305 | data_masked[260];
  assign N305 = N304 | data_masked[324];
  assign N304 = N303 | data_masked[388];
  assign N303 = N302 | data_masked[452];
  assign N302 = N301 | data_masked[516];
  assign N301 = N300 | data_masked[580];
  assign N300 = N299 | data_masked[644];
  assign N299 = N298 | data_masked[708];
  assign N298 = N297 | data_masked[772];
  assign N297 = N296 | data_masked[836];
  assign N296 = N295 | data_masked[900];
  assign N295 = N294 | data_masked[964];
  assign N294 = N293 | data_masked[1028];
  assign N293 = N292 | data_masked[1092];
  assign N292 = N291 | data_masked[1156];
  assign N291 = N290 | data_masked[1220];
  assign N290 = N289 | data_masked[1284];
  assign N289 = N288 | data_masked[1348];
  assign N288 = N287 | data_masked[1412];
  assign N287 = N286 | data_masked[1476];
  assign N286 = N285 | data_masked[1540];
  assign N285 = N284 | data_masked[1604];
  assign N284 = N283 | data_masked[1668];
  assign N283 = N282 | data_masked[1732];
  assign N282 = N281 | data_masked[1796];
  assign N281 = N280 | data_masked[1860];
  assign N280 = N279 | data_masked[1924];
  assign N279 = N278 | data_masked[1988];
  assign N278 = N277 | data_masked[2052];
  assign N277 = N276 | data_masked[2116];
  assign N276 = N275 | data_masked[2180];
  assign N275 = N274 | data_masked[2244];
  assign N274 = N273 | data_masked[2308];
  assign N273 = N272 | data_masked[2372];
  assign N272 = N271 | data_masked[2436];
  assign N271 = N270 | data_masked[2500];
  assign N270 = N269 | data_masked[2564];
  assign N269 = N268 | data_masked[2628];
  assign N268 = N267 | data_masked[2692];
  assign N267 = N266 | data_masked[2756];
  assign N266 = N265 | data_masked[2820];
  assign N265 = N264 | data_masked[2884];
  assign N264 = N263 | data_masked[2948];
  assign N263 = N262 | data_masked[3012];
  assign N262 = N261 | data_masked[3076];
  assign N261 = N260 | data_masked[3140];
  assign N260 = N259 | data_masked[3204];
  assign N259 = N258 | data_masked[3268];
  assign N258 = N257 | data_masked[3332];
  assign N257 = N256 | data_masked[3396];
  assign N256 = N255 | data_masked[3460];
  assign N255 = N254 | data_masked[3524];
  assign N254 = N253 | data_masked[3588];
  assign N253 = N252 | data_masked[3652];
  assign N252 = N251 | data_masked[3716];
  assign N251 = N250 | data_masked[3780];
  assign N250 = N249 | data_masked[3844];
  assign N249 = N248 | data_masked[3908];
  assign N248 = data_masked[4036] | data_masked[3972];
  assign data_o[5] = N371 | data_masked[5];
  assign N371 = N370 | data_masked[69];
  assign N370 = N369 | data_masked[133];
  assign N369 = N368 | data_masked[197];
  assign N368 = N367 | data_masked[261];
  assign N367 = N366 | data_masked[325];
  assign N366 = N365 | data_masked[389];
  assign N365 = N364 | data_masked[453];
  assign N364 = N363 | data_masked[517];
  assign N363 = N362 | data_masked[581];
  assign N362 = N361 | data_masked[645];
  assign N361 = N360 | data_masked[709];
  assign N360 = N359 | data_masked[773];
  assign N359 = N358 | data_masked[837];
  assign N358 = N357 | data_masked[901];
  assign N357 = N356 | data_masked[965];
  assign N356 = N355 | data_masked[1029];
  assign N355 = N354 | data_masked[1093];
  assign N354 = N353 | data_masked[1157];
  assign N353 = N352 | data_masked[1221];
  assign N352 = N351 | data_masked[1285];
  assign N351 = N350 | data_masked[1349];
  assign N350 = N349 | data_masked[1413];
  assign N349 = N348 | data_masked[1477];
  assign N348 = N347 | data_masked[1541];
  assign N347 = N346 | data_masked[1605];
  assign N346 = N345 | data_masked[1669];
  assign N345 = N344 | data_masked[1733];
  assign N344 = N343 | data_masked[1797];
  assign N343 = N342 | data_masked[1861];
  assign N342 = N341 | data_masked[1925];
  assign N341 = N340 | data_masked[1989];
  assign N340 = N339 | data_masked[2053];
  assign N339 = N338 | data_masked[2117];
  assign N338 = N337 | data_masked[2181];
  assign N337 = N336 | data_masked[2245];
  assign N336 = N335 | data_masked[2309];
  assign N335 = N334 | data_masked[2373];
  assign N334 = N333 | data_masked[2437];
  assign N333 = N332 | data_masked[2501];
  assign N332 = N331 | data_masked[2565];
  assign N331 = N330 | data_masked[2629];
  assign N330 = N329 | data_masked[2693];
  assign N329 = N328 | data_masked[2757];
  assign N328 = N327 | data_masked[2821];
  assign N327 = N326 | data_masked[2885];
  assign N326 = N325 | data_masked[2949];
  assign N325 = N324 | data_masked[3013];
  assign N324 = N323 | data_masked[3077];
  assign N323 = N322 | data_masked[3141];
  assign N322 = N321 | data_masked[3205];
  assign N321 = N320 | data_masked[3269];
  assign N320 = N319 | data_masked[3333];
  assign N319 = N318 | data_masked[3397];
  assign N318 = N317 | data_masked[3461];
  assign N317 = N316 | data_masked[3525];
  assign N316 = N315 | data_masked[3589];
  assign N315 = N314 | data_masked[3653];
  assign N314 = N313 | data_masked[3717];
  assign N313 = N312 | data_masked[3781];
  assign N312 = N311 | data_masked[3845];
  assign N311 = N310 | data_masked[3909];
  assign N310 = data_masked[4037] | data_masked[3973];
  assign data_o[6] = N433 | data_masked[6];
  assign N433 = N432 | data_masked[70];
  assign N432 = N431 | data_masked[134];
  assign N431 = N430 | data_masked[198];
  assign N430 = N429 | data_masked[262];
  assign N429 = N428 | data_masked[326];
  assign N428 = N427 | data_masked[390];
  assign N427 = N426 | data_masked[454];
  assign N426 = N425 | data_masked[518];
  assign N425 = N424 | data_masked[582];
  assign N424 = N423 | data_masked[646];
  assign N423 = N422 | data_masked[710];
  assign N422 = N421 | data_masked[774];
  assign N421 = N420 | data_masked[838];
  assign N420 = N419 | data_masked[902];
  assign N419 = N418 | data_masked[966];
  assign N418 = N417 | data_masked[1030];
  assign N417 = N416 | data_masked[1094];
  assign N416 = N415 | data_masked[1158];
  assign N415 = N414 | data_masked[1222];
  assign N414 = N413 | data_masked[1286];
  assign N413 = N412 | data_masked[1350];
  assign N412 = N411 | data_masked[1414];
  assign N411 = N410 | data_masked[1478];
  assign N410 = N409 | data_masked[1542];
  assign N409 = N408 | data_masked[1606];
  assign N408 = N407 | data_masked[1670];
  assign N407 = N406 | data_masked[1734];
  assign N406 = N405 | data_masked[1798];
  assign N405 = N404 | data_masked[1862];
  assign N404 = N403 | data_masked[1926];
  assign N403 = N402 | data_masked[1990];
  assign N402 = N401 | data_masked[2054];
  assign N401 = N400 | data_masked[2118];
  assign N400 = N399 | data_masked[2182];
  assign N399 = N398 | data_masked[2246];
  assign N398 = N397 | data_masked[2310];
  assign N397 = N396 | data_masked[2374];
  assign N396 = N395 | data_masked[2438];
  assign N395 = N394 | data_masked[2502];
  assign N394 = N393 | data_masked[2566];
  assign N393 = N392 | data_masked[2630];
  assign N392 = N391 | data_masked[2694];
  assign N391 = N390 | data_masked[2758];
  assign N390 = N389 | data_masked[2822];
  assign N389 = N388 | data_masked[2886];
  assign N388 = N387 | data_masked[2950];
  assign N387 = N386 | data_masked[3014];
  assign N386 = N385 | data_masked[3078];
  assign N385 = N384 | data_masked[3142];
  assign N384 = N383 | data_masked[3206];
  assign N383 = N382 | data_masked[3270];
  assign N382 = N381 | data_masked[3334];
  assign N381 = N380 | data_masked[3398];
  assign N380 = N379 | data_masked[3462];
  assign N379 = N378 | data_masked[3526];
  assign N378 = N377 | data_masked[3590];
  assign N377 = N376 | data_masked[3654];
  assign N376 = N375 | data_masked[3718];
  assign N375 = N374 | data_masked[3782];
  assign N374 = N373 | data_masked[3846];
  assign N373 = N372 | data_masked[3910];
  assign N372 = data_masked[4038] | data_masked[3974];
  assign data_o[7] = N495 | data_masked[7];
  assign N495 = N494 | data_masked[71];
  assign N494 = N493 | data_masked[135];
  assign N493 = N492 | data_masked[199];
  assign N492 = N491 | data_masked[263];
  assign N491 = N490 | data_masked[327];
  assign N490 = N489 | data_masked[391];
  assign N489 = N488 | data_masked[455];
  assign N488 = N487 | data_masked[519];
  assign N487 = N486 | data_masked[583];
  assign N486 = N485 | data_masked[647];
  assign N485 = N484 | data_masked[711];
  assign N484 = N483 | data_masked[775];
  assign N483 = N482 | data_masked[839];
  assign N482 = N481 | data_masked[903];
  assign N481 = N480 | data_masked[967];
  assign N480 = N479 | data_masked[1031];
  assign N479 = N478 | data_masked[1095];
  assign N478 = N477 | data_masked[1159];
  assign N477 = N476 | data_masked[1223];
  assign N476 = N475 | data_masked[1287];
  assign N475 = N474 | data_masked[1351];
  assign N474 = N473 | data_masked[1415];
  assign N473 = N472 | data_masked[1479];
  assign N472 = N471 | data_masked[1543];
  assign N471 = N470 | data_masked[1607];
  assign N470 = N469 | data_masked[1671];
  assign N469 = N468 | data_masked[1735];
  assign N468 = N467 | data_masked[1799];
  assign N467 = N466 | data_masked[1863];
  assign N466 = N465 | data_masked[1927];
  assign N465 = N464 | data_masked[1991];
  assign N464 = N463 | data_masked[2055];
  assign N463 = N462 | data_masked[2119];
  assign N462 = N461 | data_masked[2183];
  assign N461 = N460 | data_masked[2247];
  assign N460 = N459 | data_masked[2311];
  assign N459 = N458 | data_masked[2375];
  assign N458 = N457 | data_masked[2439];
  assign N457 = N456 | data_masked[2503];
  assign N456 = N455 | data_masked[2567];
  assign N455 = N454 | data_masked[2631];
  assign N454 = N453 | data_masked[2695];
  assign N453 = N452 | data_masked[2759];
  assign N452 = N451 | data_masked[2823];
  assign N451 = N450 | data_masked[2887];
  assign N450 = N449 | data_masked[2951];
  assign N449 = N448 | data_masked[3015];
  assign N448 = N447 | data_masked[3079];
  assign N447 = N446 | data_masked[3143];
  assign N446 = N445 | data_masked[3207];
  assign N445 = N444 | data_masked[3271];
  assign N444 = N443 | data_masked[3335];
  assign N443 = N442 | data_masked[3399];
  assign N442 = N441 | data_masked[3463];
  assign N441 = N440 | data_masked[3527];
  assign N440 = N439 | data_masked[3591];
  assign N439 = N438 | data_masked[3655];
  assign N438 = N437 | data_masked[3719];
  assign N437 = N436 | data_masked[3783];
  assign N436 = N435 | data_masked[3847];
  assign N435 = N434 | data_masked[3911];
  assign N434 = data_masked[4039] | data_masked[3975];
  assign data_o[8] = N557 | data_masked[8];
  assign N557 = N556 | data_masked[72];
  assign N556 = N555 | data_masked[136];
  assign N555 = N554 | data_masked[200];
  assign N554 = N553 | data_masked[264];
  assign N553 = N552 | data_masked[328];
  assign N552 = N551 | data_masked[392];
  assign N551 = N550 | data_masked[456];
  assign N550 = N549 | data_masked[520];
  assign N549 = N548 | data_masked[584];
  assign N548 = N547 | data_masked[648];
  assign N547 = N546 | data_masked[712];
  assign N546 = N545 | data_masked[776];
  assign N545 = N544 | data_masked[840];
  assign N544 = N543 | data_masked[904];
  assign N543 = N542 | data_masked[968];
  assign N542 = N541 | data_masked[1032];
  assign N541 = N540 | data_masked[1096];
  assign N540 = N539 | data_masked[1160];
  assign N539 = N538 | data_masked[1224];
  assign N538 = N537 | data_masked[1288];
  assign N537 = N536 | data_masked[1352];
  assign N536 = N535 | data_masked[1416];
  assign N535 = N534 | data_masked[1480];
  assign N534 = N533 | data_masked[1544];
  assign N533 = N532 | data_masked[1608];
  assign N532 = N531 | data_masked[1672];
  assign N531 = N530 | data_masked[1736];
  assign N530 = N529 | data_masked[1800];
  assign N529 = N528 | data_masked[1864];
  assign N528 = N527 | data_masked[1928];
  assign N527 = N526 | data_masked[1992];
  assign N526 = N525 | data_masked[2056];
  assign N525 = N524 | data_masked[2120];
  assign N524 = N523 | data_masked[2184];
  assign N523 = N522 | data_masked[2248];
  assign N522 = N521 | data_masked[2312];
  assign N521 = N520 | data_masked[2376];
  assign N520 = N519 | data_masked[2440];
  assign N519 = N518 | data_masked[2504];
  assign N518 = N517 | data_masked[2568];
  assign N517 = N516 | data_masked[2632];
  assign N516 = N515 | data_masked[2696];
  assign N515 = N514 | data_masked[2760];
  assign N514 = N513 | data_masked[2824];
  assign N513 = N512 | data_masked[2888];
  assign N512 = N511 | data_masked[2952];
  assign N511 = N510 | data_masked[3016];
  assign N510 = N509 | data_masked[3080];
  assign N509 = N508 | data_masked[3144];
  assign N508 = N507 | data_masked[3208];
  assign N507 = N506 | data_masked[3272];
  assign N506 = N505 | data_masked[3336];
  assign N505 = N504 | data_masked[3400];
  assign N504 = N503 | data_masked[3464];
  assign N503 = N502 | data_masked[3528];
  assign N502 = N501 | data_masked[3592];
  assign N501 = N500 | data_masked[3656];
  assign N500 = N499 | data_masked[3720];
  assign N499 = N498 | data_masked[3784];
  assign N498 = N497 | data_masked[3848];
  assign N497 = N496 | data_masked[3912];
  assign N496 = data_masked[4040] | data_masked[3976];
  assign data_o[9] = N619 | data_masked[9];
  assign N619 = N618 | data_masked[73];
  assign N618 = N617 | data_masked[137];
  assign N617 = N616 | data_masked[201];
  assign N616 = N615 | data_masked[265];
  assign N615 = N614 | data_masked[329];
  assign N614 = N613 | data_masked[393];
  assign N613 = N612 | data_masked[457];
  assign N612 = N611 | data_masked[521];
  assign N611 = N610 | data_masked[585];
  assign N610 = N609 | data_masked[649];
  assign N609 = N608 | data_masked[713];
  assign N608 = N607 | data_masked[777];
  assign N607 = N606 | data_masked[841];
  assign N606 = N605 | data_masked[905];
  assign N605 = N604 | data_masked[969];
  assign N604 = N603 | data_masked[1033];
  assign N603 = N602 | data_masked[1097];
  assign N602 = N601 | data_masked[1161];
  assign N601 = N600 | data_masked[1225];
  assign N600 = N599 | data_masked[1289];
  assign N599 = N598 | data_masked[1353];
  assign N598 = N597 | data_masked[1417];
  assign N597 = N596 | data_masked[1481];
  assign N596 = N595 | data_masked[1545];
  assign N595 = N594 | data_masked[1609];
  assign N594 = N593 | data_masked[1673];
  assign N593 = N592 | data_masked[1737];
  assign N592 = N591 | data_masked[1801];
  assign N591 = N590 | data_masked[1865];
  assign N590 = N589 | data_masked[1929];
  assign N589 = N588 | data_masked[1993];
  assign N588 = N587 | data_masked[2057];
  assign N587 = N586 | data_masked[2121];
  assign N586 = N585 | data_masked[2185];
  assign N585 = N584 | data_masked[2249];
  assign N584 = N583 | data_masked[2313];
  assign N583 = N582 | data_masked[2377];
  assign N582 = N581 | data_masked[2441];
  assign N581 = N580 | data_masked[2505];
  assign N580 = N579 | data_masked[2569];
  assign N579 = N578 | data_masked[2633];
  assign N578 = N577 | data_masked[2697];
  assign N577 = N576 | data_masked[2761];
  assign N576 = N575 | data_masked[2825];
  assign N575 = N574 | data_masked[2889];
  assign N574 = N573 | data_masked[2953];
  assign N573 = N572 | data_masked[3017];
  assign N572 = N571 | data_masked[3081];
  assign N571 = N570 | data_masked[3145];
  assign N570 = N569 | data_masked[3209];
  assign N569 = N568 | data_masked[3273];
  assign N568 = N567 | data_masked[3337];
  assign N567 = N566 | data_masked[3401];
  assign N566 = N565 | data_masked[3465];
  assign N565 = N564 | data_masked[3529];
  assign N564 = N563 | data_masked[3593];
  assign N563 = N562 | data_masked[3657];
  assign N562 = N561 | data_masked[3721];
  assign N561 = N560 | data_masked[3785];
  assign N560 = N559 | data_masked[3849];
  assign N559 = N558 | data_masked[3913];
  assign N558 = data_masked[4041] | data_masked[3977];
  assign data_o[10] = N681 | data_masked[10];
  assign N681 = N680 | data_masked[74];
  assign N680 = N679 | data_masked[138];
  assign N679 = N678 | data_masked[202];
  assign N678 = N677 | data_masked[266];
  assign N677 = N676 | data_masked[330];
  assign N676 = N675 | data_masked[394];
  assign N675 = N674 | data_masked[458];
  assign N674 = N673 | data_masked[522];
  assign N673 = N672 | data_masked[586];
  assign N672 = N671 | data_masked[650];
  assign N671 = N670 | data_masked[714];
  assign N670 = N669 | data_masked[778];
  assign N669 = N668 | data_masked[842];
  assign N668 = N667 | data_masked[906];
  assign N667 = N666 | data_masked[970];
  assign N666 = N665 | data_masked[1034];
  assign N665 = N664 | data_masked[1098];
  assign N664 = N663 | data_masked[1162];
  assign N663 = N662 | data_masked[1226];
  assign N662 = N661 | data_masked[1290];
  assign N661 = N660 | data_masked[1354];
  assign N660 = N659 | data_masked[1418];
  assign N659 = N658 | data_masked[1482];
  assign N658 = N657 | data_masked[1546];
  assign N657 = N656 | data_masked[1610];
  assign N656 = N655 | data_masked[1674];
  assign N655 = N654 | data_masked[1738];
  assign N654 = N653 | data_masked[1802];
  assign N653 = N652 | data_masked[1866];
  assign N652 = N651 | data_masked[1930];
  assign N651 = N650 | data_masked[1994];
  assign N650 = N649 | data_masked[2058];
  assign N649 = N648 | data_masked[2122];
  assign N648 = N647 | data_masked[2186];
  assign N647 = N646 | data_masked[2250];
  assign N646 = N645 | data_masked[2314];
  assign N645 = N644 | data_masked[2378];
  assign N644 = N643 | data_masked[2442];
  assign N643 = N642 | data_masked[2506];
  assign N642 = N641 | data_masked[2570];
  assign N641 = N640 | data_masked[2634];
  assign N640 = N639 | data_masked[2698];
  assign N639 = N638 | data_masked[2762];
  assign N638 = N637 | data_masked[2826];
  assign N637 = N636 | data_masked[2890];
  assign N636 = N635 | data_masked[2954];
  assign N635 = N634 | data_masked[3018];
  assign N634 = N633 | data_masked[3082];
  assign N633 = N632 | data_masked[3146];
  assign N632 = N631 | data_masked[3210];
  assign N631 = N630 | data_masked[3274];
  assign N630 = N629 | data_masked[3338];
  assign N629 = N628 | data_masked[3402];
  assign N628 = N627 | data_masked[3466];
  assign N627 = N626 | data_masked[3530];
  assign N626 = N625 | data_masked[3594];
  assign N625 = N624 | data_masked[3658];
  assign N624 = N623 | data_masked[3722];
  assign N623 = N622 | data_masked[3786];
  assign N622 = N621 | data_masked[3850];
  assign N621 = N620 | data_masked[3914];
  assign N620 = data_masked[4042] | data_masked[3978];
  assign data_o[11] = N743 | data_masked[11];
  assign N743 = N742 | data_masked[75];
  assign N742 = N741 | data_masked[139];
  assign N741 = N740 | data_masked[203];
  assign N740 = N739 | data_masked[267];
  assign N739 = N738 | data_masked[331];
  assign N738 = N737 | data_masked[395];
  assign N737 = N736 | data_masked[459];
  assign N736 = N735 | data_masked[523];
  assign N735 = N734 | data_masked[587];
  assign N734 = N733 | data_masked[651];
  assign N733 = N732 | data_masked[715];
  assign N732 = N731 | data_masked[779];
  assign N731 = N730 | data_masked[843];
  assign N730 = N729 | data_masked[907];
  assign N729 = N728 | data_masked[971];
  assign N728 = N727 | data_masked[1035];
  assign N727 = N726 | data_masked[1099];
  assign N726 = N725 | data_masked[1163];
  assign N725 = N724 | data_masked[1227];
  assign N724 = N723 | data_masked[1291];
  assign N723 = N722 | data_masked[1355];
  assign N722 = N721 | data_masked[1419];
  assign N721 = N720 | data_masked[1483];
  assign N720 = N719 | data_masked[1547];
  assign N719 = N718 | data_masked[1611];
  assign N718 = N717 | data_masked[1675];
  assign N717 = N716 | data_masked[1739];
  assign N716 = N715 | data_masked[1803];
  assign N715 = N714 | data_masked[1867];
  assign N714 = N713 | data_masked[1931];
  assign N713 = N712 | data_masked[1995];
  assign N712 = N711 | data_masked[2059];
  assign N711 = N710 | data_masked[2123];
  assign N710 = N709 | data_masked[2187];
  assign N709 = N708 | data_masked[2251];
  assign N708 = N707 | data_masked[2315];
  assign N707 = N706 | data_masked[2379];
  assign N706 = N705 | data_masked[2443];
  assign N705 = N704 | data_masked[2507];
  assign N704 = N703 | data_masked[2571];
  assign N703 = N702 | data_masked[2635];
  assign N702 = N701 | data_masked[2699];
  assign N701 = N700 | data_masked[2763];
  assign N700 = N699 | data_masked[2827];
  assign N699 = N698 | data_masked[2891];
  assign N698 = N697 | data_masked[2955];
  assign N697 = N696 | data_masked[3019];
  assign N696 = N695 | data_masked[3083];
  assign N695 = N694 | data_masked[3147];
  assign N694 = N693 | data_masked[3211];
  assign N693 = N692 | data_masked[3275];
  assign N692 = N691 | data_masked[3339];
  assign N691 = N690 | data_masked[3403];
  assign N690 = N689 | data_masked[3467];
  assign N689 = N688 | data_masked[3531];
  assign N688 = N687 | data_masked[3595];
  assign N687 = N686 | data_masked[3659];
  assign N686 = N685 | data_masked[3723];
  assign N685 = N684 | data_masked[3787];
  assign N684 = N683 | data_masked[3851];
  assign N683 = N682 | data_masked[3915];
  assign N682 = data_masked[4043] | data_masked[3979];
  assign data_o[12] = N805 | data_masked[12];
  assign N805 = N804 | data_masked[76];
  assign N804 = N803 | data_masked[140];
  assign N803 = N802 | data_masked[204];
  assign N802 = N801 | data_masked[268];
  assign N801 = N800 | data_masked[332];
  assign N800 = N799 | data_masked[396];
  assign N799 = N798 | data_masked[460];
  assign N798 = N797 | data_masked[524];
  assign N797 = N796 | data_masked[588];
  assign N796 = N795 | data_masked[652];
  assign N795 = N794 | data_masked[716];
  assign N794 = N793 | data_masked[780];
  assign N793 = N792 | data_masked[844];
  assign N792 = N791 | data_masked[908];
  assign N791 = N790 | data_masked[972];
  assign N790 = N789 | data_masked[1036];
  assign N789 = N788 | data_masked[1100];
  assign N788 = N787 | data_masked[1164];
  assign N787 = N786 | data_masked[1228];
  assign N786 = N785 | data_masked[1292];
  assign N785 = N784 | data_masked[1356];
  assign N784 = N783 | data_masked[1420];
  assign N783 = N782 | data_masked[1484];
  assign N782 = N781 | data_masked[1548];
  assign N781 = N780 | data_masked[1612];
  assign N780 = N779 | data_masked[1676];
  assign N779 = N778 | data_masked[1740];
  assign N778 = N777 | data_masked[1804];
  assign N777 = N776 | data_masked[1868];
  assign N776 = N775 | data_masked[1932];
  assign N775 = N774 | data_masked[1996];
  assign N774 = N773 | data_masked[2060];
  assign N773 = N772 | data_masked[2124];
  assign N772 = N771 | data_masked[2188];
  assign N771 = N770 | data_masked[2252];
  assign N770 = N769 | data_masked[2316];
  assign N769 = N768 | data_masked[2380];
  assign N768 = N767 | data_masked[2444];
  assign N767 = N766 | data_masked[2508];
  assign N766 = N765 | data_masked[2572];
  assign N765 = N764 | data_masked[2636];
  assign N764 = N763 | data_masked[2700];
  assign N763 = N762 | data_masked[2764];
  assign N762 = N761 | data_masked[2828];
  assign N761 = N760 | data_masked[2892];
  assign N760 = N759 | data_masked[2956];
  assign N759 = N758 | data_masked[3020];
  assign N758 = N757 | data_masked[3084];
  assign N757 = N756 | data_masked[3148];
  assign N756 = N755 | data_masked[3212];
  assign N755 = N754 | data_masked[3276];
  assign N754 = N753 | data_masked[3340];
  assign N753 = N752 | data_masked[3404];
  assign N752 = N751 | data_masked[3468];
  assign N751 = N750 | data_masked[3532];
  assign N750 = N749 | data_masked[3596];
  assign N749 = N748 | data_masked[3660];
  assign N748 = N747 | data_masked[3724];
  assign N747 = N746 | data_masked[3788];
  assign N746 = N745 | data_masked[3852];
  assign N745 = N744 | data_masked[3916];
  assign N744 = data_masked[4044] | data_masked[3980];
  assign data_o[13] = N867 | data_masked[13];
  assign N867 = N866 | data_masked[77];
  assign N866 = N865 | data_masked[141];
  assign N865 = N864 | data_masked[205];
  assign N864 = N863 | data_masked[269];
  assign N863 = N862 | data_masked[333];
  assign N862 = N861 | data_masked[397];
  assign N861 = N860 | data_masked[461];
  assign N860 = N859 | data_masked[525];
  assign N859 = N858 | data_masked[589];
  assign N858 = N857 | data_masked[653];
  assign N857 = N856 | data_masked[717];
  assign N856 = N855 | data_masked[781];
  assign N855 = N854 | data_masked[845];
  assign N854 = N853 | data_masked[909];
  assign N853 = N852 | data_masked[973];
  assign N852 = N851 | data_masked[1037];
  assign N851 = N850 | data_masked[1101];
  assign N850 = N849 | data_masked[1165];
  assign N849 = N848 | data_masked[1229];
  assign N848 = N847 | data_masked[1293];
  assign N847 = N846 | data_masked[1357];
  assign N846 = N845 | data_masked[1421];
  assign N845 = N844 | data_masked[1485];
  assign N844 = N843 | data_masked[1549];
  assign N843 = N842 | data_masked[1613];
  assign N842 = N841 | data_masked[1677];
  assign N841 = N840 | data_masked[1741];
  assign N840 = N839 | data_masked[1805];
  assign N839 = N838 | data_masked[1869];
  assign N838 = N837 | data_masked[1933];
  assign N837 = N836 | data_masked[1997];
  assign N836 = N835 | data_masked[2061];
  assign N835 = N834 | data_masked[2125];
  assign N834 = N833 | data_masked[2189];
  assign N833 = N832 | data_masked[2253];
  assign N832 = N831 | data_masked[2317];
  assign N831 = N830 | data_masked[2381];
  assign N830 = N829 | data_masked[2445];
  assign N829 = N828 | data_masked[2509];
  assign N828 = N827 | data_masked[2573];
  assign N827 = N826 | data_masked[2637];
  assign N826 = N825 | data_masked[2701];
  assign N825 = N824 | data_masked[2765];
  assign N824 = N823 | data_masked[2829];
  assign N823 = N822 | data_masked[2893];
  assign N822 = N821 | data_masked[2957];
  assign N821 = N820 | data_masked[3021];
  assign N820 = N819 | data_masked[3085];
  assign N819 = N818 | data_masked[3149];
  assign N818 = N817 | data_masked[3213];
  assign N817 = N816 | data_masked[3277];
  assign N816 = N815 | data_masked[3341];
  assign N815 = N814 | data_masked[3405];
  assign N814 = N813 | data_masked[3469];
  assign N813 = N812 | data_masked[3533];
  assign N812 = N811 | data_masked[3597];
  assign N811 = N810 | data_masked[3661];
  assign N810 = N809 | data_masked[3725];
  assign N809 = N808 | data_masked[3789];
  assign N808 = N807 | data_masked[3853];
  assign N807 = N806 | data_masked[3917];
  assign N806 = data_masked[4045] | data_masked[3981];
  assign data_o[14] = N929 | data_masked[14];
  assign N929 = N928 | data_masked[78];
  assign N928 = N927 | data_masked[142];
  assign N927 = N926 | data_masked[206];
  assign N926 = N925 | data_masked[270];
  assign N925 = N924 | data_masked[334];
  assign N924 = N923 | data_masked[398];
  assign N923 = N922 | data_masked[462];
  assign N922 = N921 | data_masked[526];
  assign N921 = N920 | data_masked[590];
  assign N920 = N919 | data_masked[654];
  assign N919 = N918 | data_masked[718];
  assign N918 = N917 | data_masked[782];
  assign N917 = N916 | data_masked[846];
  assign N916 = N915 | data_masked[910];
  assign N915 = N914 | data_masked[974];
  assign N914 = N913 | data_masked[1038];
  assign N913 = N912 | data_masked[1102];
  assign N912 = N911 | data_masked[1166];
  assign N911 = N910 | data_masked[1230];
  assign N910 = N909 | data_masked[1294];
  assign N909 = N908 | data_masked[1358];
  assign N908 = N907 | data_masked[1422];
  assign N907 = N906 | data_masked[1486];
  assign N906 = N905 | data_masked[1550];
  assign N905 = N904 | data_masked[1614];
  assign N904 = N903 | data_masked[1678];
  assign N903 = N902 | data_masked[1742];
  assign N902 = N901 | data_masked[1806];
  assign N901 = N900 | data_masked[1870];
  assign N900 = N899 | data_masked[1934];
  assign N899 = N898 | data_masked[1998];
  assign N898 = N897 | data_masked[2062];
  assign N897 = N896 | data_masked[2126];
  assign N896 = N895 | data_masked[2190];
  assign N895 = N894 | data_masked[2254];
  assign N894 = N893 | data_masked[2318];
  assign N893 = N892 | data_masked[2382];
  assign N892 = N891 | data_masked[2446];
  assign N891 = N890 | data_masked[2510];
  assign N890 = N889 | data_masked[2574];
  assign N889 = N888 | data_masked[2638];
  assign N888 = N887 | data_masked[2702];
  assign N887 = N886 | data_masked[2766];
  assign N886 = N885 | data_masked[2830];
  assign N885 = N884 | data_masked[2894];
  assign N884 = N883 | data_masked[2958];
  assign N883 = N882 | data_masked[3022];
  assign N882 = N881 | data_masked[3086];
  assign N881 = N880 | data_masked[3150];
  assign N880 = N879 | data_masked[3214];
  assign N879 = N878 | data_masked[3278];
  assign N878 = N877 | data_masked[3342];
  assign N877 = N876 | data_masked[3406];
  assign N876 = N875 | data_masked[3470];
  assign N875 = N874 | data_masked[3534];
  assign N874 = N873 | data_masked[3598];
  assign N873 = N872 | data_masked[3662];
  assign N872 = N871 | data_masked[3726];
  assign N871 = N870 | data_masked[3790];
  assign N870 = N869 | data_masked[3854];
  assign N869 = N868 | data_masked[3918];
  assign N868 = data_masked[4046] | data_masked[3982];
  assign data_o[15] = N991 | data_masked[15];
  assign N991 = N990 | data_masked[79];
  assign N990 = N989 | data_masked[143];
  assign N989 = N988 | data_masked[207];
  assign N988 = N987 | data_masked[271];
  assign N987 = N986 | data_masked[335];
  assign N986 = N985 | data_masked[399];
  assign N985 = N984 | data_masked[463];
  assign N984 = N983 | data_masked[527];
  assign N983 = N982 | data_masked[591];
  assign N982 = N981 | data_masked[655];
  assign N981 = N980 | data_masked[719];
  assign N980 = N979 | data_masked[783];
  assign N979 = N978 | data_masked[847];
  assign N978 = N977 | data_masked[911];
  assign N977 = N976 | data_masked[975];
  assign N976 = N975 | data_masked[1039];
  assign N975 = N974 | data_masked[1103];
  assign N974 = N973 | data_masked[1167];
  assign N973 = N972 | data_masked[1231];
  assign N972 = N971 | data_masked[1295];
  assign N971 = N970 | data_masked[1359];
  assign N970 = N969 | data_masked[1423];
  assign N969 = N968 | data_masked[1487];
  assign N968 = N967 | data_masked[1551];
  assign N967 = N966 | data_masked[1615];
  assign N966 = N965 | data_masked[1679];
  assign N965 = N964 | data_masked[1743];
  assign N964 = N963 | data_masked[1807];
  assign N963 = N962 | data_masked[1871];
  assign N962 = N961 | data_masked[1935];
  assign N961 = N960 | data_masked[1999];
  assign N960 = N959 | data_masked[2063];
  assign N959 = N958 | data_masked[2127];
  assign N958 = N957 | data_masked[2191];
  assign N957 = N956 | data_masked[2255];
  assign N956 = N955 | data_masked[2319];
  assign N955 = N954 | data_masked[2383];
  assign N954 = N953 | data_masked[2447];
  assign N953 = N952 | data_masked[2511];
  assign N952 = N951 | data_masked[2575];
  assign N951 = N950 | data_masked[2639];
  assign N950 = N949 | data_masked[2703];
  assign N949 = N948 | data_masked[2767];
  assign N948 = N947 | data_masked[2831];
  assign N947 = N946 | data_masked[2895];
  assign N946 = N945 | data_masked[2959];
  assign N945 = N944 | data_masked[3023];
  assign N944 = N943 | data_masked[3087];
  assign N943 = N942 | data_masked[3151];
  assign N942 = N941 | data_masked[3215];
  assign N941 = N940 | data_masked[3279];
  assign N940 = N939 | data_masked[3343];
  assign N939 = N938 | data_masked[3407];
  assign N938 = N937 | data_masked[3471];
  assign N937 = N936 | data_masked[3535];
  assign N936 = N935 | data_masked[3599];
  assign N935 = N934 | data_masked[3663];
  assign N934 = N933 | data_masked[3727];
  assign N933 = N932 | data_masked[3791];
  assign N932 = N931 | data_masked[3855];
  assign N931 = N930 | data_masked[3919];
  assign N930 = data_masked[4047] | data_masked[3983];
  assign data_o[16] = N1053 | data_masked[16];
  assign N1053 = N1052 | data_masked[80];
  assign N1052 = N1051 | data_masked[144];
  assign N1051 = N1050 | data_masked[208];
  assign N1050 = N1049 | data_masked[272];
  assign N1049 = N1048 | data_masked[336];
  assign N1048 = N1047 | data_masked[400];
  assign N1047 = N1046 | data_masked[464];
  assign N1046 = N1045 | data_masked[528];
  assign N1045 = N1044 | data_masked[592];
  assign N1044 = N1043 | data_masked[656];
  assign N1043 = N1042 | data_masked[720];
  assign N1042 = N1041 | data_masked[784];
  assign N1041 = N1040 | data_masked[848];
  assign N1040 = N1039 | data_masked[912];
  assign N1039 = N1038 | data_masked[976];
  assign N1038 = N1037 | data_masked[1040];
  assign N1037 = N1036 | data_masked[1104];
  assign N1036 = N1035 | data_masked[1168];
  assign N1035 = N1034 | data_masked[1232];
  assign N1034 = N1033 | data_masked[1296];
  assign N1033 = N1032 | data_masked[1360];
  assign N1032 = N1031 | data_masked[1424];
  assign N1031 = N1030 | data_masked[1488];
  assign N1030 = N1029 | data_masked[1552];
  assign N1029 = N1028 | data_masked[1616];
  assign N1028 = N1027 | data_masked[1680];
  assign N1027 = N1026 | data_masked[1744];
  assign N1026 = N1025 | data_masked[1808];
  assign N1025 = N1024 | data_masked[1872];
  assign N1024 = N1023 | data_masked[1936];
  assign N1023 = N1022 | data_masked[2000];
  assign N1022 = N1021 | data_masked[2064];
  assign N1021 = N1020 | data_masked[2128];
  assign N1020 = N1019 | data_masked[2192];
  assign N1019 = N1018 | data_masked[2256];
  assign N1018 = N1017 | data_masked[2320];
  assign N1017 = N1016 | data_masked[2384];
  assign N1016 = N1015 | data_masked[2448];
  assign N1015 = N1014 | data_masked[2512];
  assign N1014 = N1013 | data_masked[2576];
  assign N1013 = N1012 | data_masked[2640];
  assign N1012 = N1011 | data_masked[2704];
  assign N1011 = N1010 | data_masked[2768];
  assign N1010 = N1009 | data_masked[2832];
  assign N1009 = N1008 | data_masked[2896];
  assign N1008 = N1007 | data_masked[2960];
  assign N1007 = N1006 | data_masked[3024];
  assign N1006 = N1005 | data_masked[3088];
  assign N1005 = N1004 | data_masked[3152];
  assign N1004 = N1003 | data_masked[3216];
  assign N1003 = N1002 | data_masked[3280];
  assign N1002 = N1001 | data_masked[3344];
  assign N1001 = N1000 | data_masked[3408];
  assign N1000 = N999 | data_masked[3472];
  assign N999 = N998 | data_masked[3536];
  assign N998 = N997 | data_masked[3600];
  assign N997 = N996 | data_masked[3664];
  assign N996 = N995 | data_masked[3728];
  assign N995 = N994 | data_masked[3792];
  assign N994 = N993 | data_masked[3856];
  assign N993 = N992 | data_masked[3920];
  assign N992 = data_masked[4048] | data_masked[3984];
  assign data_o[17] = N1115 | data_masked[17];
  assign N1115 = N1114 | data_masked[81];
  assign N1114 = N1113 | data_masked[145];
  assign N1113 = N1112 | data_masked[209];
  assign N1112 = N1111 | data_masked[273];
  assign N1111 = N1110 | data_masked[337];
  assign N1110 = N1109 | data_masked[401];
  assign N1109 = N1108 | data_masked[465];
  assign N1108 = N1107 | data_masked[529];
  assign N1107 = N1106 | data_masked[593];
  assign N1106 = N1105 | data_masked[657];
  assign N1105 = N1104 | data_masked[721];
  assign N1104 = N1103 | data_masked[785];
  assign N1103 = N1102 | data_masked[849];
  assign N1102 = N1101 | data_masked[913];
  assign N1101 = N1100 | data_masked[977];
  assign N1100 = N1099 | data_masked[1041];
  assign N1099 = N1098 | data_masked[1105];
  assign N1098 = N1097 | data_masked[1169];
  assign N1097 = N1096 | data_masked[1233];
  assign N1096 = N1095 | data_masked[1297];
  assign N1095 = N1094 | data_masked[1361];
  assign N1094 = N1093 | data_masked[1425];
  assign N1093 = N1092 | data_masked[1489];
  assign N1092 = N1091 | data_masked[1553];
  assign N1091 = N1090 | data_masked[1617];
  assign N1090 = N1089 | data_masked[1681];
  assign N1089 = N1088 | data_masked[1745];
  assign N1088 = N1087 | data_masked[1809];
  assign N1087 = N1086 | data_masked[1873];
  assign N1086 = N1085 | data_masked[1937];
  assign N1085 = N1084 | data_masked[2001];
  assign N1084 = N1083 | data_masked[2065];
  assign N1083 = N1082 | data_masked[2129];
  assign N1082 = N1081 | data_masked[2193];
  assign N1081 = N1080 | data_masked[2257];
  assign N1080 = N1079 | data_masked[2321];
  assign N1079 = N1078 | data_masked[2385];
  assign N1078 = N1077 | data_masked[2449];
  assign N1077 = N1076 | data_masked[2513];
  assign N1076 = N1075 | data_masked[2577];
  assign N1075 = N1074 | data_masked[2641];
  assign N1074 = N1073 | data_masked[2705];
  assign N1073 = N1072 | data_masked[2769];
  assign N1072 = N1071 | data_masked[2833];
  assign N1071 = N1070 | data_masked[2897];
  assign N1070 = N1069 | data_masked[2961];
  assign N1069 = N1068 | data_masked[3025];
  assign N1068 = N1067 | data_masked[3089];
  assign N1067 = N1066 | data_masked[3153];
  assign N1066 = N1065 | data_masked[3217];
  assign N1065 = N1064 | data_masked[3281];
  assign N1064 = N1063 | data_masked[3345];
  assign N1063 = N1062 | data_masked[3409];
  assign N1062 = N1061 | data_masked[3473];
  assign N1061 = N1060 | data_masked[3537];
  assign N1060 = N1059 | data_masked[3601];
  assign N1059 = N1058 | data_masked[3665];
  assign N1058 = N1057 | data_masked[3729];
  assign N1057 = N1056 | data_masked[3793];
  assign N1056 = N1055 | data_masked[3857];
  assign N1055 = N1054 | data_masked[3921];
  assign N1054 = data_masked[4049] | data_masked[3985];
  assign data_o[18] = N1177 | data_masked[18];
  assign N1177 = N1176 | data_masked[82];
  assign N1176 = N1175 | data_masked[146];
  assign N1175 = N1174 | data_masked[210];
  assign N1174 = N1173 | data_masked[274];
  assign N1173 = N1172 | data_masked[338];
  assign N1172 = N1171 | data_masked[402];
  assign N1171 = N1170 | data_masked[466];
  assign N1170 = N1169 | data_masked[530];
  assign N1169 = N1168 | data_masked[594];
  assign N1168 = N1167 | data_masked[658];
  assign N1167 = N1166 | data_masked[722];
  assign N1166 = N1165 | data_masked[786];
  assign N1165 = N1164 | data_masked[850];
  assign N1164 = N1163 | data_masked[914];
  assign N1163 = N1162 | data_masked[978];
  assign N1162 = N1161 | data_masked[1042];
  assign N1161 = N1160 | data_masked[1106];
  assign N1160 = N1159 | data_masked[1170];
  assign N1159 = N1158 | data_masked[1234];
  assign N1158 = N1157 | data_masked[1298];
  assign N1157 = N1156 | data_masked[1362];
  assign N1156 = N1155 | data_masked[1426];
  assign N1155 = N1154 | data_masked[1490];
  assign N1154 = N1153 | data_masked[1554];
  assign N1153 = N1152 | data_masked[1618];
  assign N1152 = N1151 | data_masked[1682];
  assign N1151 = N1150 | data_masked[1746];
  assign N1150 = N1149 | data_masked[1810];
  assign N1149 = N1148 | data_masked[1874];
  assign N1148 = N1147 | data_masked[1938];
  assign N1147 = N1146 | data_masked[2002];
  assign N1146 = N1145 | data_masked[2066];
  assign N1145 = N1144 | data_masked[2130];
  assign N1144 = N1143 | data_masked[2194];
  assign N1143 = N1142 | data_masked[2258];
  assign N1142 = N1141 | data_masked[2322];
  assign N1141 = N1140 | data_masked[2386];
  assign N1140 = N1139 | data_masked[2450];
  assign N1139 = N1138 | data_masked[2514];
  assign N1138 = N1137 | data_masked[2578];
  assign N1137 = N1136 | data_masked[2642];
  assign N1136 = N1135 | data_masked[2706];
  assign N1135 = N1134 | data_masked[2770];
  assign N1134 = N1133 | data_masked[2834];
  assign N1133 = N1132 | data_masked[2898];
  assign N1132 = N1131 | data_masked[2962];
  assign N1131 = N1130 | data_masked[3026];
  assign N1130 = N1129 | data_masked[3090];
  assign N1129 = N1128 | data_masked[3154];
  assign N1128 = N1127 | data_masked[3218];
  assign N1127 = N1126 | data_masked[3282];
  assign N1126 = N1125 | data_masked[3346];
  assign N1125 = N1124 | data_masked[3410];
  assign N1124 = N1123 | data_masked[3474];
  assign N1123 = N1122 | data_masked[3538];
  assign N1122 = N1121 | data_masked[3602];
  assign N1121 = N1120 | data_masked[3666];
  assign N1120 = N1119 | data_masked[3730];
  assign N1119 = N1118 | data_masked[3794];
  assign N1118 = N1117 | data_masked[3858];
  assign N1117 = N1116 | data_masked[3922];
  assign N1116 = data_masked[4050] | data_masked[3986];
  assign data_o[19] = N1239 | data_masked[19];
  assign N1239 = N1238 | data_masked[83];
  assign N1238 = N1237 | data_masked[147];
  assign N1237 = N1236 | data_masked[211];
  assign N1236 = N1235 | data_masked[275];
  assign N1235 = N1234 | data_masked[339];
  assign N1234 = N1233 | data_masked[403];
  assign N1233 = N1232 | data_masked[467];
  assign N1232 = N1231 | data_masked[531];
  assign N1231 = N1230 | data_masked[595];
  assign N1230 = N1229 | data_masked[659];
  assign N1229 = N1228 | data_masked[723];
  assign N1228 = N1227 | data_masked[787];
  assign N1227 = N1226 | data_masked[851];
  assign N1226 = N1225 | data_masked[915];
  assign N1225 = N1224 | data_masked[979];
  assign N1224 = N1223 | data_masked[1043];
  assign N1223 = N1222 | data_masked[1107];
  assign N1222 = N1221 | data_masked[1171];
  assign N1221 = N1220 | data_masked[1235];
  assign N1220 = N1219 | data_masked[1299];
  assign N1219 = N1218 | data_masked[1363];
  assign N1218 = N1217 | data_masked[1427];
  assign N1217 = N1216 | data_masked[1491];
  assign N1216 = N1215 | data_masked[1555];
  assign N1215 = N1214 | data_masked[1619];
  assign N1214 = N1213 | data_masked[1683];
  assign N1213 = N1212 | data_masked[1747];
  assign N1212 = N1211 | data_masked[1811];
  assign N1211 = N1210 | data_masked[1875];
  assign N1210 = N1209 | data_masked[1939];
  assign N1209 = N1208 | data_masked[2003];
  assign N1208 = N1207 | data_masked[2067];
  assign N1207 = N1206 | data_masked[2131];
  assign N1206 = N1205 | data_masked[2195];
  assign N1205 = N1204 | data_masked[2259];
  assign N1204 = N1203 | data_masked[2323];
  assign N1203 = N1202 | data_masked[2387];
  assign N1202 = N1201 | data_masked[2451];
  assign N1201 = N1200 | data_masked[2515];
  assign N1200 = N1199 | data_masked[2579];
  assign N1199 = N1198 | data_masked[2643];
  assign N1198 = N1197 | data_masked[2707];
  assign N1197 = N1196 | data_masked[2771];
  assign N1196 = N1195 | data_masked[2835];
  assign N1195 = N1194 | data_masked[2899];
  assign N1194 = N1193 | data_masked[2963];
  assign N1193 = N1192 | data_masked[3027];
  assign N1192 = N1191 | data_masked[3091];
  assign N1191 = N1190 | data_masked[3155];
  assign N1190 = N1189 | data_masked[3219];
  assign N1189 = N1188 | data_masked[3283];
  assign N1188 = N1187 | data_masked[3347];
  assign N1187 = N1186 | data_masked[3411];
  assign N1186 = N1185 | data_masked[3475];
  assign N1185 = N1184 | data_masked[3539];
  assign N1184 = N1183 | data_masked[3603];
  assign N1183 = N1182 | data_masked[3667];
  assign N1182 = N1181 | data_masked[3731];
  assign N1181 = N1180 | data_masked[3795];
  assign N1180 = N1179 | data_masked[3859];
  assign N1179 = N1178 | data_masked[3923];
  assign N1178 = data_masked[4051] | data_masked[3987];
  assign data_o[20] = N1301 | data_masked[20];
  assign N1301 = N1300 | data_masked[84];
  assign N1300 = N1299 | data_masked[148];
  assign N1299 = N1298 | data_masked[212];
  assign N1298 = N1297 | data_masked[276];
  assign N1297 = N1296 | data_masked[340];
  assign N1296 = N1295 | data_masked[404];
  assign N1295 = N1294 | data_masked[468];
  assign N1294 = N1293 | data_masked[532];
  assign N1293 = N1292 | data_masked[596];
  assign N1292 = N1291 | data_masked[660];
  assign N1291 = N1290 | data_masked[724];
  assign N1290 = N1289 | data_masked[788];
  assign N1289 = N1288 | data_masked[852];
  assign N1288 = N1287 | data_masked[916];
  assign N1287 = N1286 | data_masked[980];
  assign N1286 = N1285 | data_masked[1044];
  assign N1285 = N1284 | data_masked[1108];
  assign N1284 = N1283 | data_masked[1172];
  assign N1283 = N1282 | data_masked[1236];
  assign N1282 = N1281 | data_masked[1300];
  assign N1281 = N1280 | data_masked[1364];
  assign N1280 = N1279 | data_masked[1428];
  assign N1279 = N1278 | data_masked[1492];
  assign N1278 = N1277 | data_masked[1556];
  assign N1277 = N1276 | data_masked[1620];
  assign N1276 = N1275 | data_masked[1684];
  assign N1275 = N1274 | data_masked[1748];
  assign N1274 = N1273 | data_masked[1812];
  assign N1273 = N1272 | data_masked[1876];
  assign N1272 = N1271 | data_masked[1940];
  assign N1271 = N1270 | data_masked[2004];
  assign N1270 = N1269 | data_masked[2068];
  assign N1269 = N1268 | data_masked[2132];
  assign N1268 = N1267 | data_masked[2196];
  assign N1267 = N1266 | data_masked[2260];
  assign N1266 = N1265 | data_masked[2324];
  assign N1265 = N1264 | data_masked[2388];
  assign N1264 = N1263 | data_masked[2452];
  assign N1263 = N1262 | data_masked[2516];
  assign N1262 = N1261 | data_masked[2580];
  assign N1261 = N1260 | data_masked[2644];
  assign N1260 = N1259 | data_masked[2708];
  assign N1259 = N1258 | data_masked[2772];
  assign N1258 = N1257 | data_masked[2836];
  assign N1257 = N1256 | data_masked[2900];
  assign N1256 = N1255 | data_masked[2964];
  assign N1255 = N1254 | data_masked[3028];
  assign N1254 = N1253 | data_masked[3092];
  assign N1253 = N1252 | data_masked[3156];
  assign N1252 = N1251 | data_masked[3220];
  assign N1251 = N1250 | data_masked[3284];
  assign N1250 = N1249 | data_masked[3348];
  assign N1249 = N1248 | data_masked[3412];
  assign N1248 = N1247 | data_masked[3476];
  assign N1247 = N1246 | data_masked[3540];
  assign N1246 = N1245 | data_masked[3604];
  assign N1245 = N1244 | data_masked[3668];
  assign N1244 = N1243 | data_masked[3732];
  assign N1243 = N1242 | data_masked[3796];
  assign N1242 = N1241 | data_masked[3860];
  assign N1241 = N1240 | data_masked[3924];
  assign N1240 = data_masked[4052] | data_masked[3988];
  assign data_o[21] = N1363 | data_masked[21];
  assign N1363 = N1362 | data_masked[85];
  assign N1362 = N1361 | data_masked[149];
  assign N1361 = N1360 | data_masked[213];
  assign N1360 = N1359 | data_masked[277];
  assign N1359 = N1358 | data_masked[341];
  assign N1358 = N1357 | data_masked[405];
  assign N1357 = N1356 | data_masked[469];
  assign N1356 = N1355 | data_masked[533];
  assign N1355 = N1354 | data_masked[597];
  assign N1354 = N1353 | data_masked[661];
  assign N1353 = N1352 | data_masked[725];
  assign N1352 = N1351 | data_masked[789];
  assign N1351 = N1350 | data_masked[853];
  assign N1350 = N1349 | data_masked[917];
  assign N1349 = N1348 | data_masked[981];
  assign N1348 = N1347 | data_masked[1045];
  assign N1347 = N1346 | data_masked[1109];
  assign N1346 = N1345 | data_masked[1173];
  assign N1345 = N1344 | data_masked[1237];
  assign N1344 = N1343 | data_masked[1301];
  assign N1343 = N1342 | data_masked[1365];
  assign N1342 = N1341 | data_masked[1429];
  assign N1341 = N1340 | data_masked[1493];
  assign N1340 = N1339 | data_masked[1557];
  assign N1339 = N1338 | data_masked[1621];
  assign N1338 = N1337 | data_masked[1685];
  assign N1337 = N1336 | data_masked[1749];
  assign N1336 = N1335 | data_masked[1813];
  assign N1335 = N1334 | data_masked[1877];
  assign N1334 = N1333 | data_masked[1941];
  assign N1333 = N1332 | data_masked[2005];
  assign N1332 = N1331 | data_masked[2069];
  assign N1331 = N1330 | data_masked[2133];
  assign N1330 = N1329 | data_masked[2197];
  assign N1329 = N1328 | data_masked[2261];
  assign N1328 = N1327 | data_masked[2325];
  assign N1327 = N1326 | data_masked[2389];
  assign N1326 = N1325 | data_masked[2453];
  assign N1325 = N1324 | data_masked[2517];
  assign N1324 = N1323 | data_masked[2581];
  assign N1323 = N1322 | data_masked[2645];
  assign N1322 = N1321 | data_masked[2709];
  assign N1321 = N1320 | data_masked[2773];
  assign N1320 = N1319 | data_masked[2837];
  assign N1319 = N1318 | data_masked[2901];
  assign N1318 = N1317 | data_masked[2965];
  assign N1317 = N1316 | data_masked[3029];
  assign N1316 = N1315 | data_masked[3093];
  assign N1315 = N1314 | data_masked[3157];
  assign N1314 = N1313 | data_masked[3221];
  assign N1313 = N1312 | data_masked[3285];
  assign N1312 = N1311 | data_masked[3349];
  assign N1311 = N1310 | data_masked[3413];
  assign N1310 = N1309 | data_masked[3477];
  assign N1309 = N1308 | data_masked[3541];
  assign N1308 = N1307 | data_masked[3605];
  assign N1307 = N1306 | data_masked[3669];
  assign N1306 = N1305 | data_masked[3733];
  assign N1305 = N1304 | data_masked[3797];
  assign N1304 = N1303 | data_masked[3861];
  assign N1303 = N1302 | data_masked[3925];
  assign N1302 = data_masked[4053] | data_masked[3989];
  assign data_o[22] = N1425 | data_masked[22];
  assign N1425 = N1424 | data_masked[86];
  assign N1424 = N1423 | data_masked[150];
  assign N1423 = N1422 | data_masked[214];
  assign N1422 = N1421 | data_masked[278];
  assign N1421 = N1420 | data_masked[342];
  assign N1420 = N1419 | data_masked[406];
  assign N1419 = N1418 | data_masked[470];
  assign N1418 = N1417 | data_masked[534];
  assign N1417 = N1416 | data_masked[598];
  assign N1416 = N1415 | data_masked[662];
  assign N1415 = N1414 | data_masked[726];
  assign N1414 = N1413 | data_masked[790];
  assign N1413 = N1412 | data_masked[854];
  assign N1412 = N1411 | data_masked[918];
  assign N1411 = N1410 | data_masked[982];
  assign N1410 = N1409 | data_masked[1046];
  assign N1409 = N1408 | data_masked[1110];
  assign N1408 = N1407 | data_masked[1174];
  assign N1407 = N1406 | data_masked[1238];
  assign N1406 = N1405 | data_masked[1302];
  assign N1405 = N1404 | data_masked[1366];
  assign N1404 = N1403 | data_masked[1430];
  assign N1403 = N1402 | data_masked[1494];
  assign N1402 = N1401 | data_masked[1558];
  assign N1401 = N1400 | data_masked[1622];
  assign N1400 = N1399 | data_masked[1686];
  assign N1399 = N1398 | data_masked[1750];
  assign N1398 = N1397 | data_masked[1814];
  assign N1397 = N1396 | data_masked[1878];
  assign N1396 = N1395 | data_masked[1942];
  assign N1395 = N1394 | data_masked[2006];
  assign N1394 = N1393 | data_masked[2070];
  assign N1393 = N1392 | data_masked[2134];
  assign N1392 = N1391 | data_masked[2198];
  assign N1391 = N1390 | data_masked[2262];
  assign N1390 = N1389 | data_masked[2326];
  assign N1389 = N1388 | data_masked[2390];
  assign N1388 = N1387 | data_masked[2454];
  assign N1387 = N1386 | data_masked[2518];
  assign N1386 = N1385 | data_masked[2582];
  assign N1385 = N1384 | data_masked[2646];
  assign N1384 = N1383 | data_masked[2710];
  assign N1383 = N1382 | data_masked[2774];
  assign N1382 = N1381 | data_masked[2838];
  assign N1381 = N1380 | data_masked[2902];
  assign N1380 = N1379 | data_masked[2966];
  assign N1379 = N1378 | data_masked[3030];
  assign N1378 = N1377 | data_masked[3094];
  assign N1377 = N1376 | data_masked[3158];
  assign N1376 = N1375 | data_masked[3222];
  assign N1375 = N1374 | data_masked[3286];
  assign N1374 = N1373 | data_masked[3350];
  assign N1373 = N1372 | data_masked[3414];
  assign N1372 = N1371 | data_masked[3478];
  assign N1371 = N1370 | data_masked[3542];
  assign N1370 = N1369 | data_masked[3606];
  assign N1369 = N1368 | data_masked[3670];
  assign N1368 = N1367 | data_masked[3734];
  assign N1367 = N1366 | data_masked[3798];
  assign N1366 = N1365 | data_masked[3862];
  assign N1365 = N1364 | data_masked[3926];
  assign N1364 = data_masked[4054] | data_masked[3990];
  assign data_o[23] = N1487 | data_masked[23];
  assign N1487 = N1486 | data_masked[87];
  assign N1486 = N1485 | data_masked[151];
  assign N1485 = N1484 | data_masked[215];
  assign N1484 = N1483 | data_masked[279];
  assign N1483 = N1482 | data_masked[343];
  assign N1482 = N1481 | data_masked[407];
  assign N1481 = N1480 | data_masked[471];
  assign N1480 = N1479 | data_masked[535];
  assign N1479 = N1478 | data_masked[599];
  assign N1478 = N1477 | data_masked[663];
  assign N1477 = N1476 | data_masked[727];
  assign N1476 = N1475 | data_masked[791];
  assign N1475 = N1474 | data_masked[855];
  assign N1474 = N1473 | data_masked[919];
  assign N1473 = N1472 | data_masked[983];
  assign N1472 = N1471 | data_masked[1047];
  assign N1471 = N1470 | data_masked[1111];
  assign N1470 = N1469 | data_masked[1175];
  assign N1469 = N1468 | data_masked[1239];
  assign N1468 = N1467 | data_masked[1303];
  assign N1467 = N1466 | data_masked[1367];
  assign N1466 = N1465 | data_masked[1431];
  assign N1465 = N1464 | data_masked[1495];
  assign N1464 = N1463 | data_masked[1559];
  assign N1463 = N1462 | data_masked[1623];
  assign N1462 = N1461 | data_masked[1687];
  assign N1461 = N1460 | data_masked[1751];
  assign N1460 = N1459 | data_masked[1815];
  assign N1459 = N1458 | data_masked[1879];
  assign N1458 = N1457 | data_masked[1943];
  assign N1457 = N1456 | data_masked[2007];
  assign N1456 = N1455 | data_masked[2071];
  assign N1455 = N1454 | data_masked[2135];
  assign N1454 = N1453 | data_masked[2199];
  assign N1453 = N1452 | data_masked[2263];
  assign N1452 = N1451 | data_masked[2327];
  assign N1451 = N1450 | data_masked[2391];
  assign N1450 = N1449 | data_masked[2455];
  assign N1449 = N1448 | data_masked[2519];
  assign N1448 = N1447 | data_masked[2583];
  assign N1447 = N1446 | data_masked[2647];
  assign N1446 = N1445 | data_masked[2711];
  assign N1445 = N1444 | data_masked[2775];
  assign N1444 = N1443 | data_masked[2839];
  assign N1443 = N1442 | data_masked[2903];
  assign N1442 = N1441 | data_masked[2967];
  assign N1441 = N1440 | data_masked[3031];
  assign N1440 = N1439 | data_masked[3095];
  assign N1439 = N1438 | data_masked[3159];
  assign N1438 = N1437 | data_masked[3223];
  assign N1437 = N1436 | data_masked[3287];
  assign N1436 = N1435 | data_masked[3351];
  assign N1435 = N1434 | data_masked[3415];
  assign N1434 = N1433 | data_masked[3479];
  assign N1433 = N1432 | data_masked[3543];
  assign N1432 = N1431 | data_masked[3607];
  assign N1431 = N1430 | data_masked[3671];
  assign N1430 = N1429 | data_masked[3735];
  assign N1429 = N1428 | data_masked[3799];
  assign N1428 = N1427 | data_masked[3863];
  assign N1427 = N1426 | data_masked[3927];
  assign N1426 = data_masked[4055] | data_masked[3991];
  assign data_o[24] = N1549 | data_masked[24];
  assign N1549 = N1548 | data_masked[88];
  assign N1548 = N1547 | data_masked[152];
  assign N1547 = N1546 | data_masked[216];
  assign N1546 = N1545 | data_masked[280];
  assign N1545 = N1544 | data_masked[344];
  assign N1544 = N1543 | data_masked[408];
  assign N1543 = N1542 | data_masked[472];
  assign N1542 = N1541 | data_masked[536];
  assign N1541 = N1540 | data_masked[600];
  assign N1540 = N1539 | data_masked[664];
  assign N1539 = N1538 | data_masked[728];
  assign N1538 = N1537 | data_masked[792];
  assign N1537 = N1536 | data_masked[856];
  assign N1536 = N1535 | data_masked[920];
  assign N1535 = N1534 | data_masked[984];
  assign N1534 = N1533 | data_masked[1048];
  assign N1533 = N1532 | data_masked[1112];
  assign N1532 = N1531 | data_masked[1176];
  assign N1531 = N1530 | data_masked[1240];
  assign N1530 = N1529 | data_masked[1304];
  assign N1529 = N1528 | data_masked[1368];
  assign N1528 = N1527 | data_masked[1432];
  assign N1527 = N1526 | data_masked[1496];
  assign N1526 = N1525 | data_masked[1560];
  assign N1525 = N1524 | data_masked[1624];
  assign N1524 = N1523 | data_masked[1688];
  assign N1523 = N1522 | data_masked[1752];
  assign N1522 = N1521 | data_masked[1816];
  assign N1521 = N1520 | data_masked[1880];
  assign N1520 = N1519 | data_masked[1944];
  assign N1519 = N1518 | data_masked[2008];
  assign N1518 = N1517 | data_masked[2072];
  assign N1517 = N1516 | data_masked[2136];
  assign N1516 = N1515 | data_masked[2200];
  assign N1515 = N1514 | data_masked[2264];
  assign N1514 = N1513 | data_masked[2328];
  assign N1513 = N1512 | data_masked[2392];
  assign N1512 = N1511 | data_masked[2456];
  assign N1511 = N1510 | data_masked[2520];
  assign N1510 = N1509 | data_masked[2584];
  assign N1509 = N1508 | data_masked[2648];
  assign N1508 = N1507 | data_masked[2712];
  assign N1507 = N1506 | data_masked[2776];
  assign N1506 = N1505 | data_masked[2840];
  assign N1505 = N1504 | data_masked[2904];
  assign N1504 = N1503 | data_masked[2968];
  assign N1503 = N1502 | data_masked[3032];
  assign N1502 = N1501 | data_masked[3096];
  assign N1501 = N1500 | data_masked[3160];
  assign N1500 = N1499 | data_masked[3224];
  assign N1499 = N1498 | data_masked[3288];
  assign N1498 = N1497 | data_masked[3352];
  assign N1497 = N1496 | data_masked[3416];
  assign N1496 = N1495 | data_masked[3480];
  assign N1495 = N1494 | data_masked[3544];
  assign N1494 = N1493 | data_masked[3608];
  assign N1493 = N1492 | data_masked[3672];
  assign N1492 = N1491 | data_masked[3736];
  assign N1491 = N1490 | data_masked[3800];
  assign N1490 = N1489 | data_masked[3864];
  assign N1489 = N1488 | data_masked[3928];
  assign N1488 = data_masked[4056] | data_masked[3992];
  assign data_o[25] = N1611 | data_masked[25];
  assign N1611 = N1610 | data_masked[89];
  assign N1610 = N1609 | data_masked[153];
  assign N1609 = N1608 | data_masked[217];
  assign N1608 = N1607 | data_masked[281];
  assign N1607 = N1606 | data_masked[345];
  assign N1606 = N1605 | data_masked[409];
  assign N1605 = N1604 | data_masked[473];
  assign N1604 = N1603 | data_masked[537];
  assign N1603 = N1602 | data_masked[601];
  assign N1602 = N1601 | data_masked[665];
  assign N1601 = N1600 | data_masked[729];
  assign N1600 = N1599 | data_masked[793];
  assign N1599 = N1598 | data_masked[857];
  assign N1598 = N1597 | data_masked[921];
  assign N1597 = N1596 | data_masked[985];
  assign N1596 = N1595 | data_masked[1049];
  assign N1595 = N1594 | data_masked[1113];
  assign N1594 = N1593 | data_masked[1177];
  assign N1593 = N1592 | data_masked[1241];
  assign N1592 = N1591 | data_masked[1305];
  assign N1591 = N1590 | data_masked[1369];
  assign N1590 = N1589 | data_masked[1433];
  assign N1589 = N1588 | data_masked[1497];
  assign N1588 = N1587 | data_masked[1561];
  assign N1587 = N1586 | data_masked[1625];
  assign N1586 = N1585 | data_masked[1689];
  assign N1585 = N1584 | data_masked[1753];
  assign N1584 = N1583 | data_masked[1817];
  assign N1583 = N1582 | data_masked[1881];
  assign N1582 = N1581 | data_masked[1945];
  assign N1581 = N1580 | data_masked[2009];
  assign N1580 = N1579 | data_masked[2073];
  assign N1579 = N1578 | data_masked[2137];
  assign N1578 = N1577 | data_masked[2201];
  assign N1577 = N1576 | data_masked[2265];
  assign N1576 = N1575 | data_masked[2329];
  assign N1575 = N1574 | data_masked[2393];
  assign N1574 = N1573 | data_masked[2457];
  assign N1573 = N1572 | data_masked[2521];
  assign N1572 = N1571 | data_masked[2585];
  assign N1571 = N1570 | data_masked[2649];
  assign N1570 = N1569 | data_masked[2713];
  assign N1569 = N1568 | data_masked[2777];
  assign N1568 = N1567 | data_masked[2841];
  assign N1567 = N1566 | data_masked[2905];
  assign N1566 = N1565 | data_masked[2969];
  assign N1565 = N1564 | data_masked[3033];
  assign N1564 = N1563 | data_masked[3097];
  assign N1563 = N1562 | data_masked[3161];
  assign N1562 = N1561 | data_masked[3225];
  assign N1561 = N1560 | data_masked[3289];
  assign N1560 = N1559 | data_masked[3353];
  assign N1559 = N1558 | data_masked[3417];
  assign N1558 = N1557 | data_masked[3481];
  assign N1557 = N1556 | data_masked[3545];
  assign N1556 = N1555 | data_masked[3609];
  assign N1555 = N1554 | data_masked[3673];
  assign N1554 = N1553 | data_masked[3737];
  assign N1553 = N1552 | data_masked[3801];
  assign N1552 = N1551 | data_masked[3865];
  assign N1551 = N1550 | data_masked[3929];
  assign N1550 = data_masked[4057] | data_masked[3993];
  assign data_o[26] = N1673 | data_masked[26];
  assign N1673 = N1672 | data_masked[90];
  assign N1672 = N1671 | data_masked[154];
  assign N1671 = N1670 | data_masked[218];
  assign N1670 = N1669 | data_masked[282];
  assign N1669 = N1668 | data_masked[346];
  assign N1668 = N1667 | data_masked[410];
  assign N1667 = N1666 | data_masked[474];
  assign N1666 = N1665 | data_masked[538];
  assign N1665 = N1664 | data_masked[602];
  assign N1664 = N1663 | data_masked[666];
  assign N1663 = N1662 | data_masked[730];
  assign N1662 = N1661 | data_masked[794];
  assign N1661 = N1660 | data_masked[858];
  assign N1660 = N1659 | data_masked[922];
  assign N1659 = N1658 | data_masked[986];
  assign N1658 = N1657 | data_masked[1050];
  assign N1657 = N1656 | data_masked[1114];
  assign N1656 = N1655 | data_masked[1178];
  assign N1655 = N1654 | data_masked[1242];
  assign N1654 = N1653 | data_masked[1306];
  assign N1653 = N1652 | data_masked[1370];
  assign N1652 = N1651 | data_masked[1434];
  assign N1651 = N1650 | data_masked[1498];
  assign N1650 = N1649 | data_masked[1562];
  assign N1649 = N1648 | data_masked[1626];
  assign N1648 = N1647 | data_masked[1690];
  assign N1647 = N1646 | data_masked[1754];
  assign N1646 = N1645 | data_masked[1818];
  assign N1645 = N1644 | data_masked[1882];
  assign N1644 = N1643 | data_masked[1946];
  assign N1643 = N1642 | data_masked[2010];
  assign N1642 = N1641 | data_masked[2074];
  assign N1641 = N1640 | data_masked[2138];
  assign N1640 = N1639 | data_masked[2202];
  assign N1639 = N1638 | data_masked[2266];
  assign N1638 = N1637 | data_masked[2330];
  assign N1637 = N1636 | data_masked[2394];
  assign N1636 = N1635 | data_masked[2458];
  assign N1635 = N1634 | data_masked[2522];
  assign N1634 = N1633 | data_masked[2586];
  assign N1633 = N1632 | data_masked[2650];
  assign N1632 = N1631 | data_masked[2714];
  assign N1631 = N1630 | data_masked[2778];
  assign N1630 = N1629 | data_masked[2842];
  assign N1629 = N1628 | data_masked[2906];
  assign N1628 = N1627 | data_masked[2970];
  assign N1627 = N1626 | data_masked[3034];
  assign N1626 = N1625 | data_masked[3098];
  assign N1625 = N1624 | data_masked[3162];
  assign N1624 = N1623 | data_masked[3226];
  assign N1623 = N1622 | data_masked[3290];
  assign N1622 = N1621 | data_masked[3354];
  assign N1621 = N1620 | data_masked[3418];
  assign N1620 = N1619 | data_masked[3482];
  assign N1619 = N1618 | data_masked[3546];
  assign N1618 = N1617 | data_masked[3610];
  assign N1617 = N1616 | data_masked[3674];
  assign N1616 = N1615 | data_masked[3738];
  assign N1615 = N1614 | data_masked[3802];
  assign N1614 = N1613 | data_masked[3866];
  assign N1613 = N1612 | data_masked[3930];
  assign N1612 = data_masked[4058] | data_masked[3994];
  assign data_o[27] = N1735 | data_masked[27];
  assign N1735 = N1734 | data_masked[91];
  assign N1734 = N1733 | data_masked[155];
  assign N1733 = N1732 | data_masked[219];
  assign N1732 = N1731 | data_masked[283];
  assign N1731 = N1730 | data_masked[347];
  assign N1730 = N1729 | data_masked[411];
  assign N1729 = N1728 | data_masked[475];
  assign N1728 = N1727 | data_masked[539];
  assign N1727 = N1726 | data_masked[603];
  assign N1726 = N1725 | data_masked[667];
  assign N1725 = N1724 | data_masked[731];
  assign N1724 = N1723 | data_masked[795];
  assign N1723 = N1722 | data_masked[859];
  assign N1722 = N1721 | data_masked[923];
  assign N1721 = N1720 | data_masked[987];
  assign N1720 = N1719 | data_masked[1051];
  assign N1719 = N1718 | data_masked[1115];
  assign N1718 = N1717 | data_masked[1179];
  assign N1717 = N1716 | data_masked[1243];
  assign N1716 = N1715 | data_masked[1307];
  assign N1715 = N1714 | data_masked[1371];
  assign N1714 = N1713 | data_masked[1435];
  assign N1713 = N1712 | data_masked[1499];
  assign N1712 = N1711 | data_masked[1563];
  assign N1711 = N1710 | data_masked[1627];
  assign N1710 = N1709 | data_masked[1691];
  assign N1709 = N1708 | data_masked[1755];
  assign N1708 = N1707 | data_masked[1819];
  assign N1707 = N1706 | data_masked[1883];
  assign N1706 = N1705 | data_masked[1947];
  assign N1705 = N1704 | data_masked[2011];
  assign N1704 = N1703 | data_masked[2075];
  assign N1703 = N1702 | data_masked[2139];
  assign N1702 = N1701 | data_masked[2203];
  assign N1701 = N1700 | data_masked[2267];
  assign N1700 = N1699 | data_masked[2331];
  assign N1699 = N1698 | data_masked[2395];
  assign N1698 = N1697 | data_masked[2459];
  assign N1697 = N1696 | data_masked[2523];
  assign N1696 = N1695 | data_masked[2587];
  assign N1695 = N1694 | data_masked[2651];
  assign N1694 = N1693 | data_masked[2715];
  assign N1693 = N1692 | data_masked[2779];
  assign N1692 = N1691 | data_masked[2843];
  assign N1691 = N1690 | data_masked[2907];
  assign N1690 = N1689 | data_masked[2971];
  assign N1689 = N1688 | data_masked[3035];
  assign N1688 = N1687 | data_masked[3099];
  assign N1687 = N1686 | data_masked[3163];
  assign N1686 = N1685 | data_masked[3227];
  assign N1685 = N1684 | data_masked[3291];
  assign N1684 = N1683 | data_masked[3355];
  assign N1683 = N1682 | data_masked[3419];
  assign N1682 = N1681 | data_masked[3483];
  assign N1681 = N1680 | data_masked[3547];
  assign N1680 = N1679 | data_masked[3611];
  assign N1679 = N1678 | data_masked[3675];
  assign N1678 = N1677 | data_masked[3739];
  assign N1677 = N1676 | data_masked[3803];
  assign N1676 = N1675 | data_masked[3867];
  assign N1675 = N1674 | data_masked[3931];
  assign N1674 = data_masked[4059] | data_masked[3995];
  assign data_o[28] = N1797 | data_masked[28];
  assign N1797 = N1796 | data_masked[92];
  assign N1796 = N1795 | data_masked[156];
  assign N1795 = N1794 | data_masked[220];
  assign N1794 = N1793 | data_masked[284];
  assign N1793 = N1792 | data_masked[348];
  assign N1792 = N1791 | data_masked[412];
  assign N1791 = N1790 | data_masked[476];
  assign N1790 = N1789 | data_masked[540];
  assign N1789 = N1788 | data_masked[604];
  assign N1788 = N1787 | data_masked[668];
  assign N1787 = N1786 | data_masked[732];
  assign N1786 = N1785 | data_masked[796];
  assign N1785 = N1784 | data_masked[860];
  assign N1784 = N1783 | data_masked[924];
  assign N1783 = N1782 | data_masked[988];
  assign N1782 = N1781 | data_masked[1052];
  assign N1781 = N1780 | data_masked[1116];
  assign N1780 = N1779 | data_masked[1180];
  assign N1779 = N1778 | data_masked[1244];
  assign N1778 = N1777 | data_masked[1308];
  assign N1777 = N1776 | data_masked[1372];
  assign N1776 = N1775 | data_masked[1436];
  assign N1775 = N1774 | data_masked[1500];
  assign N1774 = N1773 | data_masked[1564];
  assign N1773 = N1772 | data_masked[1628];
  assign N1772 = N1771 | data_masked[1692];
  assign N1771 = N1770 | data_masked[1756];
  assign N1770 = N1769 | data_masked[1820];
  assign N1769 = N1768 | data_masked[1884];
  assign N1768 = N1767 | data_masked[1948];
  assign N1767 = N1766 | data_masked[2012];
  assign N1766 = N1765 | data_masked[2076];
  assign N1765 = N1764 | data_masked[2140];
  assign N1764 = N1763 | data_masked[2204];
  assign N1763 = N1762 | data_masked[2268];
  assign N1762 = N1761 | data_masked[2332];
  assign N1761 = N1760 | data_masked[2396];
  assign N1760 = N1759 | data_masked[2460];
  assign N1759 = N1758 | data_masked[2524];
  assign N1758 = N1757 | data_masked[2588];
  assign N1757 = N1756 | data_masked[2652];
  assign N1756 = N1755 | data_masked[2716];
  assign N1755 = N1754 | data_masked[2780];
  assign N1754 = N1753 | data_masked[2844];
  assign N1753 = N1752 | data_masked[2908];
  assign N1752 = N1751 | data_masked[2972];
  assign N1751 = N1750 | data_masked[3036];
  assign N1750 = N1749 | data_masked[3100];
  assign N1749 = N1748 | data_masked[3164];
  assign N1748 = N1747 | data_masked[3228];
  assign N1747 = N1746 | data_masked[3292];
  assign N1746 = N1745 | data_masked[3356];
  assign N1745 = N1744 | data_masked[3420];
  assign N1744 = N1743 | data_masked[3484];
  assign N1743 = N1742 | data_masked[3548];
  assign N1742 = N1741 | data_masked[3612];
  assign N1741 = N1740 | data_masked[3676];
  assign N1740 = N1739 | data_masked[3740];
  assign N1739 = N1738 | data_masked[3804];
  assign N1738 = N1737 | data_masked[3868];
  assign N1737 = N1736 | data_masked[3932];
  assign N1736 = data_masked[4060] | data_masked[3996];
  assign data_o[29] = N1859 | data_masked[29];
  assign N1859 = N1858 | data_masked[93];
  assign N1858 = N1857 | data_masked[157];
  assign N1857 = N1856 | data_masked[221];
  assign N1856 = N1855 | data_masked[285];
  assign N1855 = N1854 | data_masked[349];
  assign N1854 = N1853 | data_masked[413];
  assign N1853 = N1852 | data_masked[477];
  assign N1852 = N1851 | data_masked[541];
  assign N1851 = N1850 | data_masked[605];
  assign N1850 = N1849 | data_masked[669];
  assign N1849 = N1848 | data_masked[733];
  assign N1848 = N1847 | data_masked[797];
  assign N1847 = N1846 | data_masked[861];
  assign N1846 = N1845 | data_masked[925];
  assign N1845 = N1844 | data_masked[989];
  assign N1844 = N1843 | data_masked[1053];
  assign N1843 = N1842 | data_masked[1117];
  assign N1842 = N1841 | data_masked[1181];
  assign N1841 = N1840 | data_masked[1245];
  assign N1840 = N1839 | data_masked[1309];
  assign N1839 = N1838 | data_masked[1373];
  assign N1838 = N1837 | data_masked[1437];
  assign N1837 = N1836 | data_masked[1501];
  assign N1836 = N1835 | data_masked[1565];
  assign N1835 = N1834 | data_masked[1629];
  assign N1834 = N1833 | data_masked[1693];
  assign N1833 = N1832 | data_masked[1757];
  assign N1832 = N1831 | data_masked[1821];
  assign N1831 = N1830 | data_masked[1885];
  assign N1830 = N1829 | data_masked[1949];
  assign N1829 = N1828 | data_masked[2013];
  assign N1828 = N1827 | data_masked[2077];
  assign N1827 = N1826 | data_masked[2141];
  assign N1826 = N1825 | data_masked[2205];
  assign N1825 = N1824 | data_masked[2269];
  assign N1824 = N1823 | data_masked[2333];
  assign N1823 = N1822 | data_masked[2397];
  assign N1822 = N1821 | data_masked[2461];
  assign N1821 = N1820 | data_masked[2525];
  assign N1820 = N1819 | data_masked[2589];
  assign N1819 = N1818 | data_masked[2653];
  assign N1818 = N1817 | data_masked[2717];
  assign N1817 = N1816 | data_masked[2781];
  assign N1816 = N1815 | data_masked[2845];
  assign N1815 = N1814 | data_masked[2909];
  assign N1814 = N1813 | data_masked[2973];
  assign N1813 = N1812 | data_masked[3037];
  assign N1812 = N1811 | data_masked[3101];
  assign N1811 = N1810 | data_masked[3165];
  assign N1810 = N1809 | data_masked[3229];
  assign N1809 = N1808 | data_masked[3293];
  assign N1808 = N1807 | data_masked[3357];
  assign N1807 = N1806 | data_masked[3421];
  assign N1806 = N1805 | data_masked[3485];
  assign N1805 = N1804 | data_masked[3549];
  assign N1804 = N1803 | data_masked[3613];
  assign N1803 = N1802 | data_masked[3677];
  assign N1802 = N1801 | data_masked[3741];
  assign N1801 = N1800 | data_masked[3805];
  assign N1800 = N1799 | data_masked[3869];
  assign N1799 = N1798 | data_masked[3933];
  assign N1798 = data_masked[4061] | data_masked[3997];
  assign data_o[30] = N1921 | data_masked[30];
  assign N1921 = N1920 | data_masked[94];
  assign N1920 = N1919 | data_masked[158];
  assign N1919 = N1918 | data_masked[222];
  assign N1918 = N1917 | data_masked[286];
  assign N1917 = N1916 | data_masked[350];
  assign N1916 = N1915 | data_masked[414];
  assign N1915 = N1914 | data_masked[478];
  assign N1914 = N1913 | data_masked[542];
  assign N1913 = N1912 | data_masked[606];
  assign N1912 = N1911 | data_masked[670];
  assign N1911 = N1910 | data_masked[734];
  assign N1910 = N1909 | data_masked[798];
  assign N1909 = N1908 | data_masked[862];
  assign N1908 = N1907 | data_masked[926];
  assign N1907 = N1906 | data_masked[990];
  assign N1906 = N1905 | data_masked[1054];
  assign N1905 = N1904 | data_masked[1118];
  assign N1904 = N1903 | data_masked[1182];
  assign N1903 = N1902 | data_masked[1246];
  assign N1902 = N1901 | data_masked[1310];
  assign N1901 = N1900 | data_masked[1374];
  assign N1900 = N1899 | data_masked[1438];
  assign N1899 = N1898 | data_masked[1502];
  assign N1898 = N1897 | data_masked[1566];
  assign N1897 = N1896 | data_masked[1630];
  assign N1896 = N1895 | data_masked[1694];
  assign N1895 = N1894 | data_masked[1758];
  assign N1894 = N1893 | data_masked[1822];
  assign N1893 = N1892 | data_masked[1886];
  assign N1892 = N1891 | data_masked[1950];
  assign N1891 = N1890 | data_masked[2014];
  assign N1890 = N1889 | data_masked[2078];
  assign N1889 = N1888 | data_masked[2142];
  assign N1888 = N1887 | data_masked[2206];
  assign N1887 = N1886 | data_masked[2270];
  assign N1886 = N1885 | data_masked[2334];
  assign N1885 = N1884 | data_masked[2398];
  assign N1884 = N1883 | data_masked[2462];
  assign N1883 = N1882 | data_masked[2526];
  assign N1882 = N1881 | data_masked[2590];
  assign N1881 = N1880 | data_masked[2654];
  assign N1880 = N1879 | data_masked[2718];
  assign N1879 = N1878 | data_masked[2782];
  assign N1878 = N1877 | data_masked[2846];
  assign N1877 = N1876 | data_masked[2910];
  assign N1876 = N1875 | data_masked[2974];
  assign N1875 = N1874 | data_masked[3038];
  assign N1874 = N1873 | data_masked[3102];
  assign N1873 = N1872 | data_masked[3166];
  assign N1872 = N1871 | data_masked[3230];
  assign N1871 = N1870 | data_masked[3294];
  assign N1870 = N1869 | data_masked[3358];
  assign N1869 = N1868 | data_masked[3422];
  assign N1868 = N1867 | data_masked[3486];
  assign N1867 = N1866 | data_masked[3550];
  assign N1866 = N1865 | data_masked[3614];
  assign N1865 = N1864 | data_masked[3678];
  assign N1864 = N1863 | data_masked[3742];
  assign N1863 = N1862 | data_masked[3806];
  assign N1862 = N1861 | data_masked[3870];
  assign N1861 = N1860 | data_masked[3934];
  assign N1860 = data_masked[4062] | data_masked[3998];
  assign data_o[31] = N1983 | data_masked[31];
  assign N1983 = N1982 | data_masked[95];
  assign N1982 = N1981 | data_masked[159];
  assign N1981 = N1980 | data_masked[223];
  assign N1980 = N1979 | data_masked[287];
  assign N1979 = N1978 | data_masked[351];
  assign N1978 = N1977 | data_masked[415];
  assign N1977 = N1976 | data_masked[479];
  assign N1976 = N1975 | data_masked[543];
  assign N1975 = N1974 | data_masked[607];
  assign N1974 = N1973 | data_masked[671];
  assign N1973 = N1972 | data_masked[735];
  assign N1972 = N1971 | data_masked[799];
  assign N1971 = N1970 | data_masked[863];
  assign N1970 = N1969 | data_masked[927];
  assign N1969 = N1968 | data_masked[991];
  assign N1968 = N1967 | data_masked[1055];
  assign N1967 = N1966 | data_masked[1119];
  assign N1966 = N1965 | data_masked[1183];
  assign N1965 = N1964 | data_masked[1247];
  assign N1964 = N1963 | data_masked[1311];
  assign N1963 = N1962 | data_masked[1375];
  assign N1962 = N1961 | data_masked[1439];
  assign N1961 = N1960 | data_masked[1503];
  assign N1960 = N1959 | data_masked[1567];
  assign N1959 = N1958 | data_masked[1631];
  assign N1958 = N1957 | data_masked[1695];
  assign N1957 = N1956 | data_masked[1759];
  assign N1956 = N1955 | data_masked[1823];
  assign N1955 = N1954 | data_masked[1887];
  assign N1954 = N1953 | data_masked[1951];
  assign N1953 = N1952 | data_masked[2015];
  assign N1952 = N1951 | data_masked[2079];
  assign N1951 = N1950 | data_masked[2143];
  assign N1950 = N1949 | data_masked[2207];
  assign N1949 = N1948 | data_masked[2271];
  assign N1948 = N1947 | data_masked[2335];
  assign N1947 = N1946 | data_masked[2399];
  assign N1946 = N1945 | data_masked[2463];
  assign N1945 = N1944 | data_masked[2527];
  assign N1944 = N1943 | data_masked[2591];
  assign N1943 = N1942 | data_masked[2655];
  assign N1942 = N1941 | data_masked[2719];
  assign N1941 = N1940 | data_masked[2783];
  assign N1940 = N1939 | data_masked[2847];
  assign N1939 = N1938 | data_masked[2911];
  assign N1938 = N1937 | data_masked[2975];
  assign N1937 = N1936 | data_masked[3039];
  assign N1936 = N1935 | data_masked[3103];
  assign N1935 = N1934 | data_masked[3167];
  assign N1934 = N1933 | data_masked[3231];
  assign N1933 = N1932 | data_masked[3295];
  assign N1932 = N1931 | data_masked[3359];
  assign N1931 = N1930 | data_masked[3423];
  assign N1930 = N1929 | data_masked[3487];
  assign N1929 = N1928 | data_masked[3551];
  assign N1928 = N1927 | data_masked[3615];
  assign N1927 = N1926 | data_masked[3679];
  assign N1926 = N1925 | data_masked[3743];
  assign N1925 = N1924 | data_masked[3807];
  assign N1924 = N1923 | data_masked[3871];
  assign N1923 = N1922 | data_masked[3935];
  assign N1922 = data_masked[4063] | data_masked[3999];
  assign data_o[32] = N2045 | data_masked[32];
  assign N2045 = N2044 | data_masked[96];
  assign N2044 = N2043 | data_masked[160];
  assign N2043 = N2042 | data_masked[224];
  assign N2042 = N2041 | data_masked[288];
  assign N2041 = N2040 | data_masked[352];
  assign N2040 = N2039 | data_masked[416];
  assign N2039 = N2038 | data_masked[480];
  assign N2038 = N2037 | data_masked[544];
  assign N2037 = N2036 | data_masked[608];
  assign N2036 = N2035 | data_masked[672];
  assign N2035 = N2034 | data_masked[736];
  assign N2034 = N2033 | data_masked[800];
  assign N2033 = N2032 | data_masked[864];
  assign N2032 = N2031 | data_masked[928];
  assign N2031 = N2030 | data_masked[992];
  assign N2030 = N2029 | data_masked[1056];
  assign N2029 = N2028 | data_masked[1120];
  assign N2028 = N2027 | data_masked[1184];
  assign N2027 = N2026 | data_masked[1248];
  assign N2026 = N2025 | data_masked[1312];
  assign N2025 = N2024 | data_masked[1376];
  assign N2024 = N2023 | data_masked[1440];
  assign N2023 = N2022 | data_masked[1504];
  assign N2022 = N2021 | data_masked[1568];
  assign N2021 = N2020 | data_masked[1632];
  assign N2020 = N2019 | data_masked[1696];
  assign N2019 = N2018 | data_masked[1760];
  assign N2018 = N2017 | data_masked[1824];
  assign N2017 = N2016 | data_masked[1888];
  assign N2016 = N2015 | data_masked[1952];
  assign N2015 = N2014 | data_masked[2016];
  assign N2014 = N2013 | data_masked[2080];
  assign N2013 = N2012 | data_masked[2144];
  assign N2012 = N2011 | data_masked[2208];
  assign N2011 = N2010 | data_masked[2272];
  assign N2010 = N2009 | data_masked[2336];
  assign N2009 = N2008 | data_masked[2400];
  assign N2008 = N2007 | data_masked[2464];
  assign N2007 = N2006 | data_masked[2528];
  assign N2006 = N2005 | data_masked[2592];
  assign N2005 = N2004 | data_masked[2656];
  assign N2004 = N2003 | data_masked[2720];
  assign N2003 = N2002 | data_masked[2784];
  assign N2002 = N2001 | data_masked[2848];
  assign N2001 = N2000 | data_masked[2912];
  assign N2000 = N1999 | data_masked[2976];
  assign N1999 = N1998 | data_masked[3040];
  assign N1998 = N1997 | data_masked[3104];
  assign N1997 = N1996 | data_masked[3168];
  assign N1996 = N1995 | data_masked[3232];
  assign N1995 = N1994 | data_masked[3296];
  assign N1994 = N1993 | data_masked[3360];
  assign N1993 = N1992 | data_masked[3424];
  assign N1992 = N1991 | data_masked[3488];
  assign N1991 = N1990 | data_masked[3552];
  assign N1990 = N1989 | data_masked[3616];
  assign N1989 = N1988 | data_masked[3680];
  assign N1988 = N1987 | data_masked[3744];
  assign N1987 = N1986 | data_masked[3808];
  assign N1986 = N1985 | data_masked[3872];
  assign N1985 = N1984 | data_masked[3936];
  assign N1984 = data_masked[4064] | data_masked[4000];
  assign data_o[33] = N2107 | data_masked[33];
  assign N2107 = N2106 | data_masked[97];
  assign N2106 = N2105 | data_masked[161];
  assign N2105 = N2104 | data_masked[225];
  assign N2104 = N2103 | data_masked[289];
  assign N2103 = N2102 | data_masked[353];
  assign N2102 = N2101 | data_masked[417];
  assign N2101 = N2100 | data_masked[481];
  assign N2100 = N2099 | data_masked[545];
  assign N2099 = N2098 | data_masked[609];
  assign N2098 = N2097 | data_masked[673];
  assign N2097 = N2096 | data_masked[737];
  assign N2096 = N2095 | data_masked[801];
  assign N2095 = N2094 | data_masked[865];
  assign N2094 = N2093 | data_masked[929];
  assign N2093 = N2092 | data_masked[993];
  assign N2092 = N2091 | data_masked[1057];
  assign N2091 = N2090 | data_masked[1121];
  assign N2090 = N2089 | data_masked[1185];
  assign N2089 = N2088 | data_masked[1249];
  assign N2088 = N2087 | data_masked[1313];
  assign N2087 = N2086 | data_masked[1377];
  assign N2086 = N2085 | data_masked[1441];
  assign N2085 = N2084 | data_masked[1505];
  assign N2084 = N2083 | data_masked[1569];
  assign N2083 = N2082 | data_masked[1633];
  assign N2082 = N2081 | data_masked[1697];
  assign N2081 = N2080 | data_masked[1761];
  assign N2080 = N2079 | data_masked[1825];
  assign N2079 = N2078 | data_masked[1889];
  assign N2078 = N2077 | data_masked[1953];
  assign N2077 = N2076 | data_masked[2017];
  assign N2076 = N2075 | data_masked[2081];
  assign N2075 = N2074 | data_masked[2145];
  assign N2074 = N2073 | data_masked[2209];
  assign N2073 = N2072 | data_masked[2273];
  assign N2072 = N2071 | data_masked[2337];
  assign N2071 = N2070 | data_masked[2401];
  assign N2070 = N2069 | data_masked[2465];
  assign N2069 = N2068 | data_masked[2529];
  assign N2068 = N2067 | data_masked[2593];
  assign N2067 = N2066 | data_masked[2657];
  assign N2066 = N2065 | data_masked[2721];
  assign N2065 = N2064 | data_masked[2785];
  assign N2064 = N2063 | data_masked[2849];
  assign N2063 = N2062 | data_masked[2913];
  assign N2062 = N2061 | data_masked[2977];
  assign N2061 = N2060 | data_masked[3041];
  assign N2060 = N2059 | data_masked[3105];
  assign N2059 = N2058 | data_masked[3169];
  assign N2058 = N2057 | data_masked[3233];
  assign N2057 = N2056 | data_masked[3297];
  assign N2056 = N2055 | data_masked[3361];
  assign N2055 = N2054 | data_masked[3425];
  assign N2054 = N2053 | data_masked[3489];
  assign N2053 = N2052 | data_masked[3553];
  assign N2052 = N2051 | data_masked[3617];
  assign N2051 = N2050 | data_masked[3681];
  assign N2050 = N2049 | data_masked[3745];
  assign N2049 = N2048 | data_masked[3809];
  assign N2048 = N2047 | data_masked[3873];
  assign N2047 = N2046 | data_masked[3937];
  assign N2046 = data_masked[4065] | data_masked[4001];
  assign data_o[34] = N2169 | data_masked[34];
  assign N2169 = N2168 | data_masked[98];
  assign N2168 = N2167 | data_masked[162];
  assign N2167 = N2166 | data_masked[226];
  assign N2166 = N2165 | data_masked[290];
  assign N2165 = N2164 | data_masked[354];
  assign N2164 = N2163 | data_masked[418];
  assign N2163 = N2162 | data_masked[482];
  assign N2162 = N2161 | data_masked[546];
  assign N2161 = N2160 | data_masked[610];
  assign N2160 = N2159 | data_masked[674];
  assign N2159 = N2158 | data_masked[738];
  assign N2158 = N2157 | data_masked[802];
  assign N2157 = N2156 | data_masked[866];
  assign N2156 = N2155 | data_masked[930];
  assign N2155 = N2154 | data_masked[994];
  assign N2154 = N2153 | data_masked[1058];
  assign N2153 = N2152 | data_masked[1122];
  assign N2152 = N2151 | data_masked[1186];
  assign N2151 = N2150 | data_masked[1250];
  assign N2150 = N2149 | data_masked[1314];
  assign N2149 = N2148 | data_masked[1378];
  assign N2148 = N2147 | data_masked[1442];
  assign N2147 = N2146 | data_masked[1506];
  assign N2146 = N2145 | data_masked[1570];
  assign N2145 = N2144 | data_masked[1634];
  assign N2144 = N2143 | data_masked[1698];
  assign N2143 = N2142 | data_masked[1762];
  assign N2142 = N2141 | data_masked[1826];
  assign N2141 = N2140 | data_masked[1890];
  assign N2140 = N2139 | data_masked[1954];
  assign N2139 = N2138 | data_masked[2018];
  assign N2138 = N2137 | data_masked[2082];
  assign N2137 = N2136 | data_masked[2146];
  assign N2136 = N2135 | data_masked[2210];
  assign N2135 = N2134 | data_masked[2274];
  assign N2134 = N2133 | data_masked[2338];
  assign N2133 = N2132 | data_masked[2402];
  assign N2132 = N2131 | data_masked[2466];
  assign N2131 = N2130 | data_masked[2530];
  assign N2130 = N2129 | data_masked[2594];
  assign N2129 = N2128 | data_masked[2658];
  assign N2128 = N2127 | data_masked[2722];
  assign N2127 = N2126 | data_masked[2786];
  assign N2126 = N2125 | data_masked[2850];
  assign N2125 = N2124 | data_masked[2914];
  assign N2124 = N2123 | data_masked[2978];
  assign N2123 = N2122 | data_masked[3042];
  assign N2122 = N2121 | data_masked[3106];
  assign N2121 = N2120 | data_masked[3170];
  assign N2120 = N2119 | data_masked[3234];
  assign N2119 = N2118 | data_masked[3298];
  assign N2118 = N2117 | data_masked[3362];
  assign N2117 = N2116 | data_masked[3426];
  assign N2116 = N2115 | data_masked[3490];
  assign N2115 = N2114 | data_masked[3554];
  assign N2114 = N2113 | data_masked[3618];
  assign N2113 = N2112 | data_masked[3682];
  assign N2112 = N2111 | data_masked[3746];
  assign N2111 = N2110 | data_masked[3810];
  assign N2110 = N2109 | data_masked[3874];
  assign N2109 = N2108 | data_masked[3938];
  assign N2108 = data_masked[4066] | data_masked[4002];
  assign data_o[35] = N2231 | data_masked[35];
  assign N2231 = N2230 | data_masked[99];
  assign N2230 = N2229 | data_masked[163];
  assign N2229 = N2228 | data_masked[227];
  assign N2228 = N2227 | data_masked[291];
  assign N2227 = N2226 | data_masked[355];
  assign N2226 = N2225 | data_masked[419];
  assign N2225 = N2224 | data_masked[483];
  assign N2224 = N2223 | data_masked[547];
  assign N2223 = N2222 | data_masked[611];
  assign N2222 = N2221 | data_masked[675];
  assign N2221 = N2220 | data_masked[739];
  assign N2220 = N2219 | data_masked[803];
  assign N2219 = N2218 | data_masked[867];
  assign N2218 = N2217 | data_masked[931];
  assign N2217 = N2216 | data_masked[995];
  assign N2216 = N2215 | data_masked[1059];
  assign N2215 = N2214 | data_masked[1123];
  assign N2214 = N2213 | data_masked[1187];
  assign N2213 = N2212 | data_masked[1251];
  assign N2212 = N2211 | data_masked[1315];
  assign N2211 = N2210 | data_masked[1379];
  assign N2210 = N2209 | data_masked[1443];
  assign N2209 = N2208 | data_masked[1507];
  assign N2208 = N2207 | data_masked[1571];
  assign N2207 = N2206 | data_masked[1635];
  assign N2206 = N2205 | data_masked[1699];
  assign N2205 = N2204 | data_masked[1763];
  assign N2204 = N2203 | data_masked[1827];
  assign N2203 = N2202 | data_masked[1891];
  assign N2202 = N2201 | data_masked[1955];
  assign N2201 = N2200 | data_masked[2019];
  assign N2200 = N2199 | data_masked[2083];
  assign N2199 = N2198 | data_masked[2147];
  assign N2198 = N2197 | data_masked[2211];
  assign N2197 = N2196 | data_masked[2275];
  assign N2196 = N2195 | data_masked[2339];
  assign N2195 = N2194 | data_masked[2403];
  assign N2194 = N2193 | data_masked[2467];
  assign N2193 = N2192 | data_masked[2531];
  assign N2192 = N2191 | data_masked[2595];
  assign N2191 = N2190 | data_masked[2659];
  assign N2190 = N2189 | data_masked[2723];
  assign N2189 = N2188 | data_masked[2787];
  assign N2188 = N2187 | data_masked[2851];
  assign N2187 = N2186 | data_masked[2915];
  assign N2186 = N2185 | data_masked[2979];
  assign N2185 = N2184 | data_masked[3043];
  assign N2184 = N2183 | data_masked[3107];
  assign N2183 = N2182 | data_masked[3171];
  assign N2182 = N2181 | data_masked[3235];
  assign N2181 = N2180 | data_masked[3299];
  assign N2180 = N2179 | data_masked[3363];
  assign N2179 = N2178 | data_masked[3427];
  assign N2178 = N2177 | data_masked[3491];
  assign N2177 = N2176 | data_masked[3555];
  assign N2176 = N2175 | data_masked[3619];
  assign N2175 = N2174 | data_masked[3683];
  assign N2174 = N2173 | data_masked[3747];
  assign N2173 = N2172 | data_masked[3811];
  assign N2172 = N2171 | data_masked[3875];
  assign N2171 = N2170 | data_masked[3939];
  assign N2170 = data_masked[4067] | data_masked[4003];
  assign data_o[36] = N2293 | data_masked[36];
  assign N2293 = N2292 | data_masked[100];
  assign N2292 = N2291 | data_masked[164];
  assign N2291 = N2290 | data_masked[228];
  assign N2290 = N2289 | data_masked[292];
  assign N2289 = N2288 | data_masked[356];
  assign N2288 = N2287 | data_masked[420];
  assign N2287 = N2286 | data_masked[484];
  assign N2286 = N2285 | data_masked[548];
  assign N2285 = N2284 | data_masked[612];
  assign N2284 = N2283 | data_masked[676];
  assign N2283 = N2282 | data_masked[740];
  assign N2282 = N2281 | data_masked[804];
  assign N2281 = N2280 | data_masked[868];
  assign N2280 = N2279 | data_masked[932];
  assign N2279 = N2278 | data_masked[996];
  assign N2278 = N2277 | data_masked[1060];
  assign N2277 = N2276 | data_masked[1124];
  assign N2276 = N2275 | data_masked[1188];
  assign N2275 = N2274 | data_masked[1252];
  assign N2274 = N2273 | data_masked[1316];
  assign N2273 = N2272 | data_masked[1380];
  assign N2272 = N2271 | data_masked[1444];
  assign N2271 = N2270 | data_masked[1508];
  assign N2270 = N2269 | data_masked[1572];
  assign N2269 = N2268 | data_masked[1636];
  assign N2268 = N2267 | data_masked[1700];
  assign N2267 = N2266 | data_masked[1764];
  assign N2266 = N2265 | data_masked[1828];
  assign N2265 = N2264 | data_masked[1892];
  assign N2264 = N2263 | data_masked[1956];
  assign N2263 = N2262 | data_masked[2020];
  assign N2262 = N2261 | data_masked[2084];
  assign N2261 = N2260 | data_masked[2148];
  assign N2260 = N2259 | data_masked[2212];
  assign N2259 = N2258 | data_masked[2276];
  assign N2258 = N2257 | data_masked[2340];
  assign N2257 = N2256 | data_masked[2404];
  assign N2256 = N2255 | data_masked[2468];
  assign N2255 = N2254 | data_masked[2532];
  assign N2254 = N2253 | data_masked[2596];
  assign N2253 = N2252 | data_masked[2660];
  assign N2252 = N2251 | data_masked[2724];
  assign N2251 = N2250 | data_masked[2788];
  assign N2250 = N2249 | data_masked[2852];
  assign N2249 = N2248 | data_masked[2916];
  assign N2248 = N2247 | data_masked[2980];
  assign N2247 = N2246 | data_masked[3044];
  assign N2246 = N2245 | data_masked[3108];
  assign N2245 = N2244 | data_masked[3172];
  assign N2244 = N2243 | data_masked[3236];
  assign N2243 = N2242 | data_masked[3300];
  assign N2242 = N2241 | data_masked[3364];
  assign N2241 = N2240 | data_masked[3428];
  assign N2240 = N2239 | data_masked[3492];
  assign N2239 = N2238 | data_masked[3556];
  assign N2238 = N2237 | data_masked[3620];
  assign N2237 = N2236 | data_masked[3684];
  assign N2236 = N2235 | data_masked[3748];
  assign N2235 = N2234 | data_masked[3812];
  assign N2234 = N2233 | data_masked[3876];
  assign N2233 = N2232 | data_masked[3940];
  assign N2232 = data_masked[4068] | data_masked[4004];
  assign data_o[37] = N2355 | data_masked[37];
  assign N2355 = N2354 | data_masked[101];
  assign N2354 = N2353 | data_masked[165];
  assign N2353 = N2352 | data_masked[229];
  assign N2352 = N2351 | data_masked[293];
  assign N2351 = N2350 | data_masked[357];
  assign N2350 = N2349 | data_masked[421];
  assign N2349 = N2348 | data_masked[485];
  assign N2348 = N2347 | data_masked[549];
  assign N2347 = N2346 | data_masked[613];
  assign N2346 = N2345 | data_masked[677];
  assign N2345 = N2344 | data_masked[741];
  assign N2344 = N2343 | data_masked[805];
  assign N2343 = N2342 | data_masked[869];
  assign N2342 = N2341 | data_masked[933];
  assign N2341 = N2340 | data_masked[997];
  assign N2340 = N2339 | data_masked[1061];
  assign N2339 = N2338 | data_masked[1125];
  assign N2338 = N2337 | data_masked[1189];
  assign N2337 = N2336 | data_masked[1253];
  assign N2336 = N2335 | data_masked[1317];
  assign N2335 = N2334 | data_masked[1381];
  assign N2334 = N2333 | data_masked[1445];
  assign N2333 = N2332 | data_masked[1509];
  assign N2332 = N2331 | data_masked[1573];
  assign N2331 = N2330 | data_masked[1637];
  assign N2330 = N2329 | data_masked[1701];
  assign N2329 = N2328 | data_masked[1765];
  assign N2328 = N2327 | data_masked[1829];
  assign N2327 = N2326 | data_masked[1893];
  assign N2326 = N2325 | data_masked[1957];
  assign N2325 = N2324 | data_masked[2021];
  assign N2324 = N2323 | data_masked[2085];
  assign N2323 = N2322 | data_masked[2149];
  assign N2322 = N2321 | data_masked[2213];
  assign N2321 = N2320 | data_masked[2277];
  assign N2320 = N2319 | data_masked[2341];
  assign N2319 = N2318 | data_masked[2405];
  assign N2318 = N2317 | data_masked[2469];
  assign N2317 = N2316 | data_masked[2533];
  assign N2316 = N2315 | data_masked[2597];
  assign N2315 = N2314 | data_masked[2661];
  assign N2314 = N2313 | data_masked[2725];
  assign N2313 = N2312 | data_masked[2789];
  assign N2312 = N2311 | data_masked[2853];
  assign N2311 = N2310 | data_masked[2917];
  assign N2310 = N2309 | data_masked[2981];
  assign N2309 = N2308 | data_masked[3045];
  assign N2308 = N2307 | data_masked[3109];
  assign N2307 = N2306 | data_masked[3173];
  assign N2306 = N2305 | data_masked[3237];
  assign N2305 = N2304 | data_masked[3301];
  assign N2304 = N2303 | data_masked[3365];
  assign N2303 = N2302 | data_masked[3429];
  assign N2302 = N2301 | data_masked[3493];
  assign N2301 = N2300 | data_masked[3557];
  assign N2300 = N2299 | data_masked[3621];
  assign N2299 = N2298 | data_masked[3685];
  assign N2298 = N2297 | data_masked[3749];
  assign N2297 = N2296 | data_masked[3813];
  assign N2296 = N2295 | data_masked[3877];
  assign N2295 = N2294 | data_masked[3941];
  assign N2294 = data_masked[4069] | data_masked[4005];
  assign data_o[38] = N2417 | data_masked[38];
  assign N2417 = N2416 | data_masked[102];
  assign N2416 = N2415 | data_masked[166];
  assign N2415 = N2414 | data_masked[230];
  assign N2414 = N2413 | data_masked[294];
  assign N2413 = N2412 | data_masked[358];
  assign N2412 = N2411 | data_masked[422];
  assign N2411 = N2410 | data_masked[486];
  assign N2410 = N2409 | data_masked[550];
  assign N2409 = N2408 | data_masked[614];
  assign N2408 = N2407 | data_masked[678];
  assign N2407 = N2406 | data_masked[742];
  assign N2406 = N2405 | data_masked[806];
  assign N2405 = N2404 | data_masked[870];
  assign N2404 = N2403 | data_masked[934];
  assign N2403 = N2402 | data_masked[998];
  assign N2402 = N2401 | data_masked[1062];
  assign N2401 = N2400 | data_masked[1126];
  assign N2400 = N2399 | data_masked[1190];
  assign N2399 = N2398 | data_masked[1254];
  assign N2398 = N2397 | data_masked[1318];
  assign N2397 = N2396 | data_masked[1382];
  assign N2396 = N2395 | data_masked[1446];
  assign N2395 = N2394 | data_masked[1510];
  assign N2394 = N2393 | data_masked[1574];
  assign N2393 = N2392 | data_masked[1638];
  assign N2392 = N2391 | data_masked[1702];
  assign N2391 = N2390 | data_masked[1766];
  assign N2390 = N2389 | data_masked[1830];
  assign N2389 = N2388 | data_masked[1894];
  assign N2388 = N2387 | data_masked[1958];
  assign N2387 = N2386 | data_masked[2022];
  assign N2386 = N2385 | data_masked[2086];
  assign N2385 = N2384 | data_masked[2150];
  assign N2384 = N2383 | data_masked[2214];
  assign N2383 = N2382 | data_masked[2278];
  assign N2382 = N2381 | data_masked[2342];
  assign N2381 = N2380 | data_masked[2406];
  assign N2380 = N2379 | data_masked[2470];
  assign N2379 = N2378 | data_masked[2534];
  assign N2378 = N2377 | data_masked[2598];
  assign N2377 = N2376 | data_masked[2662];
  assign N2376 = N2375 | data_masked[2726];
  assign N2375 = N2374 | data_masked[2790];
  assign N2374 = N2373 | data_masked[2854];
  assign N2373 = N2372 | data_masked[2918];
  assign N2372 = N2371 | data_masked[2982];
  assign N2371 = N2370 | data_masked[3046];
  assign N2370 = N2369 | data_masked[3110];
  assign N2369 = N2368 | data_masked[3174];
  assign N2368 = N2367 | data_masked[3238];
  assign N2367 = N2366 | data_masked[3302];
  assign N2366 = N2365 | data_masked[3366];
  assign N2365 = N2364 | data_masked[3430];
  assign N2364 = N2363 | data_masked[3494];
  assign N2363 = N2362 | data_masked[3558];
  assign N2362 = N2361 | data_masked[3622];
  assign N2361 = N2360 | data_masked[3686];
  assign N2360 = N2359 | data_masked[3750];
  assign N2359 = N2358 | data_masked[3814];
  assign N2358 = N2357 | data_masked[3878];
  assign N2357 = N2356 | data_masked[3942];
  assign N2356 = data_masked[4070] | data_masked[4006];
  assign data_o[39] = N2479 | data_masked[39];
  assign N2479 = N2478 | data_masked[103];
  assign N2478 = N2477 | data_masked[167];
  assign N2477 = N2476 | data_masked[231];
  assign N2476 = N2475 | data_masked[295];
  assign N2475 = N2474 | data_masked[359];
  assign N2474 = N2473 | data_masked[423];
  assign N2473 = N2472 | data_masked[487];
  assign N2472 = N2471 | data_masked[551];
  assign N2471 = N2470 | data_masked[615];
  assign N2470 = N2469 | data_masked[679];
  assign N2469 = N2468 | data_masked[743];
  assign N2468 = N2467 | data_masked[807];
  assign N2467 = N2466 | data_masked[871];
  assign N2466 = N2465 | data_masked[935];
  assign N2465 = N2464 | data_masked[999];
  assign N2464 = N2463 | data_masked[1063];
  assign N2463 = N2462 | data_masked[1127];
  assign N2462 = N2461 | data_masked[1191];
  assign N2461 = N2460 | data_masked[1255];
  assign N2460 = N2459 | data_masked[1319];
  assign N2459 = N2458 | data_masked[1383];
  assign N2458 = N2457 | data_masked[1447];
  assign N2457 = N2456 | data_masked[1511];
  assign N2456 = N2455 | data_masked[1575];
  assign N2455 = N2454 | data_masked[1639];
  assign N2454 = N2453 | data_masked[1703];
  assign N2453 = N2452 | data_masked[1767];
  assign N2452 = N2451 | data_masked[1831];
  assign N2451 = N2450 | data_masked[1895];
  assign N2450 = N2449 | data_masked[1959];
  assign N2449 = N2448 | data_masked[2023];
  assign N2448 = N2447 | data_masked[2087];
  assign N2447 = N2446 | data_masked[2151];
  assign N2446 = N2445 | data_masked[2215];
  assign N2445 = N2444 | data_masked[2279];
  assign N2444 = N2443 | data_masked[2343];
  assign N2443 = N2442 | data_masked[2407];
  assign N2442 = N2441 | data_masked[2471];
  assign N2441 = N2440 | data_masked[2535];
  assign N2440 = N2439 | data_masked[2599];
  assign N2439 = N2438 | data_masked[2663];
  assign N2438 = N2437 | data_masked[2727];
  assign N2437 = N2436 | data_masked[2791];
  assign N2436 = N2435 | data_masked[2855];
  assign N2435 = N2434 | data_masked[2919];
  assign N2434 = N2433 | data_masked[2983];
  assign N2433 = N2432 | data_masked[3047];
  assign N2432 = N2431 | data_masked[3111];
  assign N2431 = N2430 | data_masked[3175];
  assign N2430 = N2429 | data_masked[3239];
  assign N2429 = N2428 | data_masked[3303];
  assign N2428 = N2427 | data_masked[3367];
  assign N2427 = N2426 | data_masked[3431];
  assign N2426 = N2425 | data_masked[3495];
  assign N2425 = N2424 | data_masked[3559];
  assign N2424 = N2423 | data_masked[3623];
  assign N2423 = N2422 | data_masked[3687];
  assign N2422 = N2421 | data_masked[3751];
  assign N2421 = N2420 | data_masked[3815];
  assign N2420 = N2419 | data_masked[3879];
  assign N2419 = N2418 | data_masked[3943];
  assign N2418 = data_masked[4071] | data_masked[4007];
  assign data_o[40] = N2541 | data_masked[40];
  assign N2541 = N2540 | data_masked[104];
  assign N2540 = N2539 | data_masked[168];
  assign N2539 = N2538 | data_masked[232];
  assign N2538 = N2537 | data_masked[296];
  assign N2537 = N2536 | data_masked[360];
  assign N2536 = N2535 | data_masked[424];
  assign N2535 = N2534 | data_masked[488];
  assign N2534 = N2533 | data_masked[552];
  assign N2533 = N2532 | data_masked[616];
  assign N2532 = N2531 | data_masked[680];
  assign N2531 = N2530 | data_masked[744];
  assign N2530 = N2529 | data_masked[808];
  assign N2529 = N2528 | data_masked[872];
  assign N2528 = N2527 | data_masked[936];
  assign N2527 = N2526 | data_masked[1000];
  assign N2526 = N2525 | data_masked[1064];
  assign N2525 = N2524 | data_masked[1128];
  assign N2524 = N2523 | data_masked[1192];
  assign N2523 = N2522 | data_masked[1256];
  assign N2522 = N2521 | data_masked[1320];
  assign N2521 = N2520 | data_masked[1384];
  assign N2520 = N2519 | data_masked[1448];
  assign N2519 = N2518 | data_masked[1512];
  assign N2518 = N2517 | data_masked[1576];
  assign N2517 = N2516 | data_masked[1640];
  assign N2516 = N2515 | data_masked[1704];
  assign N2515 = N2514 | data_masked[1768];
  assign N2514 = N2513 | data_masked[1832];
  assign N2513 = N2512 | data_masked[1896];
  assign N2512 = N2511 | data_masked[1960];
  assign N2511 = N2510 | data_masked[2024];
  assign N2510 = N2509 | data_masked[2088];
  assign N2509 = N2508 | data_masked[2152];
  assign N2508 = N2507 | data_masked[2216];
  assign N2507 = N2506 | data_masked[2280];
  assign N2506 = N2505 | data_masked[2344];
  assign N2505 = N2504 | data_masked[2408];
  assign N2504 = N2503 | data_masked[2472];
  assign N2503 = N2502 | data_masked[2536];
  assign N2502 = N2501 | data_masked[2600];
  assign N2501 = N2500 | data_masked[2664];
  assign N2500 = N2499 | data_masked[2728];
  assign N2499 = N2498 | data_masked[2792];
  assign N2498 = N2497 | data_masked[2856];
  assign N2497 = N2496 | data_masked[2920];
  assign N2496 = N2495 | data_masked[2984];
  assign N2495 = N2494 | data_masked[3048];
  assign N2494 = N2493 | data_masked[3112];
  assign N2493 = N2492 | data_masked[3176];
  assign N2492 = N2491 | data_masked[3240];
  assign N2491 = N2490 | data_masked[3304];
  assign N2490 = N2489 | data_masked[3368];
  assign N2489 = N2488 | data_masked[3432];
  assign N2488 = N2487 | data_masked[3496];
  assign N2487 = N2486 | data_masked[3560];
  assign N2486 = N2485 | data_masked[3624];
  assign N2485 = N2484 | data_masked[3688];
  assign N2484 = N2483 | data_masked[3752];
  assign N2483 = N2482 | data_masked[3816];
  assign N2482 = N2481 | data_masked[3880];
  assign N2481 = N2480 | data_masked[3944];
  assign N2480 = data_masked[4072] | data_masked[4008];
  assign data_o[41] = N2603 | data_masked[41];
  assign N2603 = N2602 | data_masked[105];
  assign N2602 = N2601 | data_masked[169];
  assign N2601 = N2600 | data_masked[233];
  assign N2600 = N2599 | data_masked[297];
  assign N2599 = N2598 | data_masked[361];
  assign N2598 = N2597 | data_masked[425];
  assign N2597 = N2596 | data_masked[489];
  assign N2596 = N2595 | data_masked[553];
  assign N2595 = N2594 | data_masked[617];
  assign N2594 = N2593 | data_masked[681];
  assign N2593 = N2592 | data_masked[745];
  assign N2592 = N2591 | data_masked[809];
  assign N2591 = N2590 | data_masked[873];
  assign N2590 = N2589 | data_masked[937];
  assign N2589 = N2588 | data_masked[1001];
  assign N2588 = N2587 | data_masked[1065];
  assign N2587 = N2586 | data_masked[1129];
  assign N2586 = N2585 | data_masked[1193];
  assign N2585 = N2584 | data_masked[1257];
  assign N2584 = N2583 | data_masked[1321];
  assign N2583 = N2582 | data_masked[1385];
  assign N2582 = N2581 | data_masked[1449];
  assign N2581 = N2580 | data_masked[1513];
  assign N2580 = N2579 | data_masked[1577];
  assign N2579 = N2578 | data_masked[1641];
  assign N2578 = N2577 | data_masked[1705];
  assign N2577 = N2576 | data_masked[1769];
  assign N2576 = N2575 | data_masked[1833];
  assign N2575 = N2574 | data_masked[1897];
  assign N2574 = N2573 | data_masked[1961];
  assign N2573 = N2572 | data_masked[2025];
  assign N2572 = N2571 | data_masked[2089];
  assign N2571 = N2570 | data_masked[2153];
  assign N2570 = N2569 | data_masked[2217];
  assign N2569 = N2568 | data_masked[2281];
  assign N2568 = N2567 | data_masked[2345];
  assign N2567 = N2566 | data_masked[2409];
  assign N2566 = N2565 | data_masked[2473];
  assign N2565 = N2564 | data_masked[2537];
  assign N2564 = N2563 | data_masked[2601];
  assign N2563 = N2562 | data_masked[2665];
  assign N2562 = N2561 | data_masked[2729];
  assign N2561 = N2560 | data_masked[2793];
  assign N2560 = N2559 | data_masked[2857];
  assign N2559 = N2558 | data_masked[2921];
  assign N2558 = N2557 | data_masked[2985];
  assign N2557 = N2556 | data_masked[3049];
  assign N2556 = N2555 | data_masked[3113];
  assign N2555 = N2554 | data_masked[3177];
  assign N2554 = N2553 | data_masked[3241];
  assign N2553 = N2552 | data_masked[3305];
  assign N2552 = N2551 | data_masked[3369];
  assign N2551 = N2550 | data_masked[3433];
  assign N2550 = N2549 | data_masked[3497];
  assign N2549 = N2548 | data_masked[3561];
  assign N2548 = N2547 | data_masked[3625];
  assign N2547 = N2546 | data_masked[3689];
  assign N2546 = N2545 | data_masked[3753];
  assign N2545 = N2544 | data_masked[3817];
  assign N2544 = N2543 | data_masked[3881];
  assign N2543 = N2542 | data_masked[3945];
  assign N2542 = data_masked[4073] | data_masked[4009];
  assign data_o[42] = N2665 | data_masked[42];
  assign N2665 = N2664 | data_masked[106];
  assign N2664 = N2663 | data_masked[170];
  assign N2663 = N2662 | data_masked[234];
  assign N2662 = N2661 | data_masked[298];
  assign N2661 = N2660 | data_masked[362];
  assign N2660 = N2659 | data_masked[426];
  assign N2659 = N2658 | data_masked[490];
  assign N2658 = N2657 | data_masked[554];
  assign N2657 = N2656 | data_masked[618];
  assign N2656 = N2655 | data_masked[682];
  assign N2655 = N2654 | data_masked[746];
  assign N2654 = N2653 | data_masked[810];
  assign N2653 = N2652 | data_masked[874];
  assign N2652 = N2651 | data_masked[938];
  assign N2651 = N2650 | data_masked[1002];
  assign N2650 = N2649 | data_masked[1066];
  assign N2649 = N2648 | data_masked[1130];
  assign N2648 = N2647 | data_masked[1194];
  assign N2647 = N2646 | data_masked[1258];
  assign N2646 = N2645 | data_masked[1322];
  assign N2645 = N2644 | data_masked[1386];
  assign N2644 = N2643 | data_masked[1450];
  assign N2643 = N2642 | data_masked[1514];
  assign N2642 = N2641 | data_masked[1578];
  assign N2641 = N2640 | data_masked[1642];
  assign N2640 = N2639 | data_masked[1706];
  assign N2639 = N2638 | data_masked[1770];
  assign N2638 = N2637 | data_masked[1834];
  assign N2637 = N2636 | data_masked[1898];
  assign N2636 = N2635 | data_masked[1962];
  assign N2635 = N2634 | data_masked[2026];
  assign N2634 = N2633 | data_masked[2090];
  assign N2633 = N2632 | data_masked[2154];
  assign N2632 = N2631 | data_masked[2218];
  assign N2631 = N2630 | data_masked[2282];
  assign N2630 = N2629 | data_masked[2346];
  assign N2629 = N2628 | data_masked[2410];
  assign N2628 = N2627 | data_masked[2474];
  assign N2627 = N2626 | data_masked[2538];
  assign N2626 = N2625 | data_masked[2602];
  assign N2625 = N2624 | data_masked[2666];
  assign N2624 = N2623 | data_masked[2730];
  assign N2623 = N2622 | data_masked[2794];
  assign N2622 = N2621 | data_masked[2858];
  assign N2621 = N2620 | data_masked[2922];
  assign N2620 = N2619 | data_masked[2986];
  assign N2619 = N2618 | data_masked[3050];
  assign N2618 = N2617 | data_masked[3114];
  assign N2617 = N2616 | data_masked[3178];
  assign N2616 = N2615 | data_masked[3242];
  assign N2615 = N2614 | data_masked[3306];
  assign N2614 = N2613 | data_masked[3370];
  assign N2613 = N2612 | data_masked[3434];
  assign N2612 = N2611 | data_masked[3498];
  assign N2611 = N2610 | data_masked[3562];
  assign N2610 = N2609 | data_masked[3626];
  assign N2609 = N2608 | data_masked[3690];
  assign N2608 = N2607 | data_masked[3754];
  assign N2607 = N2606 | data_masked[3818];
  assign N2606 = N2605 | data_masked[3882];
  assign N2605 = N2604 | data_masked[3946];
  assign N2604 = data_masked[4074] | data_masked[4010];
  assign data_o[43] = N2727 | data_masked[43];
  assign N2727 = N2726 | data_masked[107];
  assign N2726 = N2725 | data_masked[171];
  assign N2725 = N2724 | data_masked[235];
  assign N2724 = N2723 | data_masked[299];
  assign N2723 = N2722 | data_masked[363];
  assign N2722 = N2721 | data_masked[427];
  assign N2721 = N2720 | data_masked[491];
  assign N2720 = N2719 | data_masked[555];
  assign N2719 = N2718 | data_masked[619];
  assign N2718 = N2717 | data_masked[683];
  assign N2717 = N2716 | data_masked[747];
  assign N2716 = N2715 | data_masked[811];
  assign N2715 = N2714 | data_masked[875];
  assign N2714 = N2713 | data_masked[939];
  assign N2713 = N2712 | data_masked[1003];
  assign N2712 = N2711 | data_masked[1067];
  assign N2711 = N2710 | data_masked[1131];
  assign N2710 = N2709 | data_masked[1195];
  assign N2709 = N2708 | data_masked[1259];
  assign N2708 = N2707 | data_masked[1323];
  assign N2707 = N2706 | data_masked[1387];
  assign N2706 = N2705 | data_masked[1451];
  assign N2705 = N2704 | data_masked[1515];
  assign N2704 = N2703 | data_masked[1579];
  assign N2703 = N2702 | data_masked[1643];
  assign N2702 = N2701 | data_masked[1707];
  assign N2701 = N2700 | data_masked[1771];
  assign N2700 = N2699 | data_masked[1835];
  assign N2699 = N2698 | data_masked[1899];
  assign N2698 = N2697 | data_masked[1963];
  assign N2697 = N2696 | data_masked[2027];
  assign N2696 = N2695 | data_masked[2091];
  assign N2695 = N2694 | data_masked[2155];
  assign N2694 = N2693 | data_masked[2219];
  assign N2693 = N2692 | data_masked[2283];
  assign N2692 = N2691 | data_masked[2347];
  assign N2691 = N2690 | data_masked[2411];
  assign N2690 = N2689 | data_masked[2475];
  assign N2689 = N2688 | data_masked[2539];
  assign N2688 = N2687 | data_masked[2603];
  assign N2687 = N2686 | data_masked[2667];
  assign N2686 = N2685 | data_masked[2731];
  assign N2685 = N2684 | data_masked[2795];
  assign N2684 = N2683 | data_masked[2859];
  assign N2683 = N2682 | data_masked[2923];
  assign N2682 = N2681 | data_masked[2987];
  assign N2681 = N2680 | data_masked[3051];
  assign N2680 = N2679 | data_masked[3115];
  assign N2679 = N2678 | data_masked[3179];
  assign N2678 = N2677 | data_masked[3243];
  assign N2677 = N2676 | data_masked[3307];
  assign N2676 = N2675 | data_masked[3371];
  assign N2675 = N2674 | data_masked[3435];
  assign N2674 = N2673 | data_masked[3499];
  assign N2673 = N2672 | data_masked[3563];
  assign N2672 = N2671 | data_masked[3627];
  assign N2671 = N2670 | data_masked[3691];
  assign N2670 = N2669 | data_masked[3755];
  assign N2669 = N2668 | data_masked[3819];
  assign N2668 = N2667 | data_masked[3883];
  assign N2667 = N2666 | data_masked[3947];
  assign N2666 = data_masked[4075] | data_masked[4011];
  assign data_o[44] = N2789 | data_masked[44];
  assign N2789 = N2788 | data_masked[108];
  assign N2788 = N2787 | data_masked[172];
  assign N2787 = N2786 | data_masked[236];
  assign N2786 = N2785 | data_masked[300];
  assign N2785 = N2784 | data_masked[364];
  assign N2784 = N2783 | data_masked[428];
  assign N2783 = N2782 | data_masked[492];
  assign N2782 = N2781 | data_masked[556];
  assign N2781 = N2780 | data_masked[620];
  assign N2780 = N2779 | data_masked[684];
  assign N2779 = N2778 | data_masked[748];
  assign N2778 = N2777 | data_masked[812];
  assign N2777 = N2776 | data_masked[876];
  assign N2776 = N2775 | data_masked[940];
  assign N2775 = N2774 | data_masked[1004];
  assign N2774 = N2773 | data_masked[1068];
  assign N2773 = N2772 | data_masked[1132];
  assign N2772 = N2771 | data_masked[1196];
  assign N2771 = N2770 | data_masked[1260];
  assign N2770 = N2769 | data_masked[1324];
  assign N2769 = N2768 | data_masked[1388];
  assign N2768 = N2767 | data_masked[1452];
  assign N2767 = N2766 | data_masked[1516];
  assign N2766 = N2765 | data_masked[1580];
  assign N2765 = N2764 | data_masked[1644];
  assign N2764 = N2763 | data_masked[1708];
  assign N2763 = N2762 | data_masked[1772];
  assign N2762 = N2761 | data_masked[1836];
  assign N2761 = N2760 | data_masked[1900];
  assign N2760 = N2759 | data_masked[1964];
  assign N2759 = N2758 | data_masked[2028];
  assign N2758 = N2757 | data_masked[2092];
  assign N2757 = N2756 | data_masked[2156];
  assign N2756 = N2755 | data_masked[2220];
  assign N2755 = N2754 | data_masked[2284];
  assign N2754 = N2753 | data_masked[2348];
  assign N2753 = N2752 | data_masked[2412];
  assign N2752 = N2751 | data_masked[2476];
  assign N2751 = N2750 | data_masked[2540];
  assign N2750 = N2749 | data_masked[2604];
  assign N2749 = N2748 | data_masked[2668];
  assign N2748 = N2747 | data_masked[2732];
  assign N2747 = N2746 | data_masked[2796];
  assign N2746 = N2745 | data_masked[2860];
  assign N2745 = N2744 | data_masked[2924];
  assign N2744 = N2743 | data_masked[2988];
  assign N2743 = N2742 | data_masked[3052];
  assign N2742 = N2741 | data_masked[3116];
  assign N2741 = N2740 | data_masked[3180];
  assign N2740 = N2739 | data_masked[3244];
  assign N2739 = N2738 | data_masked[3308];
  assign N2738 = N2737 | data_masked[3372];
  assign N2737 = N2736 | data_masked[3436];
  assign N2736 = N2735 | data_masked[3500];
  assign N2735 = N2734 | data_masked[3564];
  assign N2734 = N2733 | data_masked[3628];
  assign N2733 = N2732 | data_masked[3692];
  assign N2732 = N2731 | data_masked[3756];
  assign N2731 = N2730 | data_masked[3820];
  assign N2730 = N2729 | data_masked[3884];
  assign N2729 = N2728 | data_masked[3948];
  assign N2728 = data_masked[4076] | data_masked[4012];
  assign data_o[45] = N2851 | data_masked[45];
  assign N2851 = N2850 | data_masked[109];
  assign N2850 = N2849 | data_masked[173];
  assign N2849 = N2848 | data_masked[237];
  assign N2848 = N2847 | data_masked[301];
  assign N2847 = N2846 | data_masked[365];
  assign N2846 = N2845 | data_masked[429];
  assign N2845 = N2844 | data_masked[493];
  assign N2844 = N2843 | data_masked[557];
  assign N2843 = N2842 | data_masked[621];
  assign N2842 = N2841 | data_masked[685];
  assign N2841 = N2840 | data_masked[749];
  assign N2840 = N2839 | data_masked[813];
  assign N2839 = N2838 | data_masked[877];
  assign N2838 = N2837 | data_masked[941];
  assign N2837 = N2836 | data_masked[1005];
  assign N2836 = N2835 | data_masked[1069];
  assign N2835 = N2834 | data_masked[1133];
  assign N2834 = N2833 | data_masked[1197];
  assign N2833 = N2832 | data_masked[1261];
  assign N2832 = N2831 | data_masked[1325];
  assign N2831 = N2830 | data_masked[1389];
  assign N2830 = N2829 | data_masked[1453];
  assign N2829 = N2828 | data_masked[1517];
  assign N2828 = N2827 | data_masked[1581];
  assign N2827 = N2826 | data_masked[1645];
  assign N2826 = N2825 | data_masked[1709];
  assign N2825 = N2824 | data_masked[1773];
  assign N2824 = N2823 | data_masked[1837];
  assign N2823 = N2822 | data_masked[1901];
  assign N2822 = N2821 | data_masked[1965];
  assign N2821 = N2820 | data_masked[2029];
  assign N2820 = N2819 | data_masked[2093];
  assign N2819 = N2818 | data_masked[2157];
  assign N2818 = N2817 | data_masked[2221];
  assign N2817 = N2816 | data_masked[2285];
  assign N2816 = N2815 | data_masked[2349];
  assign N2815 = N2814 | data_masked[2413];
  assign N2814 = N2813 | data_masked[2477];
  assign N2813 = N2812 | data_masked[2541];
  assign N2812 = N2811 | data_masked[2605];
  assign N2811 = N2810 | data_masked[2669];
  assign N2810 = N2809 | data_masked[2733];
  assign N2809 = N2808 | data_masked[2797];
  assign N2808 = N2807 | data_masked[2861];
  assign N2807 = N2806 | data_masked[2925];
  assign N2806 = N2805 | data_masked[2989];
  assign N2805 = N2804 | data_masked[3053];
  assign N2804 = N2803 | data_masked[3117];
  assign N2803 = N2802 | data_masked[3181];
  assign N2802 = N2801 | data_masked[3245];
  assign N2801 = N2800 | data_masked[3309];
  assign N2800 = N2799 | data_masked[3373];
  assign N2799 = N2798 | data_masked[3437];
  assign N2798 = N2797 | data_masked[3501];
  assign N2797 = N2796 | data_masked[3565];
  assign N2796 = N2795 | data_masked[3629];
  assign N2795 = N2794 | data_masked[3693];
  assign N2794 = N2793 | data_masked[3757];
  assign N2793 = N2792 | data_masked[3821];
  assign N2792 = N2791 | data_masked[3885];
  assign N2791 = N2790 | data_masked[3949];
  assign N2790 = data_masked[4077] | data_masked[4013];
  assign data_o[46] = N2913 | data_masked[46];
  assign N2913 = N2912 | data_masked[110];
  assign N2912 = N2911 | data_masked[174];
  assign N2911 = N2910 | data_masked[238];
  assign N2910 = N2909 | data_masked[302];
  assign N2909 = N2908 | data_masked[366];
  assign N2908 = N2907 | data_masked[430];
  assign N2907 = N2906 | data_masked[494];
  assign N2906 = N2905 | data_masked[558];
  assign N2905 = N2904 | data_masked[622];
  assign N2904 = N2903 | data_masked[686];
  assign N2903 = N2902 | data_masked[750];
  assign N2902 = N2901 | data_masked[814];
  assign N2901 = N2900 | data_masked[878];
  assign N2900 = N2899 | data_masked[942];
  assign N2899 = N2898 | data_masked[1006];
  assign N2898 = N2897 | data_masked[1070];
  assign N2897 = N2896 | data_masked[1134];
  assign N2896 = N2895 | data_masked[1198];
  assign N2895 = N2894 | data_masked[1262];
  assign N2894 = N2893 | data_masked[1326];
  assign N2893 = N2892 | data_masked[1390];
  assign N2892 = N2891 | data_masked[1454];
  assign N2891 = N2890 | data_masked[1518];
  assign N2890 = N2889 | data_masked[1582];
  assign N2889 = N2888 | data_masked[1646];
  assign N2888 = N2887 | data_masked[1710];
  assign N2887 = N2886 | data_masked[1774];
  assign N2886 = N2885 | data_masked[1838];
  assign N2885 = N2884 | data_masked[1902];
  assign N2884 = N2883 | data_masked[1966];
  assign N2883 = N2882 | data_masked[2030];
  assign N2882 = N2881 | data_masked[2094];
  assign N2881 = N2880 | data_masked[2158];
  assign N2880 = N2879 | data_masked[2222];
  assign N2879 = N2878 | data_masked[2286];
  assign N2878 = N2877 | data_masked[2350];
  assign N2877 = N2876 | data_masked[2414];
  assign N2876 = N2875 | data_masked[2478];
  assign N2875 = N2874 | data_masked[2542];
  assign N2874 = N2873 | data_masked[2606];
  assign N2873 = N2872 | data_masked[2670];
  assign N2872 = N2871 | data_masked[2734];
  assign N2871 = N2870 | data_masked[2798];
  assign N2870 = N2869 | data_masked[2862];
  assign N2869 = N2868 | data_masked[2926];
  assign N2868 = N2867 | data_masked[2990];
  assign N2867 = N2866 | data_masked[3054];
  assign N2866 = N2865 | data_masked[3118];
  assign N2865 = N2864 | data_masked[3182];
  assign N2864 = N2863 | data_masked[3246];
  assign N2863 = N2862 | data_masked[3310];
  assign N2862 = N2861 | data_masked[3374];
  assign N2861 = N2860 | data_masked[3438];
  assign N2860 = N2859 | data_masked[3502];
  assign N2859 = N2858 | data_masked[3566];
  assign N2858 = N2857 | data_masked[3630];
  assign N2857 = N2856 | data_masked[3694];
  assign N2856 = N2855 | data_masked[3758];
  assign N2855 = N2854 | data_masked[3822];
  assign N2854 = N2853 | data_masked[3886];
  assign N2853 = N2852 | data_masked[3950];
  assign N2852 = data_masked[4078] | data_masked[4014];
  assign data_o[47] = N2975 | data_masked[47];
  assign N2975 = N2974 | data_masked[111];
  assign N2974 = N2973 | data_masked[175];
  assign N2973 = N2972 | data_masked[239];
  assign N2972 = N2971 | data_masked[303];
  assign N2971 = N2970 | data_masked[367];
  assign N2970 = N2969 | data_masked[431];
  assign N2969 = N2968 | data_masked[495];
  assign N2968 = N2967 | data_masked[559];
  assign N2967 = N2966 | data_masked[623];
  assign N2966 = N2965 | data_masked[687];
  assign N2965 = N2964 | data_masked[751];
  assign N2964 = N2963 | data_masked[815];
  assign N2963 = N2962 | data_masked[879];
  assign N2962 = N2961 | data_masked[943];
  assign N2961 = N2960 | data_masked[1007];
  assign N2960 = N2959 | data_masked[1071];
  assign N2959 = N2958 | data_masked[1135];
  assign N2958 = N2957 | data_masked[1199];
  assign N2957 = N2956 | data_masked[1263];
  assign N2956 = N2955 | data_masked[1327];
  assign N2955 = N2954 | data_masked[1391];
  assign N2954 = N2953 | data_masked[1455];
  assign N2953 = N2952 | data_masked[1519];
  assign N2952 = N2951 | data_masked[1583];
  assign N2951 = N2950 | data_masked[1647];
  assign N2950 = N2949 | data_masked[1711];
  assign N2949 = N2948 | data_masked[1775];
  assign N2948 = N2947 | data_masked[1839];
  assign N2947 = N2946 | data_masked[1903];
  assign N2946 = N2945 | data_masked[1967];
  assign N2945 = N2944 | data_masked[2031];
  assign N2944 = N2943 | data_masked[2095];
  assign N2943 = N2942 | data_masked[2159];
  assign N2942 = N2941 | data_masked[2223];
  assign N2941 = N2940 | data_masked[2287];
  assign N2940 = N2939 | data_masked[2351];
  assign N2939 = N2938 | data_masked[2415];
  assign N2938 = N2937 | data_masked[2479];
  assign N2937 = N2936 | data_masked[2543];
  assign N2936 = N2935 | data_masked[2607];
  assign N2935 = N2934 | data_masked[2671];
  assign N2934 = N2933 | data_masked[2735];
  assign N2933 = N2932 | data_masked[2799];
  assign N2932 = N2931 | data_masked[2863];
  assign N2931 = N2930 | data_masked[2927];
  assign N2930 = N2929 | data_masked[2991];
  assign N2929 = N2928 | data_masked[3055];
  assign N2928 = N2927 | data_masked[3119];
  assign N2927 = N2926 | data_masked[3183];
  assign N2926 = N2925 | data_masked[3247];
  assign N2925 = N2924 | data_masked[3311];
  assign N2924 = N2923 | data_masked[3375];
  assign N2923 = N2922 | data_masked[3439];
  assign N2922 = N2921 | data_masked[3503];
  assign N2921 = N2920 | data_masked[3567];
  assign N2920 = N2919 | data_masked[3631];
  assign N2919 = N2918 | data_masked[3695];
  assign N2918 = N2917 | data_masked[3759];
  assign N2917 = N2916 | data_masked[3823];
  assign N2916 = N2915 | data_masked[3887];
  assign N2915 = N2914 | data_masked[3951];
  assign N2914 = data_masked[4079] | data_masked[4015];
  assign data_o[48] = N3037 | data_masked[48];
  assign N3037 = N3036 | data_masked[112];
  assign N3036 = N3035 | data_masked[176];
  assign N3035 = N3034 | data_masked[240];
  assign N3034 = N3033 | data_masked[304];
  assign N3033 = N3032 | data_masked[368];
  assign N3032 = N3031 | data_masked[432];
  assign N3031 = N3030 | data_masked[496];
  assign N3030 = N3029 | data_masked[560];
  assign N3029 = N3028 | data_masked[624];
  assign N3028 = N3027 | data_masked[688];
  assign N3027 = N3026 | data_masked[752];
  assign N3026 = N3025 | data_masked[816];
  assign N3025 = N3024 | data_masked[880];
  assign N3024 = N3023 | data_masked[944];
  assign N3023 = N3022 | data_masked[1008];
  assign N3022 = N3021 | data_masked[1072];
  assign N3021 = N3020 | data_masked[1136];
  assign N3020 = N3019 | data_masked[1200];
  assign N3019 = N3018 | data_masked[1264];
  assign N3018 = N3017 | data_masked[1328];
  assign N3017 = N3016 | data_masked[1392];
  assign N3016 = N3015 | data_masked[1456];
  assign N3015 = N3014 | data_masked[1520];
  assign N3014 = N3013 | data_masked[1584];
  assign N3013 = N3012 | data_masked[1648];
  assign N3012 = N3011 | data_masked[1712];
  assign N3011 = N3010 | data_masked[1776];
  assign N3010 = N3009 | data_masked[1840];
  assign N3009 = N3008 | data_masked[1904];
  assign N3008 = N3007 | data_masked[1968];
  assign N3007 = N3006 | data_masked[2032];
  assign N3006 = N3005 | data_masked[2096];
  assign N3005 = N3004 | data_masked[2160];
  assign N3004 = N3003 | data_masked[2224];
  assign N3003 = N3002 | data_masked[2288];
  assign N3002 = N3001 | data_masked[2352];
  assign N3001 = N3000 | data_masked[2416];
  assign N3000 = N2999 | data_masked[2480];
  assign N2999 = N2998 | data_masked[2544];
  assign N2998 = N2997 | data_masked[2608];
  assign N2997 = N2996 | data_masked[2672];
  assign N2996 = N2995 | data_masked[2736];
  assign N2995 = N2994 | data_masked[2800];
  assign N2994 = N2993 | data_masked[2864];
  assign N2993 = N2992 | data_masked[2928];
  assign N2992 = N2991 | data_masked[2992];
  assign N2991 = N2990 | data_masked[3056];
  assign N2990 = N2989 | data_masked[3120];
  assign N2989 = N2988 | data_masked[3184];
  assign N2988 = N2987 | data_masked[3248];
  assign N2987 = N2986 | data_masked[3312];
  assign N2986 = N2985 | data_masked[3376];
  assign N2985 = N2984 | data_masked[3440];
  assign N2984 = N2983 | data_masked[3504];
  assign N2983 = N2982 | data_masked[3568];
  assign N2982 = N2981 | data_masked[3632];
  assign N2981 = N2980 | data_masked[3696];
  assign N2980 = N2979 | data_masked[3760];
  assign N2979 = N2978 | data_masked[3824];
  assign N2978 = N2977 | data_masked[3888];
  assign N2977 = N2976 | data_masked[3952];
  assign N2976 = data_masked[4080] | data_masked[4016];
  assign data_o[49] = N3099 | data_masked[49];
  assign N3099 = N3098 | data_masked[113];
  assign N3098 = N3097 | data_masked[177];
  assign N3097 = N3096 | data_masked[241];
  assign N3096 = N3095 | data_masked[305];
  assign N3095 = N3094 | data_masked[369];
  assign N3094 = N3093 | data_masked[433];
  assign N3093 = N3092 | data_masked[497];
  assign N3092 = N3091 | data_masked[561];
  assign N3091 = N3090 | data_masked[625];
  assign N3090 = N3089 | data_masked[689];
  assign N3089 = N3088 | data_masked[753];
  assign N3088 = N3087 | data_masked[817];
  assign N3087 = N3086 | data_masked[881];
  assign N3086 = N3085 | data_masked[945];
  assign N3085 = N3084 | data_masked[1009];
  assign N3084 = N3083 | data_masked[1073];
  assign N3083 = N3082 | data_masked[1137];
  assign N3082 = N3081 | data_masked[1201];
  assign N3081 = N3080 | data_masked[1265];
  assign N3080 = N3079 | data_masked[1329];
  assign N3079 = N3078 | data_masked[1393];
  assign N3078 = N3077 | data_masked[1457];
  assign N3077 = N3076 | data_masked[1521];
  assign N3076 = N3075 | data_masked[1585];
  assign N3075 = N3074 | data_masked[1649];
  assign N3074 = N3073 | data_masked[1713];
  assign N3073 = N3072 | data_masked[1777];
  assign N3072 = N3071 | data_masked[1841];
  assign N3071 = N3070 | data_masked[1905];
  assign N3070 = N3069 | data_masked[1969];
  assign N3069 = N3068 | data_masked[2033];
  assign N3068 = N3067 | data_masked[2097];
  assign N3067 = N3066 | data_masked[2161];
  assign N3066 = N3065 | data_masked[2225];
  assign N3065 = N3064 | data_masked[2289];
  assign N3064 = N3063 | data_masked[2353];
  assign N3063 = N3062 | data_masked[2417];
  assign N3062 = N3061 | data_masked[2481];
  assign N3061 = N3060 | data_masked[2545];
  assign N3060 = N3059 | data_masked[2609];
  assign N3059 = N3058 | data_masked[2673];
  assign N3058 = N3057 | data_masked[2737];
  assign N3057 = N3056 | data_masked[2801];
  assign N3056 = N3055 | data_masked[2865];
  assign N3055 = N3054 | data_masked[2929];
  assign N3054 = N3053 | data_masked[2993];
  assign N3053 = N3052 | data_masked[3057];
  assign N3052 = N3051 | data_masked[3121];
  assign N3051 = N3050 | data_masked[3185];
  assign N3050 = N3049 | data_masked[3249];
  assign N3049 = N3048 | data_masked[3313];
  assign N3048 = N3047 | data_masked[3377];
  assign N3047 = N3046 | data_masked[3441];
  assign N3046 = N3045 | data_masked[3505];
  assign N3045 = N3044 | data_masked[3569];
  assign N3044 = N3043 | data_masked[3633];
  assign N3043 = N3042 | data_masked[3697];
  assign N3042 = N3041 | data_masked[3761];
  assign N3041 = N3040 | data_masked[3825];
  assign N3040 = N3039 | data_masked[3889];
  assign N3039 = N3038 | data_masked[3953];
  assign N3038 = data_masked[4081] | data_masked[4017];
  assign data_o[50] = N3161 | data_masked[50];
  assign N3161 = N3160 | data_masked[114];
  assign N3160 = N3159 | data_masked[178];
  assign N3159 = N3158 | data_masked[242];
  assign N3158 = N3157 | data_masked[306];
  assign N3157 = N3156 | data_masked[370];
  assign N3156 = N3155 | data_masked[434];
  assign N3155 = N3154 | data_masked[498];
  assign N3154 = N3153 | data_masked[562];
  assign N3153 = N3152 | data_masked[626];
  assign N3152 = N3151 | data_masked[690];
  assign N3151 = N3150 | data_masked[754];
  assign N3150 = N3149 | data_masked[818];
  assign N3149 = N3148 | data_masked[882];
  assign N3148 = N3147 | data_masked[946];
  assign N3147 = N3146 | data_masked[1010];
  assign N3146 = N3145 | data_masked[1074];
  assign N3145 = N3144 | data_masked[1138];
  assign N3144 = N3143 | data_masked[1202];
  assign N3143 = N3142 | data_masked[1266];
  assign N3142 = N3141 | data_masked[1330];
  assign N3141 = N3140 | data_masked[1394];
  assign N3140 = N3139 | data_masked[1458];
  assign N3139 = N3138 | data_masked[1522];
  assign N3138 = N3137 | data_masked[1586];
  assign N3137 = N3136 | data_masked[1650];
  assign N3136 = N3135 | data_masked[1714];
  assign N3135 = N3134 | data_masked[1778];
  assign N3134 = N3133 | data_masked[1842];
  assign N3133 = N3132 | data_masked[1906];
  assign N3132 = N3131 | data_masked[1970];
  assign N3131 = N3130 | data_masked[2034];
  assign N3130 = N3129 | data_masked[2098];
  assign N3129 = N3128 | data_masked[2162];
  assign N3128 = N3127 | data_masked[2226];
  assign N3127 = N3126 | data_masked[2290];
  assign N3126 = N3125 | data_masked[2354];
  assign N3125 = N3124 | data_masked[2418];
  assign N3124 = N3123 | data_masked[2482];
  assign N3123 = N3122 | data_masked[2546];
  assign N3122 = N3121 | data_masked[2610];
  assign N3121 = N3120 | data_masked[2674];
  assign N3120 = N3119 | data_masked[2738];
  assign N3119 = N3118 | data_masked[2802];
  assign N3118 = N3117 | data_masked[2866];
  assign N3117 = N3116 | data_masked[2930];
  assign N3116 = N3115 | data_masked[2994];
  assign N3115 = N3114 | data_masked[3058];
  assign N3114 = N3113 | data_masked[3122];
  assign N3113 = N3112 | data_masked[3186];
  assign N3112 = N3111 | data_masked[3250];
  assign N3111 = N3110 | data_masked[3314];
  assign N3110 = N3109 | data_masked[3378];
  assign N3109 = N3108 | data_masked[3442];
  assign N3108 = N3107 | data_masked[3506];
  assign N3107 = N3106 | data_masked[3570];
  assign N3106 = N3105 | data_masked[3634];
  assign N3105 = N3104 | data_masked[3698];
  assign N3104 = N3103 | data_masked[3762];
  assign N3103 = N3102 | data_masked[3826];
  assign N3102 = N3101 | data_masked[3890];
  assign N3101 = N3100 | data_masked[3954];
  assign N3100 = data_masked[4082] | data_masked[4018];
  assign data_o[51] = N3223 | data_masked[51];
  assign N3223 = N3222 | data_masked[115];
  assign N3222 = N3221 | data_masked[179];
  assign N3221 = N3220 | data_masked[243];
  assign N3220 = N3219 | data_masked[307];
  assign N3219 = N3218 | data_masked[371];
  assign N3218 = N3217 | data_masked[435];
  assign N3217 = N3216 | data_masked[499];
  assign N3216 = N3215 | data_masked[563];
  assign N3215 = N3214 | data_masked[627];
  assign N3214 = N3213 | data_masked[691];
  assign N3213 = N3212 | data_masked[755];
  assign N3212 = N3211 | data_masked[819];
  assign N3211 = N3210 | data_masked[883];
  assign N3210 = N3209 | data_masked[947];
  assign N3209 = N3208 | data_masked[1011];
  assign N3208 = N3207 | data_masked[1075];
  assign N3207 = N3206 | data_masked[1139];
  assign N3206 = N3205 | data_masked[1203];
  assign N3205 = N3204 | data_masked[1267];
  assign N3204 = N3203 | data_masked[1331];
  assign N3203 = N3202 | data_masked[1395];
  assign N3202 = N3201 | data_masked[1459];
  assign N3201 = N3200 | data_masked[1523];
  assign N3200 = N3199 | data_masked[1587];
  assign N3199 = N3198 | data_masked[1651];
  assign N3198 = N3197 | data_masked[1715];
  assign N3197 = N3196 | data_masked[1779];
  assign N3196 = N3195 | data_masked[1843];
  assign N3195 = N3194 | data_masked[1907];
  assign N3194 = N3193 | data_masked[1971];
  assign N3193 = N3192 | data_masked[2035];
  assign N3192 = N3191 | data_masked[2099];
  assign N3191 = N3190 | data_masked[2163];
  assign N3190 = N3189 | data_masked[2227];
  assign N3189 = N3188 | data_masked[2291];
  assign N3188 = N3187 | data_masked[2355];
  assign N3187 = N3186 | data_masked[2419];
  assign N3186 = N3185 | data_masked[2483];
  assign N3185 = N3184 | data_masked[2547];
  assign N3184 = N3183 | data_masked[2611];
  assign N3183 = N3182 | data_masked[2675];
  assign N3182 = N3181 | data_masked[2739];
  assign N3181 = N3180 | data_masked[2803];
  assign N3180 = N3179 | data_masked[2867];
  assign N3179 = N3178 | data_masked[2931];
  assign N3178 = N3177 | data_masked[2995];
  assign N3177 = N3176 | data_masked[3059];
  assign N3176 = N3175 | data_masked[3123];
  assign N3175 = N3174 | data_masked[3187];
  assign N3174 = N3173 | data_masked[3251];
  assign N3173 = N3172 | data_masked[3315];
  assign N3172 = N3171 | data_masked[3379];
  assign N3171 = N3170 | data_masked[3443];
  assign N3170 = N3169 | data_masked[3507];
  assign N3169 = N3168 | data_masked[3571];
  assign N3168 = N3167 | data_masked[3635];
  assign N3167 = N3166 | data_masked[3699];
  assign N3166 = N3165 | data_masked[3763];
  assign N3165 = N3164 | data_masked[3827];
  assign N3164 = N3163 | data_masked[3891];
  assign N3163 = N3162 | data_masked[3955];
  assign N3162 = data_masked[4083] | data_masked[4019];
  assign data_o[52] = N3285 | data_masked[52];
  assign N3285 = N3284 | data_masked[116];
  assign N3284 = N3283 | data_masked[180];
  assign N3283 = N3282 | data_masked[244];
  assign N3282 = N3281 | data_masked[308];
  assign N3281 = N3280 | data_masked[372];
  assign N3280 = N3279 | data_masked[436];
  assign N3279 = N3278 | data_masked[500];
  assign N3278 = N3277 | data_masked[564];
  assign N3277 = N3276 | data_masked[628];
  assign N3276 = N3275 | data_masked[692];
  assign N3275 = N3274 | data_masked[756];
  assign N3274 = N3273 | data_masked[820];
  assign N3273 = N3272 | data_masked[884];
  assign N3272 = N3271 | data_masked[948];
  assign N3271 = N3270 | data_masked[1012];
  assign N3270 = N3269 | data_masked[1076];
  assign N3269 = N3268 | data_masked[1140];
  assign N3268 = N3267 | data_masked[1204];
  assign N3267 = N3266 | data_masked[1268];
  assign N3266 = N3265 | data_masked[1332];
  assign N3265 = N3264 | data_masked[1396];
  assign N3264 = N3263 | data_masked[1460];
  assign N3263 = N3262 | data_masked[1524];
  assign N3262 = N3261 | data_masked[1588];
  assign N3261 = N3260 | data_masked[1652];
  assign N3260 = N3259 | data_masked[1716];
  assign N3259 = N3258 | data_masked[1780];
  assign N3258 = N3257 | data_masked[1844];
  assign N3257 = N3256 | data_masked[1908];
  assign N3256 = N3255 | data_masked[1972];
  assign N3255 = N3254 | data_masked[2036];
  assign N3254 = N3253 | data_masked[2100];
  assign N3253 = N3252 | data_masked[2164];
  assign N3252 = N3251 | data_masked[2228];
  assign N3251 = N3250 | data_masked[2292];
  assign N3250 = N3249 | data_masked[2356];
  assign N3249 = N3248 | data_masked[2420];
  assign N3248 = N3247 | data_masked[2484];
  assign N3247 = N3246 | data_masked[2548];
  assign N3246 = N3245 | data_masked[2612];
  assign N3245 = N3244 | data_masked[2676];
  assign N3244 = N3243 | data_masked[2740];
  assign N3243 = N3242 | data_masked[2804];
  assign N3242 = N3241 | data_masked[2868];
  assign N3241 = N3240 | data_masked[2932];
  assign N3240 = N3239 | data_masked[2996];
  assign N3239 = N3238 | data_masked[3060];
  assign N3238 = N3237 | data_masked[3124];
  assign N3237 = N3236 | data_masked[3188];
  assign N3236 = N3235 | data_masked[3252];
  assign N3235 = N3234 | data_masked[3316];
  assign N3234 = N3233 | data_masked[3380];
  assign N3233 = N3232 | data_masked[3444];
  assign N3232 = N3231 | data_masked[3508];
  assign N3231 = N3230 | data_masked[3572];
  assign N3230 = N3229 | data_masked[3636];
  assign N3229 = N3228 | data_masked[3700];
  assign N3228 = N3227 | data_masked[3764];
  assign N3227 = N3226 | data_masked[3828];
  assign N3226 = N3225 | data_masked[3892];
  assign N3225 = N3224 | data_masked[3956];
  assign N3224 = data_masked[4084] | data_masked[4020];
  assign data_o[53] = N3347 | data_masked[53];
  assign N3347 = N3346 | data_masked[117];
  assign N3346 = N3345 | data_masked[181];
  assign N3345 = N3344 | data_masked[245];
  assign N3344 = N3343 | data_masked[309];
  assign N3343 = N3342 | data_masked[373];
  assign N3342 = N3341 | data_masked[437];
  assign N3341 = N3340 | data_masked[501];
  assign N3340 = N3339 | data_masked[565];
  assign N3339 = N3338 | data_masked[629];
  assign N3338 = N3337 | data_masked[693];
  assign N3337 = N3336 | data_masked[757];
  assign N3336 = N3335 | data_masked[821];
  assign N3335 = N3334 | data_masked[885];
  assign N3334 = N3333 | data_masked[949];
  assign N3333 = N3332 | data_masked[1013];
  assign N3332 = N3331 | data_masked[1077];
  assign N3331 = N3330 | data_masked[1141];
  assign N3330 = N3329 | data_masked[1205];
  assign N3329 = N3328 | data_masked[1269];
  assign N3328 = N3327 | data_masked[1333];
  assign N3327 = N3326 | data_masked[1397];
  assign N3326 = N3325 | data_masked[1461];
  assign N3325 = N3324 | data_masked[1525];
  assign N3324 = N3323 | data_masked[1589];
  assign N3323 = N3322 | data_masked[1653];
  assign N3322 = N3321 | data_masked[1717];
  assign N3321 = N3320 | data_masked[1781];
  assign N3320 = N3319 | data_masked[1845];
  assign N3319 = N3318 | data_masked[1909];
  assign N3318 = N3317 | data_masked[1973];
  assign N3317 = N3316 | data_masked[2037];
  assign N3316 = N3315 | data_masked[2101];
  assign N3315 = N3314 | data_masked[2165];
  assign N3314 = N3313 | data_masked[2229];
  assign N3313 = N3312 | data_masked[2293];
  assign N3312 = N3311 | data_masked[2357];
  assign N3311 = N3310 | data_masked[2421];
  assign N3310 = N3309 | data_masked[2485];
  assign N3309 = N3308 | data_masked[2549];
  assign N3308 = N3307 | data_masked[2613];
  assign N3307 = N3306 | data_masked[2677];
  assign N3306 = N3305 | data_masked[2741];
  assign N3305 = N3304 | data_masked[2805];
  assign N3304 = N3303 | data_masked[2869];
  assign N3303 = N3302 | data_masked[2933];
  assign N3302 = N3301 | data_masked[2997];
  assign N3301 = N3300 | data_masked[3061];
  assign N3300 = N3299 | data_masked[3125];
  assign N3299 = N3298 | data_masked[3189];
  assign N3298 = N3297 | data_masked[3253];
  assign N3297 = N3296 | data_masked[3317];
  assign N3296 = N3295 | data_masked[3381];
  assign N3295 = N3294 | data_masked[3445];
  assign N3294 = N3293 | data_masked[3509];
  assign N3293 = N3292 | data_masked[3573];
  assign N3292 = N3291 | data_masked[3637];
  assign N3291 = N3290 | data_masked[3701];
  assign N3290 = N3289 | data_masked[3765];
  assign N3289 = N3288 | data_masked[3829];
  assign N3288 = N3287 | data_masked[3893];
  assign N3287 = N3286 | data_masked[3957];
  assign N3286 = data_masked[4085] | data_masked[4021];
  assign data_o[54] = N3409 | data_masked[54];
  assign N3409 = N3408 | data_masked[118];
  assign N3408 = N3407 | data_masked[182];
  assign N3407 = N3406 | data_masked[246];
  assign N3406 = N3405 | data_masked[310];
  assign N3405 = N3404 | data_masked[374];
  assign N3404 = N3403 | data_masked[438];
  assign N3403 = N3402 | data_masked[502];
  assign N3402 = N3401 | data_masked[566];
  assign N3401 = N3400 | data_masked[630];
  assign N3400 = N3399 | data_masked[694];
  assign N3399 = N3398 | data_masked[758];
  assign N3398 = N3397 | data_masked[822];
  assign N3397 = N3396 | data_masked[886];
  assign N3396 = N3395 | data_masked[950];
  assign N3395 = N3394 | data_masked[1014];
  assign N3394 = N3393 | data_masked[1078];
  assign N3393 = N3392 | data_masked[1142];
  assign N3392 = N3391 | data_masked[1206];
  assign N3391 = N3390 | data_masked[1270];
  assign N3390 = N3389 | data_masked[1334];
  assign N3389 = N3388 | data_masked[1398];
  assign N3388 = N3387 | data_masked[1462];
  assign N3387 = N3386 | data_masked[1526];
  assign N3386 = N3385 | data_masked[1590];
  assign N3385 = N3384 | data_masked[1654];
  assign N3384 = N3383 | data_masked[1718];
  assign N3383 = N3382 | data_masked[1782];
  assign N3382 = N3381 | data_masked[1846];
  assign N3381 = N3380 | data_masked[1910];
  assign N3380 = N3379 | data_masked[1974];
  assign N3379 = N3378 | data_masked[2038];
  assign N3378 = N3377 | data_masked[2102];
  assign N3377 = N3376 | data_masked[2166];
  assign N3376 = N3375 | data_masked[2230];
  assign N3375 = N3374 | data_masked[2294];
  assign N3374 = N3373 | data_masked[2358];
  assign N3373 = N3372 | data_masked[2422];
  assign N3372 = N3371 | data_masked[2486];
  assign N3371 = N3370 | data_masked[2550];
  assign N3370 = N3369 | data_masked[2614];
  assign N3369 = N3368 | data_masked[2678];
  assign N3368 = N3367 | data_masked[2742];
  assign N3367 = N3366 | data_masked[2806];
  assign N3366 = N3365 | data_masked[2870];
  assign N3365 = N3364 | data_masked[2934];
  assign N3364 = N3363 | data_masked[2998];
  assign N3363 = N3362 | data_masked[3062];
  assign N3362 = N3361 | data_masked[3126];
  assign N3361 = N3360 | data_masked[3190];
  assign N3360 = N3359 | data_masked[3254];
  assign N3359 = N3358 | data_masked[3318];
  assign N3358 = N3357 | data_masked[3382];
  assign N3357 = N3356 | data_masked[3446];
  assign N3356 = N3355 | data_masked[3510];
  assign N3355 = N3354 | data_masked[3574];
  assign N3354 = N3353 | data_masked[3638];
  assign N3353 = N3352 | data_masked[3702];
  assign N3352 = N3351 | data_masked[3766];
  assign N3351 = N3350 | data_masked[3830];
  assign N3350 = N3349 | data_masked[3894];
  assign N3349 = N3348 | data_masked[3958];
  assign N3348 = data_masked[4086] | data_masked[4022];
  assign data_o[55] = N3471 | data_masked[55];
  assign N3471 = N3470 | data_masked[119];
  assign N3470 = N3469 | data_masked[183];
  assign N3469 = N3468 | data_masked[247];
  assign N3468 = N3467 | data_masked[311];
  assign N3467 = N3466 | data_masked[375];
  assign N3466 = N3465 | data_masked[439];
  assign N3465 = N3464 | data_masked[503];
  assign N3464 = N3463 | data_masked[567];
  assign N3463 = N3462 | data_masked[631];
  assign N3462 = N3461 | data_masked[695];
  assign N3461 = N3460 | data_masked[759];
  assign N3460 = N3459 | data_masked[823];
  assign N3459 = N3458 | data_masked[887];
  assign N3458 = N3457 | data_masked[951];
  assign N3457 = N3456 | data_masked[1015];
  assign N3456 = N3455 | data_masked[1079];
  assign N3455 = N3454 | data_masked[1143];
  assign N3454 = N3453 | data_masked[1207];
  assign N3453 = N3452 | data_masked[1271];
  assign N3452 = N3451 | data_masked[1335];
  assign N3451 = N3450 | data_masked[1399];
  assign N3450 = N3449 | data_masked[1463];
  assign N3449 = N3448 | data_masked[1527];
  assign N3448 = N3447 | data_masked[1591];
  assign N3447 = N3446 | data_masked[1655];
  assign N3446 = N3445 | data_masked[1719];
  assign N3445 = N3444 | data_masked[1783];
  assign N3444 = N3443 | data_masked[1847];
  assign N3443 = N3442 | data_masked[1911];
  assign N3442 = N3441 | data_masked[1975];
  assign N3441 = N3440 | data_masked[2039];
  assign N3440 = N3439 | data_masked[2103];
  assign N3439 = N3438 | data_masked[2167];
  assign N3438 = N3437 | data_masked[2231];
  assign N3437 = N3436 | data_masked[2295];
  assign N3436 = N3435 | data_masked[2359];
  assign N3435 = N3434 | data_masked[2423];
  assign N3434 = N3433 | data_masked[2487];
  assign N3433 = N3432 | data_masked[2551];
  assign N3432 = N3431 | data_masked[2615];
  assign N3431 = N3430 | data_masked[2679];
  assign N3430 = N3429 | data_masked[2743];
  assign N3429 = N3428 | data_masked[2807];
  assign N3428 = N3427 | data_masked[2871];
  assign N3427 = N3426 | data_masked[2935];
  assign N3426 = N3425 | data_masked[2999];
  assign N3425 = N3424 | data_masked[3063];
  assign N3424 = N3423 | data_masked[3127];
  assign N3423 = N3422 | data_masked[3191];
  assign N3422 = N3421 | data_masked[3255];
  assign N3421 = N3420 | data_masked[3319];
  assign N3420 = N3419 | data_masked[3383];
  assign N3419 = N3418 | data_masked[3447];
  assign N3418 = N3417 | data_masked[3511];
  assign N3417 = N3416 | data_masked[3575];
  assign N3416 = N3415 | data_masked[3639];
  assign N3415 = N3414 | data_masked[3703];
  assign N3414 = N3413 | data_masked[3767];
  assign N3413 = N3412 | data_masked[3831];
  assign N3412 = N3411 | data_masked[3895];
  assign N3411 = N3410 | data_masked[3959];
  assign N3410 = data_masked[4087] | data_masked[4023];
  assign data_o[56] = N3533 | data_masked[56];
  assign N3533 = N3532 | data_masked[120];
  assign N3532 = N3531 | data_masked[184];
  assign N3531 = N3530 | data_masked[248];
  assign N3530 = N3529 | data_masked[312];
  assign N3529 = N3528 | data_masked[376];
  assign N3528 = N3527 | data_masked[440];
  assign N3527 = N3526 | data_masked[504];
  assign N3526 = N3525 | data_masked[568];
  assign N3525 = N3524 | data_masked[632];
  assign N3524 = N3523 | data_masked[696];
  assign N3523 = N3522 | data_masked[760];
  assign N3522 = N3521 | data_masked[824];
  assign N3521 = N3520 | data_masked[888];
  assign N3520 = N3519 | data_masked[952];
  assign N3519 = N3518 | data_masked[1016];
  assign N3518 = N3517 | data_masked[1080];
  assign N3517 = N3516 | data_masked[1144];
  assign N3516 = N3515 | data_masked[1208];
  assign N3515 = N3514 | data_masked[1272];
  assign N3514 = N3513 | data_masked[1336];
  assign N3513 = N3512 | data_masked[1400];
  assign N3512 = N3511 | data_masked[1464];
  assign N3511 = N3510 | data_masked[1528];
  assign N3510 = N3509 | data_masked[1592];
  assign N3509 = N3508 | data_masked[1656];
  assign N3508 = N3507 | data_masked[1720];
  assign N3507 = N3506 | data_masked[1784];
  assign N3506 = N3505 | data_masked[1848];
  assign N3505 = N3504 | data_masked[1912];
  assign N3504 = N3503 | data_masked[1976];
  assign N3503 = N3502 | data_masked[2040];
  assign N3502 = N3501 | data_masked[2104];
  assign N3501 = N3500 | data_masked[2168];
  assign N3500 = N3499 | data_masked[2232];
  assign N3499 = N3498 | data_masked[2296];
  assign N3498 = N3497 | data_masked[2360];
  assign N3497 = N3496 | data_masked[2424];
  assign N3496 = N3495 | data_masked[2488];
  assign N3495 = N3494 | data_masked[2552];
  assign N3494 = N3493 | data_masked[2616];
  assign N3493 = N3492 | data_masked[2680];
  assign N3492 = N3491 | data_masked[2744];
  assign N3491 = N3490 | data_masked[2808];
  assign N3490 = N3489 | data_masked[2872];
  assign N3489 = N3488 | data_masked[2936];
  assign N3488 = N3487 | data_masked[3000];
  assign N3487 = N3486 | data_masked[3064];
  assign N3486 = N3485 | data_masked[3128];
  assign N3485 = N3484 | data_masked[3192];
  assign N3484 = N3483 | data_masked[3256];
  assign N3483 = N3482 | data_masked[3320];
  assign N3482 = N3481 | data_masked[3384];
  assign N3481 = N3480 | data_masked[3448];
  assign N3480 = N3479 | data_masked[3512];
  assign N3479 = N3478 | data_masked[3576];
  assign N3478 = N3477 | data_masked[3640];
  assign N3477 = N3476 | data_masked[3704];
  assign N3476 = N3475 | data_masked[3768];
  assign N3475 = N3474 | data_masked[3832];
  assign N3474 = N3473 | data_masked[3896];
  assign N3473 = N3472 | data_masked[3960];
  assign N3472 = data_masked[4088] | data_masked[4024];
  assign data_o[57] = N3595 | data_masked[57];
  assign N3595 = N3594 | data_masked[121];
  assign N3594 = N3593 | data_masked[185];
  assign N3593 = N3592 | data_masked[249];
  assign N3592 = N3591 | data_masked[313];
  assign N3591 = N3590 | data_masked[377];
  assign N3590 = N3589 | data_masked[441];
  assign N3589 = N3588 | data_masked[505];
  assign N3588 = N3587 | data_masked[569];
  assign N3587 = N3586 | data_masked[633];
  assign N3586 = N3585 | data_masked[697];
  assign N3585 = N3584 | data_masked[761];
  assign N3584 = N3583 | data_masked[825];
  assign N3583 = N3582 | data_masked[889];
  assign N3582 = N3581 | data_masked[953];
  assign N3581 = N3580 | data_masked[1017];
  assign N3580 = N3579 | data_masked[1081];
  assign N3579 = N3578 | data_masked[1145];
  assign N3578 = N3577 | data_masked[1209];
  assign N3577 = N3576 | data_masked[1273];
  assign N3576 = N3575 | data_masked[1337];
  assign N3575 = N3574 | data_masked[1401];
  assign N3574 = N3573 | data_masked[1465];
  assign N3573 = N3572 | data_masked[1529];
  assign N3572 = N3571 | data_masked[1593];
  assign N3571 = N3570 | data_masked[1657];
  assign N3570 = N3569 | data_masked[1721];
  assign N3569 = N3568 | data_masked[1785];
  assign N3568 = N3567 | data_masked[1849];
  assign N3567 = N3566 | data_masked[1913];
  assign N3566 = N3565 | data_masked[1977];
  assign N3565 = N3564 | data_masked[2041];
  assign N3564 = N3563 | data_masked[2105];
  assign N3563 = N3562 | data_masked[2169];
  assign N3562 = N3561 | data_masked[2233];
  assign N3561 = N3560 | data_masked[2297];
  assign N3560 = N3559 | data_masked[2361];
  assign N3559 = N3558 | data_masked[2425];
  assign N3558 = N3557 | data_masked[2489];
  assign N3557 = N3556 | data_masked[2553];
  assign N3556 = N3555 | data_masked[2617];
  assign N3555 = N3554 | data_masked[2681];
  assign N3554 = N3553 | data_masked[2745];
  assign N3553 = N3552 | data_masked[2809];
  assign N3552 = N3551 | data_masked[2873];
  assign N3551 = N3550 | data_masked[2937];
  assign N3550 = N3549 | data_masked[3001];
  assign N3549 = N3548 | data_masked[3065];
  assign N3548 = N3547 | data_masked[3129];
  assign N3547 = N3546 | data_masked[3193];
  assign N3546 = N3545 | data_masked[3257];
  assign N3545 = N3544 | data_masked[3321];
  assign N3544 = N3543 | data_masked[3385];
  assign N3543 = N3542 | data_masked[3449];
  assign N3542 = N3541 | data_masked[3513];
  assign N3541 = N3540 | data_masked[3577];
  assign N3540 = N3539 | data_masked[3641];
  assign N3539 = N3538 | data_masked[3705];
  assign N3538 = N3537 | data_masked[3769];
  assign N3537 = N3536 | data_masked[3833];
  assign N3536 = N3535 | data_masked[3897];
  assign N3535 = N3534 | data_masked[3961];
  assign N3534 = data_masked[4089] | data_masked[4025];
  assign data_o[58] = N3657 | data_masked[58];
  assign N3657 = N3656 | data_masked[122];
  assign N3656 = N3655 | data_masked[186];
  assign N3655 = N3654 | data_masked[250];
  assign N3654 = N3653 | data_masked[314];
  assign N3653 = N3652 | data_masked[378];
  assign N3652 = N3651 | data_masked[442];
  assign N3651 = N3650 | data_masked[506];
  assign N3650 = N3649 | data_masked[570];
  assign N3649 = N3648 | data_masked[634];
  assign N3648 = N3647 | data_masked[698];
  assign N3647 = N3646 | data_masked[762];
  assign N3646 = N3645 | data_masked[826];
  assign N3645 = N3644 | data_masked[890];
  assign N3644 = N3643 | data_masked[954];
  assign N3643 = N3642 | data_masked[1018];
  assign N3642 = N3641 | data_masked[1082];
  assign N3641 = N3640 | data_masked[1146];
  assign N3640 = N3639 | data_masked[1210];
  assign N3639 = N3638 | data_masked[1274];
  assign N3638 = N3637 | data_masked[1338];
  assign N3637 = N3636 | data_masked[1402];
  assign N3636 = N3635 | data_masked[1466];
  assign N3635 = N3634 | data_masked[1530];
  assign N3634 = N3633 | data_masked[1594];
  assign N3633 = N3632 | data_masked[1658];
  assign N3632 = N3631 | data_masked[1722];
  assign N3631 = N3630 | data_masked[1786];
  assign N3630 = N3629 | data_masked[1850];
  assign N3629 = N3628 | data_masked[1914];
  assign N3628 = N3627 | data_masked[1978];
  assign N3627 = N3626 | data_masked[2042];
  assign N3626 = N3625 | data_masked[2106];
  assign N3625 = N3624 | data_masked[2170];
  assign N3624 = N3623 | data_masked[2234];
  assign N3623 = N3622 | data_masked[2298];
  assign N3622 = N3621 | data_masked[2362];
  assign N3621 = N3620 | data_masked[2426];
  assign N3620 = N3619 | data_masked[2490];
  assign N3619 = N3618 | data_masked[2554];
  assign N3618 = N3617 | data_masked[2618];
  assign N3617 = N3616 | data_masked[2682];
  assign N3616 = N3615 | data_masked[2746];
  assign N3615 = N3614 | data_masked[2810];
  assign N3614 = N3613 | data_masked[2874];
  assign N3613 = N3612 | data_masked[2938];
  assign N3612 = N3611 | data_masked[3002];
  assign N3611 = N3610 | data_masked[3066];
  assign N3610 = N3609 | data_masked[3130];
  assign N3609 = N3608 | data_masked[3194];
  assign N3608 = N3607 | data_masked[3258];
  assign N3607 = N3606 | data_masked[3322];
  assign N3606 = N3605 | data_masked[3386];
  assign N3605 = N3604 | data_masked[3450];
  assign N3604 = N3603 | data_masked[3514];
  assign N3603 = N3602 | data_masked[3578];
  assign N3602 = N3601 | data_masked[3642];
  assign N3601 = N3600 | data_masked[3706];
  assign N3600 = N3599 | data_masked[3770];
  assign N3599 = N3598 | data_masked[3834];
  assign N3598 = N3597 | data_masked[3898];
  assign N3597 = N3596 | data_masked[3962];
  assign N3596 = data_masked[4090] | data_masked[4026];
  assign data_o[59] = N3719 | data_masked[59];
  assign N3719 = N3718 | data_masked[123];
  assign N3718 = N3717 | data_masked[187];
  assign N3717 = N3716 | data_masked[251];
  assign N3716 = N3715 | data_masked[315];
  assign N3715 = N3714 | data_masked[379];
  assign N3714 = N3713 | data_masked[443];
  assign N3713 = N3712 | data_masked[507];
  assign N3712 = N3711 | data_masked[571];
  assign N3711 = N3710 | data_masked[635];
  assign N3710 = N3709 | data_masked[699];
  assign N3709 = N3708 | data_masked[763];
  assign N3708 = N3707 | data_masked[827];
  assign N3707 = N3706 | data_masked[891];
  assign N3706 = N3705 | data_masked[955];
  assign N3705 = N3704 | data_masked[1019];
  assign N3704 = N3703 | data_masked[1083];
  assign N3703 = N3702 | data_masked[1147];
  assign N3702 = N3701 | data_masked[1211];
  assign N3701 = N3700 | data_masked[1275];
  assign N3700 = N3699 | data_masked[1339];
  assign N3699 = N3698 | data_masked[1403];
  assign N3698 = N3697 | data_masked[1467];
  assign N3697 = N3696 | data_masked[1531];
  assign N3696 = N3695 | data_masked[1595];
  assign N3695 = N3694 | data_masked[1659];
  assign N3694 = N3693 | data_masked[1723];
  assign N3693 = N3692 | data_masked[1787];
  assign N3692 = N3691 | data_masked[1851];
  assign N3691 = N3690 | data_masked[1915];
  assign N3690 = N3689 | data_masked[1979];
  assign N3689 = N3688 | data_masked[2043];
  assign N3688 = N3687 | data_masked[2107];
  assign N3687 = N3686 | data_masked[2171];
  assign N3686 = N3685 | data_masked[2235];
  assign N3685 = N3684 | data_masked[2299];
  assign N3684 = N3683 | data_masked[2363];
  assign N3683 = N3682 | data_masked[2427];
  assign N3682 = N3681 | data_masked[2491];
  assign N3681 = N3680 | data_masked[2555];
  assign N3680 = N3679 | data_masked[2619];
  assign N3679 = N3678 | data_masked[2683];
  assign N3678 = N3677 | data_masked[2747];
  assign N3677 = N3676 | data_masked[2811];
  assign N3676 = N3675 | data_masked[2875];
  assign N3675 = N3674 | data_masked[2939];
  assign N3674 = N3673 | data_masked[3003];
  assign N3673 = N3672 | data_masked[3067];
  assign N3672 = N3671 | data_masked[3131];
  assign N3671 = N3670 | data_masked[3195];
  assign N3670 = N3669 | data_masked[3259];
  assign N3669 = N3668 | data_masked[3323];
  assign N3668 = N3667 | data_masked[3387];
  assign N3667 = N3666 | data_masked[3451];
  assign N3666 = N3665 | data_masked[3515];
  assign N3665 = N3664 | data_masked[3579];
  assign N3664 = N3663 | data_masked[3643];
  assign N3663 = N3662 | data_masked[3707];
  assign N3662 = N3661 | data_masked[3771];
  assign N3661 = N3660 | data_masked[3835];
  assign N3660 = N3659 | data_masked[3899];
  assign N3659 = N3658 | data_masked[3963];
  assign N3658 = data_masked[4091] | data_masked[4027];
  assign data_o[60] = N3781 | data_masked[60];
  assign N3781 = N3780 | data_masked[124];
  assign N3780 = N3779 | data_masked[188];
  assign N3779 = N3778 | data_masked[252];
  assign N3778 = N3777 | data_masked[316];
  assign N3777 = N3776 | data_masked[380];
  assign N3776 = N3775 | data_masked[444];
  assign N3775 = N3774 | data_masked[508];
  assign N3774 = N3773 | data_masked[572];
  assign N3773 = N3772 | data_masked[636];
  assign N3772 = N3771 | data_masked[700];
  assign N3771 = N3770 | data_masked[764];
  assign N3770 = N3769 | data_masked[828];
  assign N3769 = N3768 | data_masked[892];
  assign N3768 = N3767 | data_masked[956];
  assign N3767 = N3766 | data_masked[1020];
  assign N3766 = N3765 | data_masked[1084];
  assign N3765 = N3764 | data_masked[1148];
  assign N3764 = N3763 | data_masked[1212];
  assign N3763 = N3762 | data_masked[1276];
  assign N3762 = N3761 | data_masked[1340];
  assign N3761 = N3760 | data_masked[1404];
  assign N3760 = N3759 | data_masked[1468];
  assign N3759 = N3758 | data_masked[1532];
  assign N3758 = N3757 | data_masked[1596];
  assign N3757 = N3756 | data_masked[1660];
  assign N3756 = N3755 | data_masked[1724];
  assign N3755 = N3754 | data_masked[1788];
  assign N3754 = N3753 | data_masked[1852];
  assign N3753 = N3752 | data_masked[1916];
  assign N3752 = N3751 | data_masked[1980];
  assign N3751 = N3750 | data_masked[2044];
  assign N3750 = N3749 | data_masked[2108];
  assign N3749 = N3748 | data_masked[2172];
  assign N3748 = N3747 | data_masked[2236];
  assign N3747 = N3746 | data_masked[2300];
  assign N3746 = N3745 | data_masked[2364];
  assign N3745 = N3744 | data_masked[2428];
  assign N3744 = N3743 | data_masked[2492];
  assign N3743 = N3742 | data_masked[2556];
  assign N3742 = N3741 | data_masked[2620];
  assign N3741 = N3740 | data_masked[2684];
  assign N3740 = N3739 | data_masked[2748];
  assign N3739 = N3738 | data_masked[2812];
  assign N3738 = N3737 | data_masked[2876];
  assign N3737 = N3736 | data_masked[2940];
  assign N3736 = N3735 | data_masked[3004];
  assign N3735 = N3734 | data_masked[3068];
  assign N3734 = N3733 | data_masked[3132];
  assign N3733 = N3732 | data_masked[3196];
  assign N3732 = N3731 | data_masked[3260];
  assign N3731 = N3730 | data_masked[3324];
  assign N3730 = N3729 | data_masked[3388];
  assign N3729 = N3728 | data_masked[3452];
  assign N3728 = N3727 | data_masked[3516];
  assign N3727 = N3726 | data_masked[3580];
  assign N3726 = N3725 | data_masked[3644];
  assign N3725 = N3724 | data_masked[3708];
  assign N3724 = N3723 | data_masked[3772];
  assign N3723 = N3722 | data_masked[3836];
  assign N3722 = N3721 | data_masked[3900];
  assign N3721 = N3720 | data_masked[3964];
  assign N3720 = data_masked[4092] | data_masked[4028];
  assign data_o[61] = N3843 | data_masked[61];
  assign N3843 = N3842 | data_masked[125];
  assign N3842 = N3841 | data_masked[189];
  assign N3841 = N3840 | data_masked[253];
  assign N3840 = N3839 | data_masked[317];
  assign N3839 = N3838 | data_masked[381];
  assign N3838 = N3837 | data_masked[445];
  assign N3837 = N3836 | data_masked[509];
  assign N3836 = N3835 | data_masked[573];
  assign N3835 = N3834 | data_masked[637];
  assign N3834 = N3833 | data_masked[701];
  assign N3833 = N3832 | data_masked[765];
  assign N3832 = N3831 | data_masked[829];
  assign N3831 = N3830 | data_masked[893];
  assign N3830 = N3829 | data_masked[957];
  assign N3829 = N3828 | data_masked[1021];
  assign N3828 = N3827 | data_masked[1085];
  assign N3827 = N3826 | data_masked[1149];
  assign N3826 = N3825 | data_masked[1213];
  assign N3825 = N3824 | data_masked[1277];
  assign N3824 = N3823 | data_masked[1341];
  assign N3823 = N3822 | data_masked[1405];
  assign N3822 = N3821 | data_masked[1469];
  assign N3821 = N3820 | data_masked[1533];
  assign N3820 = N3819 | data_masked[1597];
  assign N3819 = N3818 | data_masked[1661];
  assign N3818 = N3817 | data_masked[1725];
  assign N3817 = N3816 | data_masked[1789];
  assign N3816 = N3815 | data_masked[1853];
  assign N3815 = N3814 | data_masked[1917];
  assign N3814 = N3813 | data_masked[1981];
  assign N3813 = N3812 | data_masked[2045];
  assign N3812 = N3811 | data_masked[2109];
  assign N3811 = N3810 | data_masked[2173];
  assign N3810 = N3809 | data_masked[2237];
  assign N3809 = N3808 | data_masked[2301];
  assign N3808 = N3807 | data_masked[2365];
  assign N3807 = N3806 | data_masked[2429];
  assign N3806 = N3805 | data_masked[2493];
  assign N3805 = N3804 | data_masked[2557];
  assign N3804 = N3803 | data_masked[2621];
  assign N3803 = N3802 | data_masked[2685];
  assign N3802 = N3801 | data_masked[2749];
  assign N3801 = N3800 | data_masked[2813];
  assign N3800 = N3799 | data_masked[2877];
  assign N3799 = N3798 | data_masked[2941];
  assign N3798 = N3797 | data_masked[3005];
  assign N3797 = N3796 | data_masked[3069];
  assign N3796 = N3795 | data_masked[3133];
  assign N3795 = N3794 | data_masked[3197];
  assign N3794 = N3793 | data_masked[3261];
  assign N3793 = N3792 | data_masked[3325];
  assign N3792 = N3791 | data_masked[3389];
  assign N3791 = N3790 | data_masked[3453];
  assign N3790 = N3789 | data_masked[3517];
  assign N3789 = N3788 | data_masked[3581];
  assign N3788 = N3787 | data_masked[3645];
  assign N3787 = N3786 | data_masked[3709];
  assign N3786 = N3785 | data_masked[3773];
  assign N3785 = N3784 | data_masked[3837];
  assign N3784 = N3783 | data_masked[3901];
  assign N3783 = N3782 | data_masked[3965];
  assign N3782 = data_masked[4093] | data_masked[4029];
  assign data_o[62] = N3905 | data_masked[62];
  assign N3905 = N3904 | data_masked[126];
  assign N3904 = N3903 | data_masked[190];
  assign N3903 = N3902 | data_masked[254];
  assign N3902 = N3901 | data_masked[318];
  assign N3901 = N3900 | data_masked[382];
  assign N3900 = N3899 | data_masked[446];
  assign N3899 = N3898 | data_masked[510];
  assign N3898 = N3897 | data_masked[574];
  assign N3897 = N3896 | data_masked[638];
  assign N3896 = N3895 | data_masked[702];
  assign N3895 = N3894 | data_masked[766];
  assign N3894 = N3893 | data_masked[830];
  assign N3893 = N3892 | data_masked[894];
  assign N3892 = N3891 | data_masked[958];
  assign N3891 = N3890 | data_masked[1022];
  assign N3890 = N3889 | data_masked[1086];
  assign N3889 = N3888 | data_masked[1150];
  assign N3888 = N3887 | data_masked[1214];
  assign N3887 = N3886 | data_masked[1278];
  assign N3886 = N3885 | data_masked[1342];
  assign N3885 = N3884 | data_masked[1406];
  assign N3884 = N3883 | data_masked[1470];
  assign N3883 = N3882 | data_masked[1534];
  assign N3882 = N3881 | data_masked[1598];
  assign N3881 = N3880 | data_masked[1662];
  assign N3880 = N3879 | data_masked[1726];
  assign N3879 = N3878 | data_masked[1790];
  assign N3878 = N3877 | data_masked[1854];
  assign N3877 = N3876 | data_masked[1918];
  assign N3876 = N3875 | data_masked[1982];
  assign N3875 = N3874 | data_masked[2046];
  assign N3874 = N3873 | data_masked[2110];
  assign N3873 = N3872 | data_masked[2174];
  assign N3872 = N3871 | data_masked[2238];
  assign N3871 = N3870 | data_masked[2302];
  assign N3870 = N3869 | data_masked[2366];
  assign N3869 = N3868 | data_masked[2430];
  assign N3868 = N3867 | data_masked[2494];
  assign N3867 = N3866 | data_masked[2558];
  assign N3866 = N3865 | data_masked[2622];
  assign N3865 = N3864 | data_masked[2686];
  assign N3864 = N3863 | data_masked[2750];
  assign N3863 = N3862 | data_masked[2814];
  assign N3862 = N3861 | data_masked[2878];
  assign N3861 = N3860 | data_masked[2942];
  assign N3860 = N3859 | data_masked[3006];
  assign N3859 = N3858 | data_masked[3070];
  assign N3858 = N3857 | data_masked[3134];
  assign N3857 = N3856 | data_masked[3198];
  assign N3856 = N3855 | data_masked[3262];
  assign N3855 = N3854 | data_masked[3326];
  assign N3854 = N3853 | data_masked[3390];
  assign N3853 = N3852 | data_masked[3454];
  assign N3852 = N3851 | data_masked[3518];
  assign N3851 = N3850 | data_masked[3582];
  assign N3850 = N3849 | data_masked[3646];
  assign N3849 = N3848 | data_masked[3710];
  assign N3848 = N3847 | data_masked[3774];
  assign N3847 = N3846 | data_masked[3838];
  assign N3846 = N3845 | data_masked[3902];
  assign N3845 = N3844 | data_masked[3966];
  assign N3844 = data_masked[4094] | data_masked[4030];
  assign data_o[63] = N3967 | data_masked[63];
  assign N3967 = N3966 | data_masked[127];
  assign N3966 = N3965 | data_masked[191];
  assign N3965 = N3964 | data_masked[255];
  assign N3964 = N3963 | data_masked[319];
  assign N3963 = N3962 | data_masked[383];
  assign N3962 = N3961 | data_masked[447];
  assign N3961 = N3960 | data_masked[511];
  assign N3960 = N3959 | data_masked[575];
  assign N3959 = N3958 | data_masked[639];
  assign N3958 = N3957 | data_masked[703];
  assign N3957 = N3956 | data_masked[767];
  assign N3956 = N3955 | data_masked[831];
  assign N3955 = N3954 | data_masked[895];
  assign N3954 = N3953 | data_masked[959];
  assign N3953 = N3952 | data_masked[1023];
  assign N3952 = N3951 | data_masked[1087];
  assign N3951 = N3950 | data_masked[1151];
  assign N3950 = N3949 | data_masked[1215];
  assign N3949 = N3948 | data_masked[1279];
  assign N3948 = N3947 | data_masked[1343];
  assign N3947 = N3946 | data_masked[1407];
  assign N3946 = N3945 | data_masked[1471];
  assign N3945 = N3944 | data_masked[1535];
  assign N3944 = N3943 | data_masked[1599];
  assign N3943 = N3942 | data_masked[1663];
  assign N3942 = N3941 | data_masked[1727];
  assign N3941 = N3940 | data_masked[1791];
  assign N3940 = N3939 | data_masked[1855];
  assign N3939 = N3938 | data_masked[1919];
  assign N3938 = N3937 | data_masked[1983];
  assign N3937 = N3936 | data_masked[2047];
  assign N3936 = N3935 | data_masked[2111];
  assign N3935 = N3934 | data_masked[2175];
  assign N3934 = N3933 | data_masked[2239];
  assign N3933 = N3932 | data_masked[2303];
  assign N3932 = N3931 | data_masked[2367];
  assign N3931 = N3930 | data_masked[2431];
  assign N3930 = N3929 | data_masked[2495];
  assign N3929 = N3928 | data_masked[2559];
  assign N3928 = N3927 | data_masked[2623];
  assign N3927 = N3926 | data_masked[2687];
  assign N3926 = N3925 | data_masked[2751];
  assign N3925 = N3924 | data_masked[2815];
  assign N3924 = N3923 | data_masked[2879];
  assign N3923 = N3922 | data_masked[2943];
  assign N3922 = N3921 | data_masked[3007];
  assign N3921 = N3920 | data_masked[3071];
  assign N3920 = N3919 | data_masked[3135];
  assign N3919 = N3918 | data_masked[3199];
  assign N3918 = N3917 | data_masked[3263];
  assign N3917 = N3916 | data_masked[3327];
  assign N3916 = N3915 | data_masked[3391];
  assign N3915 = N3914 | data_masked[3455];
  assign N3914 = N3913 | data_masked[3519];
  assign N3913 = N3912 | data_masked[3583];
  assign N3912 = N3911 | data_masked[3647];
  assign N3911 = N3910 | data_masked[3711];
  assign N3910 = N3909 | data_masked[3775];
  assign N3909 = N3908 | data_masked[3839];
  assign N3908 = N3907 | data_masked[3903];
  assign N3907 = N3906 | data_masked[3967];
  assign N3906 = data_masked[4095] | data_masked[4031];

endmodule



module bsg_crossbar_o_by_i
(
  i,
  sel_oi_one_hot_i,
  o
);

  input [4095:0] i;
  input [4095:0] sel_oi_one_hot_i;
  output [4095:0] o;
  wire [4095:0] o;

  bsg_mux_one_hot_width_p64_els_p64
  genblk1_0__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[63:0]),
    .data_o(o[63:0])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_1__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[127:64]),
    .data_o(o[127:64])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_2__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[191:128]),
    .data_o(o[191:128])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_3__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[255:192]),
    .data_o(o[255:192])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_4__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[319:256]),
    .data_o(o[319:256])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_5__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[383:320]),
    .data_o(o[383:320])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_6__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[447:384]),
    .data_o(o[447:384])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_7__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[511:448]),
    .data_o(o[511:448])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_8__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[575:512]),
    .data_o(o[575:512])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_9__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[639:576]),
    .data_o(o[639:576])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_10__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[703:640]),
    .data_o(o[703:640])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_11__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[767:704]),
    .data_o(o[767:704])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_12__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[831:768]),
    .data_o(o[831:768])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_13__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[895:832]),
    .data_o(o[895:832])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_14__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[959:896]),
    .data_o(o[959:896])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_15__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1023:960]),
    .data_o(o[1023:960])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_16__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1087:1024]),
    .data_o(o[1087:1024])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_17__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1151:1088]),
    .data_o(o[1151:1088])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_18__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1215:1152]),
    .data_o(o[1215:1152])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_19__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1279:1216]),
    .data_o(o[1279:1216])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_20__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1343:1280]),
    .data_o(o[1343:1280])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_21__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1407:1344]),
    .data_o(o[1407:1344])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_22__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1471:1408]),
    .data_o(o[1471:1408])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_23__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1535:1472]),
    .data_o(o[1535:1472])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_24__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1599:1536]),
    .data_o(o[1599:1536])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_25__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1663:1600]),
    .data_o(o[1663:1600])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_26__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1727:1664]),
    .data_o(o[1727:1664])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_27__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1791:1728]),
    .data_o(o[1791:1728])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_28__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1855:1792]),
    .data_o(o[1855:1792])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_29__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1919:1856]),
    .data_o(o[1919:1856])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_30__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1983:1920]),
    .data_o(o[1983:1920])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_31__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2047:1984]),
    .data_o(o[2047:1984])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_32__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2111:2048]),
    .data_o(o[2111:2048])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_33__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2175:2112]),
    .data_o(o[2175:2112])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_34__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2239:2176]),
    .data_o(o[2239:2176])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_35__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2303:2240]),
    .data_o(o[2303:2240])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_36__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2367:2304]),
    .data_o(o[2367:2304])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_37__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2431:2368]),
    .data_o(o[2431:2368])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_38__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2495:2432]),
    .data_o(o[2495:2432])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_39__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2559:2496]),
    .data_o(o[2559:2496])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_40__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2623:2560]),
    .data_o(o[2623:2560])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_41__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2687:2624]),
    .data_o(o[2687:2624])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_42__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2751:2688]),
    .data_o(o[2751:2688])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_43__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2815:2752]),
    .data_o(o[2815:2752])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_44__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2879:2816]),
    .data_o(o[2879:2816])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_45__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[2943:2880]),
    .data_o(o[2943:2880])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_46__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3007:2944]),
    .data_o(o[3007:2944])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_47__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3071:3008]),
    .data_o(o[3071:3008])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_48__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3135:3072]),
    .data_o(o[3135:3072])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_49__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3199:3136]),
    .data_o(o[3199:3136])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_50__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3263:3200]),
    .data_o(o[3263:3200])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_51__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3327:3264]),
    .data_o(o[3327:3264])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_52__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3391:3328]),
    .data_o(o[3391:3328])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_53__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3455:3392]),
    .data_o(o[3455:3392])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_54__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3519:3456]),
    .data_o(o[3519:3456])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_55__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3583:3520]),
    .data_o(o[3583:3520])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_56__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3647:3584]),
    .data_o(o[3647:3584])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_57__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3711:3648]),
    .data_o(o[3711:3648])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_58__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3775:3712]),
    .data_o(o[3775:3712])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_59__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3839:3776]),
    .data_o(o[3839:3776])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_60__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3903:3840]),
    .data_o(o[3903:3840])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_61__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[3967:3904]),
    .data_o(o[3967:3904])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_62__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[4031:3968]),
    .data_o(o[4031:3968])
  );


  bsg_mux_one_hot_width_p64_els_p64
  genblk1_63__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[4095:4032]),
    .data_o(o[4095:4032])
  );


endmodule

