

module top
(
  i,
  o
);

  input [63:0] i;
  output [63:0] o;

  bsg_inv
  wrapper
  (
    .i(i),
    .o(o)
  );


endmodule



module bsg_inv
(
  i,
  o
);

  input [63:0] i;
  output [63:0] o;
  wire [63:0] o;
  assign o[63] = ~i[63];
  assign o[62] = ~i[62];
  assign o[61] = ~i[61];
  assign o[60] = ~i[60];
  assign o[59] = ~i[59];
  assign o[58] = ~i[58];
  assign o[57] = ~i[57];
  assign o[56] = ~i[56];
  assign o[55] = ~i[55];
  assign o[54] = ~i[54];
  assign o[53] = ~i[53];
  assign o[52] = ~i[52];
  assign o[51] = ~i[51];
  assign o[50] = ~i[50];
  assign o[49] = ~i[49];
  assign o[48] = ~i[48];
  assign o[47] = ~i[47];
  assign o[46] = ~i[46];
  assign o[45] = ~i[45];
  assign o[44] = ~i[44];
  assign o[43] = ~i[43];
  assign o[42] = ~i[42];
  assign o[41] = ~i[41];
  assign o[40] = ~i[40];
  assign o[39] = ~i[39];
  assign o[38] = ~i[38];
  assign o[37] = ~i[37];
  assign o[36] = ~i[36];
  assign o[35] = ~i[35];
  assign o[34] = ~i[34];
  assign o[33] = ~i[33];
  assign o[32] = ~i[32];
  assign o[31] = ~i[31];
  assign o[30] = ~i[30];
  assign o[29] = ~i[29];
  assign o[28] = ~i[28];
  assign o[27] = ~i[27];
  assign o[26] = ~i[26];
  assign o[25] = ~i[25];
  assign o[24] = ~i[24];
  assign o[23] = ~i[23];
  assign o[22] = ~i[22];
  assign o[21] = ~i[21];
  assign o[20] = ~i[20];
  assign o[19] = ~i[19];
  assign o[18] = ~i[18];
  assign o[17] = ~i[17];
  assign o[16] = ~i[16];
  assign o[15] = ~i[15];
  assign o[14] = ~i[14];
  assign o[13] = ~i[13];
  assign o[12] = ~i[12];
  assign o[11] = ~i[11];
  assign o[10] = ~i[10];
  assign o[9] = ~i[9];
  assign o[8] = ~i[8];
  assign o[7] = ~i[7];
  assign o[6] = ~i[6];
  assign o[5] = ~i[5];
  assign o[4] = ~i[4];
  assign o[3] = ~i[3];
  assign o[2] = ~i[2];
  assign o[1] = ~i[1];
  assign o[0] = ~i[0];

endmodule

