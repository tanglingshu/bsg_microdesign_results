

module top
(
  clk_i,
  data_i,
  sel_i,
  data_o
);

  input [15:0] data_i;
  input [127:0] sel_i;
  output [15:0] data_o;
  input clk_i;

  bsg_fifo_shift_datapath
  wrapper
  (
    .data_i(data_i),
    .sel_i(sel_i),
    .data_o(data_o),
    .clk_i(clk_i)
  );


endmodule



module bsg_fifo_shift_datapath
(
  clk_i,
  data_i,
  sel_i,
  data_o
);

  input [15:0] data_i;
  input [127:0] sel_i;
  output [15:0] data_o;
  input clk_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,
  r_n_0__15_,r_n_0__14_,r_n_0__13_,r_n_0__12_,r_n_0__11_,r_n_0__10_,r_n_0__9_,
  r_n_0__8_,r_n_0__7_,r_n_0__6_,r_n_0__5_,r_n_0__4_,r_n_0__3_,r_n_0__2_,r_n_0__1_,
  r_n_0__0_,r_n_32__15_,r_n_32__14_,r_n_32__13_,r_n_32__12_,r_n_32__11_,r_n_32__10_,
  r_n_32__9_,r_n_32__8_,r_n_32__7_,r_n_32__6_,r_n_32__5_,r_n_32__4_,r_n_32__3_,
  r_n_32__2_,r_n_32__1_,r_n_32__0_,r_n_31__15_,r_n_31__14_,r_n_31__13_,r_n_31__12_,
  r_n_31__11_,r_n_31__10_,r_n_31__9_,r_n_31__8_,r_n_31__7_,r_n_31__6_,r_n_31__5_,
  r_n_31__4_,r_n_31__3_,r_n_31__2_,r_n_31__1_,r_n_31__0_,r_n_30__15_,r_n_30__14_,
  r_n_30__13_,r_n_30__12_,r_n_30__11_,r_n_30__10_,r_n_30__9_,r_n_30__8_,r_n_30__7_,
  r_n_30__6_,r_n_30__5_,r_n_30__4_,r_n_30__3_,r_n_30__2_,r_n_30__1_,r_n_30__0_,r_n_29__15_,
  r_n_29__14_,r_n_29__13_,r_n_29__12_,r_n_29__11_,r_n_29__10_,r_n_29__9_,
  r_n_29__8_,r_n_29__7_,r_n_29__6_,r_n_29__5_,r_n_29__4_,r_n_29__3_,r_n_29__2_,r_n_29__1_,
  r_n_29__0_,r_n_28__15_,r_n_28__14_,r_n_28__13_,r_n_28__12_,r_n_28__11_,
  r_n_28__10_,r_n_28__9_,r_n_28__8_,r_n_28__7_,r_n_28__6_,r_n_28__5_,r_n_28__4_,r_n_28__3_,
  r_n_28__2_,r_n_28__1_,r_n_28__0_,r_n_27__15_,r_n_27__14_,r_n_27__13_,r_n_27__12_,
  r_n_27__11_,r_n_27__10_,r_n_27__9_,r_n_27__8_,r_n_27__7_,r_n_27__6_,r_n_27__5_,
  r_n_27__4_,r_n_27__3_,r_n_27__2_,r_n_27__1_,r_n_27__0_,r_n_26__15_,r_n_26__14_,
  r_n_26__13_,r_n_26__12_,r_n_26__11_,r_n_26__10_,r_n_26__9_,r_n_26__8_,r_n_26__7_,
  r_n_26__6_,r_n_26__5_,r_n_26__4_,r_n_26__3_,r_n_26__2_,r_n_26__1_,r_n_26__0_,
  r_n_25__15_,r_n_25__14_,r_n_25__13_,r_n_25__12_,r_n_25__11_,r_n_25__10_,r_n_25__9_,
  r_n_25__8_,r_n_25__7_,r_n_25__6_,r_n_25__5_,r_n_25__4_,r_n_25__3_,r_n_25__2_,
  r_n_25__1_,r_n_25__0_,r_n_24__15_,r_n_24__14_,r_n_24__13_,r_n_24__12_,r_n_24__11_,
  r_n_24__10_,r_n_24__9_,r_n_24__8_,r_n_24__7_,r_n_24__6_,r_n_24__5_,r_n_24__4_,
  r_n_24__3_,r_n_24__2_,r_n_24__1_,r_n_24__0_,r_n_23__15_,r_n_23__14_,r_n_23__13_,
  r_n_23__12_,r_n_23__11_,r_n_23__10_,r_n_23__9_,r_n_23__8_,r_n_23__7_,r_n_23__6_,
  r_n_23__5_,r_n_23__4_,r_n_23__3_,r_n_23__2_,r_n_23__1_,r_n_23__0_,r_n_22__15_,
  r_n_22__14_,r_n_22__13_,r_n_22__12_,r_n_22__11_,r_n_22__10_,r_n_22__9_,r_n_22__8_,
  r_n_22__7_,r_n_22__6_,r_n_22__5_,r_n_22__4_,r_n_22__3_,r_n_22__2_,r_n_22__1_,
  r_n_22__0_,r_n_21__15_,r_n_21__14_,r_n_21__13_,r_n_21__12_,r_n_21__11_,r_n_21__10_,
  r_n_21__9_,r_n_21__8_,r_n_21__7_,r_n_21__6_,r_n_21__5_,r_n_21__4_,r_n_21__3_,
  r_n_21__2_,r_n_21__1_,r_n_21__0_,r_n_20__15_,r_n_20__14_,r_n_20__13_,r_n_20__12_,
  r_n_20__11_,r_n_20__10_,r_n_20__9_,r_n_20__8_,r_n_20__7_,r_n_20__6_,r_n_20__5_,
  r_n_20__4_,r_n_20__3_,r_n_20__2_,r_n_20__1_,r_n_20__0_,r_n_19__15_,r_n_19__14_,
  r_n_19__13_,r_n_19__12_,r_n_19__11_,r_n_19__10_,r_n_19__9_,r_n_19__8_,r_n_19__7_,
  r_n_19__6_,r_n_19__5_,r_n_19__4_,r_n_19__3_,r_n_19__2_,r_n_19__1_,r_n_19__0_,
  r_n_18__15_,r_n_18__14_,r_n_18__13_,r_n_18__12_,r_n_18__11_,r_n_18__10_,r_n_18__9_,
  r_n_18__8_,r_n_18__7_,r_n_18__6_,r_n_18__5_,r_n_18__4_,r_n_18__3_,r_n_18__2_,r_n_18__1_,
  r_n_18__0_,r_n_17__15_,r_n_17__14_,r_n_17__13_,r_n_17__12_,r_n_17__11_,
  r_n_17__10_,r_n_17__9_,r_n_17__8_,r_n_17__7_,r_n_17__6_,r_n_17__5_,r_n_17__4_,r_n_17__3_,
  r_n_17__2_,r_n_17__1_,r_n_17__0_,r_n_16__15_,r_n_16__14_,r_n_16__13_,
  r_n_16__12_,r_n_16__11_,r_n_16__10_,r_n_16__9_,r_n_16__8_,r_n_16__7_,r_n_16__6_,r_n_16__5_,
  r_n_16__4_,r_n_16__3_,r_n_16__2_,r_n_16__1_,r_n_16__0_,r_n_15__15_,r_n_15__14_,
  r_n_15__13_,r_n_15__12_,r_n_15__11_,r_n_15__10_,r_n_15__9_,r_n_15__8_,r_n_15__7_,
  r_n_15__6_,r_n_15__5_,r_n_15__4_,r_n_15__3_,r_n_15__2_,r_n_15__1_,r_n_15__0_,
  r_n_14__15_,r_n_14__14_,r_n_14__13_,r_n_14__12_,r_n_14__11_,r_n_14__10_,r_n_14__9_,
  r_n_14__8_,r_n_14__7_,r_n_14__6_,r_n_14__5_,r_n_14__4_,r_n_14__3_,r_n_14__2_,
  r_n_14__1_,r_n_14__0_,r_n_13__15_,r_n_13__14_,r_n_13__13_,r_n_13__12_,r_n_13__11_,
  r_n_13__10_,r_n_13__9_,r_n_13__8_,r_n_13__7_,r_n_13__6_,r_n_13__5_,r_n_13__4_,
  r_n_13__3_,r_n_13__2_,r_n_13__1_,r_n_13__0_,r_n_12__15_,r_n_12__14_,r_n_12__13_,
  r_n_12__12_,r_n_12__11_,r_n_12__10_,r_n_12__9_,r_n_12__8_,r_n_12__7_,r_n_12__6_,
  r_n_12__5_,r_n_12__4_,r_n_12__3_,r_n_12__2_,r_n_12__1_,r_n_12__0_,r_n_11__15_,
  r_n_11__14_,r_n_11__13_,r_n_11__12_,r_n_11__11_,r_n_11__10_,r_n_11__9_,r_n_11__8_,
  r_n_11__7_,r_n_11__6_,r_n_11__5_,r_n_11__4_,r_n_11__3_,r_n_11__2_,r_n_11__1_,
  r_n_11__0_,r_n_10__15_,r_n_10__14_,r_n_10__13_,r_n_10__12_,r_n_10__11_,r_n_10__10_,
  r_n_10__9_,r_n_10__8_,r_n_10__7_,r_n_10__6_,r_n_10__5_,r_n_10__4_,r_n_10__3_,
  r_n_10__2_,r_n_10__1_,r_n_10__0_,r_n_9__15_,r_n_9__14_,r_n_9__13_,r_n_9__12_,
  r_n_9__11_,r_n_9__10_,r_n_9__9_,r_n_9__8_,r_n_9__7_,r_n_9__6_,r_n_9__5_,r_n_9__4_,
  r_n_9__3_,r_n_9__2_,r_n_9__1_,r_n_9__0_,r_n_8__15_,r_n_8__14_,r_n_8__13_,r_n_8__12_,
  r_n_8__11_,r_n_8__10_,r_n_8__9_,r_n_8__8_,r_n_8__7_,r_n_8__6_,r_n_8__5_,r_n_8__4_,
  r_n_8__3_,r_n_8__2_,r_n_8__1_,r_n_8__0_,r_n_7__15_,r_n_7__14_,r_n_7__13_,
  r_n_7__12_,r_n_7__11_,r_n_7__10_,r_n_7__9_,r_n_7__8_,r_n_7__7_,r_n_7__6_,r_n_7__5_,
  r_n_7__4_,r_n_7__3_,r_n_7__2_,r_n_7__1_,r_n_7__0_,r_n_6__15_,r_n_6__14_,r_n_6__13_,
  r_n_6__12_,r_n_6__11_,r_n_6__10_,r_n_6__9_,r_n_6__8_,r_n_6__7_,r_n_6__6_,
  r_n_6__5_,r_n_6__4_,r_n_6__3_,r_n_6__2_,r_n_6__1_,r_n_6__0_,r_n_5__15_,r_n_5__14_,
  r_n_5__13_,r_n_5__12_,r_n_5__11_,r_n_5__10_,r_n_5__9_,r_n_5__8_,r_n_5__7_,r_n_5__6_,
  r_n_5__5_,r_n_5__4_,r_n_5__3_,r_n_5__2_,r_n_5__1_,r_n_5__0_,r_n_4__15_,r_n_4__14_,
  r_n_4__13_,r_n_4__12_,r_n_4__11_,r_n_4__10_,r_n_4__9_,r_n_4__8_,r_n_4__7_,
  r_n_4__6_,r_n_4__5_,r_n_4__4_,r_n_4__3_,r_n_4__2_,r_n_4__1_,r_n_4__0_,r_n_3__15_,
  r_n_3__14_,r_n_3__13_,r_n_3__12_,r_n_3__11_,r_n_3__10_,r_n_3__9_,r_n_3__8_,r_n_3__7_,
  r_n_3__6_,r_n_3__5_,r_n_3__4_,r_n_3__3_,r_n_3__2_,r_n_3__1_,r_n_3__0_,r_n_2__15_,
  r_n_2__14_,r_n_2__13_,r_n_2__12_,r_n_2__11_,r_n_2__10_,r_n_2__9_,r_n_2__8_,
  r_n_2__7_,r_n_2__6_,r_n_2__5_,r_n_2__4_,r_n_2__3_,r_n_2__2_,r_n_2__1_,r_n_2__0_,
  r_n_1__15_,r_n_1__14_,r_n_1__13_,r_n_1__12_,r_n_1__11_,r_n_1__10_,r_n_1__9_,
  r_n_1__8_,r_n_1__7_,r_n_1__6_,r_n_1__5_,r_n_1__4_,r_n_1__3_,r_n_1__2_,r_n_1__1_,
  r_n_1__0_,r_n_63__15_,r_n_63__14_,r_n_63__13_,r_n_63__12_,r_n_63__11_,r_n_63__10_,
  r_n_63__9_,r_n_63__8_,r_n_63__7_,r_n_63__6_,r_n_63__5_,r_n_63__4_,r_n_63__3_,
  r_n_63__2_,r_n_63__1_,r_n_63__0_,r_n_62__15_,r_n_62__14_,r_n_62__13_,r_n_62__12_,
  r_n_62__11_,r_n_62__10_,r_n_62__9_,r_n_62__8_,r_n_62__7_,r_n_62__6_,r_n_62__5_,
  r_n_62__4_,r_n_62__3_,r_n_62__2_,r_n_62__1_,r_n_62__0_,r_n_61__15_,r_n_61__14_,
  r_n_61__13_,r_n_61__12_,r_n_61__11_,r_n_61__10_,r_n_61__9_,r_n_61__8_,r_n_61__7_,
  r_n_61__6_,r_n_61__5_,r_n_61__4_,r_n_61__3_,r_n_61__2_,r_n_61__1_,r_n_61__0_,r_n_60__15_,
  r_n_60__14_,r_n_60__13_,r_n_60__12_,r_n_60__11_,r_n_60__10_,r_n_60__9_,
  r_n_60__8_,r_n_60__7_,r_n_60__6_,r_n_60__5_,r_n_60__4_,r_n_60__3_,r_n_60__2_,r_n_60__1_,
  r_n_60__0_,r_n_59__15_,r_n_59__14_,r_n_59__13_,r_n_59__12_,r_n_59__11_,
  r_n_59__10_,r_n_59__9_,r_n_59__8_,r_n_59__7_,r_n_59__6_,r_n_59__5_,r_n_59__4_,r_n_59__3_,
  r_n_59__2_,r_n_59__1_,r_n_59__0_,r_n_58__15_,r_n_58__14_,r_n_58__13_,r_n_58__12_,
  r_n_58__11_,r_n_58__10_,r_n_58__9_,r_n_58__8_,r_n_58__7_,r_n_58__6_,r_n_58__5_,
  r_n_58__4_,r_n_58__3_,r_n_58__2_,r_n_58__1_,r_n_58__0_,r_n_57__15_,r_n_57__14_,
  r_n_57__13_,r_n_57__12_,r_n_57__11_,r_n_57__10_,r_n_57__9_,r_n_57__8_,r_n_57__7_,
  r_n_57__6_,r_n_57__5_,r_n_57__4_,r_n_57__3_,r_n_57__2_,r_n_57__1_,r_n_57__0_,
  r_n_56__15_,r_n_56__14_,r_n_56__13_,r_n_56__12_,r_n_56__11_,r_n_56__10_,r_n_56__9_,
  r_n_56__8_,r_n_56__7_,r_n_56__6_,r_n_56__5_,r_n_56__4_,r_n_56__3_,r_n_56__2_,
  r_n_56__1_,r_n_56__0_,r_n_55__15_,r_n_55__14_,r_n_55__13_,r_n_55__12_,r_n_55__11_,
  r_n_55__10_,r_n_55__9_,r_n_55__8_,r_n_55__7_,r_n_55__6_,r_n_55__5_,r_n_55__4_,
  r_n_55__3_,r_n_55__2_,r_n_55__1_,r_n_55__0_,r_n_54__15_,r_n_54__14_,r_n_54__13_,
  r_n_54__12_,r_n_54__11_,r_n_54__10_,r_n_54__9_,r_n_54__8_,r_n_54__7_,r_n_54__6_,
  r_n_54__5_,r_n_54__4_,r_n_54__3_,r_n_54__2_,r_n_54__1_,r_n_54__0_,r_n_53__15_,
  r_n_53__14_,r_n_53__13_,r_n_53__12_,r_n_53__11_,r_n_53__10_,r_n_53__9_,r_n_53__8_,
  r_n_53__7_,r_n_53__6_,r_n_53__5_,r_n_53__4_,r_n_53__3_,r_n_53__2_,r_n_53__1_,
  r_n_53__0_,r_n_52__15_,r_n_52__14_,r_n_52__13_,r_n_52__12_,r_n_52__11_,r_n_52__10_,
  r_n_52__9_,r_n_52__8_,r_n_52__7_,r_n_52__6_,r_n_52__5_,r_n_52__4_,r_n_52__3_,
  r_n_52__2_,r_n_52__1_,r_n_52__0_,r_n_51__15_,r_n_51__14_,r_n_51__13_,r_n_51__12_,
  r_n_51__11_,r_n_51__10_,r_n_51__9_,r_n_51__8_,r_n_51__7_,r_n_51__6_,r_n_51__5_,
  r_n_51__4_,r_n_51__3_,r_n_51__2_,r_n_51__1_,r_n_51__0_,r_n_50__15_,r_n_50__14_,
  r_n_50__13_,r_n_50__12_,r_n_50__11_,r_n_50__10_,r_n_50__9_,r_n_50__8_,r_n_50__7_,
  r_n_50__6_,r_n_50__5_,r_n_50__4_,r_n_50__3_,r_n_50__2_,r_n_50__1_,r_n_50__0_,
  r_n_49__15_,r_n_49__14_,r_n_49__13_,r_n_49__12_,r_n_49__11_,r_n_49__10_,r_n_49__9_,
  r_n_49__8_,r_n_49__7_,r_n_49__6_,r_n_49__5_,r_n_49__4_,r_n_49__3_,r_n_49__2_,r_n_49__1_,
  r_n_49__0_,r_n_48__15_,r_n_48__14_,r_n_48__13_,r_n_48__12_,r_n_48__11_,
  r_n_48__10_,r_n_48__9_,r_n_48__8_,r_n_48__7_,r_n_48__6_,r_n_48__5_,r_n_48__4_,r_n_48__3_,
  r_n_48__2_,r_n_48__1_,r_n_48__0_,r_n_47__15_,r_n_47__14_,r_n_47__13_,
  r_n_47__12_,r_n_47__11_,r_n_47__10_,r_n_47__9_,r_n_47__8_,r_n_47__7_,r_n_47__6_,r_n_47__5_,
  r_n_47__4_,r_n_47__3_,r_n_47__2_,r_n_47__1_,r_n_47__0_,r_n_46__15_,r_n_46__14_,
  r_n_46__13_,r_n_46__12_,r_n_46__11_,r_n_46__10_,r_n_46__9_,r_n_46__8_,r_n_46__7_,
  r_n_46__6_,r_n_46__5_,r_n_46__4_,r_n_46__3_,r_n_46__2_,r_n_46__1_,r_n_46__0_,
  r_n_45__15_,r_n_45__14_,r_n_45__13_,r_n_45__12_,r_n_45__11_,r_n_45__10_,r_n_45__9_,
  r_n_45__8_,r_n_45__7_,r_n_45__6_,r_n_45__5_,r_n_45__4_,r_n_45__3_,r_n_45__2_,
  r_n_45__1_,r_n_45__0_,r_n_44__15_,r_n_44__14_,r_n_44__13_,r_n_44__12_,r_n_44__11_,
  r_n_44__10_,r_n_44__9_,r_n_44__8_,r_n_44__7_,r_n_44__6_,r_n_44__5_,r_n_44__4_,
  r_n_44__3_,r_n_44__2_,r_n_44__1_,r_n_44__0_,r_n_43__15_,r_n_43__14_,r_n_43__13_,
  r_n_43__12_,r_n_43__11_,r_n_43__10_,r_n_43__9_,r_n_43__8_,r_n_43__7_,r_n_43__6_,
  r_n_43__5_,r_n_43__4_,r_n_43__3_,r_n_43__2_,r_n_43__1_,r_n_43__0_,r_n_42__15_,
  r_n_42__14_,r_n_42__13_,r_n_42__12_,r_n_42__11_,r_n_42__10_,r_n_42__9_,r_n_42__8_,
  r_n_42__7_,r_n_42__6_,r_n_42__5_,r_n_42__4_,r_n_42__3_,r_n_42__2_,r_n_42__1_,
  r_n_42__0_,r_n_41__15_,r_n_41__14_,r_n_41__13_,r_n_41__12_,r_n_41__11_,r_n_41__10_,
  r_n_41__9_,r_n_41__8_,r_n_41__7_,r_n_41__6_,r_n_41__5_,r_n_41__4_,r_n_41__3_,
  r_n_41__2_,r_n_41__1_,r_n_41__0_,r_n_40__15_,r_n_40__14_,r_n_40__13_,r_n_40__12_,
  r_n_40__11_,r_n_40__10_,r_n_40__9_,r_n_40__8_,r_n_40__7_,r_n_40__6_,r_n_40__5_,
  r_n_40__4_,r_n_40__3_,r_n_40__2_,r_n_40__1_,r_n_40__0_,r_n_39__15_,r_n_39__14_,
  r_n_39__13_,r_n_39__12_,r_n_39__11_,r_n_39__10_,r_n_39__9_,r_n_39__8_,r_n_39__7_,
  r_n_39__6_,r_n_39__5_,r_n_39__4_,r_n_39__3_,r_n_39__2_,r_n_39__1_,r_n_39__0_,
  r_n_38__15_,r_n_38__14_,r_n_38__13_,r_n_38__12_,r_n_38__11_,r_n_38__10_,r_n_38__9_,
  r_n_38__8_,r_n_38__7_,r_n_38__6_,r_n_38__5_,r_n_38__4_,r_n_38__3_,r_n_38__2_,
  r_n_38__1_,r_n_38__0_,r_n_37__15_,r_n_37__14_,r_n_37__13_,r_n_37__12_,r_n_37__11_,
  r_n_37__10_,r_n_37__9_,r_n_37__8_,r_n_37__7_,r_n_37__6_,r_n_37__5_,r_n_37__4_,
  r_n_37__3_,r_n_37__2_,r_n_37__1_,r_n_37__0_,r_n_36__15_,r_n_36__14_,r_n_36__13_,
  r_n_36__12_,r_n_36__11_,r_n_36__10_,r_n_36__9_,r_n_36__8_,r_n_36__7_,r_n_36__6_,
  r_n_36__5_,r_n_36__4_,r_n_36__3_,r_n_36__2_,r_n_36__1_,r_n_36__0_,r_n_35__15_,
  r_n_35__14_,r_n_35__13_,r_n_35__12_,r_n_35__11_,r_n_35__10_,r_n_35__9_,r_n_35__8_,
  r_n_35__7_,r_n_35__6_,r_n_35__5_,r_n_35__4_,r_n_35__3_,r_n_35__2_,r_n_35__1_,r_n_35__0_,
  r_n_34__15_,r_n_34__14_,r_n_34__13_,r_n_34__12_,r_n_34__11_,r_n_34__10_,
  r_n_34__9_,r_n_34__8_,r_n_34__7_,r_n_34__6_,r_n_34__5_,r_n_34__4_,r_n_34__3_,r_n_34__2_,
  r_n_34__1_,r_n_34__0_,r_n_33__15_,r_n_33__14_,r_n_33__13_,r_n_33__12_,
  r_n_33__11_,r_n_33__10_,r_n_33__9_,r_n_33__8_,r_n_33__7_,r_n_33__6_,r_n_33__5_,r_n_33__4_,
  r_n_33__3_,r_n_33__2_,r_n_33__1_,r_n_33__0_,N133,N134,N135,N136,N137,N138,N139,
  N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,
  N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,
  N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,
  N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,
  N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,
  N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,
  N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,
  N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,
  N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,
  N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,
  N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,
  N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,
  N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,
  N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,
  N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,
  N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,
  N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,
  N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,
  N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,
  N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,
  N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,
  N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,
  N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,
  N508,N509,N510,N511;
  reg [15:0] data_o;
  reg r_1__15_,r_1__14_,r_1__13_,r_1__12_,r_1__11_,r_1__10_,r_1__9_,r_1__8_,r_1__7_,
  r_1__6_,r_1__5_,r_1__4_,r_1__3_,r_1__2_,r_1__1_,r_1__0_,r_2__15_,r_2__14_,
  r_2__13_,r_2__12_,r_2__11_,r_2__10_,r_2__9_,r_2__8_,r_2__7_,r_2__6_,r_2__5_,r_2__4_,
  r_2__3_,r_2__2_,r_2__1_,r_2__0_,r_3__15_,r_3__14_,r_3__13_,r_3__12_,r_3__11_,
  r_3__10_,r_3__9_,r_3__8_,r_3__7_,r_3__6_,r_3__5_,r_3__4_,r_3__3_,r_3__2_,r_3__1_,
  r_3__0_,r_4__15_,r_4__14_,r_4__13_,r_4__12_,r_4__11_,r_4__10_,r_4__9_,r_4__8_,r_4__7_,
  r_4__6_,r_4__5_,r_4__4_,r_4__3_,r_4__2_,r_4__1_,r_4__0_,r_5__15_,r_5__14_,
  r_5__13_,r_5__12_,r_5__11_,r_5__10_,r_5__9_,r_5__8_,r_5__7_,r_5__6_,r_5__5_,r_5__4_,
  r_5__3_,r_5__2_,r_5__1_,r_5__0_,r_6__15_,r_6__14_,r_6__13_,r_6__12_,r_6__11_,
  r_6__10_,r_6__9_,r_6__8_,r_6__7_,r_6__6_,r_6__5_,r_6__4_,r_6__3_,r_6__2_,r_6__1_,
  r_6__0_,r_7__15_,r_7__14_,r_7__13_,r_7__12_,r_7__11_,r_7__10_,r_7__9_,r_7__8_,
  r_7__7_,r_7__6_,r_7__5_,r_7__4_,r_7__3_,r_7__2_,r_7__1_,r_7__0_,r_8__15_,r_8__14_,
  r_8__13_,r_8__12_,r_8__11_,r_8__10_,r_8__9_,r_8__8_,r_8__7_,r_8__6_,r_8__5_,r_8__4_,
  r_8__3_,r_8__2_,r_8__1_,r_8__0_,r_9__15_,r_9__14_,r_9__13_,r_9__12_,r_9__11_,
  r_9__10_,r_9__9_,r_9__8_,r_9__7_,r_9__6_,r_9__5_,r_9__4_,r_9__3_,r_9__2_,r_9__1_,
  r_9__0_,r_10__15_,r_10__14_,r_10__13_,r_10__12_,r_10__11_,r_10__10_,r_10__9_,
  r_10__8_,r_10__7_,r_10__6_,r_10__5_,r_10__4_,r_10__3_,r_10__2_,r_10__1_,r_10__0_,
  r_11__15_,r_11__14_,r_11__13_,r_11__12_,r_11__11_,r_11__10_,r_11__9_,r_11__8_,
  r_11__7_,r_11__6_,r_11__5_,r_11__4_,r_11__3_,r_11__2_,r_11__1_,r_11__0_,r_12__15_,
  r_12__14_,r_12__13_,r_12__12_,r_12__11_,r_12__10_,r_12__9_,r_12__8_,r_12__7_,
  r_12__6_,r_12__5_,r_12__4_,r_12__3_,r_12__2_,r_12__1_,r_12__0_,r_13__15_,r_13__14_,
  r_13__13_,r_13__12_,r_13__11_,r_13__10_,r_13__9_,r_13__8_,r_13__7_,r_13__6_,
  r_13__5_,r_13__4_,r_13__3_,r_13__2_,r_13__1_,r_13__0_,r_14__15_,r_14__14_,r_14__13_,
  r_14__12_,r_14__11_,r_14__10_,r_14__9_,r_14__8_,r_14__7_,r_14__6_,r_14__5_,r_14__4_,
  r_14__3_,r_14__2_,r_14__1_,r_14__0_,r_15__15_,r_15__14_,r_15__13_,r_15__12_,
  r_15__11_,r_15__10_,r_15__9_,r_15__8_,r_15__7_,r_15__6_,r_15__5_,r_15__4_,r_15__3_,
  r_15__2_,r_15__1_,r_15__0_,r_16__15_,r_16__14_,r_16__13_,r_16__12_,r_16__11_,
  r_16__10_,r_16__9_,r_16__8_,r_16__7_,r_16__6_,r_16__5_,r_16__4_,r_16__3_,r_16__2_,
  r_16__1_,r_16__0_,r_17__15_,r_17__14_,r_17__13_,r_17__12_,r_17__11_,r_17__10_,
  r_17__9_,r_17__8_,r_17__7_,r_17__6_,r_17__5_,r_17__4_,r_17__3_,r_17__2_,r_17__1_,
  r_17__0_,r_18__15_,r_18__14_,r_18__13_,r_18__12_,r_18__11_,r_18__10_,r_18__9_,
  r_18__8_,r_18__7_,r_18__6_,r_18__5_,r_18__4_,r_18__3_,r_18__2_,r_18__1_,r_18__0_,
  r_19__15_,r_19__14_,r_19__13_,r_19__12_,r_19__11_,r_19__10_,r_19__9_,r_19__8_,
  r_19__7_,r_19__6_,r_19__5_,r_19__4_,r_19__3_,r_19__2_,r_19__1_,r_19__0_,r_20__15_,
  r_20__14_,r_20__13_,r_20__12_,r_20__11_,r_20__10_,r_20__9_,r_20__8_,r_20__7_,
  r_20__6_,r_20__5_,r_20__4_,r_20__3_,r_20__2_,r_20__1_,r_20__0_,r_21__15_,r_21__14_,
  r_21__13_,r_21__12_,r_21__11_,r_21__10_,r_21__9_,r_21__8_,r_21__7_,r_21__6_,
  r_21__5_,r_21__4_,r_21__3_,r_21__2_,r_21__1_,r_21__0_,r_22__15_,r_22__14_,r_22__13_,
  r_22__12_,r_22__11_,r_22__10_,r_22__9_,r_22__8_,r_22__7_,r_22__6_,r_22__5_,r_22__4_,
  r_22__3_,r_22__2_,r_22__1_,r_22__0_,r_23__15_,r_23__14_,r_23__13_,r_23__12_,
  r_23__11_,r_23__10_,r_23__9_,r_23__8_,r_23__7_,r_23__6_,r_23__5_,r_23__4_,r_23__3_,
  r_23__2_,r_23__1_,r_23__0_,r_24__15_,r_24__14_,r_24__13_,r_24__12_,r_24__11_,
  r_24__10_,r_24__9_,r_24__8_,r_24__7_,r_24__6_,r_24__5_,r_24__4_,r_24__3_,r_24__2_,
  r_24__1_,r_24__0_,r_25__15_,r_25__14_,r_25__13_,r_25__12_,r_25__11_,r_25__10_,
  r_25__9_,r_25__8_,r_25__7_,r_25__6_,r_25__5_,r_25__4_,r_25__3_,r_25__2_,r_25__1_,
  r_25__0_,r_26__15_,r_26__14_,r_26__13_,r_26__12_,r_26__11_,r_26__10_,r_26__9_,
  r_26__8_,r_26__7_,r_26__6_,r_26__5_,r_26__4_,r_26__3_,r_26__2_,r_26__1_,r_26__0_,
  r_27__15_,r_27__14_,r_27__13_,r_27__12_,r_27__11_,r_27__10_,r_27__9_,r_27__8_,
  r_27__7_,r_27__6_,r_27__5_,r_27__4_,r_27__3_,r_27__2_,r_27__1_,r_27__0_,r_28__15_,
  r_28__14_,r_28__13_,r_28__12_,r_28__11_,r_28__10_,r_28__9_,r_28__8_,r_28__7_,
  r_28__6_,r_28__5_,r_28__4_,r_28__3_,r_28__2_,r_28__1_,r_28__0_,r_29__15_,r_29__14_,
  r_29__13_,r_29__12_,r_29__11_,r_29__10_,r_29__9_,r_29__8_,r_29__7_,r_29__6_,
  r_29__5_,r_29__4_,r_29__3_,r_29__2_,r_29__1_,r_29__0_,r_30__15_,r_30__14_,r_30__13_,
  r_30__12_,r_30__11_,r_30__10_,r_30__9_,r_30__8_,r_30__7_,r_30__6_,r_30__5_,r_30__4_,
  r_30__3_,r_30__2_,r_30__1_,r_30__0_,r_31__15_,r_31__14_,r_31__13_,r_31__12_,
  r_31__11_,r_31__10_,r_31__9_,r_31__8_,r_31__7_,r_31__6_,r_31__5_,r_31__4_,r_31__3_,
  r_31__2_,r_31__1_,r_31__0_,r_32__15_,r_32__14_,r_32__13_,r_32__12_,r_32__11_,
  r_32__10_,r_32__9_,r_32__8_,r_32__7_,r_32__6_,r_32__5_,r_32__4_,r_32__3_,r_32__2_,
  r_32__1_,r_32__0_,r_33__15_,r_33__14_,r_33__13_,r_33__12_,r_33__11_,r_33__10_,
  r_33__9_,r_33__8_,r_33__7_,r_33__6_,r_33__5_,r_33__4_,r_33__3_,r_33__2_,r_33__1_,
  r_33__0_,r_34__15_,r_34__14_,r_34__13_,r_34__12_,r_34__11_,r_34__10_,r_34__9_,
  r_34__8_,r_34__7_,r_34__6_,r_34__5_,r_34__4_,r_34__3_,r_34__2_,r_34__1_,r_34__0_,
  r_35__15_,r_35__14_,r_35__13_,r_35__12_,r_35__11_,r_35__10_,r_35__9_,r_35__8_,
  r_35__7_,r_35__6_,r_35__5_,r_35__4_,r_35__3_,r_35__2_,r_35__1_,r_35__0_,r_36__15_,
  r_36__14_,r_36__13_,r_36__12_,r_36__11_,r_36__10_,r_36__9_,r_36__8_,r_36__7_,
  r_36__6_,r_36__5_,r_36__4_,r_36__3_,r_36__2_,r_36__1_,r_36__0_,r_37__15_,r_37__14_,
  r_37__13_,r_37__12_,r_37__11_,r_37__10_,r_37__9_,r_37__8_,r_37__7_,r_37__6_,
  r_37__5_,r_37__4_,r_37__3_,r_37__2_,r_37__1_,r_37__0_,r_38__15_,r_38__14_,r_38__13_,
  r_38__12_,r_38__11_,r_38__10_,r_38__9_,r_38__8_,r_38__7_,r_38__6_,r_38__5_,r_38__4_,
  r_38__3_,r_38__2_,r_38__1_,r_38__0_,r_39__15_,r_39__14_,r_39__13_,r_39__12_,
  r_39__11_,r_39__10_,r_39__9_,r_39__8_,r_39__7_,r_39__6_,r_39__5_,r_39__4_,r_39__3_,
  r_39__2_,r_39__1_,r_39__0_,r_40__15_,r_40__14_,r_40__13_,r_40__12_,r_40__11_,
  r_40__10_,r_40__9_,r_40__8_,r_40__7_,r_40__6_,r_40__5_,r_40__4_,r_40__3_,r_40__2_,
  r_40__1_,r_40__0_,r_41__15_,r_41__14_,r_41__13_,r_41__12_,r_41__11_,r_41__10_,
  r_41__9_,r_41__8_,r_41__7_,r_41__6_,r_41__5_,r_41__4_,r_41__3_,r_41__2_,r_41__1_,
  r_41__0_,r_42__15_,r_42__14_,r_42__13_,r_42__12_,r_42__11_,r_42__10_,r_42__9_,
  r_42__8_,r_42__7_,r_42__6_,r_42__5_,r_42__4_,r_42__3_,r_42__2_,r_42__1_,r_42__0_,
  r_43__15_,r_43__14_,r_43__13_,r_43__12_,r_43__11_,r_43__10_,r_43__9_,r_43__8_,
  r_43__7_,r_43__6_,r_43__5_,r_43__4_,r_43__3_,r_43__2_,r_43__1_,r_43__0_,r_44__15_,
  r_44__14_,r_44__13_,r_44__12_,r_44__11_,r_44__10_,r_44__9_,r_44__8_,r_44__7_,
  r_44__6_,r_44__5_,r_44__4_,r_44__3_,r_44__2_,r_44__1_,r_44__0_,r_45__15_,r_45__14_,
  r_45__13_,r_45__12_,r_45__11_,r_45__10_,r_45__9_,r_45__8_,r_45__7_,r_45__6_,
  r_45__5_,r_45__4_,r_45__3_,r_45__2_,r_45__1_,r_45__0_,r_46__15_,r_46__14_,r_46__13_,
  r_46__12_,r_46__11_,r_46__10_,r_46__9_,r_46__8_,r_46__7_,r_46__6_,r_46__5_,r_46__4_,
  r_46__3_,r_46__2_,r_46__1_,r_46__0_,r_47__15_,r_47__14_,r_47__13_,r_47__12_,
  r_47__11_,r_47__10_,r_47__9_,r_47__8_,r_47__7_,r_47__6_,r_47__5_,r_47__4_,r_47__3_,
  r_47__2_,r_47__1_,r_47__0_,r_48__15_,r_48__14_,r_48__13_,r_48__12_,r_48__11_,
  r_48__10_,r_48__9_,r_48__8_,r_48__7_,r_48__6_,r_48__5_,r_48__4_,r_48__3_,r_48__2_,
  r_48__1_,r_48__0_,r_49__15_,r_49__14_,r_49__13_,r_49__12_,r_49__11_,r_49__10_,
  r_49__9_,r_49__8_,r_49__7_,r_49__6_,r_49__5_,r_49__4_,r_49__3_,r_49__2_,r_49__1_,
  r_49__0_,r_50__15_,r_50__14_,r_50__13_,r_50__12_,r_50__11_,r_50__10_,r_50__9_,
  r_50__8_,r_50__7_,r_50__6_,r_50__5_,r_50__4_,r_50__3_,r_50__2_,r_50__1_,r_50__0_,
  r_51__15_,r_51__14_,r_51__13_,r_51__12_,r_51__11_,r_51__10_,r_51__9_,r_51__8_,
  r_51__7_,r_51__6_,r_51__5_,r_51__4_,r_51__3_,r_51__2_,r_51__1_,r_51__0_,r_52__15_,
  r_52__14_,r_52__13_,r_52__12_,r_52__11_,r_52__10_,r_52__9_,r_52__8_,r_52__7_,
  r_52__6_,r_52__5_,r_52__4_,r_52__3_,r_52__2_,r_52__1_,r_52__0_,r_53__15_,r_53__14_,
  r_53__13_,r_53__12_,r_53__11_,r_53__10_,r_53__9_,r_53__8_,r_53__7_,r_53__6_,
  r_53__5_,r_53__4_,r_53__3_,r_53__2_,r_53__1_,r_53__0_,r_54__15_,r_54__14_,r_54__13_,
  r_54__12_,r_54__11_,r_54__10_,r_54__9_,r_54__8_,r_54__7_,r_54__6_,r_54__5_,r_54__4_,
  r_54__3_,r_54__2_,r_54__1_,r_54__0_,r_55__15_,r_55__14_,r_55__13_,r_55__12_,
  r_55__11_,r_55__10_,r_55__9_,r_55__8_,r_55__7_,r_55__6_,r_55__5_,r_55__4_,r_55__3_,
  r_55__2_,r_55__1_,r_55__0_,r_56__15_,r_56__14_,r_56__13_,r_56__12_,r_56__11_,
  r_56__10_,r_56__9_,r_56__8_,r_56__7_,r_56__6_,r_56__5_,r_56__4_,r_56__3_,r_56__2_,
  r_56__1_,r_56__0_,r_57__15_,r_57__14_,r_57__13_,r_57__12_,r_57__11_,r_57__10_,
  r_57__9_,r_57__8_,r_57__7_,r_57__6_,r_57__5_,r_57__4_,r_57__3_,r_57__2_,r_57__1_,
  r_57__0_,r_58__15_,r_58__14_,r_58__13_,r_58__12_,r_58__11_,r_58__10_,r_58__9_,
  r_58__8_,r_58__7_,r_58__6_,r_58__5_,r_58__4_,r_58__3_,r_58__2_,r_58__1_,r_58__0_,
  r_59__15_,r_59__14_,r_59__13_,r_59__12_,r_59__11_,r_59__10_,r_59__9_,r_59__8_,
  r_59__7_,r_59__6_,r_59__5_,r_59__4_,r_59__3_,r_59__2_,r_59__1_,r_59__0_,r_60__15_,
  r_60__14_,r_60__13_,r_60__12_,r_60__11_,r_60__10_,r_60__9_,r_60__8_,r_60__7_,
  r_60__6_,r_60__5_,r_60__4_,r_60__3_,r_60__2_,r_60__1_,r_60__0_,r_61__15_,r_61__14_,
  r_61__13_,r_61__12_,r_61__11_,r_61__10_,r_61__9_,r_61__8_,r_61__7_,r_61__6_,
  r_61__5_,r_61__4_,r_61__3_,r_61__2_,r_61__1_,r_61__0_,r_62__15_,r_62__14_,r_62__13_,
  r_62__12_,r_62__11_,r_62__10_,r_62__9_,r_62__8_,r_62__7_,r_62__6_,r_62__5_,r_62__4_,
  r_62__3_,r_62__2_,r_62__1_,r_62__0_,r_63__15_,r_63__14_,r_63__13_,r_63__12_,
  r_63__11_,r_63__10_,r_63__9_,r_63__8_,r_63__7_,r_63__6_,r_63__5_,r_63__4_,r_63__3_,
  r_63__2_,r_63__1_,r_63__0_;
  assign N128 = sel_i[1] & sel_i[0];
  assign N130 = N129 & N132;
  assign N133 = sel_i[3] & sel_i[2];
  assign N135 = N134 & N137;
  assign N138 = sel_i[5] & sel_i[4];
  assign N140 = N139 & N142;
  assign N143 = sel_i[7] & sel_i[6];
  assign N145 = N144 & N147;
  assign N148 = sel_i[9] & sel_i[8];
  assign N150 = N149 & N152;
  assign N153 = sel_i[11] & sel_i[10];
  assign N155 = N154 & N157;
  assign N158 = sel_i[13] & sel_i[12];
  assign N160 = N159 & N162;
  assign N163 = sel_i[15] & sel_i[14];
  assign N165 = N164 & N167;
  assign N168 = sel_i[17] & sel_i[16];
  assign N170 = N169 & N172;
  assign N173 = sel_i[19] & sel_i[18];
  assign N175 = N174 & N177;
  assign N178 = sel_i[21] & sel_i[20];
  assign N180 = N179 & N182;
  assign N183 = sel_i[23] & sel_i[22];
  assign N185 = N184 & N187;
  assign N188 = sel_i[25] & sel_i[24];
  assign N190 = N189 & N192;
  assign N193 = sel_i[27] & sel_i[26];
  assign N195 = N194 & N197;
  assign N198 = sel_i[29] & sel_i[28];
  assign N200 = N199 & N202;
  assign N203 = sel_i[31] & sel_i[30];
  assign N205 = N204 & N207;
  assign N208 = sel_i[33] & sel_i[32];
  assign N210 = N209 & N212;
  assign N213 = sel_i[35] & sel_i[34];
  assign N215 = N214 & N217;
  assign N218 = sel_i[37] & sel_i[36];
  assign N220 = N219 & N222;
  assign N223 = sel_i[39] & sel_i[38];
  assign N225 = N224 & N227;
  assign N228 = sel_i[41] & sel_i[40];
  assign N230 = N229 & N232;
  assign N233 = sel_i[43] & sel_i[42];
  assign N235 = N234 & N237;
  assign N238 = sel_i[45] & sel_i[44];
  assign N240 = N239 & N242;
  assign N243 = sel_i[47] & sel_i[46];
  assign N245 = N244 & N247;
  assign N248 = sel_i[49] & sel_i[48];
  assign N250 = N249 & N252;
  assign N253 = sel_i[51] & sel_i[50];
  assign N255 = N254 & N257;
  assign N258 = sel_i[53] & sel_i[52];
  assign N260 = N259 & N262;
  assign N263 = sel_i[55] & sel_i[54];
  assign N265 = N264 & N267;
  assign N268 = sel_i[57] & sel_i[56];
  assign N270 = N269 & N272;
  assign N273 = sel_i[59] & sel_i[58];
  assign N275 = N274 & N277;
  assign N278 = sel_i[61] & sel_i[60];
  assign N280 = N279 & N282;
  assign N283 = sel_i[63] & sel_i[62];
  assign N285 = N284 & N287;
  assign N288 = sel_i[65] & sel_i[64];
  assign N290 = N289 & N292;
  assign N293 = sel_i[67] & sel_i[66];
  assign N295 = N294 & N297;
  assign N298 = sel_i[69] & sel_i[68];
  assign N300 = N299 & N302;
  assign N303 = sel_i[71] & sel_i[70];
  assign N305 = N304 & N307;
  assign N308 = sel_i[73] & sel_i[72];
  assign N310 = N309 & N312;
  assign N313 = sel_i[75] & sel_i[74];
  assign N315 = N314 & N317;
  assign N318 = sel_i[77] & sel_i[76];
  assign N320 = N319 & N322;
  assign N323 = sel_i[79] & sel_i[78];
  assign N325 = N324 & N327;
  assign N328 = sel_i[81] & sel_i[80];
  assign N330 = N329 & N332;
  assign N333 = sel_i[83] & sel_i[82];
  assign N335 = N334 & N337;
  assign N338 = sel_i[85] & sel_i[84];
  assign N340 = N339 & N342;
  assign N343 = sel_i[87] & sel_i[86];
  assign N345 = N344 & N347;
  assign N348 = sel_i[89] & sel_i[88];
  assign N350 = N349 & N352;
  assign N353 = sel_i[91] & sel_i[90];
  assign N355 = N354 & N357;
  assign N358 = sel_i[93] & sel_i[92];
  assign N360 = N359 & N362;
  assign N363 = sel_i[95] & sel_i[94];
  assign N365 = N364 & N367;
  assign N368 = sel_i[97] & sel_i[96];
  assign N370 = N369 & N372;
  assign N373 = sel_i[99] & sel_i[98];
  assign N375 = N374 & N377;
  assign N378 = sel_i[101] & sel_i[100];
  assign N380 = N379 & N382;
  assign N383 = sel_i[103] & sel_i[102];
  assign N385 = N384 & N387;
  assign N388 = sel_i[105] & sel_i[104];
  assign N390 = N389 & N392;
  assign N393 = sel_i[107] & sel_i[106];
  assign N395 = N394 & N397;
  assign N398 = sel_i[109] & sel_i[108];
  assign N400 = N399 & N402;
  assign N403 = sel_i[111] & sel_i[110];
  assign N405 = N404 & N407;
  assign N408 = sel_i[113] & sel_i[112];
  assign N410 = N409 & N412;
  assign N413 = sel_i[115] & sel_i[114];
  assign N415 = N414 & N417;
  assign N418 = sel_i[117] & sel_i[116];
  assign N420 = N419 & N422;
  assign N423 = sel_i[119] & sel_i[118];
  assign N425 = N424 & N427;
  assign N428 = sel_i[121] & sel_i[120];
  assign N430 = N429 & N432;
  assign N433 = sel_i[123] & sel_i[122];
  assign N435 = N434 & N437;
  assign N438 = sel_i[125] & sel_i[124];
  assign N440 = N439 & N442;
  assign N443 = sel_i[127] & sel_i[126];
  assign N445 = N444 & N447;
  assign N132 = ~sel_i[0];
  assign N137 = ~sel_i[2];
  assign N142 = ~sel_i[4];
  assign N147 = ~sel_i[6];
  assign N152 = ~sel_i[8];
  assign N157 = ~sel_i[10];
  assign N162 = ~sel_i[12];
  assign N167 = ~sel_i[14];
  assign N172 = ~sel_i[16];
  assign N177 = ~sel_i[18];
  assign N182 = ~sel_i[20];
  assign N187 = ~sel_i[22];
  assign N192 = ~sel_i[24];
  assign N197 = ~sel_i[26];
  assign N202 = ~sel_i[28];
  assign N207 = ~sel_i[30];
  assign N212 = ~sel_i[32];
  assign N217 = ~sel_i[34];
  assign N222 = ~sel_i[36];
  assign N227 = ~sel_i[38];
  assign N232 = ~sel_i[40];
  assign N237 = ~sel_i[42];
  assign N242 = ~sel_i[44];
  assign N247 = ~sel_i[46];
  assign N252 = ~sel_i[48];
  assign N257 = ~sel_i[50];
  assign N262 = ~sel_i[52];
  assign N267 = ~sel_i[54];
  assign N272 = ~sel_i[56];
  assign N277 = ~sel_i[58];
  assign N282 = ~sel_i[60];
  assign N287 = ~sel_i[62];
  assign N292 = ~sel_i[64];
  assign N297 = ~sel_i[66];
  assign N302 = ~sel_i[68];
  assign N307 = ~sel_i[70];
  assign N312 = ~sel_i[72];
  assign N317 = ~sel_i[74];
  assign N322 = ~sel_i[76];
  assign N327 = ~sel_i[78];
  assign N332 = ~sel_i[80];
  assign N337 = ~sel_i[82];
  assign N342 = ~sel_i[84];
  assign N347 = ~sel_i[86];
  assign N352 = ~sel_i[88];
  assign N357 = ~sel_i[90];
  assign N362 = ~sel_i[92];
  assign N367 = ~sel_i[94];
  assign N372 = ~sel_i[96];
  assign N377 = ~sel_i[98];
  assign N382 = ~sel_i[100];
  assign N387 = ~sel_i[102];
  assign N392 = ~sel_i[104];
  assign N397 = ~sel_i[106];
  assign N402 = ~sel_i[108];
  assign N407 = ~sel_i[110];
  assign N412 = ~sel_i[112];
  assign N417 = ~sel_i[114];
  assign N422 = ~sel_i[116];
  assign N427 = ~sel_i[118];
  assign N432 = ~sel_i[120];
  assign N437 = ~sel_i[122];
  assign N442 = ~sel_i[124];
  assign N447 = ~sel_i[126];
  assign { r_n_0__15_, r_n_0__14_, r_n_0__13_, r_n_0__12_, r_n_0__11_, r_n_0__10_, r_n_0__9_, r_n_0__8_, r_n_0__7_, r_n_0__6_, r_n_0__5_, r_n_0__4_, r_n_0__3_, r_n_0__2_, r_n_0__1_, r_n_0__0_ } = (N0)? { r_1__15_, r_1__14_, r_1__13_, r_1__12_, r_1__11_, r_1__10_, r_1__9_, r_1__8_, r_1__7_, r_1__6_, r_1__5_, r_1__4_, r_1__3_, r_1__2_, r_1__1_, r_1__0_ } : 
                                                                                                                                                                                                    (N1)? data_i : 1'b0;
  assign N0 = sel_i[0];
  assign N1 = N132;
  assign { r_n_1__15_, r_n_1__14_, r_n_1__13_, r_n_1__12_, r_n_1__11_, r_n_1__10_, r_n_1__9_, r_n_1__8_, r_n_1__7_, r_n_1__6_, r_n_1__5_, r_n_1__4_, r_n_1__3_, r_n_1__2_, r_n_1__1_, r_n_1__0_ } = (N2)? { r_2__15_, r_2__14_, r_2__13_, r_2__12_, r_2__11_, r_2__10_, r_2__9_, r_2__8_, r_2__7_, r_2__6_, r_2__5_, r_2__4_, r_2__3_, r_2__2_, r_2__1_, r_2__0_ } : 
                                                                                                                                                                                                    (N3)? data_i : 1'b0;
  assign N2 = sel_i[2];
  assign N3 = N137;
  assign { r_n_2__15_, r_n_2__14_, r_n_2__13_, r_n_2__12_, r_n_2__11_, r_n_2__10_, r_n_2__9_, r_n_2__8_, r_n_2__7_, r_n_2__6_, r_n_2__5_, r_n_2__4_, r_n_2__3_, r_n_2__2_, r_n_2__1_, r_n_2__0_ } = (N4)? { r_3__15_, r_3__14_, r_3__13_, r_3__12_, r_3__11_, r_3__10_, r_3__9_, r_3__8_, r_3__7_, r_3__6_, r_3__5_, r_3__4_, r_3__3_, r_3__2_, r_3__1_, r_3__0_ } : 
                                                                                                                                                                                                    (N5)? data_i : 1'b0;
  assign N4 = sel_i[4];
  assign N5 = N142;
  assign { r_n_3__15_, r_n_3__14_, r_n_3__13_, r_n_3__12_, r_n_3__11_, r_n_3__10_, r_n_3__9_, r_n_3__8_, r_n_3__7_, r_n_3__6_, r_n_3__5_, r_n_3__4_, r_n_3__3_, r_n_3__2_, r_n_3__1_, r_n_3__0_ } = (N6)? { r_4__15_, r_4__14_, r_4__13_, r_4__12_, r_4__11_, r_4__10_, r_4__9_, r_4__8_, r_4__7_, r_4__6_, r_4__5_, r_4__4_, r_4__3_, r_4__2_, r_4__1_, r_4__0_ } : 
                                                                                                                                                                                                    (N7)? data_i : 1'b0;
  assign N6 = sel_i[6];
  assign N7 = N147;
  assign { r_n_4__15_, r_n_4__14_, r_n_4__13_, r_n_4__12_, r_n_4__11_, r_n_4__10_, r_n_4__9_, r_n_4__8_, r_n_4__7_, r_n_4__6_, r_n_4__5_, r_n_4__4_, r_n_4__3_, r_n_4__2_, r_n_4__1_, r_n_4__0_ } = (N8)? { r_5__15_, r_5__14_, r_5__13_, r_5__12_, r_5__11_, r_5__10_, r_5__9_, r_5__8_, r_5__7_, r_5__6_, r_5__5_, r_5__4_, r_5__3_, r_5__2_, r_5__1_, r_5__0_ } : 
                                                                                                                                                                                                    (N9)? data_i : 1'b0;
  assign N8 = sel_i[8];
  assign N9 = N152;
  assign { r_n_5__15_, r_n_5__14_, r_n_5__13_, r_n_5__12_, r_n_5__11_, r_n_5__10_, r_n_5__9_, r_n_5__8_, r_n_5__7_, r_n_5__6_, r_n_5__5_, r_n_5__4_, r_n_5__3_, r_n_5__2_, r_n_5__1_, r_n_5__0_ } = (N10)? { r_6__15_, r_6__14_, r_6__13_, r_6__12_, r_6__11_, r_6__10_, r_6__9_, r_6__8_, r_6__7_, r_6__6_, r_6__5_, r_6__4_, r_6__3_, r_6__2_, r_6__1_, r_6__0_ } : 
                                                                                                                                                                                                    (N11)? data_i : 1'b0;
  assign N10 = sel_i[10];
  assign N11 = N157;
  assign { r_n_6__15_, r_n_6__14_, r_n_6__13_, r_n_6__12_, r_n_6__11_, r_n_6__10_, r_n_6__9_, r_n_6__8_, r_n_6__7_, r_n_6__6_, r_n_6__5_, r_n_6__4_, r_n_6__3_, r_n_6__2_, r_n_6__1_, r_n_6__0_ } = (N12)? { r_7__15_, r_7__14_, r_7__13_, r_7__12_, r_7__11_, r_7__10_, r_7__9_, r_7__8_, r_7__7_, r_7__6_, r_7__5_, r_7__4_, r_7__3_, r_7__2_, r_7__1_, r_7__0_ } : 
                                                                                                                                                                                                    (N13)? data_i : 1'b0;
  assign N12 = sel_i[12];
  assign N13 = N162;
  assign { r_n_7__15_, r_n_7__14_, r_n_7__13_, r_n_7__12_, r_n_7__11_, r_n_7__10_, r_n_7__9_, r_n_7__8_, r_n_7__7_, r_n_7__6_, r_n_7__5_, r_n_7__4_, r_n_7__3_, r_n_7__2_, r_n_7__1_, r_n_7__0_ } = (N14)? { r_8__15_, r_8__14_, r_8__13_, r_8__12_, r_8__11_, r_8__10_, r_8__9_, r_8__8_, r_8__7_, r_8__6_, r_8__5_, r_8__4_, r_8__3_, r_8__2_, r_8__1_, r_8__0_ } : 
                                                                                                                                                                                                    (N15)? data_i : 1'b0;
  assign N14 = sel_i[14];
  assign N15 = N167;
  assign { r_n_8__15_, r_n_8__14_, r_n_8__13_, r_n_8__12_, r_n_8__11_, r_n_8__10_, r_n_8__9_, r_n_8__8_, r_n_8__7_, r_n_8__6_, r_n_8__5_, r_n_8__4_, r_n_8__3_, r_n_8__2_, r_n_8__1_, r_n_8__0_ } = (N16)? { r_9__15_, r_9__14_, r_9__13_, r_9__12_, r_9__11_, r_9__10_, r_9__9_, r_9__8_, r_9__7_, r_9__6_, r_9__5_, r_9__4_, r_9__3_, r_9__2_, r_9__1_, r_9__0_ } : 
                                                                                                                                                                                                    (N17)? data_i : 1'b0;
  assign N16 = sel_i[16];
  assign N17 = N172;
  assign { r_n_9__15_, r_n_9__14_, r_n_9__13_, r_n_9__12_, r_n_9__11_, r_n_9__10_, r_n_9__9_, r_n_9__8_, r_n_9__7_, r_n_9__6_, r_n_9__5_, r_n_9__4_, r_n_9__3_, r_n_9__2_, r_n_9__1_, r_n_9__0_ } = (N18)? { r_10__15_, r_10__14_, r_10__13_, r_10__12_, r_10__11_, r_10__10_, r_10__9_, r_10__8_, r_10__7_, r_10__6_, r_10__5_, r_10__4_, r_10__3_, r_10__2_, r_10__1_, r_10__0_ } : 
                                                                                                                                                                                                    (N19)? data_i : 1'b0;
  assign N18 = sel_i[18];
  assign N19 = N177;
  assign { r_n_10__15_, r_n_10__14_, r_n_10__13_, r_n_10__12_, r_n_10__11_, r_n_10__10_, r_n_10__9_, r_n_10__8_, r_n_10__7_, r_n_10__6_, r_n_10__5_, r_n_10__4_, r_n_10__3_, r_n_10__2_, r_n_10__1_, r_n_10__0_ } = (N20)? { r_11__15_, r_11__14_, r_11__13_, r_11__12_, r_11__11_, r_11__10_, r_11__9_, r_11__8_, r_11__7_, r_11__6_, r_11__5_, r_11__4_, r_11__3_, r_11__2_, r_11__1_, r_11__0_ } : 
                                                                                                                                                                                                                    (N21)? data_i : 1'b0;
  assign N20 = sel_i[20];
  assign N21 = N182;
  assign { r_n_11__15_, r_n_11__14_, r_n_11__13_, r_n_11__12_, r_n_11__11_, r_n_11__10_, r_n_11__9_, r_n_11__8_, r_n_11__7_, r_n_11__6_, r_n_11__5_, r_n_11__4_, r_n_11__3_, r_n_11__2_, r_n_11__1_, r_n_11__0_ } = (N22)? { r_12__15_, r_12__14_, r_12__13_, r_12__12_, r_12__11_, r_12__10_, r_12__9_, r_12__8_, r_12__7_, r_12__6_, r_12__5_, r_12__4_, r_12__3_, r_12__2_, r_12__1_, r_12__0_ } : 
                                                                                                                                                                                                                    (N23)? data_i : 1'b0;
  assign N22 = sel_i[22];
  assign N23 = N187;
  assign { r_n_12__15_, r_n_12__14_, r_n_12__13_, r_n_12__12_, r_n_12__11_, r_n_12__10_, r_n_12__9_, r_n_12__8_, r_n_12__7_, r_n_12__6_, r_n_12__5_, r_n_12__4_, r_n_12__3_, r_n_12__2_, r_n_12__1_, r_n_12__0_ } = (N24)? { r_13__15_, r_13__14_, r_13__13_, r_13__12_, r_13__11_, r_13__10_, r_13__9_, r_13__8_, r_13__7_, r_13__6_, r_13__5_, r_13__4_, r_13__3_, r_13__2_, r_13__1_, r_13__0_ } : 
                                                                                                                                                                                                                    (N25)? data_i : 1'b0;
  assign N24 = sel_i[24];
  assign N25 = N192;
  assign { r_n_13__15_, r_n_13__14_, r_n_13__13_, r_n_13__12_, r_n_13__11_, r_n_13__10_, r_n_13__9_, r_n_13__8_, r_n_13__7_, r_n_13__6_, r_n_13__5_, r_n_13__4_, r_n_13__3_, r_n_13__2_, r_n_13__1_, r_n_13__0_ } = (N26)? { r_14__15_, r_14__14_, r_14__13_, r_14__12_, r_14__11_, r_14__10_, r_14__9_, r_14__8_, r_14__7_, r_14__6_, r_14__5_, r_14__4_, r_14__3_, r_14__2_, r_14__1_, r_14__0_ } : 
                                                                                                                                                                                                                    (N27)? data_i : 1'b0;
  assign N26 = sel_i[26];
  assign N27 = N197;
  assign { r_n_14__15_, r_n_14__14_, r_n_14__13_, r_n_14__12_, r_n_14__11_, r_n_14__10_, r_n_14__9_, r_n_14__8_, r_n_14__7_, r_n_14__6_, r_n_14__5_, r_n_14__4_, r_n_14__3_, r_n_14__2_, r_n_14__1_, r_n_14__0_ } = (N28)? { r_15__15_, r_15__14_, r_15__13_, r_15__12_, r_15__11_, r_15__10_, r_15__9_, r_15__8_, r_15__7_, r_15__6_, r_15__5_, r_15__4_, r_15__3_, r_15__2_, r_15__1_, r_15__0_ } : 
                                                                                                                                                                                                                    (N29)? data_i : 1'b0;
  assign N28 = sel_i[28];
  assign N29 = N202;
  assign { r_n_15__15_, r_n_15__14_, r_n_15__13_, r_n_15__12_, r_n_15__11_, r_n_15__10_, r_n_15__9_, r_n_15__8_, r_n_15__7_, r_n_15__6_, r_n_15__5_, r_n_15__4_, r_n_15__3_, r_n_15__2_, r_n_15__1_, r_n_15__0_ } = (N30)? { r_16__15_, r_16__14_, r_16__13_, r_16__12_, r_16__11_, r_16__10_, r_16__9_, r_16__8_, r_16__7_, r_16__6_, r_16__5_, r_16__4_, r_16__3_, r_16__2_, r_16__1_, r_16__0_ } : 
                                                                                                                                                                                                                    (N31)? data_i : 1'b0;
  assign N30 = sel_i[30];
  assign N31 = N207;
  assign { r_n_16__15_, r_n_16__14_, r_n_16__13_, r_n_16__12_, r_n_16__11_, r_n_16__10_, r_n_16__9_, r_n_16__8_, r_n_16__7_, r_n_16__6_, r_n_16__5_, r_n_16__4_, r_n_16__3_, r_n_16__2_, r_n_16__1_, r_n_16__0_ } = (N32)? { r_17__15_, r_17__14_, r_17__13_, r_17__12_, r_17__11_, r_17__10_, r_17__9_, r_17__8_, r_17__7_, r_17__6_, r_17__5_, r_17__4_, r_17__3_, r_17__2_, r_17__1_, r_17__0_ } : 
                                                                                                                                                                                                                    (N33)? data_i : 1'b0;
  assign N32 = sel_i[32];
  assign N33 = N212;
  assign { r_n_17__15_, r_n_17__14_, r_n_17__13_, r_n_17__12_, r_n_17__11_, r_n_17__10_, r_n_17__9_, r_n_17__8_, r_n_17__7_, r_n_17__6_, r_n_17__5_, r_n_17__4_, r_n_17__3_, r_n_17__2_, r_n_17__1_, r_n_17__0_ } = (N34)? { r_18__15_, r_18__14_, r_18__13_, r_18__12_, r_18__11_, r_18__10_, r_18__9_, r_18__8_, r_18__7_, r_18__6_, r_18__5_, r_18__4_, r_18__3_, r_18__2_, r_18__1_, r_18__0_ } : 
                                                                                                                                                                                                                    (N35)? data_i : 1'b0;
  assign N34 = sel_i[34];
  assign N35 = N217;
  assign { r_n_18__15_, r_n_18__14_, r_n_18__13_, r_n_18__12_, r_n_18__11_, r_n_18__10_, r_n_18__9_, r_n_18__8_, r_n_18__7_, r_n_18__6_, r_n_18__5_, r_n_18__4_, r_n_18__3_, r_n_18__2_, r_n_18__1_, r_n_18__0_ } = (N36)? { r_19__15_, r_19__14_, r_19__13_, r_19__12_, r_19__11_, r_19__10_, r_19__9_, r_19__8_, r_19__7_, r_19__6_, r_19__5_, r_19__4_, r_19__3_, r_19__2_, r_19__1_, r_19__0_ } : 
                                                                                                                                                                                                                    (N37)? data_i : 1'b0;
  assign N36 = sel_i[36];
  assign N37 = N222;
  assign { r_n_19__15_, r_n_19__14_, r_n_19__13_, r_n_19__12_, r_n_19__11_, r_n_19__10_, r_n_19__9_, r_n_19__8_, r_n_19__7_, r_n_19__6_, r_n_19__5_, r_n_19__4_, r_n_19__3_, r_n_19__2_, r_n_19__1_, r_n_19__0_ } = (N38)? { r_20__15_, r_20__14_, r_20__13_, r_20__12_, r_20__11_, r_20__10_, r_20__9_, r_20__8_, r_20__7_, r_20__6_, r_20__5_, r_20__4_, r_20__3_, r_20__2_, r_20__1_, r_20__0_ } : 
                                                                                                                                                                                                                    (N39)? data_i : 1'b0;
  assign N38 = sel_i[38];
  assign N39 = N227;
  assign { r_n_20__15_, r_n_20__14_, r_n_20__13_, r_n_20__12_, r_n_20__11_, r_n_20__10_, r_n_20__9_, r_n_20__8_, r_n_20__7_, r_n_20__6_, r_n_20__5_, r_n_20__4_, r_n_20__3_, r_n_20__2_, r_n_20__1_, r_n_20__0_ } = (N40)? { r_21__15_, r_21__14_, r_21__13_, r_21__12_, r_21__11_, r_21__10_, r_21__9_, r_21__8_, r_21__7_, r_21__6_, r_21__5_, r_21__4_, r_21__3_, r_21__2_, r_21__1_, r_21__0_ } : 
                                                                                                                                                                                                                    (N41)? data_i : 1'b0;
  assign N40 = sel_i[40];
  assign N41 = N232;
  assign { r_n_21__15_, r_n_21__14_, r_n_21__13_, r_n_21__12_, r_n_21__11_, r_n_21__10_, r_n_21__9_, r_n_21__8_, r_n_21__7_, r_n_21__6_, r_n_21__5_, r_n_21__4_, r_n_21__3_, r_n_21__2_, r_n_21__1_, r_n_21__0_ } = (N42)? { r_22__15_, r_22__14_, r_22__13_, r_22__12_, r_22__11_, r_22__10_, r_22__9_, r_22__8_, r_22__7_, r_22__6_, r_22__5_, r_22__4_, r_22__3_, r_22__2_, r_22__1_, r_22__0_ } : 
                                                                                                                                                                                                                    (N43)? data_i : 1'b0;
  assign N42 = sel_i[42];
  assign N43 = N237;
  assign { r_n_22__15_, r_n_22__14_, r_n_22__13_, r_n_22__12_, r_n_22__11_, r_n_22__10_, r_n_22__9_, r_n_22__8_, r_n_22__7_, r_n_22__6_, r_n_22__5_, r_n_22__4_, r_n_22__3_, r_n_22__2_, r_n_22__1_, r_n_22__0_ } = (N44)? { r_23__15_, r_23__14_, r_23__13_, r_23__12_, r_23__11_, r_23__10_, r_23__9_, r_23__8_, r_23__7_, r_23__6_, r_23__5_, r_23__4_, r_23__3_, r_23__2_, r_23__1_, r_23__0_ } : 
                                                                                                                                                                                                                    (N45)? data_i : 1'b0;
  assign N44 = sel_i[44];
  assign N45 = N242;
  assign { r_n_23__15_, r_n_23__14_, r_n_23__13_, r_n_23__12_, r_n_23__11_, r_n_23__10_, r_n_23__9_, r_n_23__8_, r_n_23__7_, r_n_23__6_, r_n_23__5_, r_n_23__4_, r_n_23__3_, r_n_23__2_, r_n_23__1_, r_n_23__0_ } = (N46)? { r_24__15_, r_24__14_, r_24__13_, r_24__12_, r_24__11_, r_24__10_, r_24__9_, r_24__8_, r_24__7_, r_24__6_, r_24__5_, r_24__4_, r_24__3_, r_24__2_, r_24__1_, r_24__0_ } : 
                                                                                                                                                                                                                    (N47)? data_i : 1'b0;
  assign N46 = sel_i[46];
  assign N47 = N247;
  assign { r_n_24__15_, r_n_24__14_, r_n_24__13_, r_n_24__12_, r_n_24__11_, r_n_24__10_, r_n_24__9_, r_n_24__8_, r_n_24__7_, r_n_24__6_, r_n_24__5_, r_n_24__4_, r_n_24__3_, r_n_24__2_, r_n_24__1_, r_n_24__0_ } = (N48)? { r_25__15_, r_25__14_, r_25__13_, r_25__12_, r_25__11_, r_25__10_, r_25__9_, r_25__8_, r_25__7_, r_25__6_, r_25__5_, r_25__4_, r_25__3_, r_25__2_, r_25__1_, r_25__0_ } : 
                                                                                                                                                                                                                    (N49)? data_i : 1'b0;
  assign N48 = sel_i[48];
  assign N49 = N252;
  assign { r_n_25__15_, r_n_25__14_, r_n_25__13_, r_n_25__12_, r_n_25__11_, r_n_25__10_, r_n_25__9_, r_n_25__8_, r_n_25__7_, r_n_25__6_, r_n_25__5_, r_n_25__4_, r_n_25__3_, r_n_25__2_, r_n_25__1_, r_n_25__0_ } = (N50)? { r_26__15_, r_26__14_, r_26__13_, r_26__12_, r_26__11_, r_26__10_, r_26__9_, r_26__8_, r_26__7_, r_26__6_, r_26__5_, r_26__4_, r_26__3_, r_26__2_, r_26__1_, r_26__0_ } : 
                                                                                                                                                                                                                    (N51)? data_i : 1'b0;
  assign N50 = sel_i[50];
  assign N51 = N257;
  assign { r_n_26__15_, r_n_26__14_, r_n_26__13_, r_n_26__12_, r_n_26__11_, r_n_26__10_, r_n_26__9_, r_n_26__8_, r_n_26__7_, r_n_26__6_, r_n_26__5_, r_n_26__4_, r_n_26__3_, r_n_26__2_, r_n_26__1_, r_n_26__0_ } = (N52)? { r_27__15_, r_27__14_, r_27__13_, r_27__12_, r_27__11_, r_27__10_, r_27__9_, r_27__8_, r_27__7_, r_27__6_, r_27__5_, r_27__4_, r_27__3_, r_27__2_, r_27__1_, r_27__0_ } : 
                                                                                                                                                                                                                    (N53)? data_i : 1'b0;
  assign N52 = sel_i[52];
  assign N53 = N262;
  assign { r_n_27__15_, r_n_27__14_, r_n_27__13_, r_n_27__12_, r_n_27__11_, r_n_27__10_, r_n_27__9_, r_n_27__8_, r_n_27__7_, r_n_27__6_, r_n_27__5_, r_n_27__4_, r_n_27__3_, r_n_27__2_, r_n_27__1_, r_n_27__0_ } = (N54)? { r_28__15_, r_28__14_, r_28__13_, r_28__12_, r_28__11_, r_28__10_, r_28__9_, r_28__8_, r_28__7_, r_28__6_, r_28__5_, r_28__4_, r_28__3_, r_28__2_, r_28__1_, r_28__0_ } : 
                                                                                                                                                                                                                    (N55)? data_i : 1'b0;
  assign N54 = sel_i[54];
  assign N55 = N267;
  assign { r_n_28__15_, r_n_28__14_, r_n_28__13_, r_n_28__12_, r_n_28__11_, r_n_28__10_, r_n_28__9_, r_n_28__8_, r_n_28__7_, r_n_28__6_, r_n_28__5_, r_n_28__4_, r_n_28__3_, r_n_28__2_, r_n_28__1_, r_n_28__0_ } = (N56)? { r_29__15_, r_29__14_, r_29__13_, r_29__12_, r_29__11_, r_29__10_, r_29__9_, r_29__8_, r_29__7_, r_29__6_, r_29__5_, r_29__4_, r_29__3_, r_29__2_, r_29__1_, r_29__0_ } : 
                                                                                                                                                                                                                    (N57)? data_i : 1'b0;
  assign N56 = sel_i[56];
  assign N57 = N272;
  assign { r_n_29__15_, r_n_29__14_, r_n_29__13_, r_n_29__12_, r_n_29__11_, r_n_29__10_, r_n_29__9_, r_n_29__8_, r_n_29__7_, r_n_29__6_, r_n_29__5_, r_n_29__4_, r_n_29__3_, r_n_29__2_, r_n_29__1_, r_n_29__0_ } = (N58)? { r_30__15_, r_30__14_, r_30__13_, r_30__12_, r_30__11_, r_30__10_, r_30__9_, r_30__8_, r_30__7_, r_30__6_, r_30__5_, r_30__4_, r_30__3_, r_30__2_, r_30__1_, r_30__0_ } : 
                                                                                                                                                                                                                    (N59)? data_i : 1'b0;
  assign N58 = sel_i[58];
  assign N59 = N277;
  assign { r_n_30__15_, r_n_30__14_, r_n_30__13_, r_n_30__12_, r_n_30__11_, r_n_30__10_, r_n_30__9_, r_n_30__8_, r_n_30__7_, r_n_30__6_, r_n_30__5_, r_n_30__4_, r_n_30__3_, r_n_30__2_, r_n_30__1_, r_n_30__0_ } = (N60)? { r_31__15_, r_31__14_, r_31__13_, r_31__12_, r_31__11_, r_31__10_, r_31__9_, r_31__8_, r_31__7_, r_31__6_, r_31__5_, r_31__4_, r_31__3_, r_31__2_, r_31__1_, r_31__0_ } : 
                                                                                                                                                                                                                    (N61)? data_i : 1'b0;
  assign N60 = sel_i[60];
  assign N61 = N282;
  assign { r_n_31__15_, r_n_31__14_, r_n_31__13_, r_n_31__12_, r_n_31__11_, r_n_31__10_, r_n_31__9_, r_n_31__8_, r_n_31__7_, r_n_31__6_, r_n_31__5_, r_n_31__4_, r_n_31__3_, r_n_31__2_, r_n_31__1_, r_n_31__0_ } = (N62)? { r_32__15_, r_32__14_, r_32__13_, r_32__12_, r_32__11_, r_32__10_, r_32__9_, r_32__8_, r_32__7_, r_32__6_, r_32__5_, r_32__4_, r_32__3_, r_32__2_, r_32__1_, r_32__0_ } : 
                                                                                                                                                                                                                    (N63)? data_i : 1'b0;
  assign N62 = sel_i[62];
  assign N63 = N287;
  assign { r_n_32__15_, r_n_32__14_, r_n_32__13_, r_n_32__12_, r_n_32__11_, r_n_32__10_, r_n_32__9_, r_n_32__8_, r_n_32__7_, r_n_32__6_, r_n_32__5_, r_n_32__4_, r_n_32__3_, r_n_32__2_, r_n_32__1_, r_n_32__0_ } = (N64)? { r_33__15_, r_33__14_, r_33__13_, r_33__12_, r_33__11_, r_33__10_, r_33__9_, r_33__8_, r_33__7_, r_33__6_, r_33__5_, r_33__4_, r_33__3_, r_33__2_, r_33__1_, r_33__0_ } : 
                                                                                                                                                                                                                    (N65)? data_i : 1'b0;
  assign N64 = sel_i[64];
  assign N65 = N292;
  assign { r_n_33__15_, r_n_33__14_, r_n_33__13_, r_n_33__12_, r_n_33__11_, r_n_33__10_, r_n_33__9_, r_n_33__8_, r_n_33__7_, r_n_33__6_, r_n_33__5_, r_n_33__4_, r_n_33__3_, r_n_33__2_, r_n_33__1_, r_n_33__0_ } = (N66)? { r_34__15_, r_34__14_, r_34__13_, r_34__12_, r_34__11_, r_34__10_, r_34__9_, r_34__8_, r_34__7_, r_34__6_, r_34__5_, r_34__4_, r_34__3_, r_34__2_, r_34__1_, r_34__0_ } : 
                                                                                                                                                                                                                    (N67)? data_i : 1'b0;
  assign N66 = sel_i[66];
  assign N67 = N297;
  assign { r_n_34__15_, r_n_34__14_, r_n_34__13_, r_n_34__12_, r_n_34__11_, r_n_34__10_, r_n_34__9_, r_n_34__8_, r_n_34__7_, r_n_34__6_, r_n_34__5_, r_n_34__4_, r_n_34__3_, r_n_34__2_, r_n_34__1_, r_n_34__0_ } = (N68)? { r_35__15_, r_35__14_, r_35__13_, r_35__12_, r_35__11_, r_35__10_, r_35__9_, r_35__8_, r_35__7_, r_35__6_, r_35__5_, r_35__4_, r_35__3_, r_35__2_, r_35__1_, r_35__0_ } : 
                                                                                                                                                                                                                    (N69)? data_i : 1'b0;
  assign N68 = sel_i[68];
  assign N69 = N302;
  assign { r_n_35__15_, r_n_35__14_, r_n_35__13_, r_n_35__12_, r_n_35__11_, r_n_35__10_, r_n_35__9_, r_n_35__8_, r_n_35__7_, r_n_35__6_, r_n_35__5_, r_n_35__4_, r_n_35__3_, r_n_35__2_, r_n_35__1_, r_n_35__0_ } = (N70)? { r_36__15_, r_36__14_, r_36__13_, r_36__12_, r_36__11_, r_36__10_, r_36__9_, r_36__8_, r_36__7_, r_36__6_, r_36__5_, r_36__4_, r_36__3_, r_36__2_, r_36__1_, r_36__0_ } : 
                                                                                                                                                                                                                    (N71)? data_i : 1'b0;
  assign N70 = sel_i[70];
  assign N71 = N307;
  assign { r_n_36__15_, r_n_36__14_, r_n_36__13_, r_n_36__12_, r_n_36__11_, r_n_36__10_, r_n_36__9_, r_n_36__8_, r_n_36__7_, r_n_36__6_, r_n_36__5_, r_n_36__4_, r_n_36__3_, r_n_36__2_, r_n_36__1_, r_n_36__0_ } = (N72)? { r_37__15_, r_37__14_, r_37__13_, r_37__12_, r_37__11_, r_37__10_, r_37__9_, r_37__8_, r_37__7_, r_37__6_, r_37__5_, r_37__4_, r_37__3_, r_37__2_, r_37__1_, r_37__0_ } : 
                                                                                                                                                                                                                    (N73)? data_i : 1'b0;
  assign N72 = sel_i[72];
  assign N73 = N312;
  assign { r_n_37__15_, r_n_37__14_, r_n_37__13_, r_n_37__12_, r_n_37__11_, r_n_37__10_, r_n_37__9_, r_n_37__8_, r_n_37__7_, r_n_37__6_, r_n_37__5_, r_n_37__4_, r_n_37__3_, r_n_37__2_, r_n_37__1_, r_n_37__0_ } = (N74)? { r_38__15_, r_38__14_, r_38__13_, r_38__12_, r_38__11_, r_38__10_, r_38__9_, r_38__8_, r_38__7_, r_38__6_, r_38__5_, r_38__4_, r_38__3_, r_38__2_, r_38__1_, r_38__0_ } : 
                                                                                                                                                                                                                    (N75)? data_i : 1'b0;
  assign N74 = sel_i[74];
  assign N75 = N317;
  assign { r_n_38__15_, r_n_38__14_, r_n_38__13_, r_n_38__12_, r_n_38__11_, r_n_38__10_, r_n_38__9_, r_n_38__8_, r_n_38__7_, r_n_38__6_, r_n_38__5_, r_n_38__4_, r_n_38__3_, r_n_38__2_, r_n_38__1_, r_n_38__0_ } = (N76)? { r_39__15_, r_39__14_, r_39__13_, r_39__12_, r_39__11_, r_39__10_, r_39__9_, r_39__8_, r_39__7_, r_39__6_, r_39__5_, r_39__4_, r_39__3_, r_39__2_, r_39__1_, r_39__0_ } : 
                                                                                                                                                                                                                    (N77)? data_i : 1'b0;
  assign N76 = sel_i[76];
  assign N77 = N322;
  assign { r_n_39__15_, r_n_39__14_, r_n_39__13_, r_n_39__12_, r_n_39__11_, r_n_39__10_, r_n_39__9_, r_n_39__8_, r_n_39__7_, r_n_39__6_, r_n_39__5_, r_n_39__4_, r_n_39__3_, r_n_39__2_, r_n_39__1_, r_n_39__0_ } = (N78)? { r_40__15_, r_40__14_, r_40__13_, r_40__12_, r_40__11_, r_40__10_, r_40__9_, r_40__8_, r_40__7_, r_40__6_, r_40__5_, r_40__4_, r_40__3_, r_40__2_, r_40__1_, r_40__0_ } : 
                                                                                                                                                                                                                    (N79)? data_i : 1'b0;
  assign N78 = sel_i[78];
  assign N79 = N327;
  assign { r_n_40__15_, r_n_40__14_, r_n_40__13_, r_n_40__12_, r_n_40__11_, r_n_40__10_, r_n_40__9_, r_n_40__8_, r_n_40__7_, r_n_40__6_, r_n_40__5_, r_n_40__4_, r_n_40__3_, r_n_40__2_, r_n_40__1_, r_n_40__0_ } = (N80)? { r_41__15_, r_41__14_, r_41__13_, r_41__12_, r_41__11_, r_41__10_, r_41__9_, r_41__8_, r_41__7_, r_41__6_, r_41__5_, r_41__4_, r_41__3_, r_41__2_, r_41__1_, r_41__0_ } : 
                                                                                                                                                                                                                    (N81)? data_i : 1'b0;
  assign N80 = sel_i[80];
  assign N81 = N332;
  assign { r_n_41__15_, r_n_41__14_, r_n_41__13_, r_n_41__12_, r_n_41__11_, r_n_41__10_, r_n_41__9_, r_n_41__8_, r_n_41__7_, r_n_41__6_, r_n_41__5_, r_n_41__4_, r_n_41__3_, r_n_41__2_, r_n_41__1_, r_n_41__0_ } = (N82)? { r_42__15_, r_42__14_, r_42__13_, r_42__12_, r_42__11_, r_42__10_, r_42__9_, r_42__8_, r_42__7_, r_42__6_, r_42__5_, r_42__4_, r_42__3_, r_42__2_, r_42__1_, r_42__0_ } : 
                                                                                                                                                                                                                    (N83)? data_i : 1'b0;
  assign N82 = sel_i[82];
  assign N83 = N337;
  assign { r_n_42__15_, r_n_42__14_, r_n_42__13_, r_n_42__12_, r_n_42__11_, r_n_42__10_, r_n_42__9_, r_n_42__8_, r_n_42__7_, r_n_42__6_, r_n_42__5_, r_n_42__4_, r_n_42__3_, r_n_42__2_, r_n_42__1_, r_n_42__0_ } = (N84)? { r_43__15_, r_43__14_, r_43__13_, r_43__12_, r_43__11_, r_43__10_, r_43__9_, r_43__8_, r_43__7_, r_43__6_, r_43__5_, r_43__4_, r_43__3_, r_43__2_, r_43__1_, r_43__0_ } : 
                                                                                                                                                                                                                    (N85)? data_i : 1'b0;
  assign N84 = sel_i[84];
  assign N85 = N342;
  assign { r_n_43__15_, r_n_43__14_, r_n_43__13_, r_n_43__12_, r_n_43__11_, r_n_43__10_, r_n_43__9_, r_n_43__8_, r_n_43__7_, r_n_43__6_, r_n_43__5_, r_n_43__4_, r_n_43__3_, r_n_43__2_, r_n_43__1_, r_n_43__0_ } = (N86)? { r_44__15_, r_44__14_, r_44__13_, r_44__12_, r_44__11_, r_44__10_, r_44__9_, r_44__8_, r_44__7_, r_44__6_, r_44__5_, r_44__4_, r_44__3_, r_44__2_, r_44__1_, r_44__0_ } : 
                                                                                                                                                                                                                    (N87)? data_i : 1'b0;
  assign N86 = sel_i[86];
  assign N87 = N347;
  assign { r_n_44__15_, r_n_44__14_, r_n_44__13_, r_n_44__12_, r_n_44__11_, r_n_44__10_, r_n_44__9_, r_n_44__8_, r_n_44__7_, r_n_44__6_, r_n_44__5_, r_n_44__4_, r_n_44__3_, r_n_44__2_, r_n_44__1_, r_n_44__0_ } = (N88)? { r_45__15_, r_45__14_, r_45__13_, r_45__12_, r_45__11_, r_45__10_, r_45__9_, r_45__8_, r_45__7_, r_45__6_, r_45__5_, r_45__4_, r_45__3_, r_45__2_, r_45__1_, r_45__0_ } : 
                                                                                                                                                                                                                    (N89)? data_i : 1'b0;
  assign N88 = sel_i[88];
  assign N89 = N352;
  assign { r_n_45__15_, r_n_45__14_, r_n_45__13_, r_n_45__12_, r_n_45__11_, r_n_45__10_, r_n_45__9_, r_n_45__8_, r_n_45__7_, r_n_45__6_, r_n_45__5_, r_n_45__4_, r_n_45__3_, r_n_45__2_, r_n_45__1_, r_n_45__0_ } = (N90)? { r_46__15_, r_46__14_, r_46__13_, r_46__12_, r_46__11_, r_46__10_, r_46__9_, r_46__8_, r_46__7_, r_46__6_, r_46__5_, r_46__4_, r_46__3_, r_46__2_, r_46__1_, r_46__0_ } : 
                                                                                                                                                                                                                    (N91)? data_i : 1'b0;
  assign N90 = sel_i[90];
  assign N91 = N357;
  assign { r_n_46__15_, r_n_46__14_, r_n_46__13_, r_n_46__12_, r_n_46__11_, r_n_46__10_, r_n_46__9_, r_n_46__8_, r_n_46__7_, r_n_46__6_, r_n_46__5_, r_n_46__4_, r_n_46__3_, r_n_46__2_, r_n_46__1_, r_n_46__0_ } = (N92)? { r_47__15_, r_47__14_, r_47__13_, r_47__12_, r_47__11_, r_47__10_, r_47__9_, r_47__8_, r_47__7_, r_47__6_, r_47__5_, r_47__4_, r_47__3_, r_47__2_, r_47__1_, r_47__0_ } : 
                                                                                                                                                                                                                    (N93)? data_i : 1'b0;
  assign N92 = sel_i[92];
  assign N93 = N362;
  assign { r_n_47__15_, r_n_47__14_, r_n_47__13_, r_n_47__12_, r_n_47__11_, r_n_47__10_, r_n_47__9_, r_n_47__8_, r_n_47__7_, r_n_47__6_, r_n_47__5_, r_n_47__4_, r_n_47__3_, r_n_47__2_, r_n_47__1_, r_n_47__0_ } = (N94)? { r_48__15_, r_48__14_, r_48__13_, r_48__12_, r_48__11_, r_48__10_, r_48__9_, r_48__8_, r_48__7_, r_48__6_, r_48__5_, r_48__4_, r_48__3_, r_48__2_, r_48__1_, r_48__0_ } : 
                                                                                                                                                                                                                    (N95)? data_i : 1'b0;
  assign N94 = sel_i[94];
  assign N95 = N367;
  assign { r_n_48__15_, r_n_48__14_, r_n_48__13_, r_n_48__12_, r_n_48__11_, r_n_48__10_, r_n_48__9_, r_n_48__8_, r_n_48__7_, r_n_48__6_, r_n_48__5_, r_n_48__4_, r_n_48__3_, r_n_48__2_, r_n_48__1_, r_n_48__0_ } = (N96)? { r_49__15_, r_49__14_, r_49__13_, r_49__12_, r_49__11_, r_49__10_, r_49__9_, r_49__8_, r_49__7_, r_49__6_, r_49__5_, r_49__4_, r_49__3_, r_49__2_, r_49__1_, r_49__0_ } : 
                                                                                                                                                                                                                    (N97)? data_i : 1'b0;
  assign N96 = sel_i[96];
  assign N97 = N372;
  assign { r_n_49__15_, r_n_49__14_, r_n_49__13_, r_n_49__12_, r_n_49__11_, r_n_49__10_, r_n_49__9_, r_n_49__8_, r_n_49__7_, r_n_49__6_, r_n_49__5_, r_n_49__4_, r_n_49__3_, r_n_49__2_, r_n_49__1_, r_n_49__0_ } = (N98)? { r_50__15_, r_50__14_, r_50__13_, r_50__12_, r_50__11_, r_50__10_, r_50__9_, r_50__8_, r_50__7_, r_50__6_, r_50__5_, r_50__4_, r_50__3_, r_50__2_, r_50__1_, r_50__0_ } : 
                                                                                                                                                                                                                    (N99)? data_i : 1'b0;
  assign N98 = sel_i[98];
  assign N99 = N377;
  assign { r_n_50__15_, r_n_50__14_, r_n_50__13_, r_n_50__12_, r_n_50__11_, r_n_50__10_, r_n_50__9_, r_n_50__8_, r_n_50__7_, r_n_50__6_, r_n_50__5_, r_n_50__4_, r_n_50__3_, r_n_50__2_, r_n_50__1_, r_n_50__0_ } = (N100)? { r_51__15_, r_51__14_, r_51__13_, r_51__12_, r_51__11_, r_51__10_, r_51__9_, r_51__8_, r_51__7_, r_51__6_, r_51__5_, r_51__4_, r_51__3_, r_51__2_, r_51__1_, r_51__0_ } : 
                                                                                                                                                                                                                    (N101)? data_i : 1'b0;
  assign N100 = sel_i[100];
  assign N101 = N382;
  assign { r_n_51__15_, r_n_51__14_, r_n_51__13_, r_n_51__12_, r_n_51__11_, r_n_51__10_, r_n_51__9_, r_n_51__8_, r_n_51__7_, r_n_51__6_, r_n_51__5_, r_n_51__4_, r_n_51__3_, r_n_51__2_, r_n_51__1_, r_n_51__0_ } = (N102)? { r_52__15_, r_52__14_, r_52__13_, r_52__12_, r_52__11_, r_52__10_, r_52__9_, r_52__8_, r_52__7_, r_52__6_, r_52__5_, r_52__4_, r_52__3_, r_52__2_, r_52__1_, r_52__0_ } : 
                                                                                                                                                                                                                    (N103)? data_i : 1'b0;
  assign N102 = sel_i[102];
  assign N103 = N387;
  assign { r_n_52__15_, r_n_52__14_, r_n_52__13_, r_n_52__12_, r_n_52__11_, r_n_52__10_, r_n_52__9_, r_n_52__8_, r_n_52__7_, r_n_52__6_, r_n_52__5_, r_n_52__4_, r_n_52__3_, r_n_52__2_, r_n_52__1_, r_n_52__0_ } = (N104)? { r_53__15_, r_53__14_, r_53__13_, r_53__12_, r_53__11_, r_53__10_, r_53__9_, r_53__8_, r_53__7_, r_53__6_, r_53__5_, r_53__4_, r_53__3_, r_53__2_, r_53__1_, r_53__0_ } : 
                                                                                                                                                                                                                    (N105)? data_i : 1'b0;
  assign N104 = sel_i[104];
  assign N105 = N392;
  assign { r_n_53__15_, r_n_53__14_, r_n_53__13_, r_n_53__12_, r_n_53__11_, r_n_53__10_, r_n_53__9_, r_n_53__8_, r_n_53__7_, r_n_53__6_, r_n_53__5_, r_n_53__4_, r_n_53__3_, r_n_53__2_, r_n_53__1_, r_n_53__0_ } = (N106)? { r_54__15_, r_54__14_, r_54__13_, r_54__12_, r_54__11_, r_54__10_, r_54__9_, r_54__8_, r_54__7_, r_54__6_, r_54__5_, r_54__4_, r_54__3_, r_54__2_, r_54__1_, r_54__0_ } : 
                                                                                                                                                                                                                    (N107)? data_i : 1'b0;
  assign N106 = sel_i[106];
  assign N107 = N397;
  assign { r_n_54__15_, r_n_54__14_, r_n_54__13_, r_n_54__12_, r_n_54__11_, r_n_54__10_, r_n_54__9_, r_n_54__8_, r_n_54__7_, r_n_54__6_, r_n_54__5_, r_n_54__4_, r_n_54__3_, r_n_54__2_, r_n_54__1_, r_n_54__0_ } = (N108)? { r_55__15_, r_55__14_, r_55__13_, r_55__12_, r_55__11_, r_55__10_, r_55__9_, r_55__8_, r_55__7_, r_55__6_, r_55__5_, r_55__4_, r_55__3_, r_55__2_, r_55__1_, r_55__0_ } : 
                                                                                                                                                                                                                    (N109)? data_i : 1'b0;
  assign N108 = sel_i[108];
  assign N109 = N402;
  assign { r_n_55__15_, r_n_55__14_, r_n_55__13_, r_n_55__12_, r_n_55__11_, r_n_55__10_, r_n_55__9_, r_n_55__8_, r_n_55__7_, r_n_55__6_, r_n_55__5_, r_n_55__4_, r_n_55__3_, r_n_55__2_, r_n_55__1_, r_n_55__0_ } = (N110)? { r_56__15_, r_56__14_, r_56__13_, r_56__12_, r_56__11_, r_56__10_, r_56__9_, r_56__8_, r_56__7_, r_56__6_, r_56__5_, r_56__4_, r_56__3_, r_56__2_, r_56__1_, r_56__0_ } : 
                                                                                                                                                                                                                    (N111)? data_i : 1'b0;
  assign N110 = sel_i[110];
  assign N111 = N407;
  assign { r_n_56__15_, r_n_56__14_, r_n_56__13_, r_n_56__12_, r_n_56__11_, r_n_56__10_, r_n_56__9_, r_n_56__8_, r_n_56__7_, r_n_56__6_, r_n_56__5_, r_n_56__4_, r_n_56__3_, r_n_56__2_, r_n_56__1_, r_n_56__0_ } = (N112)? { r_57__15_, r_57__14_, r_57__13_, r_57__12_, r_57__11_, r_57__10_, r_57__9_, r_57__8_, r_57__7_, r_57__6_, r_57__5_, r_57__4_, r_57__3_, r_57__2_, r_57__1_, r_57__0_ } : 
                                                                                                                                                                                                                    (N113)? data_i : 1'b0;
  assign N112 = sel_i[112];
  assign N113 = N412;
  assign { r_n_57__15_, r_n_57__14_, r_n_57__13_, r_n_57__12_, r_n_57__11_, r_n_57__10_, r_n_57__9_, r_n_57__8_, r_n_57__7_, r_n_57__6_, r_n_57__5_, r_n_57__4_, r_n_57__3_, r_n_57__2_, r_n_57__1_, r_n_57__0_ } = (N114)? { r_58__15_, r_58__14_, r_58__13_, r_58__12_, r_58__11_, r_58__10_, r_58__9_, r_58__8_, r_58__7_, r_58__6_, r_58__5_, r_58__4_, r_58__3_, r_58__2_, r_58__1_, r_58__0_ } : 
                                                                                                                                                                                                                    (N115)? data_i : 1'b0;
  assign N114 = sel_i[114];
  assign N115 = N417;
  assign { r_n_58__15_, r_n_58__14_, r_n_58__13_, r_n_58__12_, r_n_58__11_, r_n_58__10_, r_n_58__9_, r_n_58__8_, r_n_58__7_, r_n_58__6_, r_n_58__5_, r_n_58__4_, r_n_58__3_, r_n_58__2_, r_n_58__1_, r_n_58__0_ } = (N116)? { r_59__15_, r_59__14_, r_59__13_, r_59__12_, r_59__11_, r_59__10_, r_59__9_, r_59__8_, r_59__7_, r_59__6_, r_59__5_, r_59__4_, r_59__3_, r_59__2_, r_59__1_, r_59__0_ } : 
                                                                                                                                                                                                                    (N117)? data_i : 1'b0;
  assign N116 = sel_i[116];
  assign N117 = N422;
  assign { r_n_59__15_, r_n_59__14_, r_n_59__13_, r_n_59__12_, r_n_59__11_, r_n_59__10_, r_n_59__9_, r_n_59__8_, r_n_59__7_, r_n_59__6_, r_n_59__5_, r_n_59__4_, r_n_59__3_, r_n_59__2_, r_n_59__1_, r_n_59__0_ } = (N118)? { r_60__15_, r_60__14_, r_60__13_, r_60__12_, r_60__11_, r_60__10_, r_60__9_, r_60__8_, r_60__7_, r_60__6_, r_60__5_, r_60__4_, r_60__3_, r_60__2_, r_60__1_, r_60__0_ } : 
                                                                                                                                                                                                                    (N119)? data_i : 1'b0;
  assign N118 = sel_i[118];
  assign N119 = N427;
  assign { r_n_60__15_, r_n_60__14_, r_n_60__13_, r_n_60__12_, r_n_60__11_, r_n_60__10_, r_n_60__9_, r_n_60__8_, r_n_60__7_, r_n_60__6_, r_n_60__5_, r_n_60__4_, r_n_60__3_, r_n_60__2_, r_n_60__1_, r_n_60__0_ } = (N120)? { r_61__15_, r_61__14_, r_61__13_, r_61__12_, r_61__11_, r_61__10_, r_61__9_, r_61__8_, r_61__7_, r_61__6_, r_61__5_, r_61__4_, r_61__3_, r_61__2_, r_61__1_, r_61__0_ } : 
                                                                                                                                                                                                                    (N121)? data_i : 1'b0;
  assign N120 = sel_i[120];
  assign N121 = N432;
  assign { r_n_61__15_, r_n_61__14_, r_n_61__13_, r_n_61__12_, r_n_61__11_, r_n_61__10_, r_n_61__9_, r_n_61__8_, r_n_61__7_, r_n_61__6_, r_n_61__5_, r_n_61__4_, r_n_61__3_, r_n_61__2_, r_n_61__1_, r_n_61__0_ } = (N122)? { r_62__15_, r_62__14_, r_62__13_, r_62__12_, r_62__11_, r_62__10_, r_62__9_, r_62__8_, r_62__7_, r_62__6_, r_62__5_, r_62__4_, r_62__3_, r_62__2_, r_62__1_, r_62__0_ } : 
                                                                                                                                                                                                                    (N123)? data_i : 1'b0;
  assign N122 = sel_i[122];
  assign N123 = N437;
  assign { r_n_62__15_, r_n_62__14_, r_n_62__13_, r_n_62__12_, r_n_62__11_, r_n_62__10_, r_n_62__9_, r_n_62__8_, r_n_62__7_, r_n_62__6_, r_n_62__5_, r_n_62__4_, r_n_62__3_, r_n_62__2_, r_n_62__1_, r_n_62__0_ } = (N124)? { r_63__15_, r_63__14_, r_63__13_, r_63__12_, r_63__11_, r_63__10_, r_63__9_, r_63__8_, r_63__7_, r_63__6_, r_63__5_, r_63__4_, r_63__3_, r_63__2_, r_63__1_, r_63__0_ } : 
                                                                                                                                                                                                                    (N125)? data_i : 1'b0;
  assign N124 = sel_i[124];
  assign N125 = N442;
  assign { r_n_63__15_, r_n_63__14_, r_n_63__13_, r_n_63__12_, r_n_63__11_, r_n_63__10_, r_n_63__9_, r_n_63__8_, r_n_63__7_, r_n_63__6_, r_n_63__5_, r_n_63__4_, r_n_63__3_, r_n_63__2_, r_n_63__1_, r_n_63__0_ } = (N126)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                    (N127)? data_i : 1'b0;
  assign N126 = sel_i[126];
  assign N127 = N447;
  assign N129 = ~sel_i[1];
  assign N131 = N128 | N130;
  assign N134 = ~sel_i[3];
  assign N136 = N133 | N135;
  assign N139 = ~sel_i[5];
  assign N141 = N138 | N140;
  assign N144 = ~sel_i[7];
  assign N146 = N143 | N145;
  assign N149 = ~sel_i[9];
  assign N151 = N148 | N150;
  assign N154 = ~sel_i[11];
  assign N156 = N153 | N155;
  assign N159 = ~sel_i[13];
  assign N161 = N158 | N160;
  assign N164 = ~sel_i[15];
  assign N166 = N163 | N165;
  assign N169 = ~sel_i[17];
  assign N171 = N168 | N170;
  assign N174 = ~sel_i[19];
  assign N176 = N173 | N175;
  assign N179 = ~sel_i[21];
  assign N181 = N178 | N180;
  assign N184 = ~sel_i[23];
  assign N186 = N183 | N185;
  assign N189 = ~sel_i[25];
  assign N191 = N188 | N190;
  assign N194 = ~sel_i[27];
  assign N196 = N193 | N195;
  assign N199 = ~sel_i[29];
  assign N201 = N198 | N200;
  assign N204 = ~sel_i[31];
  assign N206 = N203 | N205;
  assign N209 = ~sel_i[33];
  assign N211 = N208 | N210;
  assign N214 = ~sel_i[35];
  assign N216 = N213 | N215;
  assign N219 = ~sel_i[37];
  assign N221 = N218 | N220;
  assign N224 = ~sel_i[39];
  assign N226 = N223 | N225;
  assign N229 = ~sel_i[41];
  assign N231 = N228 | N230;
  assign N234 = ~sel_i[43];
  assign N236 = N233 | N235;
  assign N239 = ~sel_i[45];
  assign N241 = N238 | N240;
  assign N244 = ~sel_i[47];
  assign N246 = N243 | N245;
  assign N249 = ~sel_i[49];
  assign N251 = N248 | N250;
  assign N254 = ~sel_i[51];
  assign N256 = N253 | N255;
  assign N259 = ~sel_i[53];
  assign N261 = N258 | N260;
  assign N264 = ~sel_i[55];
  assign N266 = N263 | N265;
  assign N269 = ~sel_i[57];
  assign N271 = N268 | N270;
  assign N274 = ~sel_i[59];
  assign N276 = N273 | N275;
  assign N279 = ~sel_i[61];
  assign N281 = N278 | N280;
  assign N284 = ~sel_i[63];
  assign N286 = N283 | N285;
  assign N289 = ~sel_i[65];
  assign N291 = N288 | N290;
  assign N294 = ~sel_i[67];
  assign N296 = N293 | N295;
  assign N299 = ~sel_i[69];
  assign N301 = N298 | N300;
  assign N304 = ~sel_i[71];
  assign N306 = N303 | N305;
  assign N309 = ~sel_i[73];
  assign N311 = N308 | N310;
  assign N314 = ~sel_i[75];
  assign N316 = N313 | N315;
  assign N319 = ~sel_i[77];
  assign N321 = N318 | N320;
  assign N324 = ~sel_i[79];
  assign N326 = N323 | N325;
  assign N329 = ~sel_i[81];
  assign N331 = N328 | N330;
  assign N334 = ~sel_i[83];
  assign N336 = N333 | N335;
  assign N339 = ~sel_i[85];
  assign N341 = N338 | N340;
  assign N344 = ~sel_i[87];
  assign N346 = N343 | N345;
  assign N349 = ~sel_i[89];
  assign N351 = N348 | N350;
  assign N354 = ~sel_i[91];
  assign N356 = N353 | N355;
  assign N359 = ~sel_i[93];
  assign N361 = N358 | N360;
  assign N364 = ~sel_i[95];
  assign N366 = N363 | N365;
  assign N369 = ~sel_i[97];
  assign N371 = N368 | N370;
  assign N374 = ~sel_i[99];
  assign N376 = N373 | N375;
  assign N379 = ~sel_i[101];
  assign N381 = N378 | N380;
  assign N384 = ~sel_i[103];
  assign N386 = N383 | N385;
  assign N389 = ~sel_i[105];
  assign N391 = N388 | N390;
  assign N394 = ~sel_i[107];
  assign N396 = N393 | N395;
  assign N399 = ~sel_i[109];
  assign N401 = N398 | N400;
  assign N404 = ~sel_i[111];
  assign N406 = N403 | N405;
  assign N409 = ~sel_i[113];
  assign N411 = N408 | N410;
  assign N414 = ~sel_i[115];
  assign N416 = N413 | N415;
  assign N419 = ~sel_i[117];
  assign N421 = N418 | N420;
  assign N424 = ~sel_i[119];
  assign N426 = N423 | N425;
  assign N429 = ~sel_i[121];
  assign N431 = N428 | N430;
  assign N434 = ~sel_i[123];
  assign N436 = N433 | N435;
  assign N439 = ~sel_i[125];
  assign N441 = N438 | N440;
  assign N444 = ~sel_i[127];
  assign N446 = N443 | N445;
  assign N448 = ~N131;
  assign N449 = ~N136;
  assign N450 = ~N141;
  assign N451 = ~N146;
  assign N452 = ~N151;
  assign N453 = ~N156;
  assign N454 = ~N161;
  assign N455 = ~N166;
  assign N456 = ~N171;
  assign N457 = ~N176;
  assign N458 = ~N181;
  assign N459 = ~N186;
  assign N460 = ~N191;
  assign N461 = ~N196;
  assign N462 = ~N201;
  assign N463 = ~N206;
  assign N464 = ~N211;
  assign N465 = ~N216;
  assign N466 = ~N221;
  assign N467 = ~N226;
  assign N468 = ~N231;
  assign N469 = ~N236;
  assign N470 = ~N241;
  assign N471 = ~N246;
  assign N472 = ~N251;
  assign N473 = ~N256;
  assign N474 = ~N261;
  assign N475 = ~N266;
  assign N476 = ~N271;
  assign N477 = ~N276;
  assign N478 = ~N281;
  assign N479 = ~N286;
  assign N480 = ~N291;
  assign N481 = ~N296;
  assign N482 = ~N301;
  assign N483 = ~N306;
  assign N484 = ~N311;
  assign N485 = ~N316;
  assign N486 = ~N321;
  assign N487 = ~N326;
  assign N488 = ~N331;
  assign N489 = ~N336;
  assign N490 = ~N341;
  assign N491 = ~N346;
  assign N492 = ~N351;
  assign N493 = ~N356;
  assign N494 = ~N361;
  assign N495 = ~N366;
  assign N496 = ~N371;
  assign N497 = ~N376;
  assign N498 = ~N381;
  assign N499 = ~N386;
  assign N500 = ~N391;
  assign N501 = ~N396;
  assign N502 = ~N401;
  assign N503 = ~N406;
  assign N504 = ~N411;
  assign N505 = ~N416;
  assign N506 = ~N421;
  assign N507 = ~N426;
  assign N508 = ~N431;
  assign N509 = ~N436;
  assign N510 = ~N441;
  assign N511 = ~N446;

  always @(posedge clk_i) begin
    if(N448) begin
      { data_o[15:0] } <= { r_n_0__15_, r_n_0__14_, r_n_0__13_, r_n_0__12_, r_n_0__11_, r_n_0__10_, r_n_0__9_, r_n_0__8_, r_n_0__7_, r_n_0__6_, r_n_0__5_, r_n_0__4_, r_n_0__3_, r_n_0__2_, r_n_0__1_, r_n_0__0_ };
    end 
    if(N449) begin
      r_1__15_ <= r_n_1__15_;
      r_1__14_ <= r_n_1__14_;
      r_1__13_ <= r_n_1__13_;
      r_1__12_ <= r_n_1__12_;
      r_1__11_ <= r_n_1__11_;
      r_1__10_ <= r_n_1__10_;
      r_1__9_ <= r_n_1__9_;
      r_1__8_ <= r_n_1__8_;
      r_1__7_ <= r_n_1__7_;
      r_1__6_ <= r_n_1__6_;
      r_1__5_ <= r_n_1__5_;
      r_1__4_ <= r_n_1__4_;
      r_1__3_ <= r_n_1__3_;
      r_1__2_ <= r_n_1__2_;
      r_1__1_ <= r_n_1__1_;
      r_1__0_ <= r_n_1__0_;
    end 
    if(N450) begin
      r_2__15_ <= r_n_2__15_;
      r_2__14_ <= r_n_2__14_;
      r_2__13_ <= r_n_2__13_;
      r_2__12_ <= r_n_2__12_;
      r_2__11_ <= r_n_2__11_;
      r_2__10_ <= r_n_2__10_;
      r_2__9_ <= r_n_2__9_;
      r_2__8_ <= r_n_2__8_;
      r_2__7_ <= r_n_2__7_;
      r_2__6_ <= r_n_2__6_;
      r_2__5_ <= r_n_2__5_;
      r_2__4_ <= r_n_2__4_;
      r_2__3_ <= r_n_2__3_;
      r_2__2_ <= r_n_2__2_;
      r_2__1_ <= r_n_2__1_;
      r_2__0_ <= r_n_2__0_;
    end 
    if(N451) begin
      r_3__15_ <= r_n_3__15_;
      r_3__14_ <= r_n_3__14_;
      r_3__13_ <= r_n_3__13_;
      r_3__12_ <= r_n_3__12_;
      r_3__11_ <= r_n_3__11_;
      r_3__10_ <= r_n_3__10_;
      r_3__9_ <= r_n_3__9_;
      r_3__8_ <= r_n_3__8_;
      r_3__7_ <= r_n_3__7_;
      r_3__6_ <= r_n_3__6_;
      r_3__5_ <= r_n_3__5_;
      r_3__4_ <= r_n_3__4_;
      r_3__3_ <= r_n_3__3_;
      r_3__2_ <= r_n_3__2_;
      r_3__1_ <= r_n_3__1_;
      r_3__0_ <= r_n_3__0_;
    end 
    if(N452) begin
      r_4__15_ <= r_n_4__15_;
      r_4__14_ <= r_n_4__14_;
      r_4__13_ <= r_n_4__13_;
      r_4__12_ <= r_n_4__12_;
      r_4__11_ <= r_n_4__11_;
      r_4__10_ <= r_n_4__10_;
      r_4__9_ <= r_n_4__9_;
      r_4__8_ <= r_n_4__8_;
      r_4__7_ <= r_n_4__7_;
      r_4__6_ <= r_n_4__6_;
      r_4__5_ <= r_n_4__5_;
      r_4__4_ <= r_n_4__4_;
      r_4__3_ <= r_n_4__3_;
      r_4__2_ <= r_n_4__2_;
      r_4__1_ <= r_n_4__1_;
      r_4__0_ <= r_n_4__0_;
    end 
    if(N453) begin
      r_5__15_ <= r_n_5__15_;
      r_5__14_ <= r_n_5__14_;
      r_5__13_ <= r_n_5__13_;
      r_5__12_ <= r_n_5__12_;
      r_5__11_ <= r_n_5__11_;
      r_5__10_ <= r_n_5__10_;
      r_5__9_ <= r_n_5__9_;
      r_5__8_ <= r_n_5__8_;
      r_5__7_ <= r_n_5__7_;
      r_5__6_ <= r_n_5__6_;
      r_5__5_ <= r_n_5__5_;
      r_5__4_ <= r_n_5__4_;
      r_5__3_ <= r_n_5__3_;
      r_5__2_ <= r_n_5__2_;
      r_5__1_ <= r_n_5__1_;
      r_5__0_ <= r_n_5__0_;
    end 
    if(N454) begin
      r_6__15_ <= r_n_6__15_;
      r_6__14_ <= r_n_6__14_;
      r_6__13_ <= r_n_6__13_;
      r_6__12_ <= r_n_6__12_;
      r_6__11_ <= r_n_6__11_;
      r_6__10_ <= r_n_6__10_;
      r_6__9_ <= r_n_6__9_;
      r_6__8_ <= r_n_6__8_;
      r_6__7_ <= r_n_6__7_;
      r_6__6_ <= r_n_6__6_;
      r_6__5_ <= r_n_6__5_;
      r_6__4_ <= r_n_6__4_;
      r_6__3_ <= r_n_6__3_;
      r_6__2_ <= r_n_6__2_;
      r_6__1_ <= r_n_6__1_;
      r_6__0_ <= r_n_6__0_;
    end 
    if(N455) begin
      r_7__15_ <= r_n_7__15_;
      r_7__14_ <= r_n_7__14_;
      r_7__13_ <= r_n_7__13_;
      r_7__12_ <= r_n_7__12_;
      r_7__11_ <= r_n_7__11_;
      r_7__10_ <= r_n_7__10_;
      r_7__9_ <= r_n_7__9_;
      r_7__8_ <= r_n_7__8_;
      r_7__7_ <= r_n_7__7_;
      r_7__6_ <= r_n_7__6_;
      r_7__5_ <= r_n_7__5_;
      r_7__4_ <= r_n_7__4_;
      r_7__3_ <= r_n_7__3_;
      r_7__2_ <= r_n_7__2_;
      r_7__1_ <= r_n_7__1_;
      r_7__0_ <= r_n_7__0_;
    end 
    if(N456) begin
      r_8__15_ <= r_n_8__15_;
      r_8__14_ <= r_n_8__14_;
      r_8__13_ <= r_n_8__13_;
      r_8__12_ <= r_n_8__12_;
      r_8__11_ <= r_n_8__11_;
      r_8__10_ <= r_n_8__10_;
      r_8__9_ <= r_n_8__9_;
      r_8__8_ <= r_n_8__8_;
      r_8__7_ <= r_n_8__7_;
      r_8__6_ <= r_n_8__6_;
      r_8__5_ <= r_n_8__5_;
      r_8__4_ <= r_n_8__4_;
      r_8__3_ <= r_n_8__3_;
      r_8__2_ <= r_n_8__2_;
      r_8__1_ <= r_n_8__1_;
      r_8__0_ <= r_n_8__0_;
    end 
    if(N457) begin
      r_9__15_ <= r_n_9__15_;
      r_9__14_ <= r_n_9__14_;
      r_9__13_ <= r_n_9__13_;
      r_9__12_ <= r_n_9__12_;
      r_9__11_ <= r_n_9__11_;
      r_9__10_ <= r_n_9__10_;
      r_9__9_ <= r_n_9__9_;
      r_9__8_ <= r_n_9__8_;
      r_9__7_ <= r_n_9__7_;
      r_9__6_ <= r_n_9__6_;
      r_9__5_ <= r_n_9__5_;
      r_9__4_ <= r_n_9__4_;
      r_9__3_ <= r_n_9__3_;
      r_9__2_ <= r_n_9__2_;
      r_9__1_ <= r_n_9__1_;
      r_9__0_ <= r_n_9__0_;
    end 
    if(N458) begin
      r_10__15_ <= r_n_10__15_;
      r_10__14_ <= r_n_10__14_;
      r_10__13_ <= r_n_10__13_;
      r_10__12_ <= r_n_10__12_;
      r_10__11_ <= r_n_10__11_;
      r_10__10_ <= r_n_10__10_;
      r_10__9_ <= r_n_10__9_;
      r_10__8_ <= r_n_10__8_;
      r_10__7_ <= r_n_10__7_;
      r_10__6_ <= r_n_10__6_;
      r_10__5_ <= r_n_10__5_;
      r_10__4_ <= r_n_10__4_;
      r_10__3_ <= r_n_10__3_;
      r_10__2_ <= r_n_10__2_;
      r_10__1_ <= r_n_10__1_;
      r_10__0_ <= r_n_10__0_;
    end 
    if(N459) begin
      r_11__15_ <= r_n_11__15_;
      r_11__14_ <= r_n_11__14_;
      r_11__13_ <= r_n_11__13_;
      r_11__12_ <= r_n_11__12_;
      r_11__11_ <= r_n_11__11_;
      r_11__10_ <= r_n_11__10_;
      r_11__9_ <= r_n_11__9_;
      r_11__8_ <= r_n_11__8_;
      r_11__7_ <= r_n_11__7_;
      r_11__6_ <= r_n_11__6_;
      r_11__5_ <= r_n_11__5_;
      r_11__4_ <= r_n_11__4_;
      r_11__3_ <= r_n_11__3_;
      r_11__2_ <= r_n_11__2_;
      r_11__1_ <= r_n_11__1_;
      r_11__0_ <= r_n_11__0_;
    end 
    if(N460) begin
      r_12__15_ <= r_n_12__15_;
      r_12__14_ <= r_n_12__14_;
      r_12__13_ <= r_n_12__13_;
      r_12__12_ <= r_n_12__12_;
      r_12__11_ <= r_n_12__11_;
      r_12__10_ <= r_n_12__10_;
      r_12__9_ <= r_n_12__9_;
      r_12__8_ <= r_n_12__8_;
      r_12__7_ <= r_n_12__7_;
      r_12__6_ <= r_n_12__6_;
      r_12__5_ <= r_n_12__5_;
      r_12__4_ <= r_n_12__4_;
      r_12__3_ <= r_n_12__3_;
      r_12__2_ <= r_n_12__2_;
      r_12__1_ <= r_n_12__1_;
      r_12__0_ <= r_n_12__0_;
    end 
    if(N461) begin
      r_13__15_ <= r_n_13__15_;
      r_13__14_ <= r_n_13__14_;
      r_13__13_ <= r_n_13__13_;
      r_13__12_ <= r_n_13__12_;
      r_13__11_ <= r_n_13__11_;
      r_13__10_ <= r_n_13__10_;
      r_13__9_ <= r_n_13__9_;
      r_13__8_ <= r_n_13__8_;
      r_13__7_ <= r_n_13__7_;
      r_13__6_ <= r_n_13__6_;
      r_13__5_ <= r_n_13__5_;
      r_13__4_ <= r_n_13__4_;
      r_13__3_ <= r_n_13__3_;
      r_13__2_ <= r_n_13__2_;
      r_13__1_ <= r_n_13__1_;
      r_13__0_ <= r_n_13__0_;
    end 
    if(N462) begin
      r_14__15_ <= r_n_14__15_;
      r_14__14_ <= r_n_14__14_;
      r_14__13_ <= r_n_14__13_;
      r_14__12_ <= r_n_14__12_;
      r_14__11_ <= r_n_14__11_;
      r_14__10_ <= r_n_14__10_;
      r_14__9_ <= r_n_14__9_;
      r_14__8_ <= r_n_14__8_;
      r_14__7_ <= r_n_14__7_;
      r_14__6_ <= r_n_14__6_;
      r_14__5_ <= r_n_14__5_;
      r_14__4_ <= r_n_14__4_;
      r_14__3_ <= r_n_14__3_;
      r_14__2_ <= r_n_14__2_;
      r_14__1_ <= r_n_14__1_;
      r_14__0_ <= r_n_14__0_;
    end 
    if(N463) begin
      r_15__15_ <= r_n_15__15_;
      r_15__14_ <= r_n_15__14_;
      r_15__13_ <= r_n_15__13_;
      r_15__12_ <= r_n_15__12_;
      r_15__11_ <= r_n_15__11_;
      r_15__10_ <= r_n_15__10_;
      r_15__9_ <= r_n_15__9_;
      r_15__8_ <= r_n_15__8_;
      r_15__7_ <= r_n_15__7_;
      r_15__6_ <= r_n_15__6_;
      r_15__5_ <= r_n_15__5_;
      r_15__4_ <= r_n_15__4_;
      r_15__3_ <= r_n_15__3_;
      r_15__2_ <= r_n_15__2_;
      r_15__1_ <= r_n_15__1_;
      r_15__0_ <= r_n_15__0_;
    end 
    if(N464) begin
      r_16__15_ <= r_n_16__15_;
      r_16__14_ <= r_n_16__14_;
      r_16__13_ <= r_n_16__13_;
      r_16__12_ <= r_n_16__12_;
      r_16__11_ <= r_n_16__11_;
      r_16__10_ <= r_n_16__10_;
      r_16__9_ <= r_n_16__9_;
      r_16__8_ <= r_n_16__8_;
      r_16__7_ <= r_n_16__7_;
      r_16__6_ <= r_n_16__6_;
      r_16__5_ <= r_n_16__5_;
      r_16__4_ <= r_n_16__4_;
      r_16__3_ <= r_n_16__3_;
      r_16__2_ <= r_n_16__2_;
      r_16__1_ <= r_n_16__1_;
      r_16__0_ <= r_n_16__0_;
    end 
    if(N465) begin
      r_17__15_ <= r_n_17__15_;
      r_17__14_ <= r_n_17__14_;
      r_17__13_ <= r_n_17__13_;
      r_17__12_ <= r_n_17__12_;
      r_17__11_ <= r_n_17__11_;
      r_17__10_ <= r_n_17__10_;
      r_17__9_ <= r_n_17__9_;
      r_17__8_ <= r_n_17__8_;
      r_17__7_ <= r_n_17__7_;
      r_17__6_ <= r_n_17__6_;
      r_17__5_ <= r_n_17__5_;
      r_17__4_ <= r_n_17__4_;
      r_17__3_ <= r_n_17__3_;
      r_17__2_ <= r_n_17__2_;
      r_17__1_ <= r_n_17__1_;
      r_17__0_ <= r_n_17__0_;
    end 
    if(N466) begin
      r_18__15_ <= r_n_18__15_;
      r_18__14_ <= r_n_18__14_;
      r_18__13_ <= r_n_18__13_;
      r_18__12_ <= r_n_18__12_;
      r_18__11_ <= r_n_18__11_;
      r_18__10_ <= r_n_18__10_;
      r_18__9_ <= r_n_18__9_;
      r_18__8_ <= r_n_18__8_;
      r_18__7_ <= r_n_18__7_;
      r_18__6_ <= r_n_18__6_;
      r_18__5_ <= r_n_18__5_;
      r_18__4_ <= r_n_18__4_;
      r_18__3_ <= r_n_18__3_;
      r_18__2_ <= r_n_18__2_;
      r_18__1_ <= r_n_18__1_;
      r_18__0_ <= r_n_18__0_;
    end 
    if(N467) begin
      r_19__15_ <= r_n_19__15_;
      r_19__14_ <= r_n_19__14_;
      r_19__13_ <= r_n_19__13_;
      r_19__12_ <= r_n_19__12_;
      r_19__11_ <= r_n_19__11_;
      r_19__10_ <= r_n_19__10_;
      r_19__9_ <= r_n_19__9_;
      r_19__8_ <= r_n_19__8_;
      r_19__7_ <= r_n_19__7_;
      r_19__6_ <= r_n_19__6_;
      r_19__5_ <= r_n_19__5_;
      r_19__4_ <= r_n_19__4_;
      r_19__3_ <= r_n_19__3_;
      r_19__2_ <= r_n_19__2_;
      r_19__1_ <= r_n_19__1_;
      r_19__0_ <= r_n_19__0_;
    end 
    if(N468) begin
      r_20__15_ <= r_n_20__15_;
      r_20__14_ <= r_n_20__14_;
      r_20__13_ <= r_n_20__13_;
      r_20__12_ <= r_n_20__12_;
      r_20__11_ <= r_n_20__11_;
      r_20__10_ <= r_n_20__10_;
      r_20__9_ <= r_n_20__9_;
      r_20__8_ <= r_n_20__8_;
      r_20__7_ <= r_n_20__7_;
      r_20__6_ <= r_n_20__6_;
      r_20__5_ <= r_n_20__5_;
      r_20__4_ <= r_n_20__4_;
      r_20__3_ <= r_n_20__3_;
      r_20__2_ <= r_n_20__2_;
      r_20__1_ <= r_n_20__1_;
      r_20__0_ <= r_n_20__0_;
    end 
    if(N469) begin
      r_21__15_ <= r_n_21__15_;
      r_21__14_ <= r_n_21__14_;
      r_21__13_ <= r_n_21__13_;
      r_21__12_ <= r_n_21__12_;
      r_21__11_ <= r_n_21__11_;
      r_21__10_ <= r_n_21__10_;
      r_21__9_ <= r_n_21__9_;
      r_21__8_ <= r_n_21__8_;
      r_21__7_ <= r_n_21__7_;
      r_21__6_ <= r_n_21__6_;
      r_21__5_ <= r_n_21__5_;
      r_21__4_ <= r_n_21__4_;
      r_21__3_ <= r_n_21__3_;
      r_21__2_ <= r_n_21__2_;
      r_21__1_ <= r_n_21__1_;
      r_21__0_ <= r_n_21__0_;
    end 
    if(N470) begin
      r_22__15_ <= r_n_22__15_;
      r_22__14_ <= r_n_22__14_;
      r_22__13_ <= r_n_22__13_;
      r_22__12_ <= r_n_22__12_;
      r_22__11_ <= r_n_22__11_;
      r_22__10_ <= r_n_22__10_;
      r_22__9_ <= r_n_22__9_;
      r_22__8_ <= r_n_22__8_;
      r_22__7_ <= r_n_22__7_;
      r_22__6_ <= r_n_22__6_;
      r_22__5_ <= r_n_22__5_;
      r_22__4_ <= r_n_22__4_;
      r_22__3_ <= r_n_22__3_;
      r_22__2_ <= r_n_22__2_;
      r_22__1_ <= r_n_22__1_;
      r_22__0_ <= r_n_22__0_;
    end 
    if(N471) begin
      r_23__15_ <= r_n_23__15_;
      r_23__14_ <= r_n_23__14_;
      r_23__13_ <= r_n_23__13_;
      r_23__12_ <= r_n_23__12_;
      r_23__11_ <= r_n_23__11_;
      r_23__10_ <= r_n_23__10_;
      r_23__9_ <= r_n_23__9_;
      r_23__8_ <= r_n_23__8_;
      r_23__7_ <= r_n_23__7_;
      r_23__6_ <= r_n_23__6_;
      r_23__5_ <= r_n_23__5_;
      r_23__4_ <= r_n_23__4_;
      r_23__3_ <= r_n_23__3_;
      r_23__2_ <= r_n_23__2_;
      r_23__1_ <= r_n_23__1_;
      r_23__0_ <= r_n_23__0_;
    end 
    if(N472) begin
      r_24__15_ <= r_n_24__15_;
      r_24__14_ <= r_n_24__14_;
      r_24__13_ <= r_n_24__13_;
      r_24__12_ <= r_n_24__12_;
      r_24__11_ <= r_n_24__11_;
      r_24__10_ <= r_n_24__10_;
      r_24__9_ <= r_n_24__9_;
      r_24__8_ <= r_n_24__8_;
      r_24__7_ <= r_n_24__7_;
      r_24__6_ <= r_n_24__6_;
      r_24__5_ <= r_n_24__5_;
      r_24__4_ <= r_n_24__4_;
      r_24__3_ <= r_n_24__3_;
      r_24__2_ <= r_n_24__2_;
      r_24__1_ <= r_n_24__1_;
      r_24__0_ <= r_n_24__0_;
    end 
    if(N473) begin
      r_25__15_ <= r_n_25__15_;
      r_25__14_ <= r_n_25__14_;
      r_25__13_ <= r_n_25__13_;
      r_25__12_ <= r_n_25__12_;
      r_25__11_ <= r_n_25__11_;
      r_25__10_ <= r_n_25__10_;
      r_25__9_ <= r_n_25__9_;
      r_25__8_ <= r_n_25__8_;
      r_25__7_ <= r_n_25__7_;
      r_25__6_ <= r_n_25__6_;
      r_25__5_ <= r_n_25__5_;
      r_25__4_ <= r_n_25__4_;
      r_25__3_ <= r_n_25__3_;
      r_25__2_ <= r_n_25__2_;
      r_25__1_ <= r_n_25__1_;
      r_25__0_ <= r_n_25__0_;
    end 
    if(N474) begin
      r_26__15_ <= r_n_26__15_;
      r_26__14_ <= r_n_26__14_;
      r_26__13_ <= r_n_26__13_;
      r_26__12_ <= r_n_26__12_;
      r_26__11_ <= r_n_26__11_;
      r_26__10_ <= r_n_26__10_;
      r_26__9_ <= r_n_26__9_;
      r_26__8_ <= r_n_26__8_;
      r_26__7_ <= r_n_26__7_;
      r_26__6_ <= r_n_26__6_;
      r_26__5_ <= r_n_26__5_;
      r_26__4_ <= r_n_26__4_;
      r_26__3_ <= r_n_26__3_;
      r_26__2_ <= r_n_26__2_;
      r_26__1_ <= r_n_26__1_;
      r_26__0_ <= r_n_26__0_;
    end 
    if(N475) begin
      r_27__15_ <= r_n_27__15_;
      r_27__14_ <= r_n_27__14_;
      r_27__13_ <= r_n_27__13_;
      r_27__12_ <= r_n_27__12_;
      r_27__11_ <= r_n_27__11_;
      r_27__10_ <= r_n_27__10_;
      r_27__9_ <= r_n_27__9_;
      r_27__8_ <= r_n_27__8_;
      r_27__7_ <= r_n_27__7_;
      r_27__6_ <= r_n_27__6_;
      r_27__5_ <= r_n_27__5_;
      r_27__4_ <= r_n_27__4_;
      r_27__3_ <= r_n_27__3_;
      r_27__2_ <= r_n_27__2_;
      r_27__1_ <= r_n_27__1_;
      r_27__0_ <= r_n_27__0_;
    end 
    if(N476) begin
      r_28__15_ <= r_n_28__15_;
      r_28__14_ <= r_n_28__14_;
      r_28__13_ <= r_n_28__13_;
      r_28__12_ <= r_n_28__12_;
      r_28__11_ <= r_n_28__11_;
      r_28__10_ <= r_n_28__10_;
      r_28__9_ <= r_n_28__9_;
      r_28__8_ <= r_n_28__8_;
      r_28__7_ <= r_n_28__7_;
      r_28__6_ <= r_n_28__6_;
      r_28__5_ <= r_n_28__5_;
      r_28__4_ <= r_n_28__4_;
      r_28__3_ <= r_n_28__3_;
      r_28__2_ <= r_n_28__2_;
      r_28__1_ <= r_n_28__1_;
      r_28__0_ <= r_n_28__0_;
    end 
    if(N477) begin
      r_29__15_ <= r_n_29__15_;
      r_29__14_ <= r_n_29__14_;
      r_29__13_ <= r_n_29__13_;
      r_29__12_ <= r_n_29__12_;
      r_29__11_ <= r_n_29__11_;
      r_29__10_ <= r_n_29__10_;
      r_29__9_ <= r_n_29__9_;
      r_29__8_ <= r_n_29__8_;
      r_29__7_ <= r_n_29__7_;
      r_29__6_ <= r_n_29__6_;
      r_29__5_ <= r_n_29__5_;
      r_29__4_ <= r_n_29__4_;
      r_29__3_ <= r_n_29__3_;
      r_29__2_ <= r_n_29__2_;
      r_29__1_ <= r_n_29__1_;
      r_29__0_ <= r_n_29__0_;
    end 
    if(N478) begin
      r_30__15_ <= r_n_30__15_;
      r_30__14_ <= r_n_30__14_;
      r_30__13_ <= r_n_30__13_;
      r_30__12_ <= r_n_30__12_;
      r_30__11_ <= r_n_30__11_;
      r_30__10_ <= r_n_30__10_;
      r_30__9_ <= r_n_30__9_;
      r_30__8_ <= r_n_30__8_;
      r_30__7_ <= r_n_30__7_;
      r_30__6_ <= r_n_30__6_;
      r_30__5_ <= r_n_30__5_;
      r_30__4_ <= r_n_30__4_;
      r_30__3_ <= r_n_30__3_;
      r_30__2_ <= r_n_30__2_;
      r_30__1_ <= r_n_30__1_;
      r_30__0_ <= r_n_30__0_;
    end 
    if(N479) begin
      r_31__15_ <= r_n_31__15_;
      r_31__14_ <= r_n_31__14_;
      r_31__13_ <= r_n_31__13_;
      r_31__12_ <= r_n_31__12_;
      r_31__11_ <= r_n_31__11_;
      r_31__10_ <= r_n_31__10_;
      r_31__9_ <= r_n_31__9_;
      r_31__8_ <= r_n_31__8_;
      r_31__7_ <= r_n_31__7_;
      r_31__6_ <= r_n_31__6_;
      r_31__5_ <= r_n_31__5_;
      r_31__4_ <= r_n_31__4_;
      r_31__3_ <= r_n_31__3_;
      r_31__2_ <= r_n_31__2_;
      r_31__1_ <= r_n_31__1_;
      r_31__0_ <= r_n_31__0_;
    end 
    if(N480) begin
      r_32__15_ <= r_n_32__15_;
      r_32__14_ <= r_n_32__14_;
      r_32__13_ <= r_n_32__13_;
      r_32__12_ <= r_n_32__12_;
      r_32__11_ <= r_n_32__11_;
      r_32__10_ <= r_n_32__10_;
      r_32__9_ <= r_n_32__9_;
      r_32__8_ <= r_n_32__8_;
      r_32__7_ <= r_n_32__7_;
      r_32__6_ <= r_n_32__6_;
      r_32__5_ <= r_n_32__5_;
      r_32__4_ <= r_n_32__4_;
      r_32__3_ <= r_n_32__3_;
      r_32__2_ <= r_n_32__2_;
      r_32__1_ <= r_n_32__1_;
      r_32__0_ <= r_n_32__0_;
    end 
    if(N481) begin
      r_33__15_ <= r_n_33__15_;
      r_33__14_ <= r_n_33__14_;
      r_33__13_ <= r_n_33__13_;
      r_33__12_ <= r_n_33__12_;
      r_33__11_ <= r_n_33__11_;
      r_33__10_ <= r_n_33__10_;
      r_33__9_ <= r_n_33__9_;
      r_33__8_ <= r_n_33__8_;
      r_33__7_ <= r_n_33__7_;
      r_33__6_ <= r_n_33__6_;
      r_33__5_ <= r_n_33__5_;
      r_33__4_ <= r_n_33__4_;
      r_33__3_ <= r_n_33__3_;
      r_33__2_ <= r_n_33__2_;
      r_33__1_ <= r_n_33__1_;
      r_33__0_ <= r_n_33__0_;
    end 
    if(N482) begin
      r_34__15_ <= r_n_34__15_;
      r_34__14_ <= r_n_34__14_;
      r_34__13_ <= r_n_34__13_;
      r_34__12_ <= r_n_34__12_;
      r_34__11_ <= r_n_34__11_;
      r_34__10_ <= r_n_34__10_;
      r_34__9_ <= r_n_34__9_;
      r_34__8_ <= r_n_34__8_;
      r_34__7_ <= r_n_34__7_;
      r_34__6_ <= r_n_34__6_;
      r_34__5_ <= r_n_34__5_;
      r_34__4_ <= r_n_34__4_;
      r_34__3_ <= r_n_34__3_;
      r_34__2_ <= r_n_34__2_;
      r_34__1_ <= r_n_34__1_;
      r_34__0_ <= r_n_34__0_;
    end 
    if(N483) begin
      r_35__15_ <= r_n_35__15_;
      r_35__14_ <= r_n_35__14_;
      r_35__13_ <= r_n_35__13_;
      r_35__12_ <= r_n_35__12_;
      r_35__11_ <= r_n_35__11_;
      r_35__10_ <= r_n_35__10_;
      r_35__9_ <= r_n_35__9_;
      r_35__8_ <= r_n_35__8_;
      r_35__7_ <= r_n_35__7_;
      r_35__6_ <= r_n_35__6_;
      r_35__5_ <= r_n_35__5_;
      r_35__4_ <= r_n_35__4_;
      r_35__3_ <= r_n_35__3_;
      r_35__2_ <= r_n_35__2_;
      r_35__1_ <= r_n_35__1_;
      r_35__0_ <= r_n_35__0_;
    end 
    if(N484) begin
      r_36__15_ <= r_n_36__15_;
      r_36__14_ <= r_n_36__14_;
      r_36__13_ <= r_n_36__13_;
      r_36__12_ <= r_n_36__12_;
      r_36__11_ <= r_n_36__11_;
      r_36__10_ <= r_n_36__10_;
      r_36__9_ <= r_n_36__9_;
      r_36__8_ <= r_n_36__8_;
      r_36__7_ <= r_n_36__7_;
      r_36__6_ <= r_n_36__6_;
      r_36__5_ <= r_n_36__5_;
      r_36__4_ <= r_n_36__4_;
      r_36__3_ <= r_n_36__3_;
      r_36__2_ <= r_n_36__2_;
      r_36__1_ <= r_n_36__1_;
      r_36__0_ <= r_n_36__0_;
    end 
    if(N485) begin
      r_37__15_ <= r_n_37__15_;
      r_37__14_ <= r_n_37__14_;
      r_37__13_ <= r_n_37__13_;
      r_37__12_ <= r_n_37__12_;
      r_37__11_ <= r_n_37__11_;
      r_37__10_ <= r_n_37__10_;
      r_37__9_ <= r_n_37__9_;
      r_37__8_ <= r_n_37__8_;
      r_37__7_ <= r_n_37__7_;
      r_37__6_ <= r_n_37__6_;
      r_37__5_ <= r_n_37__5_;
      r_37__4_ <= r_n_37__4_;
      r_37__3_ <= r_n_37__3_;
      r_37__2_ <= r_n_37__2_;
      r_37__1_ <= r_n_37__1_;
      r_37__0_ <= r_n_37__0_;
    end 
    if(N486) begin
      r_38__15_ <= r_n_38__15_;
      r_38__14_ <= r_n_38__14_;
      r_38__13_ <= r_n_38__13_;
      r_38__12_ <= r_n_38__12_;
      r_38__11_ <= r_n_38__11_;
      r_38__10_ <= r_n_38__10_;
      r_38__9_ <= r_n_38__9_;
      r_38__8_ <= r_n_38__8_;
      r_38__7_ <= r_n_38__7_;
      r_38__6_ <= r_n_38__6_;
      r_38__5_ <= r_n_38__5_;
      r_38__4_ <= r_n_38__4_;
      r_38__3_ <= r_n_38__3_;
      r_38__2_ <= r_n_38__2_;
      r_38__1_ <= r_n_38__1_;
      r_38__0_ <= r_n_38__0_;
    end 
    if(N487) begin
      r_39__15_ <= r_n_39__15_;
      r_39__14_ <= r_n_39__14_;
      r_39__13_ <= r_n_39__13_;
      r_39__12_ <= r_n_39__12_;
      r_39__11_ <= r_n_39__11_;
      r_39__10_ <= r_n_39__10_;
      r_39__9_ <= r_n_39__9_;
      r_39__8_ <= r_n_39__8_;
      r_39__7_ <= r_n_39__7_;
      r_39__6_ <= r_n_39__6_;
      r_39__5_ <= r_n_39__5_;
      r_39__4_ <= r_n_39__4_;
      r_39__3_ <= r_n_39__3_;
      r_39__2_ <= r_n_39__2_;
      r_39__1_ <= r_n_39__1_;
      r_39__0_ <= r_n_39__0_;
    end 
    if(N488) begin
      r_40__15_ <= r_n_40__15_;
      r_40__14_ <= r_n_40__14_;
      r_40__13_ <= r_n_40__13_;
      r_40__12_ <= r_n_40__12_;
      r_40__11_ <= r_n_40__11_;
      r_40__10_ <= r_n_40__10_;
      r_40__9_ <= r_n_40__9_;
      r_40__8_ <= r_n_40__8_;
      r_40__7_ <= r_n_40__7_;
      r_40__6_ <= r_n_40__6_;
      r_40__5_ <= r_n_40__5_;
      r_40__4_ <= r_n_40__4_;
      r_40__3_ <= r_n_40__3_;
      r_40__2_ <= r_n_40__2_;
      r_40__1_ <= r_n_40__1_;
      r_40__0_ <= r_n_40__0_;
    end 
    if(N489) begin
      r_41__15_ <= r_n_41__15_;
      r_41__14_ <= r_n_41__14_;
      r_41__13_ <= r_n_41__13_;
      r_41__12_ <= r_n_41__12_;
      r_41__11_ <= r_n_41__11_;
      r_41__10_ <= r_n_41__10_;
      r_41__9_ <= r_n_41__9_;
      r_41__8_ <= r_n_41__8_;
      r_41__7_ <= r_n_41__7_;
      r_41__6_ <= r_n_41__6_;
      r_41__5_ <= r_n_41__5_;
      r_41__4_ <= r_n_41__4_;
      r_41__3_ <= r_n_41__3_;
      r_41__2_ <= r_n_41__2_;
      r_41__1_ <= r_n_41__1_;
      r_41__0_ <= r_n_41__0_;
    end 
    if(N490) begin
      r_42__15_ <= r_n_42__15_;
      r_42__14_ <= r_n_42__14_;
      r_42__13_ <= r_n_42__13_;
      r_42__12_ <= r_n_42__12_;
      r_42__11_ <= r_n_42__11_;
      r_42__10_ <= r_n_42__10_;
      r_42__9_ <= r_n_42__9_;
      r_42__8_ <= r_n_42__8_;
      r_42__7_ <= r_n_42__7_;
      r_42__6_ <= r_n_42__6_;
      r_42__5_ <= r_n_42__5_;
      r_42__4_ <= r_n_42__4_;
      r_42__3_ <= r_n_42__3_;
      r_42__2_ <= r_n_42__2_;
      r_42__1_ <= r_n_42__1_;
      r_42__0_ <= r_n_42__0_;
    end 
    if(N491) begin
      r_43__15_ <= r_n_43__15_;
      r_43__14_ <= r_n_43__14_;
      r_43__13_ <= r_n_43__13_;
      r_43__12_ <= r_n_43__12_;
      r_43__11_ <= r_n_43__11_;
      r_43__10_ <= r_n_43__10_;
      r_43__9_ <= r_n_43__9_;
      r_43__8_ <= r_n_43__8_;
      r_43__7_ <= r_n_43__7_;
      r_43__6_ <= r_n_43__6_;
      r_43__5_ <= r_n_43__5_;
      r_43__4_ <= r_n_43__4_;
      r_43__3_ <= r_n_43__3_;
      r_43__2_ <= r_n_43__2_;
      r_43__1_ <= r_n_43__1_;
      r_43__0_ <= r_n_43__0_;
    end 
    if(N492) begin
      r_44__15_ <= r_n_44__15_;
      r_44__14_ <= r_n_44__14_;
      r_44__13_ <= r_n_44__13_;
      r_44__12_ <= r_n_44__12_;
      r_44__11_ <= r_n_44__11_;
      r_44__10_ <= r_n_44__10_;
      r_44__9_ <= r_n_44__9_;
      r_44__8_ <= r_n_44__8_;
      r_44__7_ <= r_n_44__7_;
      r_44__6_ <= r_n_44__6_;
      r_44__5_ <= r_n_44__5_;
      r_44__4_ <= r_n_44__4_;
      r_44__3_ <= r_n_44__3_;
      r_44__2_ <= r_n_44__2_;
      r_44__1_ <= r_n_44__1_;
      r_44__0_ <= r_n_44__0_;
    end 
    if(N493) begin
      r_45__15_ <= r_n_45__15_;
      r_45__14_ <= r_n_45__14_;
      r_45__13_ <= r_n_45__13_;
      r_45__12_ <= r_n_45__12_;
      r_45__11_ <= r_n_45__11_;
      r_45__10_ <= r_n_45__10_;
      r_45__9_ <= r_n_45__9_;
      r_45__8_ <= r_n_45__8_;
      r_45__7_ <= r_n_45__7_;
      r_45__6_ <= r_n_45__6_;
      r_45__5_ <= r_n_45__5_;
      r_45__4_ <= r_n_45__4_;
      r_45__3_ <= r_n_45__3_;
      r_45__2_ <= r_n_45__2_;
      r_45__1_ <= r_n_45__1_;
      r_45__0_ <= r_n_45__0_;
    end 
    if(N494) begin
      r_46__15_ <= r_n_46__15_;
      r_46__14_ <= r_n_46__14_;
      r_46__13_ <= r_n_46__13_;
      r_46__12_ <= r_n_46__12_;
      r_46__11_ <= r_n_46__11_;
      r_46__10_ <= r_n_46__10_;
      r_46__9_ <= r_n_46__9_;
      r_46__8_ <= r_n_46__8_;
      r_46__7_ <= r_n_46__7_;
      r_46__6_ <= r_n_46__6_;
      r_46__5_ <= r_n_46__5_;
      r_46__4_ <= r_n_46__4_;
      r_46__3_ <= r_n_46__3_;
      r_46__2_ <= r_n_46__2_;
      r_46__1_ <= r_n_46__1_;
      r_46__0_ <= r_n_46__0_;
    end 
    if(N495) begin
      r_47__15_ <= r_n_47__15_;
      r_47__14_ <= r_n_47__14_;
      r_47__13_ <= r_n_47__13_;
      r_47__12_ <= r_n_47__12_;
      r_47__11_ <= r_n_47__11_;
      r_47__10_ <= r_n_47__10_;
      r_47__9_ <= r_n_47__9_;
      r_47__8_ <= r_n_47__8_;
      r_47__7_ <= r_n_47__7_;
      r_47__6_ <= r_n_47__6_;
      r_47__5_ <= r_n_47__5_;
      r_47__4_ <= r_n_47__4_;
      r_47__3_ <= r_n_47__3_;
      r_47__2_ <= r_n_47__2_;
      r_47__1_ <= r_n_47__1_;
      r_47__0_ <= r_n_47__0_;
    end 
    if(N496) begin
      r_48__15_ <= r_n_48__15_;
      r_48__14_ <= r_n_48__14_;
      r_48__13_ <= r_n_48__13_;
      r_48__12_ <= r_n_48__12_;
      r_48__11_ <= r_n_48__11_;
      r_48__10_ <= r_n_48__10_;
      r_48__9_ <= r_n_48__9_;
      r_48__8_ <= r_n_48__8_;
      r_48__7_ <= r_n_48__7_;
      r_48__6_ <= r_n_48__6_;
      r_48__5_ <= r_n_48__5_;
      r_48__4_ <= r_n_48__4_;
      r_48__3_ <= r_n_48__3_;
      r_48__2_ <= r_n_48__2_;
      r_48__1_ <= r_n_48__1_;
      r_48__0_ <= r_n_48__0_;
    end 
    if(N497) begin
      r_49__15_ <= r_n_49__15_;
      r_49__14_ <= r_n_49__14_;
      r_49__13_ <= r_n_49__13_;
      r_49__12_ <= r_n_49__12_;
      r_49__11_ <= r_n_49__11_;
      r_49__10_ <= r_n_49__10_;
      r_49__9_ <= r_n_49__9_;
      r_49__8_ <= r_n_49__8_;
      r_49__7_ <= r_n_49__7_;
      r_49__6_ <= r_n_49__6_;
      r_49__5_ <= r_n_49__5_;
      r_49__4_ <= r_n_49__4_;
      r_49__3_ <= r_n_49__3_;
      r_49__2_ <= r_n_49__2_;
      r_49__1_ <= r_n_49__1_;
      r_49__0_ <= r_n_49__0_;
    end 
    if(N498) begin
      r_50__15_ <= r_n_50__15_;
      r_50__14_ <= r_n_50__14_;
      r_50__13_ <= r_n_50__13_;
      r_50__12_ <= r_n_50__12_;
      r_50__11_ <= r_n_50__11_;
      r_50__10_ <= r_n_50__10_;
      r_50__9_ <= r_n_50__9_;
      r_50__8_ <= r_n_50__8_;
      r_50__7_ <= r_n_50__7_;
      r_50__6_ <= r_n_50__6_;
      r_50__5_ <= r_n_50__5_;
      r_50__4_ <= r_n_50__4_;
      r_50__3_ <= r_n_50__3_;
      r_50__2_ <= r_n_50__2_;
      r_50__1_ <= r_n_50__1_;
      r_50__0_ <= r_n_50__0_;
    end 
    if(N499) begin
      r_51__15_ <= r_n_51__15_;
      r_51__14_ <= r_n_51__14_;
      r_51__13_ <= r_n_51__13_;
      r_51__12_ <= r_n_51__12_;
      r_51__11_ <= r_n_51__11_;
      r_51__10_ <= r_n_51__10_;
      r_51__9_ <= r_n_51__9_;
      r_51__8_ <= r_n_51__8_;
      r_51__7_ <= r_n_51__7_;
      r_51__6_ <= r_n_51__6_;
      r_51__5_ <= r_n_51__5_;
      r_51__4_ <= r_n_51__4_;
      r_51__3_ <= r_n_51__3_;
      r_51__2_ <= r_n_51__2_;
      r_51__1_ <= r_n_51__1_;
      r_51__0_ <= r_n_51__0_;
    end 
    if(N500) begin
      r_52__15_ <= r_n_52__15_;
      r_52__14_ <= r_n_52__14_;
      r_52__13_ <= r_n_52__13_;
      r_52__12_ <= r_n_52__12_;
      r_52__11_ <= r_n_52__11_;
      r_52__10_ <= r_n_52__10_;
      r_52__9_ <= r_n_52__9_;
      r_52__8_ <= r_n_52__8_;
      r_52__7_ <= r_n_52__7_;
      r_52__6_ <= r_n_52__6_;
      r_52__5_ <= r_n_52__5_;
      r_52__4_ <= r_n_52__4_;
      r_52__3_ <= r_n_52__3_;
      r_52__2_ <= r_n_52__2_;
      r_52__1_ <= r_n_52__1_;
      r_52__0_ <= r_n_52__0_;
    end 
    if(N501) begin
      r_53__15_ <= r_n_53__15_;
      r_53__14_ <= r_n_53__14_;
      r_53__13_ <= r_n_53__13_;
      r_53__12_ <= r_n_53__12_;
      r_53__11_ <= r_n_53__11_;
      r_53__10_ <= r_n_53__10_;
      r_53__9_ <= r_n_53__9_;
      r_53__8_ <= r_n_53__8_;
      r_53__7_ <= r_n_53__7_;
      r_53__6_ <= r_n_53__6_;
      r_53__5_ <= r_n_53__5_;
      r_53__4_ <= r_n_53__4_;
      r_53__3_ <= r_n_53__3_;
      r_53__2_ <= r_n_53__2_;
      r_53__1_ <= r_n_53__1_;
      r_53__0_ <= r_n_53__0_;
    end 
    if(N502) begin
      r_54__15_ <= r_n_54__15_;
      r_54__14_ <= r_n_54__14_;
      r_54__13_ <= r_n_54__13_;
      r_54__12_ <= r_n_54__12_;
      r_54__11_ <= r_n_54__11_;
      r_54__10_ <= r_n_54__10_;
      r_54__9_ <= r_n_54__9_;
      r_54__8_ <= r_n_54__8_;
      r_54__7_ <= r_n_54__7_;
      r_54__6_ <= r_n_54__6_;
      r_54__5_ <= r_n_54__5_;
      r_54__4_ <= r_n_54__4_;
      r_54__3_ <= r_n_54__3_;
      r_54__2_ <= r_n_54__2_;
      r_54__1_ <= r_n_54__1_;
      r_54__0_ <= r_n_54__0_;
    end 
    if(N503) begin
      r_55__15_ <= r_n_55__15_;
      r_55__14_ <= r_n_55__14_;
      r_55__13_ <= r_n_55__13_;
      r_55__12_ <= r_n_55__12_;
      r_55__11_ <= r_n_55__11_;
      r_55__10_ <= r_n_55__10_;
      r_55__9_ <= r_n_55__9_;
      r_55__8_ <= r_n_55__8_;
      r_55__7_ <= r_n_55__7_;
      r_55__6_ <= r_n_55__6_;
      r_55__5_ <= r_n_55__5_;
      r_55__4_ <= r_n_55__4_;
      r_55__3_ <= r_n_55__3_;
      r_55__2_ <= r_n_55__2_;
      r_55__1_ <= r_n_55__1_;
      r_55__0_ <= r_n_55__0_;
    end 
    if(N504) begin
      r_56__15_ <= r_n_56__15_;
      r_56__14_ <= r_n_56__14_;
      r_56__13_ <= r_n_56__13_;
      r_56__12_ <= r_n_56__12_;
      r_56__11_ <= r_n_56__11_;
      r_56__10_ <= r_n_56__10_;
      r_56__9_ <= r_n_56__9_;
      r_56__8_ <= r_n_56__8_;
      r_56__7_ <= r_n_56__7_;
      r_56__6_ <= r_n_56__6_;
      r_56__5_ <= r_n_56__5_;
      r_56__4_ <= r_n_56__4_;
      r_56__3_ <= r_n_56__3_;
      r_56__2_ <= r_n_56__2_;
      r_56__1_ <= r_n_56__1_;
      r_56__0_ <= r_n_56__0_;
    end 
    if(N505) begin
      r_57__15_ <= r_n_57__15_;
      r_57__14_ <= r_n_57__14_;
      r_57__13_ <= r_n_57__13_;
      r_57__12_ <= r_n_57__12_;
      r_57__11_ <= r_n_57__11_;
      r_57__10_ <= r_n_57__10_;
      r_57__9_ <= r_n_57__9_;
      r_57__8_ <= r_n_57__8_;
      r_57__7_ <= r_n_57__7_;
      r_57__6_ <= r_n_57__6_;
      r_57__5_ <= r_n_57__5_;
      r_57__4_ <= r_n_57__4_;
      r_57__3_ <= r_n_57__3_;
      r_57__2_ <= r_n_57__2_;
      r_57__1_ <= r_n_57__1_;
      r_57__0_ <= r_n_57__0_;
    end 
    if(N506) begin
      r_58__15_ <= r_n_58__15_;
      r_58__14_ <= r_n_58__14_;
      r_58__13_ <= r_n_58__13_;
      r_58__12_ <= r_n_58__12_;
      r_58__11_ <= r_n_58__11_;
      r_58__10_ <= r_n_58__10_;
      r_58__9_ <= r_n_58__9_;
      r_58__8_ <= r_n_58__8_;
      r_58__7_ <= r_n_58__7_;
      r_58__6_ <= r_n_58__6_;
      r_58__5_ <= r_n_58__5_;
      r_58__4_ <= r_n_58__4_;
      r_58__3_ <= r_n_58__3_;
      r_58__2_ <= r_n_58__2_;
      r_58__1_ <= r_n_58__1_;
      r_58__0_ <= r_n_58__0_;
    end 
    if(N507) begin
      r_59__15_ <= r_n_59__15_;
      r_59__14_ <= r_n_59__14_;
      r_59__13_ <= r_n_59__13_;
      r_59__12_ <= r_n_59__12_;
      r_59__11_ <= r_n_59__11_;
      r_59__10_ <= r_n_59__10_;
      r_59__9_ <= r_n_59__9_;
      r_59__8_ <= r_n_59__8_;
      r_59__7_ <= r_n_59__7_;
      r_59__6_ <= r_n_59__6_;
      r_59__5_ <= r_n_59__5_;
      r_59__4_ <= r_n_59__4_;
      r_59__3_ <= r_n_59__3_;
      r_59__2_ <= r_n_59__2_;
      r_59__1_ <= r_n_59__1_;
      r_59__0_ <= r_n_59__0_;
    end 
    if(N508) begin
      r_60__15_ <= r_n_60__15_;
      r_60__14_ <= r_n_60__14_;
      r_60__13_ <= r_n_60__13_;
      r_60__12_ <= r_n_60__12_;
      r_60__11_ <= r_n_60__11_;
      r_60__10_ <= r_n_60__10_;
      r_60__9_ <= r_n_60__9_;
      r_60__8_ <= r_n_60__8_;
      r_60__7_ <= r_n_60__7_;
      r_60__6_ <= r_n_60__6_;
      r_60__5_ <= r_n_60__5_;
      r_60__4_ <= r_n_60__4_;
      r_60__3_ <= r_n_60__3_;
      r_60__2_ <= r_n_60__2_;
      r_60__1_ <= r_n_60__1_;
      r_60__0_ <= r_n_60__0_;
    end 
    if(N509) begin
      r_61__15_ <= r_n_61__15_;
      r_61__14_ <= r_n_61__14_;
      r_61__13_ <= r_n_61__13_;
      r_61__12_ <= r_n_61__12_;
      r_61__11_ <= r_n_61__11_;
      r_61__10_ <= r_n_61__10_;
      r_61__9_ <= r_n_61__9_;
      r_61__8_ <= r_n_61__8_;
      r_61__7_ <= r_n_61__7_;
      r_61__6_ <= r_n_61__6_;
      r_61__5_ <= r_n_61__5_;
      r_61__4_ <= r_n_61__4_;
      r_61__3_ <= r_n_61__3_;
      r_61__2_ <= r_n_61__2_;
      r_61__1_ <= r_n_61__1_;
      r_61__0_ <= r_n_61__0_;
    end 
    if(N510) begin
      r_62__15_ <= r_n_62__15_;
      r_62__14_ <= r_n_62__14_;
      r_62__13_ <= r_n_62__13_;
      r_62__12_ <= r_n_62__12_;
      r_62__11_ <= r_n_62__11_;
      r_62__10_ <= r_n_62__10_;
      r_62__9_ <= r_n_62__9_;
      r_62__8_ <= r_n_62__8_;
      r_62__7_ <= r_n_62__7_;
      r_62__6_ <= r_n_62__6_;
      r_62__5_ <= r_n_62__5_;
      r_62__4_ <= r_n_62__4_;
      r_62__3_ <= r_n_62__3_;
      r_62__2_ <= r_n_62__2_;
      r_62__1_ <= r_n_62__1_;
      r_62__0_ <= r_n_62__0_;
    end 
    if(N511) begin
      r_63__15_ <= r_n_63__15_;
      r_63__14_ <= r_n_63__14_;
      r_63__13_ <= r_n_63__13_;
      r_63__12_ <= r_n_63__12_;
      r_63__11_ <= r_n_63__11_;
      r_63__10_ <= r_n_63__10_;
      r_63__9_ <= r_n_63__9_;
      r_63__8_ <= r_n_63__8_;
      r_63__7_ <= r_n_63__7_;
      r_63__6_ <= r_n_63__6_;
      r_63__5_ <= r_n_63__5_;
      r_63__4_ <= r_n_63__4_;
      r_63__3_ <= r_n_63__3_;
      r_63__2_ <= r_n_63__2_;
      r_63__1_ <= r_n_63__1_;
      r_63__0_ <= r_n_63__0_;
    end 
  end


endmodule

