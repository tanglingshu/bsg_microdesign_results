

module top
(
  clk_i,
  data_i,
  data_o
);

  input [63:0] data_i;
  output [63:0] data_o;
  input clk_i;

  bsg_dff_chain
  wrapper
  (
    .data_i(data_i),
    .data_o(data_o),
    .clk_i(clk_i)
  );


endmodule



module bsg_dff_width_p64
(
  clk_i,
  data_i,
  data_o
);

  input [63:0] data_i;
  output [63:0] data_o;
  input clk_i;
  reg [63:0] data_o;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { data_o[63:0] } <= { data_i[63:0] };
    end 
  end


endmodule



module bsg_dff_chain
(
  clk_i,
  data_i,
  data_o
);

  input [63:0] data_i;
  output [63:0] data_o;
  input clk_i;
  wire [63:0] data_o;
  wire chained_data_delayed_63__63_,chained_data_delayed_63__62_,
  chained_data_delayed_63__61_,chained_data_delayed_63__60_,chained_data_delayed_63__59_,
  chained_data_delayed_63__58_,chained_data_delayed_63__57_,chained_data_delayed_63__56_,
  chained_data_delayed_63__55_,chained_data_delayed_63__54_,chained_data_delayed_63__53_,
  chained_data_delayed_63__52_,chained_data_delayed_63__51_,
  chained_data_delayed_63__50_,chained_data_delayed_63__49_,chained_data_delayed_63__48_,
  chained_data_delayed_63__47_,chained_data_delayed_63__46_,chained_data_delayed_63__45_,
  chained_data_delayed_63__44_,chained_data_delayed_63__43_,chained_data_delayed_63__42_,
  chained_data_delayed_63__41_,chained_data_delayed_63__40_,
  chained_data_delayed_63__39_,chained_data_delayed_63__38_,chained_data_delayed_63__37_,
  chained_data_delayed_63__36_,chained_data_delayed_63__35_,chained_data_delayed_63__34_,
  chained_data_delayed_63__33_,chained_data_delayed_63__32_,chained_data_delayed_63__31_,
  chained_data_delayed_63__30_,chained_data_delayed_63__29_,
  chained_data_delayed_63__28_,chained_data_delayed_63__27_,chained_data_delayed_63__26_,
  chained_data_delayed_63__25_,chained_data_delayed_63__24_,chained_data_delayed_63__23_,
  chained_data_delayed_63__22_,chained_data_delayed_63__21_,chained_data_delayed_63__20_,
  chained_data_delayed_63__19_,chained_data_delayed_63__18_,
  chained_data_delayed_63__17_,chained_data_delayed_63__16_,chained_data_delayed_63__15_,
  chained_data_delayed_63__14_,chained_data_delayed_63__13_,chained_data_delayed_63__12_,
  chained_data_delayed_63__11_,chained_data_delayed_63__10_,chained_data_delayed_63__9_,
  chained_data_delayed_63__8_,chained_data_delayed_63__7_,chained_data_delayed_63__6_,
  chained_data_delayed_63__5_,chained_data_delayed_63__4_,
  chained_data_delayed_63__3_,chained_data_delayed_63__2_,chained_data_delayed_63__1_,
  chained_data_delayed_63__0_,chained_data_delayed_62__63_,chained_data_delayed_62__62_,
  chained_data_delayed_62__61_,chained_data_delayed_62__60_,chained_data_delayed_62__59_,
  chained_data_delayed_62__58_,chained_data_delayed_62__57_,chained_data_delayed_62__56_,
  chained_data_delayed_62__55_,chained_data_delayed_62__54_,
  chained_data_delayed_62__53_,chained_data_delayed_62__52_,chained_data_delayed_62__51_,
  chained_data_delayed_62__50_,chained_data_delayed_62__49_,chained_data_delayed_62__48_,
  chained_data_delayed_62__47_,chained_data_delayed_62__46_,chained_data_delayed_62__45_,
  chained_data_delayed_62__44_,chained_data_delayed_62__43_,
  chained_data_delayed_62__42_,chained_data_delayed_62__41_,chained_data_delayed_62__40_,
  chained_data_delayed_62__39_,chained_data_delayed_62__38_,chained_data_delayed_62__37_,
  chained_data_delayed_62__36_,chained_data_delayed_62__35_,chained_data_delayed_62__34_,
  chained_data_delayed_62__33_,chained_data_delayed_62__32_,
  chained_data_delayed_62__31_,chained_data_delayed_62__30_,chained_data_delayed_62__29_,
  chained_data_delayed_62__28_,chained_data_delayed_62__27_,chained_data_delayed_62__26_,
  chained_data_delayed_62__25_,chained_data_delayed_62__24_,chained_data_delayed_62__23_,
  chained_data_delayed_62__22_,chained_data_delayed_62__21_,
  chained_data_delayed_62__20_,chained_data_delayed_62__19_,chained_data_delayed_62__18_,
  chained_data_delayed_62__17_,chained_data_delayed_62__16_,chained_data_delayed_62__15_,
  chained_data_delayed_62__14_,chained_data_delayed_62__13_,chained_data_delayed_62__12_,
  chained_data_delayed_62__11_,chained_data_delayed_62__10_,chained_data_delayed_62__9_,
  chained_data_delayed_62__8_,chained_data_delayed_62__7_,
  chained_data_delayed_62__6_,chained_data_delayed_62__5_,chained_data_delayed_62__4_,
  chained_data_delayed_62__3_,chained_data_delayed_62__2_,chained_data_delayed_62__1_,
  chained_data_delayed_62__0_,chained_data_delayed_61__63_,chained_data_delayed_61__62_,
  chained_data_delayed_61__61_,chained_data_delayed_61__60_,chained_data_delayed_61__59_,
  chained_data_delayed_61__58_,chained_data_delayed_61__57_,
  chained_data_delayed_61__56_,chained_data_delayed_61__55_,chained_data_delayed_61__54_,
  chained_data_delayed_61__53_,chained_data_delayed_61__52_,chained_data_delayed_61__51_,
  chained_data_delayed_61__50_,chained_data_delayed_61__49_,chained_data_delayed_61__48_,
  chained_data_delayed_61__47_,chained_data_delayed_61__46_,
  chained_data_delayed_61__45_,chained_data_delayed_61__44_,chained_data_delayed_61__43_,
  chained_data_delayed_61__42_,chained_data_delayed_61__41_,chained_data_delayed_61__40_,
  chained_data_delayed_61__39_,chained_data_delayed_61__38_,chained_data_delayed_61__37_,
  chained_data_delayed_61__36_,chained_data_delayed_61__35_,
  chained_data_delayed_61__34_,chained_data_delayed_61__33_,chained_data_delayed_61__32_,
  chained_data_delayed_61__31_,chained_data_delayed_61__30_,chained_data_delayed_61__29_,
  chained_data_delayed_61__28_,chained_data_delayed_61__27_,chained_data_delayed_61__26_,
  chained_data_delayed_61__25_,chained_data_delayed_61__24_,
  chained_data_delayed_61__23_,chained_data_delayed_61__22_,chained_data_delayed_61__21_,
  chained_data_delayed_61__20_,chained_data_delayed_61__19_,chained_data_delayed_61__18_,
  chained_data_delayed_61__17_,chained_data_delayed_61__16_,chained_data_delayed_61__15_,
  chained_data_delayed_61__14_,chained_data_delayed_61__13_,chained_data_delayed_61__12_,
  chained_data_delayed_61__11_,chained_data_delayed_61__10_,
  chained_data_delayed_61__9_,chained_data_delayed_61__8_,chained_data_delayed_61__7_,
  chained_data_delayed_61__6_,chained_data_delayed_61__5_,chained_data_delayed_61__4_,
  chained_data_delayed_61__3_,chained_data_delayed_61__2_,chained_data_delayed_61__1_,
  chained_data_delayed_61__0_,chained_data_delayed_60__63_,chained_data_delayed_60__62_,
  chained_data_delayed_60__61_,chained_data_delayed_60__60_,
  chained_data_delayed_60__59_,chained_data_delayed_60__58_,chained_data_delayed_60__57_,
  chained_data_delayed_60__56_,chained_data_delayed_60__55_,chained_data_delayed_60__54_,
  chained_data_delayed_60__53_,chained_data_delayed_60__52_,chained_data_delayed_60__51_,
  chained_data_delayed_60__50_,chained_data_delayed_60__49_,
  chained_data_delayed_60__48_,chained_data_delayed_60__47_,chained_data_delayed_60__46_,
  chained_data_delayed_60__45_,chained_data_delayed_60__44_,chained_data_delayed_60__43_,
  chained_data_delayed_60__42_,chained_data_delayed_60__41_,chained_data_delayed_60__40_,
  chained_data_delayed_60__39_,chained_data_delayed_60__38_,
  chained_data_delayed_60__37_,chained_data_delayed_60__36_,chained_data_delayed_60__35_,
  chained_data_delayed_60__34_,chained_data_delayed_60__33_,chained_data_delayed_60__32_,
  chained_data_delayed_60__31_,chained_data_delayed_60__30_,chained_data_delayed_60__29_,
  chained_data_delayed_60__28_,chained_data_delayed_60__27_,chained_data_delayed_60__26_,
  chained_data_delayed_60__25_,chained_data_delayed_60__24_,
  chained_data_delayed_60__23_,chained_data_delayed_60__22_,chained_data_delayed_60__21_,
  chained_data_delayed_60__20_,chained_data_delayed_60__19_,chained_data_delayed_60__18_,
  chained_data_delayed_60__17_,chained_data_delayed_60__16_,chained_data_delayed_60__15_,
  chained_data_delayed_60__14_,chained_data_delayed_60__13_,
  chained_data_delayed_60__12_,chained_data_delayed_60__11_,chained_data_delayed_60__10_,
  chained_data_delayed_60__9_,chained_data_delayed_60__8_,chained_data_delayed_60__7_,
  chained_data_delayed_60__6_,chained_data_delayed_60__5_,chained_data_delayed_60__4_,
  chained_data_delayed_60__3_,chained_data_delayed_60__2_,chained_data_delayed_60__1_,
  chained_data_delayed_60__0_,chained_data_delayed_59__63_,
  chained_data_delayed_59__62_,chained_data_delayed_59__61_,chained_data_delayed_59__60_,
  chained_data_delayed_59__59_,chained_data_delayed_59__58_,chained_data_delayed_59__57_,
  chained_data_delayed_59__56_,chained_data_delayed_59__55_,chained_data_delayed_59__54_,
  chained_data_delayed_59__53_,chained_data_delayed_59__52_,
  chained_data_delayed_59__51_,chained_data_delayed_59__50_,chained_data_delayed_59__49_,
  chained_data_delayed_59__48_,chained_data_delayed_59__47_,chained_data_delayed_59__46_,
  chained_data_delayed_59__45_,chained_data_delayed_59__44_,chained_data_delayed_59__43_,
  chained_data_delayed_59__42_,chained_data_delayed_59__41_,chained_data_delayed_59__40_,
  chained_data_delayed_59__39_,chained_data_delayed_59__38_,
  chained_data_delayed_59__37_,chained_data_delayed_59__36_,chained_data_delayed_59__35_,
  chained_data_delayed_59__34_,chained_data_delayed_59__33_,chained_data_delayed_59__32_,
  chained_data_delayed_59__31_,chained_data_delayed_59__30_,chained_data_delayed_59__29_,
  chained_data_delayed_59__28_,chained_data_delayed_59__27_,
  chained_data_delayed_59__26_,chained_data_delayed_59__25_,chained_data_delayed_59__24_,
  chained_data_delayed_59__23_,chained_data_delayed_59__22_,chained_data_delayed_59__21_,
  chained_data_delayed_59__20_,chained_data_delayed_59__19_,chained_data_delayed_59__18_,
  chained_data_delayed_59__17_,chained_data_delayed_59__16_,
  chained_data_delayed_59__15_,chained_data_delayed_59__14_,chained_data_delayed_59__13_,
  chained_data_delayed_59__12_,chained_data_delayed_59__11_,chained_data_delayed_59__10_,
  chained_data_delayed_59__9_,chained_data_delayed_59__8_,chained_data_delayed_59__7_,
  chained_data_delayed_59__6_,chained_data_delayed_59__5_,chained_data_delayed_59__4_,
  chained_data_delayed_59__3_,chained_data_delayed_59__2_,
  chained_data_delayed_59__1_,chained_data_delayed_59__0_,chained_data_delayed_58__63_,
  chained_data_delayed_58__62_,chained_data_delayed_58__61_,chained_data_delayed_58__60_,
  chained_data_delayed_58__59_,chained_data_delayed_58__58_,chained_data_delayed_58__57_,
  chained_data_delayed_58__56_,chained_data_delayed_58__55_,chained_data_delayed_58__54_,
  chained_data_delayed_58__53_,chained_data_delayed_58__52_,
  chained_data_delayed_58__51_,chained_data_delayed_58__50_,chained_data_delayed_58__49_,
  chained_data_delayed_58__48_,chained_data_delayed_58__47_,chained_data_delayed_58__46_,
  chained_data_delayed_58__45_,chained_data_delayed_58__44_,chained_data_delayed_58__43_,
  chained_data_delayed_58__42_,chained_data_delayed_58__41_,
  chained_data_delayed_58__40_,chained_data_delayed_58__39_,chained_data_delayed_58__38_,
  chained_data_delayed_58__37_,chained_data_delayed_58__36_,chained_data_delayed_58__35_,
  chained_data_delayed_58__34_,chained_data_delayed_58__33_,chained_data_delayed_58__32_,
  chained_data_delayed_58__31_,chained_data_delayed_58__30_,
  chained_data_delayed_58__29_,chained_data_delayed_58__28_,chained_data_delayed_58__27_,
  chained_data_delayed_58__26_,chained_data_delayed_58__25_,chained_data_delayed_58__24_,
  chained_data_delayed_58__23_,chained_data_delayed_58__22_,chained_data_delayed_58__21_,
  chained_data_delayed_58__20_,chained_data_delayed_58__19_,
  chained_data_delayed_58__18_,chained_data_delayed_58__17_,chained_data_delayed_58__16_,
  chained_data_delayed_58__15_,chained_data_delayed_58__14_,chained_data_delayed_58__13_,
  chained_data_delayed_58__12_,chained_data_delayed_58__11_,chained_data_delayed_58__10_,
  chained_data_delayed_58__9_,chained_data_delayed_58__8_,chained_data_delayed_58__7_,
  chained_data_delayed_58__6_,chained_data_delayed_58__5_,
  chained_data_delayed_58__4_,chained_data_delayed_58__3_,chained_data_delayed_58__2_,
  chained_data_delayed_58__1_,chained_data_delayed_58__0_,chained_data_delayed_57__63_,
  chained_data_delayed_57__62_,chained_data_delayed_57__61_,chained_data_delayed_57__60_,
  chained_data_delayed_57__59_,chained_data_delayed_57__58_,chained_data_delayed_57__57_,
  chained_data_delayed_57__56_,chained_data_delayed_57__55_,
  chained_data_delayed_57__54_,chained_data_delayed_57__53_,chained_data_delayed_57__52_,
  chained_data_delayed_57__51_,chained_data_delayed_57__50_,chained_data_delayed_57__49_,
  chained_data_delayed_57__48_,chained_data_delayed_57__47_,chained_data_delayed_57__46_,
  chained_data_delayed_57__45_,chained_data_delayed_57__44_,
  chained_data_delayed_57__43_,chained_data_delayed_57__42_,chained_data_delayed_57__41_,
  chained_data_delayed_57__40_,chained_data_delayed_57__39_,chained_data_delayed_57__38_,
  chained_data_delayed_57__37_,chained_data_delayed_57__36_,chained_data_delayed_57__35_,
  chained_data_delayed_57__34_,chained_data_delayed_57__33_,
  chained_data_delayed_57__32_,chained_data_delayed_57__31_,chained_data_delayed_57__30_,
  chained_data_delayed_57__29_,chained_data_delayed_57__28_,chained_data_delayed_57__27_,
  chained_data_delayed_57__26_,chained_data_delayed_57__25_,chained_data_delayed_57__24_,
  chained_data_delayed_57__23_,chained_data_delayed_57__22_,
  chained_data_delayed_57__21_,chained_data_delayed_57__20_,chained_data_delayed_57__19_,
  chained_data_delayed_57__18_,chained_data_delayed_57__17_,chained_data_delayed_57__16_,
  chained_data_delayed_57__15_,chained_data_delayed_57__14_,chained_data_delayed_57__13_,
  chained_data_delayed_57__12_,chained_data_delayed_57__11_,
  chained_data_delayed_57__10_,chained_data_delayed_57__9_,chained_data_delayed_57__8_,
  chained_data_delayed_57__7_,chained_data_delayed_57__6_,chained_data_delayed_57__5_,
  chained_data_delayed_57__4_,chained_data_delayed_57__3_,chained_data_delayed_57__2_,
  chained_data_delayed_57__1_,chained_data_delayed_57__0_,chained_data_delayed_8__63_,
  chained_data_delayed_8__62_,chained_data_delayed_8__61_,chained_data_delayed_8__60_,
  chained_data_delayed_8__59_,chained_data_delayed_8__58_,chained_data_delayed_8__57_,
  chained_data_delayed_8__56_,chained_data_delayed_8__55_,
  chained_data_delayed_8__54_,chained_data_delayed_8__53_,chained_data_delayed_8__52_,
  chained_data_delayed_8__51_,chained_data_delayed_8__50_,chained_data_delayed_8__49_,
  chained_data_delayed_8__48_,chained_data_delayed_8__47_,chained_data_delayed_8__46_,
  chained_data_delayed_8__45_,chained_data_delayed_8__44_,chained_data_delayed_8__43_,
  chained_data_delayed_8__42_,chained_data_delayed_8__41_,chained_data_delayed_8__40_,
  chained_data_delayed_8__39_,chained_data_delayed_8__38_,chained_data_delayed_8__37_,
  chained_data_delayed_8__36_,chained_data_delayed_8__35_,
  chained_data_delayed_8__34_,chained_data_delayed_8__33_,chained_data_delayed_8__32_,
  chained_data_delayed_8__31_,chained_data_delayed_8__30_,chained_data_delayed_8__29_,
  chained_data_delayed_8__28_,chained_data_delayed_8__27_,chained_data_delayed_8__26_,
  chained_data_delayed_8__25_,chained_data_delayed_8__24_,chained_data_delayed_8__23_,
  chained_data_delayed_8__22_,chained_data_delayed_8__21_,chained_data_delayed_8__20_,
  chained_data_delayed_8__19_,chained_data_delayed_8__18_,chained_data_delayed_8__17_,
  chained_data_delayed_8__16_,chained_data_delayed_8__15_,
  chained_data_delayed_8__14_,chained_data_delayed_8__13_,chained_data_delayed_8__12_,
  chained_data_delayed_8__11_,chained_data_delayed_8__10_,chained_data_delayed_8__9_,
  chained_data_delayed_8__8_,chained_data_delayed_8__7_,chained_data_delayed_8__6_,
  chained_data_delayed_8__5_,chained_data_delayed_8__4_,chained_data_delayed_8__3_,
  chained_data_delayed_8__2_,chained_data_delayed_8__1_,chained_data_delayed_8__0_,
  chained_data_delayed_7__63_,chained_data_delayed_7__62_,chained_data_delayed_7__61_,
  chained_data_delayed_7__60_,chained_data_delayed_7__59_,chained_data_delayed_7__58_,
  chained_data_delayed_7__57_,chained_data_delayed_7__56_,chained_data_delayed_7__55_,
  chained_data_delayed_7__54_,chained_data_delayed_7__53_,chained_data_delayed_7__52_,
  chained_data_delayed_7__51_,chained_data_delayed_7__50_,
  chained_data_delayed_7__49_,chained_data_delayed_7__48_,chained_data_delayed_7__47_,
  chained_data_delayed_7__46_,chained_data_delayed_7__45_,chained_data_delayed_7__44_,
  chained_data_delayed_7__43_,chained_data_delayed_7__42_,chained_data_delayed_7__41_,
  chained_data_delayed_7__40_,chained_data_delayed_7__39_,chained_data_delayed_7__38_,
  chained_data_delayed_7__37_,chained_data_delayed_7__36_,chained_data_delayed_7__35_,
  chained_data_delayed_7__34_,chained_data_delayed_7__33_,chained_data_delayed_7__32_,
  chained_data_delayed_7__31_,chained_data_delayed_7__30_,
  chained_data_delayed_7__29_,chained_data_delayed_7__28_,chained_data_delayed_7__27_,
  chained_data_delayed_7__26_,chained_data_delayed_7__25_,chained_data_delayed_7__24_,
  chained_data_delayed_7__23_,chained_data_delayed_7__22_,chained_data_delayed_7__21_,
  chained_data_delayed_7__20_,chained_data_delayed_7__19_,chained_data_delayed_7__18_,
  chained_data_delayed_7__17_,chained_data_delayed_7__16_,chained_data_delayed_7__15_,
  chained_data_delayed_7__14_,chained_data_delayed_7__13_,chained_data_delayed_7__12_,
  chained_data_delayed_7__11_,chained_data_delayed_7__10_,
  chained_data_delayed_7__9_,chained_data_delayed_7__8_,chained_data_delayed_7__7_,
  chained_data_delayed_7__6_,chained_data_delayed_7__5_,chained_data_delayed_7__4_,
  chained_data_delayed_7__3_,chained_data_delayed_7__2_,chained_data_delayed_7__1_,
  chained_data_delayed_7__0_,chained_data_delayed_6__63_,chained_data_delayed_6__62_,
  chained_data_delayed_6__61_,chained_data_delayed_6__60_,chained_data_delayed_6__59_,
  chained_data_delayed_6__58_,chained_data_delayed_6__57_,chained_data_delayed_6__56_,
  chained_data_delayed_6__55_,chained_data_delayed_6__54_,chained_data_delayed_6__53_,
  chained_data_delayed_6__52_,chained_data_delayed_6__51_,chained_data_delayed_6__50_,
  chained_data_delayed_6__49_,chained_data_delayed_6__48_,
  chained_data_delayed_6__47_,chained_data_delayed_6__46_,chained_data_delayed_6__45_,
  chained_data_delayed_6__44_,chained_data_delayed_6__43_,chained_data_delayed_6__42_,
  chained_data_delayed_6__41_,chained_data_delayed_6__40_,chained_data_delayed_6__39_,
  chained_data_delayed_6__38_,chained_data_delayed_6__37_,chained_data_delayed_6__36_,
  chained_data_delayed_6__35_,chained_data_delayed_6__34_,chained_data_delayed_6__33_,
  chained_data_delayed_6__32_,chained_data_delayed_6__31_,chained_data_delayed_6__30_,
  chained_data_delayed_6__29_,chained_data_delayed_6__28_,
  chained_data_delayed_6__27_,chained_data_delayed_6__26_,chained_data_delayed_6__25_,
  chained_data_delayed_6__24_,chained_data_delayed_6__23_,chained_data_delayed_6__22_,
  chained_data_delayed_6__21_,chained_data_delayed_6__20_,chained_data_delayed_6__19_,
  chained_data_delayed_6__18_,chained_data_delayed_6__17_,chained_data_delayed_6__16_,
  chained_data_delayed_6__15_,chained_data_delayed_6__14_,chained_data_delayed_6__13_,
  chained_data_delayed_6__12_,chained_data_delayed_6__11_,chained_data_delayed_6__10_,
  chained_data_delayed_6__9_,chained_data_delayed_6__8_,chained_data_delayed_6__7_,
  chained_data_delayed_6__6_,chained_data_delayed_6__5_,chained_data_delayed_6__4_,
  chained_data_delayed_6__3_,chained_data_delayed_6__2_,
  chained_data_delayed_6__1_,chained_data_delayed_6__0_,chained_data_delayed_5__63_,
  chained_data_delayed_5__62_,chained_data_delayed_5__61_,chained_data_delayed_5__60_,
  chained_data_delayed_5__59_,chained_data_delayed_5__58_,chained_data_delayed_5__57_,
  chained_data_delayed_5__56_,chained_data_delayed_5__55_,chained_data_delayed_5__54_,
  chained_data_delayed_5__53_,chained_data_delayed_5__52_,chained_data_delayed_5__51_,
  chained_data_delayed_5__50_,chained_data_delayed_5__49_,chained_data_delayed_5__48_,
  chained_data_delayed_5__47_,chained_data_delayed_5__46_,chained_data_delayed_5__45_,
  chained_data_delayed_5__44_,chained_data_delayed_5__43_,
  chained_data_delayed_5__42_,chained_data_delayed_5__41_,chained_data_delayed_5__40_,
  chained_data_delayed_5__39_,chained_data_delayed_5__38_,chained_data_delayed_5__37_,
  chained_data_delayed_5__36_,chained_data_delayed_5__35_,chained_data_delayed_5__34_,
  chained_data_delayed_5__33_,chained_data_delayed_5__32_,chained_data_delayed_5__31_,
  chained_data_delayed_5__30_,chained_data_delayed_5__29_,chained_data_delayed_5__28_,
  chained_data_delayed_5__27_,chained_data_delayed_5__26_,chained_data_delayed_5__25_,
  chained_data_delayed_5__24_,chained_data_delayed_5__23_,
  chained_data_delayed_5__22_,chained_data_delayed_5__21_,chained_data_delayed_5__20_,
  chained_data_delayed_5__19_,chained_data_delayed_5__18_,chained_data_delayed_5__17_,
  chained_data_delayed_5__16_,chained_data_delayed_5__15_,chained_data_delayed_5__14_,
  chained_data_delayed_5__13_,chained_data_delayed_5__12_,chained_data_delayed_5__11_,
  chained_data_delayed_5__10_,chained_data_delayed_5__9_,chained_data_delayed_5__8_,
  chained_data_delayed_5__7_,chained_data_delayed_5__6_,chained_data_delayed_5__5_,
  chained_data_delayed_5__4_,chained_data_delayed_5__3_,chained_data_delayed_5__2_,
  chained_data_delayed_5__1_,chained_data_delayed_5__0_,chained_data_delayed_4__63_,
  chained_data_delayed_4__62_,chained_data_delayed_4__61_,
  chained_data_delayed_4__60_,chained_data_delayed_4__59_,chained_data_delayed_4__58_,
  chained_data_delayed_4__57_,chained_data_delayed_4__56_,chained_data_delayed_4__55_,
  chained_data_delayed_4__54_,chained_data_delayed_4__53_,chained_data_delayed_4__52_,
  chained_data_delayed_4__51_,chained_data_delayed_4__50_,chained_data_delayed_4__49_,
  chained_data_delayed_4__48_,chained_data_delayed_4__47_,chained_data_delayed_4__46_,
  chained_data_delayed_4__45_,chained_data_delayed_4__44_,chained_data_delayed_4__43_,
  chained_data_delayed_4__42_,chained_data_delayed_4__41_,
  chained_data_delayed_4__40_,chained_data_delayed_4__39_,chained_data_delayed_4__38_,
  chained_data_delayed_4__37_,chained_data_delayed_4__36_,chained_data_delayed_4__35_,
  chained_data_delayed_4__34_,chained_data_delayed_4__33_,chained_data_delayed_4__32_,
  chained_data_delayed_4__31_,chained_data_delayed_4__30_,chained_data_delayed_4__29_,
  chained_data_delayed_4__28_,chained_data_delayed_4__27_,chained_data_delayed_4__26_,
  chained_data_delayed_4__25_,chained_data_delayed_4__24_,chained_data_delayed_4__23_,
  chained_data_delayed_4__22_,chained_data_delayed_4__21_,
  chained_data_delayed_4__20_,chained_data_delayed_4__19_,chained_data_delayed_4__18_,
  chained_data_delayed_4__17_,chained_data_delayed_4__16_,chained_data_delayed_4__15_,
  chained_data_delayed_4__14_,chained_data_delayed_4__13_,chained_data_delayed_4__12_,
  chained_data_delayed_4__11_,chained_data_delayed_4__10_,chained_data_delayed_4__9_,
  chained_data_delayed_4__8_,chained_data_delayed_4__7_,chained_data_delayed_4__6_,
  chained_data_delayed_4__5_,chained_data_delayed_4__4_,chained_data_delayed_4__3_,
  chained_data_delayed_4__2_,chained_data_delayed_4__1_,chained_data_delayed_4__0_,
  chained_data_delayed_3__63_,chained_data_delayed_3__62_,chained_data_delayed_3__61_,
  chained_data_delayed_3__60_,chained_data_delayed_3__59_,chained_data_delayed_3__58_,
  chained_data_delayed_3__57_,chained_data_delayed_3__56_,
  chained_data_delayed_3__55_,chained_data_delayed_3__54_,chained_data_delayed_3__53_,
  chained_data_delayed_3__52_,chained_data_delayed_3__51_,chained_data_delayed_3__50_,
  chained_data_delayed_3__49_,chained_data_delayed_3__48_,chained_data_delayed_3__47_,
  chained_data_delayed_3__46_,chained_data_delayed_3__45_,chained_data_delayed_3__44_,
  chained_data_delayed_3__43_,chained_data_delayed_3__42_,chained_data_delayed_3__41_,
  chained_data_delayed_3__40_,chained_data_delayed_3__39_,chained_data_delayed_3__38_,
  chained_data_delayed_3__37_,chained_data_delayed_3__36_,
  chained_data_delayed_3__35_,chained_data_delayed_3__34_,chained_data_delayed_3__33_,
  chained_data_delayed_3__32_,chained_data_delayed_3__31_,chained_data_delayed_3__30_,
  chained_data_delayed_3__29_,chained_data_delayed_3__28_,chained_data_delayed_3__27_,
  chained_data_delayed_3__26_,chained_data_delayed_3__25_,chained_data_delayed_3__24_,
  chained_data_delayed_3__23_,chained_data_delayed_3__22_,chained_data_delayed_3__21_,
  chained_data_delayed_3__20_,chained_data_delayed_3__19_,chained_data_delayed_3__18_,
  chained_data_delayed_3__17_,chained_data_delayed_3__16_,
  chained_data_delayed_3__15_,chained_data_delayed_3__14_,chained_data_delayed_3__13_,
  chained_data_delayed_3__12_,chained_data_delayed_3__11_,chained_data_delayed_3__10_,
  chained_data_delayed_3__9_,chained_data_delayed_3__8_,chained_data_delayed_3__7_,
  chained_data_delayed_3__6_,chained_data_delayed_3__5_,chained_data_delayed_3__4_,
  chained_data_delayed_3__3_,chained_data_delayed_3__2_,chained_data_delayed_3__1_,
  chained_data_delayed_3__0_,chained_data_delayed_2__63_,chained_data_delayed_2__62_,
  chained_data_delayed_2__61_,chained_data_delayed_2__60_,chained_data_delayed_2__59_,
  chained_data_delayed_2__58_,chained_data_delayed_2__57_,chained_data_delayed_2__56_,
  chained_data_delayed_2__55_,chained_data_delayed_2__54_,
  chained_data_delayed_2__53_,chained_data_delayed_2__52_,chained_data_delayed_2__51_,
  chained_data_delayed_2__50_,chained_data_delayed_2__49_,chained_data_delayed_2__48_,
  chained_data_delayed_2__47_,chained_data_delayed_2__46_,chained_data_delayed_2__45_,
  chained_data_delayed_2__44_,chained_data_delayed_2__43_,chained_data_delayed_2__42_,
  chained_data_delayed_2__41_,chained_data_delayed_2__40_,chained_data_delayed_2__39_,
  chained_data_delayed_2__38_,chained_data_delayed_2__37_,chained_data_delayed_2__36_,
  chained_data_delayed_2__35_,chained_data_delayed_2__34_,
  chained_data_delayed_2__33_,chained_data_delayed_2__32_,chained_data_delayed_2__31_,
  chained_data_delayed_2__30_,chained_data_delayed_2__29_,chained_data_delayed_2__28_,
  chained_data_delayed_2__27_,chained_data_delayed_2__26_,chained_data_delayed_2__25_,
  chained_data_delayed_2__24_,chained_data_delayed_2__23_,chained_data_delayed_2__22_,
  chained_data_delayed_2__21_,chained_data_delayed_2__20_,chained_data_delayed_2__19_,
  chained_data_delayed_2__18_,chained_data_delayed_2__17_,chained_data_delayed_2__16_,
  chained_data_delayed_2__15_,chained_data_delayed_2__14_,
  chained_data_delayed_2__13_,chained_data_delayed_2__12_,chained_data_delayed_2__11_,
  chained_data_delayed_2__10_,chained_data_delayed_2__9_,chained_data_delayed_2__8_,
  chained_data_delayed_2__7_,chained_data_delayed_2__6_,chained_data_delayed_2__5_,
  chained_data_delayed_2__4_,chained_data_delayed_2__3_,chained_data_delayed_2__2_,
  chained_data_delayed_2__1_,chained_data_delayed_2__0_,chained_data_delayed_1__63_,
  chained_data_delayed_1__62_,chained_data_delayed_1__61_,chained_data_delayed_1__60_,
  chained_data_delayed_1__59_,chained_data_delayed_1__58_,chained_data_delayed_1__57_,
  chained_data_delayed_1__56_,chained_data_delayed_1__55_,chained_data_delayed_1__54_,
  chained_data_delayed_1__53_,chained_data_delayed_1__52_,chained_data_delayed_1__51_,
  chained_data_delayed_1__50_,chained_data_delayed_1__49_,
  chained_data_delayed_1__48_,chained_data_delayed_1__47_,chained_data_delayed_1__46_,
  chained_data_delayed_1__45_,chained_data_delayed_1__44_,chained_data_delayed_1__43_,
  chained_data_delayed_1__42_,chained_data_delayed_1__41_,chained_data_delayed_1__40_,
  chained_data_delayed_1__39_,chained_data_delayed_1__38_,chained_data_delayed_1__37_,
  chained_data_delayed_1__36_,chained_data_delayed_1__35_,chained_data_delayed_1__34_,
  chained_data_delayed_1__33_,chained_data_delayed_1__32_,chained_data_delayed_1__31_,
  chained_data_delayed_1__30_,chained_data_delayed_1__29_,
  chained_data_delayed_1__28_,chained_data_delayed_1__27_,chained_data_delayed_1__26_,
  chained_data_delayed_1__25_,chained_data_delayed_1__24_,chained_data_delayed_1__23_,
  chained_data_delayed_1__22_,chained_data_delayed_1__21_,chained_data_delayed_1__20_,
  chained_data_delayed_1__19_,chained_data_delayed_1__18_,chained_data_delayed_1__17_,
  chained_data_delayed_1__16_,chained_data_delayed_1__15_,chained_data_delayed_1__14_,
  chained_data_delayed_1__13_,chained_data_delayed_1__12_,chained_data_delayed_1__11_,
  chained_data_delayed_1__10_,chained_data_delayed_1__9_,
  chained_data_delayed_1__8_,chained_data_delayed_1__7_,chained_data_delayed_1__6_,
  chained_data_delayed_1__5_,chained_data_delayed_1__4_,chained_data_delayed_1__3_,
  chained_data_delayed_1__2_,chained_data_delayed_1__1_,chained_data_delayed_1__0_,
  chained_data_delayed_16__63_,chained_data_delayed_16__62_,chained_data_delayed_16__61_,
  chained_data_delayed_16__60_,chained_data_delayed_16__59_,chained_data_delayed_16__58_,
  chained_data_delayed_16__57_,chained_data_delayed_16__56_,chained_data_delayed_16__55_,
  chained_data_delayed_16__54_,chained_data_delayed_16__53_,
  chained_data_delayed_16__52_,chained_data_delayed_16__51_,chained_data_delayed_16__50_,
  chained_data_delayed_16__49_,chained_data_delayed_16__48_,chained_data_delayed_16__47_,
  chained_data_delayed_16__46_,chained_data_delayed_16__45_,chained_data_delayed_16__44_,
  chained_data_delayed_16__43_,chained_data_delayed_16__42_,
  chained_data_delayed_16__41_,chained_data_delayed_16__40_,chained_data_delayed_16__39_,
  chained_data_delayed_16__38_,chained_data_delayed_16__37_,chained_data_delayed_16__36_,
  chained_data_delayed_16__35_,chained_data_delayed_16__34_,chained_data_delayed_16__33_,
  chained_data_delayed_16__32_,chained_data_delayed_16__31_,
  chained_data_delayed_16__30_,chained_data_delayed_16__29_,chained_data_delayed_16__28_,
  chained_data_delayed_16__27_,chained_data_delayed_16__26_,chained_data_delayed_16__25_,
  chained_data_delayed_16__24_,chained_data_delayed_16__23_,chained_data_delayed_16__22_,
  chained_data_delayed_16__21_,chained_data_delayed_16__20_,
  chained_data_delayed_16__19_,chained_data_delayed_16__18_,chained_data_delayed_16__17_,
  chained_data_delayed_16__16_,chained_data_delayed_16__15_,chained_data_delayed_16__14_,
  chained_data_delayed_16__13_,chained_data_delayed_16__12_,chained_data_delayed_16__11_,
  chained_data_delayed_16__10_,chained_data_delayed_16__9_,chained_data_delayed_16__8_,
  chained_data_delayed_16__7_,chained_data_delayed_16__6_,
  chained_data_delayed_16__5_,chained_data_delayed_16__4_,chained_data_delayed_16__3_,
  chained_data_delayed_16__2_,chained_data_delayed_16__1_,chained_data_delayed_16__0_,
  chained_data_delayed_15__63_,chained_data_delayed_15__62_,chained_data_delayed_15__61_,
  chained_data_delayed_15__60_,chained_data_delayed_15__59_,chained_data_delayed_15__58_,
  chained_data_delayed_15__57_,chained_data_delayed_15__56_,
  chained_data_delayed_15__55_,chained_data_delayed_15__54_,chained_data_delayed_15__53_,
  chained_data_delayed_15__52_,chained_data_delayed_15__51_,chained_data_delayed_15__50_,
  chained_data_delayed_15__49_,chained_data_delayed_15__48_,chained_data_delayed_15__47_,
  chained_data_delayed_15__46_,chained_data_delayed_15__45_,
  chained_data_delayed_15__44_,chained_data_delayed_15__43_,chained_data_delayed_15__42_,
  chained_data_delayed_15__41_,chained_data_delayed_15__40_,chained_data_delayed_15__39_,
  chained_data_delayed_15__38_,chained_data_delayed_15__37_,chained_data_delayed_15__36_,
  chained_data_delayed_15__35_,chained_data_delayed_15__34_,
  chained_data_delayed_15__33_,chained_data_delayed_15__32_,chained_data_delayed_15__31_,
  chained_data_delayed_15__30_,chained_data_delayed_15__29_,chained_data_delayed_15__28_,
  chained_data_delayed_15__27_,chained_data_delayed_15__26_,chained_data_delayed_15__25_,
  chained_data_delayed_15__24_,chained_data_delayed_15__23_,
  chained_data_delayed_15__22_,chained_data_delayed_15__21_,chained_data_delayed_15__20_,
  chained_data_delayed_15__19_,chained_data_delayed_15__18_,chained_data_delayed_15__17_,
  chained_data_delayed_15__16_,chained_data_delayed_15__15_,chained_data_delayed_15__14_,
  chained_data_delayed_15__13_,chained_data_delayed_15__12_,
  chained_data_delayed_15__11_,chained_data_delayed_15__10_,chained_data_delayed_15__9_,
  chained_data_delayed_15__8_,chained_data_delayed_15__7_,chained_data_delayed_15__6_,
  chained_data_delayed_15__5_,chained_data_delayed_15__4_,chained_data_delayed_15__3_,
  chained_data_delayed_15__2_,chained_data_delayed_15__1_,chained_data_delayed_15__0_,
  chained_data_delayed_14__63_,chained_data_delayed_14__62_,chained_data_delayed_14__61_,
  chained_data_delayed_14__60_,chained_data_delayed_14__59_,
  chained_data_delayed_14__58_,chained_data_delayed_14__57_,chained_data_delayed_14__56_,
  chained_data_delayed_14__55_,chained_data_delayed_14__54_,chained_data_delayed_14__53_,
  chained_data_delayed_14__52_,chained_data_delayed_14__51_,chained_data_delayed_14__50_,
  chained_data_delayed_14__49_,chained_data_delayed_14__48_,
  chained_data_delayed_14__47_,chained_data_delayed_14__46_,chained_data_delayed_14__45_,
  chained_data_delayed_14__44_,chained_data_delayed_14__43_,chained_data_delayed_14__42_,
  chained_data_delayed_14__41_,chained_data_delayed_14__40_,chained_data_delayed_14__39_,
  chained_data_delayed_14__38_,chained_data_delayed_14__37_,
  chained_data_delayed_14__36_,chained_data_delayed_14__35_,chained_data_delayed_14__34_,
  chained_data_delayed_14__33_,chained_data_delayed_14__32_,chained_data_delayed_14__31_,
  chained_data_delayed_14__30_,chained_data_delayed_14__29_,chained_data_delayed_14__28_,
  chained_data_delayed_14__27_,chained_data_delayed_14__26_,
  chained_data_delayed_14__25_,chained_data_delayed_14__24_,chained_data_delayed_14__23_,
  chained_data_delayed_14__22_,chained_data_delayed_14__21_,chained_data_delayed_14__20_,
  chained_data_delayed_14__19_,chained_data_delayed_14__18_,chained_data_delayed_14__17_,
  chained_data_delayed_14__16_,chained_data_delayed_14__15_,chained_data_delayed_14__14_,
  chained_data_delayed_14__13_,chained_data_delayed_14__12_,
  chained_data_delayed_14__11_,chained_data_delayed_14__10_,chained_data_delayed_14__9_,
  chained_data_delayed_14__8_,chained_data_delayed_14__7_,chained_data_delayed_14__6_,
  chained_data_delayed_14__5_,chained_data_delayed_14__4_,chained_data_delayed_14__3_,
  chained_data_delayed_14__2_,chained_data_delayed_14__1_,chained_data_delayed_14__0_,
  chained_data_delayed_13__63_,chained_data_delayed_13__62_,
  chained_data_delayed_13__61_,chained_data_delayed_13__60_,chained_data_delayed_13__59_,
  chained_data_delayed_13__58_,chained_data_delayed_13__57_,chained_data_delayed_13__56_,
  chained_data_delayed_13__55_,chained_data_delayed_13__54_,chained_data_delayed_13__53_,
  chained_data_delayed_13__52_,chained_data_delayed_13__51_,
  chained_data_delayed_13__50_,chained_data_delayed_13__49_,chained_data_delayed_13__48_,
  chained_data_delayed_13__47_,chained_data_delayed_13__46_,chained_data_delayed_13__45_,
  chained_data_delayed_13__44_,chained_data_delayed_13__43_,chained_data_delayed_13__42_,
  chained_data_delayed_13__41_,chained_data_delayed_13__40_,
  chained_data_delayed_13__39_,chained_data_delayed_13__38_,chained_data_delayed_13__37_,
  chained_data_delayed_13__36_,chained_data_delayed_13__35_,chained_data_delayed_13__34_,
  chained_data_delayed_13__33_,chained_data_delayed_13__32_,chained_data_delayed_13__31_,
  chained_data_delayed_13__30_,chained_data_delayed_13__29_,chained_data_delayed_13__28_,
  chained_data_delayed_13__27_,chained_data_delayed_13__26_,
  chained_data_delayed_13__25_,chained_data_delayed_13__24_,chained_data_delayed_13__23_,
  chained_data_delayed_13__22_,chained_data_delayed_13__21_,chained_data_delayed_13__20_,
  chained_data_delayed_13__19_,chained_data_delayed_13__18_,chained_data_delayed_13__17_,
  chained_data_delayed_13__16_,chained_data_delayed_13__15_,
  chained_data_delayed_13__14_,chained_data_delayed_13__13_,chained_data_delayed_13__12_,
  chained_data_delayed_13__11_,chained_data_delayed_13__10_,chained_data_delayed_13__9_,
  chained_data_delayed_13__8_,chained_data_delayed_13__7_,chained_data_delayed_13__6_,
  chained_data_delayed_13__5_,chained_data_delayed_13__4_,chained_data_delayed_13__3_,
  chained_data_delayed_13__2_,chained_data_delayed_13__1_,
  chained_data_delayed_13__0_,chained_data_delayed_12__63_,chained_data_delayed_12__62_,
  chained_data_delayed_12__61_,chained_data_delayed_12__60_,chained_data_delayed_12__59_,
  chained_data_delayed_12__58_,chained_data_delayed_12__57_,chained_data_delayed_12__56_,
  chained_data_delayed_12__55_,chained_data_delayed_12__54_,
  chained_data_delayed_12__53_,chained_data_delayed_12__52_,chained_data_delayed_12__51_,
  chained_data_delayed_12__50_,chained_data_delayed_12__49_,chained_data_delayed_12__48_,
  chained_data_delayed_12__47_,chained_data_delayed_12__46_,chained_data_delayed_12__45_,
  chained_data_delayed_12__44_,chained_data_delayed_12__43_,chained_data_delayed_12__42_,
  chained_data_delayed_12__41_,chained_data_delayed_12__40_,
  chained_data_delayed_12__39_,chained_data_delayed_12__38_,chained_data_delayed_12__37_,
  chained_data_delayed_12__36_,chained_data_delayed_12__35_,chained_data_delayed_12__34_,
  chained_data_delayed_12__33_,chained_data_delayed_12__32_,chained_data_delayed_12__31_,
  chained_data_delayed_12__30_,chained_data_delayed_12__29_,
  chained_data_delayed_12__28_,chained_data_delayed_12__27_,chained_data_delayed_12__26_,
  chained_data_delayed_12__25_,chained_data_delayed_12__24_,chained_data_delayed_12__23_,
  chained_data_delayed_12__22_,chained_data_delayed_12__21_,chained_data_delayed_12__20_,
  chained_data_delayed_12__19_,chained_data_delayed_12__18_,
  chained_data_delayed_12__17_,chained_data_delayed_12__16_,chained_data_delayed_12__15_,
  chained_data_delayed_12__14_,chained_data_delayed_12__13_,chained_data_delayed_12__12_,
  chained_data_delayed_12__11_,chained_data_delayed_12__10_,chained_data_delayed_12__9_,
  chained_data_delayed_12__8_,chained_data_delayed_12__7_,chained_data_delayed_12__6_,
  chained_data_delayed_12__5_,chained_data_delayed_12__4_,
  chained_data_delayed_12__3_,chained_data_delayed_12__2_,chained_data_delayed_12__1_,
  chained_data_delayed_12__0_,chained_data_delayed_11__63_,chained_data_delayed_11__62_,
  chained_data_delayed_11__61_,chained_data_delayed_11__60_,chained_data_delayed_11__59_,
  chained_data_delayed_11__58_,chained_data_delayed_11__57_,chained_data_delayed_11__56_,
  chained_data_delayed_11__55_,chained_data_delayed_11__54_,
  chained_data_delayed_11__53_,chained_data_delayed_11__52_,chained_data_delayed_11__51_,
  chained_data_delayed_11__50_,chained_data_delayed_11__49_,chained_data_delayed_11__48_,
  chained_data_delayed_11__47_,chained_data_delayed_11__46_,chained_data_delayed_11__45_,
  chained_data_delayed_11__44_,chained_data_delayed_11__43_,
  chained_data_delayed_11__42_,chained_data_delayed_11__41_,chained_data_delayed_11__40_,
  chained_data_delayed_11__39_,chained_data_delayed_11__38_,chained_data_delayed_11__37_,
  chained_data_delayed_11__36_,chained_data_delayed_11__35_,chained_data_delayed_11__34_,
  chained_data_delayed_11__33_,chained_data_delayed_11__32_,
  chained_data_delayed_11__31_,chained_data_delayed_11__30_,chained_data_delayed_11__29_,
  chained_data_delayed_11__28_,chained_data_delayed_11__27_,chained_data_delayed_11__26_,
  chained_data_delayed_11__25_,chained_data_delayed_11__24_,chained_data_delayed_11__23_,
  chained_data_delayed_11__22_,chained_data_delayed_11__21_,
  chained_data_delayed_11__20_,chained_data_delayed_11__19_,chained_data_delayed_11__18_,
  chained_data_delayed_11__17_,chained_data_delayed_11__16_,chained_data_delayed_11__15_,
  chained_data_delayed_11__14_,chained_data_delayed_11__13_,chained_data_delayed_11__12_,
  chained_data_delayed_11__11_,chained_data_delayed_11__10_,
  chained_data_delayed_11__9_,chained_data_delayed_11__8_,chained_data_delayed_11__7_,
  chained_data_delayed_11__6_,chained_data_delayed_11__5_,chained_data_delayed_11__4_,
  chained_data_delayed_11__3_,chained_data_delayed_11__2_,chained_data_delayed_11__1_,
  chained_data_delayed_11__0_,chained_data_delayed_10__63_,chained_data_delayed_10__62_,
  chained_data_delayed_10__61_,chained_data_delayed_10__60_,chained_data_delayed_10__59_,
  chained_data_delayed_10__58_,chained_data_delayed_10__57_,
  chained_data_delayed_10__56_,chained_data_delayed_10__55_,chained_data_delayed_10__54_,
  chained_data_delayed_10__53_,chained_data_delayed_10__52_,chained_data_delayed_10__51_,
  chained_data_delayed_10__50_,chained_data_delayed_10__49_,chained_data_delayed_10__48_,
  chained_data_delayed_10__47_,chained_data_delayed_10__46_,
  chained_data_delayed_10__45_,chained_data_delayed_10__44_,chained_data_delayed_10__43_,
  chained_data_delayed_10__42_,chained_data_delayed_10__41_,chained_data_delayed_10__40_,
  chained_data_delayed_10__39_,chained_data_delayed_10__38_,chained_data_delayed_10__37_,
  chained_data_delayed_10__36_,chained_data_delayed_10__35_,
  chained_data_delayed_10__34_,chained_data_delayed_10__33_,chained_data_delayed_10__32_,
  chained_data_delayed_10__31_,chained_data_delayed_10__30_,chained_data_delayed_10__29_,
  chained_data_delayed_10__28_,chained_data_delayed_10__27_,chained_data_delayed_10__26_,
  chained_data_delayed_10__25_,chained_data_delayed_10__24_,
  chained_data_delayed_10__23_,chained_data_delayed_10__22_,chained_data_delayed_10__21_,
  chained_data_delayed_10__20_,chained_data_delayed_10__19_,chained_data_delayed_10__18_,
  chained_data_delayed_10__17_,chained_data_delayed_10__16_,chained_data_delayed_10__15_,
  chained_data_delayed_10__14_,chained_data_delayed_10__13_,
  chained_data_delayed_10__12_,chained_data_delayed_10__11_,chained_data_delayed_10__10_,
  chained_data_delayed_10__9_,chained_data_delayed_10__8_,chained_data_delayed_10__7_,
  chained_data_delayed_10__6_,chained_data_delayed_10__5_,chained_data_delayed_10__4_,
  chained_data_delayed_10__3_,chained_data_delayed_10__2_,chained_data_delayed_10__1_,
  chained_data_delayed_10__0_,chained_data_delayed_9__63_,chained_data_delayed_9__62_,
  chained_data_delayed_9__61_,chained_data_delayed_9__60_,chained_data_delayed_9__59_,
  chained_data_delayed_9__58_,chained_data_delayed_9__57_,
  chained_data_delayed_9__56_,chained_data_delayed_9__55_,chained_data_delayed_9__54_,
  chained_data_delayed_9__53_,chained_data_delayed_9__52_,chained_data_delayed_9__51_,
  chained_data_delayed_9__50_,chained_data_delayed_9__49_,chained_data_delayed_9__48_,
  chained_data_delayed_9__47_,chained_data_delayed_9__46_,chained_data_delayed_9__45_,
  chained_data_delayed_9__44_,chained_data_delayed_9__43_,chained_data_delayed_9__42_,
  chained_data_delayed_9__41_,chained_data_delayed_9__40_,chained_data_delayed_9__39_,
  chained_data_delayed_9__38_,chained_data_delayed_9__37_,
  chained_data_delayed_9__36_,chained_data_delayed_9__35_,chained_data_delayed_9__34_,
  chained_data_delayed_9__33_,chained_data_delayed_9__32_,chained_data_delayed_9__31_,
  chained_data_delayed_9__30_,chained_data_delayed_9__29_,chained_data_delayed_9__28_,
  chained_data_delayed_9__27_,chained_data_delayed_9__26_,chained_data_delayed_9__25_,
  chained_data_delayed_9__24_,chained_data_delayed_9__23_,chained_data_delayed_9__22_,
  chained_data_delayed_9__21_,chained_data_delayed_9__20_,chained_data_delayed_9__19_,
  chained_data_delayed_9__18_,chained_data_delayed_9__17_,
  chained_data_delayed_9__16_,chained_data_delayed_9__15_,chained_data_delayed_9__14_,
  chained_data_delayed_9__13_,chained_data_delayed_9__12_,chained_data_delayed_9__11_,
  chained_data_delayed_9__10_,chained_data_delayed_9__9_,chained_data_delayed_9__8_,
  chained_data_delayed_9__7_,chained_data_delayed_9__6_,chained_data_delayed_9__5_,
  chained_data_delayed_9__4_,chained_data_delayed_9__3_,chained_data_delayed_9__2_,
  chained_data_delayed_9__1_,chained_data_delayed_9__0_,chained_data_delayed_24__63_,
  chained_data_delayed_24__62_,chained_data_delayed_24__61_,chained_data_delayed_24__60_,
  chained_data_delayed_24__59_,chained_data_delayed_24__58_,
  chained_data_delayed_24__57_,chained_data_delayed_24__56_,chained_data_delayed_24__55_,
  chained_data_delayed_24__54_,chained_data_delayed_24__53_,chained_data_delayed_24__52_,
  chained_data_delayed_24__51_,chained_data_delayed_24__50_,chained_data_delayed_24__49_,
  chained_data_delayed_24__48_,chained_data_delayed_24__47_,
  chained_data_delayed_24__46_,chained_data_delayed_24__45_,chained_data_delayed_24__44_,
  chained_data_delayed_24__43_,chained_data_delayed_24__42_,chained_data_delayed_24__41_,
  chained_data_delayed_24__40_,chained_data_delayed_24__39_,chained_data_delayed_24__38_,
  chained_data_delayed_24__37_,chained_data_delayed_24__36_,
  chained_data_delayed_24__35_,chained_data_delayed_24__34_,chained_data_delayed_24__33_,
  chained_data_delayed_24__32_,chained_data_delayed_24__31_,chained_data_delayed_24__30_,
  chained_data_delayed_24__29_,chained_data_delayed_24__28_,chained_data_delayed_24__27_,
  chained_data_delayed_24__26_,chained_data_delayed_24__25_,
  chained_data_delayed_24__24_,chained_data_delayed_24__23_,chained_data_delayed_24__22_,
  chained_data_delayed_24__21_,chained_data_delayed_24__20_,chained_data_delayed_24__19_,
  chained_data_delayed_24__18_,chained_data_delayed_24__17_,chained_data_delayed_24__16_,
  chained_data_delayed_24__15_,chained_data_delayed_24__14_,
  chained_data_delayed_24__13_,chained_data_delayed_24__12_,chained_data_delayed_24__11_,
  chained_data_delayed_24__10_,chained_data_delayed_24__9_,chained_data_delayed_24__8_,
  chained_data_delayed_24__7_,chained_data_delayed_24__6_,chained_data_delayed_24__5_,
  chained_data_delayed_24__4_,chained_data_delayed_24__3_,chained_data_delayed_24__2_,
  chained_data_delayed_24__1_,chained_data_delayed_24__0_,chained_data_delayed_23__63_,
  chained_data_delayed_23__62_,chained_data_delayed_23__61_,
  chained_data_delayed_23__60_,chained_data_delayed_23__59_,chained_data_delayed_23__58_,
  chained_data_delayed_23__57_,chained_data_delayed_23__56_,chained_data_delayed_23__55_,
  chained_data_delayed_23__54_,chained_data_delayed_23__53_,chained_data_delayed_23__52_,
  chained_data_delayed_23__51_,chained_data_delayed_23__50_,
  chained_data_delayed_23__49_,chained_data_delayed_23__48_,chained_data_delayed_23__47_,
  chained_data_delayed_23__46_,chained_data_delayed_23__45_,chained_data_delayed_23__44_,
  chained_data_delayed_23__43_,chained_data_delayed_23__42_,chained_data_delayed_23__41_,
  chained_data_delayed_23__40_,chained_data_delayed_23__39_,
  chained_data_delayed_23__38_,chained_data_delayed_23__37_,chained_data_delayed_23__36_,
  chained_data_delayed_23__35_,chained_data_delayed_23__34_,chained_data_delayed_23__33_,
  chained_data_delayed_23__32_,chained_data_delayed_23__31_,chained_data_delayed_23__30_,
  chained_data_delayed_23__29_,chained_data_delayed_23__28_,
  chained_data_delayed_23__27_,chained_data_delayed_23__26_,chained_data_delayed_23__25_,
  chained_data_delayed_23__24_,chained_data_delayed_23__23_,chained_data_delayed_23__22_,
  chained_data_delayed_23__21_,chained_data_delayed_23__20_,chained_data_delayed_23__19_,
  chained_data_delayed_23__18_,chained_data_delayed_23__17_,chained_data_delayed_23__16_,
  chained_data_delayed_23__15_,chained_data_delayed_23__14_,
  chained_data_delayed_23__13_,chained_data_delayed_23__12_,chained_data_delayed_23__11_,
  chained_data_delayed_23__10_,chained_data_delayed_23__9_,chained_data_delayed_23__8_,
  chained_data_delayed_23__7_,chained_data_delayed_23__6_,chained_data_delayed_23__5_,
  chained_data_delayed_23__4_,chained_data_delayed_23__3_,chained_data_delayed_23__2_,
  chained_data_delayed_23__1_,chained_data_delayed_23__0_,
  chained_data_delayed_22__63_,chained_data_delayed_22__62_,chained_data_delayed_22__61_,
  chained_data_delayed_22__60_,chained_data_delayed_22__59_,chained_data_delayed_22__58_,
  chained_data_delayed_22__57_,chained_data_delayed_22__56_,chained_data_delayed_22__55_,
  chained_data_delayed_22__54_,chained_data_delayed_22__53_,
  chained_data_delayed_22__52_,chained_data_delayed_22__51_,chained_data_delayed_22__50_,
  chained_data_delayed_22__49_,chained_data_delayed_22__48_,chained_data_delayed_22__47_,
  chained_data_delayed_22__46_,chained_data_delayed_22__45_,chained_data_delayed_22__44_,
  chained_data_delayed_22__43_,chained_data_delayed_22__42_,
  chained_data_delayed_22__41_,chained_data_delayed_22__40_,chained_data_delayed_22__39_,
  chained_data_delayed_22__38_,chained_data_delayed_22__37_,chained_data_delayed_22__36_,
  chained_data_delayed_22__35_,chained_data_delayed_22__34_,chained_data_delayed_22__33_,
  chained_data_delayed_22__32_,chained_data_delayed_22__31_,chained_data_delayed_22__30_,
  chained_data_delayed_22__29_,chained_data_delayed_22__28_,
  chained_data_delayed_22__27_,chained_data_delayed_22__26_,chained_data_delayed_22__25_,
  chained_data_delayed_22__24_,chained_data_delayed_22__23_,chained_data_delayed_22__22_,
  chained_data_delayed_22__21_,chained_data_delayed_22__20_,chained_data_delayed_22__19_,
  chained_data_delayed_22__18_,chained_data_delayed_22__17_,
  chained_data_delayed_22__16_,chained_data_delayed_22__15_,chained_data_delayed_22__14_,
  chained_data_delayed_22__13_,chained_data_delayed_22__12_,chained_data_delayed_22__11_,
  chained_data_delayed_22__10_,chained_data_delayed_22__9_,chained_data_delayed_22__8_,
  chained_data_delayed_22__7_,chained_data_delayed_22__6_,chained_data_delayed_22__5_,
  chained_data_delayed_22__4_,chained_data_delayed_22__3_,
  chained_data_delayed_22__2_,chained_data_delayed_22__1_,chained_data_delayed_22__0_,
  chained_data_delayed_21__63_,chained_data_delayed_21__62_,chained_data_delayed_21__61_,
  chained_data_delayed_21__60_,chained_data_delayed_21__59_,chained_data_delayed_21__58_,
  chained_data_delayed_21__57_,chained_data_delayed_21__56_,
  chained_data_delayed_21__55_,chained_data_delayed_21__54_,chained_data_delayed_21__53_,
  chained_data_delayed_21__52_,chained_data_delayed_21__51_,chained_data_delayed_21__50_,
  chained_data_delayed_21__49_,chained_data_delayed_21__48_,chained_data_delayed_21__47_,
  chained_data_delayed_21__46_,chained_data_delayed_21__45_,chained_data_delayed_21__44_,
  chained_data_delayed_21__43_,chained_data_delayed_21__42_,
  chained_data_delayed_21__41_,chained_data_delayed_21__40_,chained_data_delayed_21__39_,
  chained_data_delayed_21__38_,chained_data_delayed_21__37_,chained_data_delayed_21__36_,
  chained_data_delayed_21__35_,chained_data_delayed_21__34_,chained_data_delayed_21__33_,
  chained_data_delayed_21__32_,chained_data_delayed_21__31_,
  chained_data_delayed_21__30_,chained_data_delayed_21__29_,chained_data_delayed_21__28_,
  chained_data_delayed_21__27_,chained_data_delayed_21__26_,chained_data_delayed_21__25_,
  chained_data_delayed_21__24_,chained_data_delayed_21__23_,chained_data_delayed_21__22_,
  chained_data_delayed_21__21_,chained_data_delayed_21__20_,
  chained_data_delayed_21__19_,chained_data_delayed_21__18_,chained_data_delayed_21__17_,
  chained_data_delayed_21__16_,chained_data_delayed_21__15_,chained_data_delayed_21__14_,
  chained_data_delayed_21__13_,chained_data_delayed_21__12_,chained_data_delayed_21__11_,
  chained_data_delayed_21__10_,chained_data_delayed_21__9_,
  chained_data_delayed_21__8_,chained_data_delayed_21__7_,chained_data_delayed_21__6_,
  chained_data_delayed_21__5_,chained_data_delayed_21__4_,chained_data_delayed_21__3_,
  chained_data_delayed_21__2_,chained_data_delayed_21__1_,chained_data_delayed_21__0_,
  chained_data_delayed_20__63_,chained_data_delayed_20__62_,chained_data_delayed_20__61_,
  chained_data_delayed_20__60_,chained_data_delayed_20__59_,chained_data_delayed_20__58_,
  chained_data_delayed_20__57_,chained_data_delayed_20__56_,
  chained_data_delayed_20__55_,chained_data_delayed_20__54_,chained_data_delayed_20__53_,
  chained_data_delayed_20__52_,chained_data_delayed_20__51_,chained_data_delayed_20__50_,
  chained_data_delayed_20__49_,chained_data_delayed_20__48_,chained_data_delayed_20__47_,
  chained_data_delayed_20__46_,chained_data_delayed_20__45_,
  chained_data_delayed_20__44_,chained_data_delayed_20__43_,chained_data_delayed_20__42_,
  chained_data_delayed_20__41_,chained_data_delayed_20__40_,chained_data_delayed_20__39_,
  chained_data_delayed_20__38_,chained_data_delayed_20__37_,chained_data_delayed_20__36_,
  chained_data_delayed_20__35_,chained_data_delayed_20__34_,
  chained_data_delayed_20__33_,chained_data_delayed_20__32_,chained_data_delayed_20__31_,
  chained_data_delayed_20__30_,chained_data_delayed_20__29_,chained_data_delayed_20__28_,
  chained_data_delayed_20__27_,chained_data_delayed_20__26_,chained_data_delayed_20__25_,
  chained_data_delayed_20__24_,chained_data_delayed_20__23_,
  chained_data_delayed_20__22_,chained_data_delayed_20__21_,chained_data_delayed_20__20_,
  chained_data_delayed_20__19_,chained_data_delayed_20__18_,chained_data_delayed_20__17_,
  chained_data_delayed_20__16_,chained_data_delayed_20__15_,chained_data_delayed_20__14_,
  chained_data_delayed_20__13_,chained_data_delayed_20__12_,
  chained_data_delayed_20__11_,chained_data_delayed_20__10_,chained_data_delayed_20__9_,
  chained_data_delayed_20__8_,chained_data_delayed_20__7_,chained_data_delayed_20__6_,
  chained_data_delayed_20__5_,chained_data_delayed_20__4_,chained_data_delayed_20__3_,
  chained_data_delayed_20__2_,chained_data_delayed_20__1_,chained_data_delayed_20__0_,
  chained_data_delayed_19__63_,chained_data_delayed_19__62_,chained_data_delayed_19__61_,
  chained_data_delayed_19__60_,chained_data_delayed_19__59_,
  chained_data_delayed_19__58_,chained_data_delayed_19__57_,chained_data_delayed_19__56_,
  chained_data_delayed_19__55_,chained_data_delayed_19__54_,chained_data_delayed_19__53_,
  chained_data_delayed_19__52_,chained_data_delayed_19__51_,chained_data_delayed_19__50_,
  chained_data_delayed_19__49_,chained_data_delayed_19__48_,
  chained_data_delayed_19__47_,chained_data_delayed_19__46_,chained_data_delayed_19__45_,
  chained_data_delayed_19__44_,chained_data_delayed_19__43_,chained_data_delayed_19__42_,
  chained_data_delayed_19__41_,chained_data_delayed_19__40_,chained_data_delayed_19__39_,
  chained_data_delayed_19__38_,chained_data_delayed_19__37_,
  chained_data_delayed_19__36_,chained_data_delayed_19__35_,chained_data_delayed_19__34_,
  chained_data_delayed_19__33_,chained_data_delayed_19__32_,chained_data_delayed_19__31_,
  chained_data_delayed_19__30_,chained_data_delayed_19__29_,chained_data_delayed_19__28_,
  chained_data_delayed_19__27_,chained_data_delayed_19__26_,
  chained_data_delayed_19__25_,chained_data_delayed_19__24_,chained_data_delayed_19__23_,
  chained_data_delayed_19__22_,chained_data_delayed_19__21_,chained_data_delayed_19__20_,
  chained_data_delayed_19__19_,chained_data_delayed_19__18_,chained_data_delayed_19__17_,
  chained_data_delayed_19__16_,chained_data_delayed_19__15_,
  chained_data_delayed_19__14_,chained_data_delayed_19__13_,chained_data_delayed_19__12_,
  chained_data_delayed_19__11_,chained_data_delayed_19__10_,chained_data_delayed_19__9_,
  chained_data_delayed_19__8_,chained_data_delayed_19__7_,chained_data_delayed_19__6_,
  chained_data_delayed_19__5_,chained_data_delayed_19__4_,chained_data_delayed_19__3_,
  chained_data_delayed_19__2_,chained_data_delayed_19__1_,chained_data_delayed_19__0_,
  chained_data_delayed_18__63_,chained_data_delayed_18__62_,
  chained_data_delayed_18__61_,chained_data_delayed_18__60_,chained_data_delayed_18__59_,
  chained_data_delayed_18__58_,chained_data_delayed_18__57_,chained_data_delayed_18__56_,
  chained_data_delayed_18__55_,chained_data_delayed_18__54_,chained_data_delayed_18__53_,
  chained_data_delayed_18__52_,chained_data_delayed_18__51_,
  chained_data_delayed_18__50_,chained_data_delayed_18__49_,chained_data_delayed_18__48_,
  chained_data_delayed_18__47_,chained_data_delayed_18__46_,chained_data_delayed_18__45_,
  chained_data_delayed_18__44_,chained_data_delayed_18__43_,chained_data_delayed_18__42_,
  chained_data_delayed_18__41_,chained_data_delayed_18__40_,
  chained_data_delayed_18__39_,chained_data_delayed_18__38_,chained_data_delayed_18__37_,
  chained_data_delayed_18__36_,chained_data_delayed_18__35_,chained_data_delayed_18__34_,
  chained_data_delayed_18__33_,chained_data_delayed_18__32_,chained_data_delayed_18__31_,
  chained_data_delayed_18__30_,chained_data_delayed_18__29_,
  chained_data_delayed_18__28_,chained_data_delayed_18__27_,chained_data_delayed_18__26_,
  chained_data_delayed_18__25_,chained_data_delayed_18__24_,chained_data_delayed_18__23_,
  chained_data_delayed_18__22_,chained_data_delayed_18__21_,chained_data_delayed_18__20_,
  chained_data_delayed_18__19_,chained_data_delayed_18__18_,
  chained_data_delayed_18__17_,chained_data_delayed_18__16_,chained_data_delayed_18__15_,
  chained_data_delayed_18__14_,chained_data_delayed_18__13_,chained_data_delayed_18__12_,
  chained_data_delayed_18__11_,chained_data_delayed_18__10_,chained_data_delayed_18__9_,
  chained_data_delayed_18__8_,chained_data_delayed_18__7_,chained_data_delayed_18__6_,
  chained_data_delayed_18__5_,chained_data_delayed_18__4_,chained_data_delayed_18__3_,
  chained_data_delayed_18__2_,chained_data_delayed_18__1_,
  chained_data_delayed_18__0_,chained_data_delayed_17__63_,chained_data_delayed_17__62_,
  chained_data_delayed_17__61_,chained_data_delayed_17__60_,chained_data_delayed_17__59_,
  chained_data_delayed_17__58_,chained_data_delayed_17__57_,chained_data_delayed_17__56_,
  chained_data_delayed_17__55_,chained_data_delayed_17__54_,
  chained_data_delayed_17__53_,chained_data_delayed_17__52_,chained_data_delayed_17__51_,
  chained_data_delayed_17__50_,chained_data_delayed_17__49_,chained_data_delayed_17__48_,
  chained_data_delayed_17__47_,chained_data_delayed_17__46_,chained_data_delayed_17__45_,
  chained_data_delayed_17__44_,chained_data_delayed_17__43_,
  chained_data_delayed_17__42_,chained_data_delayed_17__41_,chained_data_delayed_17__40_,
  chained_data_delayed_17__39_,chained_data_delayed_17__38_,chained_data_delayed_17__37_,
  chained_data_delayed_17__36_,chained_data_delayed_17__35_,chained_data_delayed_17__34_,
  chained_data_delayed_17__33_,chained_data_delayed_17__32_,
  chained_data_delayed_17__31_,chained_data_delayed_17__30_,chained_data_delayed_17__29_,
  chained_data_delayed_17__28_,chained_data_delayed_17__27_,chained_data_delayed_17__26_,
  chained_data_delayed_17__25_,chained_data_delayed_17__24_,chained_data_delayed_17__23_,
  chained_data_delayed_17__22_,chained_data_delayed_17__21_,chained_data_delayed_17__20_,
  chained_data_delayed_17__19_,chained_data_delayed_17__18_,
  chained_data_delayed_17__17_,chained_data_delayed_17__16_,chained_data_delayed_17__15_,
  chained_data_delayed_17__14_,chained_data_delayed_17__13_,chained_data_delayed_17__12_,
  chained_data_delayed_17__11_,chained_data_delayed_17__10_,chained_data_delayed_17__9_,
  chained_data_delayed_17__8_,chained_data_delayed_17__7_,
  chained_data_delayed_17__6_,chained_data_delayed_17__5_,chained_data_delayed_17__4_,
  chained_data_delayed_17__3_,chained_data_delayed_17__2_,chained_data_delayed_17__1_,
  chained_data_delayed_17__0_,chained_data_delayed_32__63_,chained_data_delayed_32__62_,
  chained_data_delayed_32__61_,chained_data_delayed_32__60_,chained_data_delayed_32__59_,
  chained_data_delayed_32__58_,chained_data_delayed_32__57_,
  chained_data_delayed_32__56_,chained_data_delayed_32__55_,chained_data_delayed_32__54_,
  chained_data_delayed_32__53_,chained_data_delayed_32__52_,chained_data_delayed_32__51_,
  chained_data_delayed_32__50_,chained_data_delayed_32__49_,chained_data_delayed_32__48_,
  chained_data_delayed_32__47_,chained_data_delayed_32__46_,
  chained_data_delayed_32__45_,chained_data_delayed_32__44_,chained_data_delayed_32__43_,
  chained_data_delayed_32__42_,chained_data_delayed_32__41_,chained_data_delayed_32__40_,
  chained_data_delayed_32__39_,chained_data_delayed_32__38_,chained_data_delayed_32__37_,
  chained_data_delayed_32__36_,chained_data_delayed_32__35_,chained_data_delayed_32__34_,
  chained_data_delayed_32__33_,chained_data_delayed_32__32_,
  chained_data_delayed_32__31_,chained_data_delayed_32__30_,chained_data_delayed_32__29_,
  chained_data_delayed_32__28_,chained_data_delayed_32__27_,chained_data_delayed_32__26_,
  chained_data_delayed_32__25_,chained_data_delayed_32__24_,chained_data_delayed_32__23_,
  chained_data_delayed_32__22_,chained_data_delayed_32__21_,
  chained_data_delayed_32__20_,chained_data_delayed_32__19_,chained_data_delayed_32__18_,
  chained_data_delayed_32__17_,chained_data_delayed_32__16_,chained_data_delayed_32__15_,
  chained_data_delayed_32__14_,chained_data_delayed_32__13_,chained_data_delayed_32__12_,
  chained_data_delayed_32__11_,chained_data_delayed_32__10_,
  chained_data_delayed_32__9_,chained_data_delayed_32__8_,chained_data_delayed_32__7_,
  chained_data_delayed_32__6_,chained_data_delayed_32__5_,chained_data_delayed_32__4_,
  chained_data_delayed_32__3_,chained_data_delayed_32__2_,chained_data_delayed_32__1_,
  chained_data_delayed_32__0_,chained_data_delayed_31__63_,chained_data_delayed_31__62_,
  chained_data_delayed_31__61_,chained_data_delayed_31__60_,
  chained_data_delayed_31__59_,chained_data_delayed_31__58_,chained_data_delayed_31__57_,
  chained_data_delayed_31__56_,chained_data_delayed_31__55_,chained_data_delayed_31__54_,
  chained_data_delayed_31__53_,chained_data_delayed_31__52_,chained_data_delayed_31__51_,
  chained_data_delayed_31__50_,chained_data_delayed_31__49_,chained_data_delayed_31__48_,
  chained_data_delayed_31__47_,chained_data_delayed_31__46_,
  chained_data_delayed_31__45_,chained_data_delayed_31__44_,chained_data_delayed_31__43_,
  chained_data_delayed_31__42_,chained_data_delayed_31__41_,chained_data_delayed_31__40_,
  chained_data_delayed_31__39_,chained_data_delayed_31__38_,chained_data_delayed_31__37_,
  chained_data_delayed_31__36_,chained_data_delayed_31__35_,
  chained_data_delayed_31__34_,chained_data_delayed_31__33_,chained_data_delayed_31__32_,
  chained_data_delayed_31__31_,chained_data_delayed_31__30_,chained_data_delayed_31__29_,
  chained_data_delayed_31__28_,chained_data_delayed_31__27_,chained_data_delayed_31__26_,
  chained_data_delayed_31__25_,chained_data_delayed_31__24_,
  chained_data_delayed_31__23_,chained_data_delayed_31__22_,chained_data_delayed_31__21_,
  chained_data_delayed_31__20_,chained_data_delayed_31__19_,chained_data_delayed_31__18_,
  chained_data_delayed_31__17_,chained_data_delayed_31__16_,chained_data_delayed_31__15_,
  chained_data_delayed_31__14_,chained_data_delayed_31__13_,
  chained_data_delayed_31__12_,chained_data_delayed_31__11_,chained_data_delayed_31__10_,
  chained_data_delayed_31__9_,chained_data_delayed_31__8_,chained_data_delayed_31__7_,
  chained_data_delayed_31__6_,chained_data_delayed_31__5_,chained_data_delayed_31__4_,
  chained_data_delayed_31__3_,chained_data_delayed_31__2_,chained_data_delayed_31__1_,
  chained_data_delayed_31__0_,chained_data_delayed_30__63_,chained_data_delayed_30__62_,
  chained_data_delayed_30__61_,chained_data_delayed_30__60_,
  chained_data_delayed_30__59_,chained_data_delayed_30__58_,chained_data_delayed_30__57_,
  chained_data_delayed_30__56_,chained_data_delayed_30__55_,chained_data_delayed_30__54_,
  chained_data_delayed_30__53_,chained_data_delayed_30__52_,chained_data_delayed_30__51_,
  chained_data_delayed_30__50_,chained_data_delayed_30__49_,
  chained_data_delayed_30__48_,chained_data_delayed_30__47_,chained_data_delayed_30__46_,
  chained_data_delayed_30__45_,chained_data_delayed_30__44_,chained_data_delayed_30__43_,
  chained_data_delayed_30__42_,chained_data_delayed_30__41_,chained_data_delayed_30__40_,
  chained_data_delayed_30__39_,chained_data_delayed_30__38_,
  chained_data_delayed_30__37_,chained_data_delayed_30__36_,chained_data_delayed_30__35_,
  chained_data_delayed_30__34_,chained_data_delayed_30__33_,chained_data_delayed_30__32_,
  chained_data_delayed_30__31_,chained_data_delayed_30__30_,chained_data_delayed_30__29_,
  chained_data_delayed_30__28_,chained_data_delayed_30__27_,
  chained_data_delayed_30__26_,chained_data_delayed_30__25_,chained_data_delayed_30__24_,
  chained_data_delayed_30__23_,chained_data_delayed_30__22_,chained_data_delayed_30__21_,
  chained_data_delayed_30__20_,chained_data_delayed_30__19_,chained_data_delayed_30__18_,
  chained_data_delayed_30__17_,chained_data_delayed_30__16_,
  chained_data_delayed_30__15_,chained_data_delayed_30__14_,chained_data_delayed_30__13_,
  chained_data_delayed_30__12_,chained_data_delayed_30__11_,chained_data_delayed_30__10_,
  chained_data_delayed_30__9_,chained_data_delayed_30__8_,chained_data_delayed_30__7_,
  chained_data_delayed_30__6_,chained_data_delayed_30__5_,chained_data_delayed_30__4_,
  chained_data_delayed_30__3_,chained_data_delayed_30__2_,chained_data_delayed_30__1_,
  chained_data_delayed_30__0_,chained_data_delayed_29__63_,
  chained_data_delayed_29__62_,chained_data_delayed_29__61_,chained_data_delayed_29__60_,
  chained_data_delayed_29__59_,chained_data_delayed_29__58_,chained_data_delayed_29__57_,
  chained_data_delayed_29__56_,chained_data_delayed_29__55_,chained_data_delayed_29__54_,
  chained_data_delayed_29__53_,chained_data_delayed_29__52_,
  chained_data_delayed_29__51_,chained_data_delayed_29__50_,chained_data_delayed_29__49_,
  chained_data_delayed_29__48_,chained_data_delayed_29__47_,chained_data_delayed_29__46_,
  chained_data_delayed_29__45_,chained_data_delayed_29__44_,chained_data_delayed_29__43_,
  chained_data_delayed_29__42_,chained_data_delayed_29__41_,
  chained_data_delayed_29__40_,chained_data_delayed_29__39_,chained_data_delayed_29__38_,
  chained_data_delayed_29__37_,chained_data_delayed_29__36_,chained_data_delayed_29__35_,
  chained_data_delayed_29__34_,chained_data_delayed_29__33_,chained_data_delayed_29__32_,
  chained_data_delayed_29__31_,chained_data_delayed_29__30_,
  chained_data_delayed_29__29_,chained_data_delayed_29__28_,chained_data_delayed_29__27_,
  chained_data_delayed_29__26_,chained_data_delayed_29__25_,chained_data_delayed_29__24_,
  chained_data_delayed_29__23_,chained_data_delayed_29__22_,chained_data_delayed_29__21_,
  chained_data_delayed_29__20_,chained_data_delayed_29__19_,
  chained_data_delayed_29__18_,chained_data_delayed_29__17_,chained_data_delayed_29__16_,
  chained_data_delayed_29__15_,chained_data_delayed_29__14_,chained_data_delayed_29__13_,
  chained_data_delayed_29__12_,chained_data_delayed_29__11_,chained_data_delayed_29__10_,
  chained_data_delayed_29__9_,chained_data_delayed_29__8_,chained_data_delayed_29__7_,
  chained_data_delayed_29__6_,chained_data_delayed_29__5_,
  chained_data_delayed_29__4_,chained_data_delayed_29__3_,chained_data_delayed_29__2_,
  chained_data_delayed_29__1_,chained_data_delayed_29__0_,chained_data_delayed_28__63_,
  chained_data_delayed_28__62_,chained_data_delayed_28__61_,chained_data_delayed_28__60_,
  chained_data_delayed_28__59_,chained_data_delayed_28__58_,chained_data_delayed_28__57_,
  chained_data_delayed_28__56_,chained_data_delayed_28__55_,
  chained_data_delayed_28__54_,chained_data_delayed_28__53_,chained_data_delayed_28__52_,
  chained_data_delayed_28__51_,chained_data_delayed_28__50_,chained_data_delayed_28__49_,
  chained_data_delayed_28__48_,chained_data_delayed_28__47_,chained_data_delayed_28__46_,
  chained_data_delayed_28__45_,chained_data_delayed_28__44_,
  chained_data_delayed_28__43_,chained_data_delayed_28__42_,chained_data_delayed_28__41_,
  chained_data_delayed_28__40_,chained_data_delayed_28__39_,chained_data_delayed_28__38_,
  chained_data_delayed_28__37_,chained_data_delayed_28__36_,chained_data_delayed_28__35_,
  chained_data_delayed_28__34_,chained_data_delayed_28__33_,
  chained_data_delayed_28__32_,chained_data_delayed_28__31_,chained_data_delayed_28__30_,
  chained_data_delayed_28__29_,chained_data_delayed_28__28_,chained_data_delayed_28__27_,
  chained_data_delayed_28__26_,chained_data_delayed_28__25_,chained_data_delayed_28__24_,
  chained_data_delayed_28__23_,chained_data_delayed_28__22_,
  chained_data_delayed_28__21_,chained_data_delayed_28__20_,chained_data_delayed_28__19_,
  chained_data_delayed_28__18_,chained_data_delayed_28__17_,chained_data_delayed_28__16_,
  chained_data_delayed_28__15_,chained_data_delayed_28__14_,chained_data_delayed_28__13_,
  chained_data_delayed_28__12_,chained_data_delayed_28__11_,chained_data_delayed_28__10_,
  chained_data_delayed_28__9_,chained_data_delayed_28__8_,
  chained_data_delayed_28__7_,chained_data_delayed_28__6_,chained_data_delayed_28__5_,
  chained_data_delayed_28__4_,chained_data_delayed_28__3_,chained_data_delayed_28__2_,
  chained_data_delayed_28__1_,chained_data_delayed_28__0_,chained_data_delayed_27__63_,
  chained_data_delayed_27__62_,chained_data_delayed_27__61_,chained_data_delayed_27__60_,
  chained_data_delayed_27__59_,chained_data_delayed_27__58_,
  chained_data_delayed_27__57_,chained_data_delayed_27__56_,chained_data_delayed_27__55_,
  chained_data_delayed_27__54_,chained_data_delayed_27__53_,chained_data_delayed_27__52_,
  chained_data_delayed_27__51_,chained_data_delayed_27__50_,chained_data_delayed_27__49_,
  chained_data_delayed_27__48_,chained_data_delayed_27__47_,
  chained_data_delayed_27__46_,chained_data_delayed_27__45_,chained_data_delayed_27__44_,
  chained_data_delayed_27__43_,chained_data_delayed_27__42_,chained_data_delayed_27__41_,
  chained_data_delayed_27__40_,chained_data_delayed_27__39_,chained_data_delayed_27__38_,
  chained_data_delayed_27__37_,chained_data_delayed_27__36_,
  chained_data_delayed_27__35_,chained_data_delayed_27__34_,chained_data_delayed_27__33_,
  chained_data_delayed_27__32_,chained_data_delayed_27__31_,chained_data_delayed_27__30_,
  chained_data_delayed_27__29_,chained_data_delayed_27__28_,chained_data_delayed_27__27_,
  chained_data_delayed_27__26_,chained_data_delayed_27__25_,chained_data_delayed_27__24_,
  chained_data_delayed_27__23_,chained_data_delayed_27__22_,
  chained_data_delayed_27__21_,chained_data_delayed_27__20_,chained_data_delayed_27__19_,
  chained_data_delayed_27__18_,chained_data_delayed_27__17_,chained_data_delayed_27__16_,
  chained_data_delayed_27__15_,chained_data_delayed_27__14_,chained_data_delayed_27__13_,
  chained_data_delayed_27__12_,chained_data_delayed_27__11_,
  chained_data_delayed_27__10_,chained_data_delayed_27__9_,chained_data_delayed_27__8_,
  chained_data_delayed_27__7_,chained_data_delayed_27__6_,chained_data_delayed_27__5_,
  chained_data_delayed_27__4_,chained_data_delayed_27__3_,chained_data_delayed_27__2_,
  chained_data_delayed_27__1_,chained_data_delayed_27__0_,chained_data_delayed_26__63_,
  chained_data_delayed_26__62_,chained_data_delayed_26__61_,
  chained_data_delayed_26__60_,chained_data_delayed_26__59_,chained_data_delayed_26__58_,
  chained_data_delayed_26__57_,chained_data_delayed_26__56_,chained_data_delayed_26__55_,
  chained_data_delayed_26__54_,chained_data_delayed_26__53_,chained_data_delayed_26__52_,
  chained_data_delayed_26__51_,chained_data_delayed_26__50_,
  chained_data_delayed_26__49_,chained_data_delayed_26__48_,chained_data_delayed_26__47_,
  chained_data_delayed_26__46_,chained_data_delayed_26__45_,chained_data_delayed_26__44_,
  chained_data_delayed_26__43_,chained_data_delayed_26__42_,chained_data_delayed_26__41_,
  chained_data_delayed_26__40_,chained_data_delayed_26__39_,chained_data_delayed_26__38_,
  chained_data_delayed_26__37_,chained_data_delayed_26__36_,
  chained_data_delayed_26__35_,chained_data_delayed_26__34_,chained_data_delayed_26__33_,
  chained_data_delayed_26__32_,chained_data_delayed_26__31_,chained_data_delayed_26__30_,
  chained_data_delayed_26__29_,chained_data_delayed_26__28_,chained_data_delayed_26__27_,
  chained_data_delayed_26__26_,chained_data_delayed_26__25_,
  chained_data_delayed_26__24_,chained_data_delayed_26__23_,chained_data_delayed_26__22_,
  chained_data_delayed_26__21_,chained_data_delayed_26__20_,chained_data_delayed_26__19_,
  chained_data_delayed_26__18_,chained_data_delayed_26__17_,chained_data_delayed_26__16_,
  chained_data_delayed_26__15_,chained_data_delayed_26__14_,
  chained_data_delayed_26__13_,chained_data_delayed_26__12_,chained_data_delayed_26__11_,
  chained_data_delayed_26__10_,chained_data_delayed_26__9_,chained_data_delayed_26__8_,
  chained_data_delayed_26__7_,chained_data_delayed_26__6_,chained_data_delayed_26__5_,
  chained_data_delayed_26__4_,chained_data_delayed_26__3_,chained_data_delayed_26__2_,
  chained_data_delayed_26__1_,chained_data_delayed_26__0_,
  chained_data_delayed_25__63_,chained_data_delayed_25__62_,chained_data_delayed_25__61_,
  chained_data_delayed_25__60_,chained_data_delayed_25__59_,chained_data_delayed_25__58_,
  chained_data_delayed_25__57_,chained_data_delayed_25__56_,chained_data_delayed_25__55_,
  chained_data_delayed_25__54_,chained_data_delayed_25__53_,chained_data_delayed_25__52_,
  chained_data_delayed_25__51_,chained_data_delayed_25__50_,
  chained_data_delayed_25__49_,chained_data_delayed_25__48_,chained_data_delayed_25__47_,
  chained_data_delayed_25__46_,chained_data_delayed_25__45_,chained_data_delayed_25__44_,
  chained_data_delayed_25__43_,chained_data_delayed_25__42_,chained_data_delayed_25__41_,
  chained_data_delayed_25__40_,chained_data_delayed_25__39_,
  chained_data_delayed_25__38_,chained_data_delayed_25__37_,chained_data_delayed_25__36_,
  chained_data_delayed_25__35_,chained_data_delayed_25__34_,chained_data_delayed_25__33_,
  chained_data_delayed_25__32_,chained_data_delayed_25__31_,chained_data_delayed_25__30_,
  chained_data_delayed_25__29_,chained_data_delayed_25__28_,
  chained_data_delayed_25__27_,chained_data_delayed_25__26_,chained_data_delayed_25__25_,
  chained_data_delayed_25__24_,chained_data_delayed_25__23_,chained_data_delayed_25__22_,
  chained_data_delayed_25__21_,chained_data_delayed_25__20_,chained_data_delayed_25__19_,
  chained_data_delayed_25__18_,chained_data_delayed_25__17_,
  chained_data_delayed_25__16_,chained_data_delayed_25__15_,chained_data_delayed_25__14_,
  chained_data_delayed_25__13_,chained_data_delayed_25__12_,chained_data_delayed_25__11_,
  chained_data_delayed_25__10_,chained_data_delayed_25__9_,chained_data_delayed_25__8_,
  chained_data_delayed_25__7_,chained_data_delayed_25__6_,chained_data_delayed_25__5_,
  chained_data_delayed_25__4_,chained_data_delayed_25__3_,
  chained_data_delayed_25__2_,chained_data_delayed_25__1_,chained_data_delayed_25__0_,
  chained_data_delayed_40__63_,chained_data_delayed_40__62_,chained_data_delayed_40__61_,
  chained_data_delayed_40__60_,chained_data_delayed_40__59_,chained_data_delayed_40__58_,
  chained_data_delayed_40__57_,chained_data_delayed_40__56_,chained_data_delayed_40__55_,
  chained_data_delayed_40__54_,chained_data_delayed_40__53_,
  chained_data_delayed_40__52_,chained_data_delayed_40__51_,chained_data_delayed_40__50_,
  chained_data_delayed_40__49_,chained_data_delayed_40__48_,chained_data_delayed_40__47_,
  chained_data_delayed_40__46_,chained_data_delayed_40__45_,chained_data_delayed_40__44_,
  chained_data_delayed_40__43_,chained_data_delayed_40__42_,
  chained_data_delayed_40__41_,chained_data_delayed_40__40_,chained_data_delayed_40__39_,
  chained_data_delayed_40__38_,chained_data_delayed_40__37_,chained_data_delayed_40__36_,
  chained_data_delayed_40__35_,chained_data_delayed_40__34_,chained_data_delayed_40__33_,
  chained_data_delayed_40__32_,chained_data_delayed_40__31_,
  chained_data_delayed_40__30_,chained_data_delayed_40__29_,chained_data_delayed_40__28_,
  chained_data_delayed_40__27_,chained_data_delayed_40__26_,chained_data_delayed_40__25_,
  chained_data_delayed_40__24_,chained_data_delayed_40__23_,chained_data_delayed_40__22_,
  chained_data_delayed_40__21_,chained_data_delayed_40__20_,
  chained_data_delayed_40__19_,chained_data_delayed_40__18_,chained_data_delayed_40__17_,
  chained_data_delayed_40__16_,chained_data_delayed_40__15_,chained_data_delayed_40__14_,
  chained_data_delayed_40__13_,chained_data_delayed_40__12_,chained_data_delayed_40__11_,
  chained_data_delayed_40__10_,chained_data_delayed_40__9_,chained_data_delayed_40__8_,
  chained_data_delayed_40__7_,chained_data_delayed_40__6_,
  chained_data_delayed_40__5_,chained_data_delayed_40__4_,chained_data_delayed_40__3_,
  chained_data_delayed_40__2_,chained_data_delayed_40__1_,chained_data_delayed_40__0_,
  chained_data_delayed_39__63_,chained_data_delayed_39__62_,chained_data_delayed_39__61_,
  chained_data_delayed_39__60_,chained_data_delayed_39__59_,chained_data_delayed_39__58_,
  chained_data_delayed_39__57_,chained_data_delayed_39__56_,
  chained_data_delayed_39__55_,chained_data_delayed_39__54_,chained_data_delayed_39__53_,
  chained_data_delayed_39__52_,chained_data_delayed_39__51_,chained_data_delayed_39__50_,
  chained_data_delayed_39__49_,chained_data_delayed_39__48_,chained_data_delayed_39__47_,
  chained_data_delayed_39__46_,chained_data_delayed_39__45_,
  chained_data_delayed_39__44_,chained_data_delayed_39__43_,chained_data_delayed_39__42_,
  chained_data_delayed_39__41_,chained_data_delayed_39__40_,chained_data_delayed_39__39_,
  chained_data_delayed_39__38_,chained_data_delayed_39__37_,chained_data_delayed_39__36_,
  chained_data_delayed_39__35_,chained_data_delayed_39__34_,
  chained_data_delayed_39__33_,chained_data_delayed_39__32_,chained_data_delayed_39__31_,
  chained_data_delayed_39__30_,chained_data_delayed_39__29_,chained_data_delayed_39__28_,
  chained_data_delayed_39__27_,chained_data_delayed_39__26_,chained_data_delayed_39__25_,
  chained_data_delayed_39__24_,chained_data_delayed_39__23_,
  chained_data_delayed_39__22_,chained_data_delayed_39__21_,chained_data_delayed_39__20_,
  chained_data_delayed_39__19_,chained_data_delayed_39__18_,chained_data_delayed_39__17_,
  chained_data_delayed_39__16_,chained_data_delayed_39__15_,chained_data_delayed_39__14_,
  chained_data_delayed_39__13_,chained_data_delayed_39__12_,
  chained_data_delayed_39__11_,chained_data_delayed_39__10_,chained_data_delayed_39__9_,
  chained_data_delayed_39__8_,chained_data_delayed_39__7_,chained_data_delayed_39__6_,
  chained_data_delayed_39__5_,chained_data_delayed_39__4_,chained_data_delayed_39__3_,
  chained_data_delayed_39__2_,chained_data_delayed_39__1_,chained_data_delayed_39__0_,
  chained_data_delayed_38__63_,chained_data_delayed_38__62_,chained_data_delayed_38__61_,
  chained_data_delayed_38__60_,chained_data_delayed_38__59_,
  chained_data_delayed_38__58_,chained_data_delayed_38__57_,chained_data_delayed_38__56_,
  chained_data_delayed_38__55_,chained_data_delayed_38__54_,chained_data_delayed_38__53_,
  chained_data_delayed_38__52_,chained_data_delayed_38__51_,chained_data_delayed_38__50_,
  chained_data_delayed_38__49_,chained_data_delayed_38__48_,
  chained_data_delayed_38__47_,chained_data_delayed_38__46_,chained_data_delayed_38__45_,
  chained_data_delayed_38__44_,chained_data_delayed_38__43_,chained_data_delayed_38__42_,
  chained_data_delayed_38__41_,chained_data_delayed_38__40_,chained_data_delayed_38__39_,
  chained_data_delayed_38__38_,chained_data_delayed_38__37_,
  chained_data_delayed_38__36_,chained_data_delayed_38__35_,chained_data_delayed_38__34_,
  chained_data_delayed_38__33_,chained_data_delayed_38__32_,chained_data_delayed_38__31_,
  chained_data_delayed_38__30_,chained_data_delayed_38__29_,chained_data_delayed_38__28_,
  chained_data_delayed_38__27_,chained_data_delayed_38__26_,
  chained_data_delayed_38__25_,chained_data_delayed_38__24_,chained_data_delayed_38__23_,
  chained_data_delayed_38__22_,chained_data_delayed_38__21_,chained_data_delayed_38__20_,
  chained_data_delayed_38__19_,chained_data_delayed_38__18_,chained_data_delayed_38__17_,
  chained_data_delayed_38__16_,chained_data_delayed_38__15_,chained_data_delayed_38__14_,
  chained_data_delayed_38__13_,chained_data_delayed_38__12_,
  chained_data_delayed_38__11_,chained_data_delayed_38__10_,chained_data_delayed_38__9_,
  chained_data_delayed_38__8_,chained_data_delayed_38__7_,chained_data_delayed_38__6_,
  chained_data_delayed_38__5_,chained_data_delayed_38__4_,chained_data_delayed_38__3_,
  chained_data_delayed_38__2_,chained_data_delayed_38__1_,chained_data_delayed_38__0_,
  chained_data_delayed_37__63_,chained_data_delayed_37__62_,
  chained_data_delayed_37__61_,chained_data_delayed_37__60_,chained_data_delayed_37__59_,
  chained_data_delayed_37__58_,chained_data_delayed_37__57_,chained_data_delayed_37__56_,
  chained_data_delayed_37__55_,chained_data_delayed_37__54_,chained_data_delayed_37__53_,
  chained_data_delayed_37__52_,chained_data_delayed_37__51_,
  chained_data_delayed_37__50_,chained_data_delayed_37__49_,chained_data_delayed_37__48_,
  chained_data_delayed_37__47_,chained_data_delayed_37__46_,chained_data_delayed_37__45_,
  chained_data_delayed_37__44_,chained_data_delayed_37__43_,chained_data_delayed_37__42_,
  chained_data_delayed_37__41_,chained_data_delayed_37__40_,
  chained_data_delayed_37__39_,chained_data_delayed_37__38_,chained_data_delayed_37__37_,
  chained_data_delayed_37__36_,chained_data_delayed_37__35_,chained_data_delayed_37__34_,
  chained_data_delayed_37__33_,chained_data_delayed_37__32_,chained_data_delayed_37__31_,
  chained_data_delayed_37__30_,chained_data_delayed_37__29_,chained_data_delayed_37__28_,
  chained_data_delayed_37__27_,chained_data_delayed_37__26_,
  chained_data_delayed_37__25_,chained_data_delayed_37__24_,chained_data_delayed_37__23_,
  chained_data_delayed_37__22_,chained_data_delayed_37__21_,chained_data_delayed_37__20_,
  chained_data_delayed_37__19_,chained_data_delayed_37__18_,chained_data_delayed_37__17_,
  chained_data_delayed_37__16_,chained_data_delayed_37__15_,
  chained_data_delayed_37__14_,chained_data_delayed_37__13_,chained_data_delayed_37__12_,
  chained_data_delayed_37__11_,chained_data_delayed_37__10_,chained_data_delayed_37__9_,
  chained_data_delayed_37__8_,chained_data_delayed_37__7_,chained_data_delayed_37__6_,
  chained_data_delayed_37__5_,chained_data_delayed_37__4_,chained_data_delayed_37__3_,
  chained_data_delayed_37__2_,chained_data_delayed_37__1_,
  chained_data_delayed_37__0_,chained_data_delayed_36__63_,chained_data_delayed_36__62_,
  chained_data_delayed_36__61_,chained_data_delayed_36__60_,chained_data_delayed_36__59_,
  chained_data_delayed_36__58_,chained_data_delayed_36__57_,chained_data_delayed_36__56_,
  chained_data_delayed_36__55_,chained_data_delayed_36__54_,
  chained_data_delayed_36__53_,chained_data_delayed_36__52_,chained_data_delayed_36__51_,
  chained_data_delayed_36__50_,chained_data_delayed_36__49_,chained_data_delayed_36__48_,
  chained_data_delayed_36__47_,chained_data_delayed_36__46_,chained_data_delayed_36__45_,
  chained_data_delayed_36__44_,chained_data_delayed_36__43_,chained_data_delayed_36__42_,
  chained_data_delayed_36__41_,chained_data_delayed_36__40_,
  chained_data_delayed_36__39_,chained_data_delayed_36__38_,chained_data_delayed_36__37_,
  chained_data_delayed_36__36_,chained_data_delayed_36__35_,chained_data_delayed_36__34_,
  chained_data_delayed_36__33_,chained_data_delayed_36__32_,chained_data_delayed_36__31_,
  chained_data_delayed_36__30_,chained_data_delayed_36__29_,
  chained_data_delayed_36__28_,chained_data_delayed_36__27_,chained_data_delayed_36__26_,
  chained_data_delayed_36__25_,chained_data_delayed_36__24_,chained_data_delayed_36__23_,
  chained_data_delayed_36__22_,chained_data_delayed_36__21_,chained_data_delayed_36__20_,
  chained_data_delayed_36__19_,chained_data_delayed_36__18_,
  chained_data_delayed_36__17_,chained_data_delayed_36__16_,chained_data_delayed_36__15_,
  chained_data_delayed_36__14_,chained_data_delayed_36__13_,chained_data_delayed_36__12_,
  chained_data_delayed_36__11_,chained_data_delayed_36__10_,chained_data_delayed_36__9_,
  chained_data_delayed_36__8_,chained_data_delayed_36__7_,chained_data_delayed_36__6_,
  chained_data_delayed_36__5_,chained_data_delayed_36__4_,
  chained_data_delayed_36__3_,chained_data_delayed_36__2_,chained_data_delayed_36__1_,
  chained_data_delayed_36__0_,chained_data_delayed_35__63_,chained_data_delayed_35__62_,
  chained_data_delayed_35__61_,chained_data_delayed_35__60_,chained_data_delayed_35__59_,
  chained_data_delayed_35__58_,chained_data_delayed_35__57_,chained_data_delayed_35__56_,
  chained_data_delayed_35__55_,chained_data_delayed_35__54_,
  chained_data_delayed_35__53_,chained_data_delayed_35__52_,chained_data_delayed_35__51_,
  chained_data_delayed_35__50_,chained_data_delayed_35__49_,chained_data_delayed_35__48_,
  chained_data_delayed_35__47_,chained_data_delayed_35__46_,chained_data_delayed_35__45_,
  chained_data_delayed_35__44_,chained_data_delayed_35__43_,
  chained_data_delayed_35__42_,chained_data_delayed_35__41_,chained_data_delayed_35__40_,
  chained_data_delayed_35__39_,chained_data_delayed_35__38_,chained_data_delayed_35__37_,
  chained_data_delayed_35__36_,chained_data_delayed_35__35_,chained_data_delayed_35__34_,
  chained_data_delayed_35__33_,chained_data_delayed_35__32_,
  chained_data_delayed_35__31_,chained_data_delayed_35__30_,chained_data_delayed_35__29_,
  chained_data_delayed_35__28_,chained_data_delayed_35__27_,chained_data_delayed_35__26_,
  chained_data_delayed_35__25_,chained_data_delayed_35__24_,chained_data_delayed_35__23_,
  chained_data_delayed_35__22_,chained_data_delayed_35__21_,
  chained_data_delayed_35__20_,chained_data_delayed_35__19_,chained_data_delayed_35__18_,
  chained_data_delayed_35__17_,chained_data_delayed_35__16_,chained_data_delayed_35__15_,
  chained_data_delayed_35__14_,chained_data_delayed_35__13_,chained_data_delayed_35__12_,
  chained_data_delayed_35__11_,chained_data_delayed_35__10_,
  chained_data_delayed_35__9_,chained_data_delayed_35__8_,chained_data_delayed_35__7_,
  chained_data_delayed_35__6_,chained_data_delayed_35__5_,chained_data_delayed_35__4_,
  chained_data_delayed_35__3_,chained_data_delayed_35__2_,chained_data_delayed_35__1_,
  chained_data_delayed_35__0_,chained_data_delayed_34__63_,chained_data_delayed_34__62_,
  chained_data_delayed_34__61_,chained_data_delayed_34__60_,chained_data_delayed_34__59_,
  chained_data_delayed_34__58_,chained_data_delayed_34__57_,
  chained_data_delayed_34__56_,chained_data_delayed_34__55_,chained_data_delayed_34__54_,
  chained_data_delayed_34__53_,chained_data_delayed_34__52_,chained_data_delayed_34__51_,
  chained_data_delayed_34__50_,chained_data_delayed_34__49_,chained_data_delayed_34__48_,
  chained_data_delayed_34__47_,chained_data_delayed_34__46_,
  chained_data_delayed_34__45_,chained_data_delayed_34__44_,chained_data_delayed_34__43_,
  chained_data_delayed_34__42_,chained_data_delayed_34__41_,chained_data_delayed_34__40_,
  chained_data_delayed_34__39_,chained_data_delayed_34__38_,chained_data_delayed_34__37_,
  chained_data_delayed_34__36_,chained_data_delayed_34__35_,
  chained_data_delayed_34__34_,chained_data_delayed_34__33_,chained_data_delayed_34__32_,
  chained_data_delayed_34__31_,chained_data_delayed_34__30_,chained_data_delayed_34__29_,
  chained_data_delayed_34__28_,chained_data_delayed_34__27_,chained_data_delayed_34__26_,
  chained_data_delayed_34__25_,chained_data_delayed_34__24_,
  chained_data_delayed_34__23_,chained_data_delayed_34__22_,chained_data_delayed_34__21_,
  chained_data_delayed_34__20_,chained_data_delayed_34__19_,chained_data_delayed_34__18_,
  chained_data_delayed_34__17_,chained_data_delayed_34__16_,chained_data_delayed_34__15_,
  chained_data_delayed_34__14_,chained_data_delayed_34__13_,
  chained_data_delayed_34__12_,chained_data_delayed_34__11_,chained_data_delayed_34__10_,
  chained_data_delayed_34__9_,chained_data_delayed_34__8_,chained_data_delayed_34__7_,
  chained_data_delayed_34__6_,chained_data_delayed_34__5_,chained_data_delayed_34__4_,
  chained_data_delayed_34__3_,chained_data_delayed_34__2_,chained_data_delayed_34__1_,
  chained_data_delayed_34__0_,chained_data_delayed_33__63_,chained_data_delayed_33__62_,
  chained_data_delayed_33__61_,chained_data_delayed_33__60_,
  chained_data_delayed_33__59_,chained_data_delayed_33__58_,chained_data_delayed_33__57_,
  chained_data_delayed_33__56_,chained_data_delayed_33__55_,chained_data_delayed_33__54_,
  chained_data_delayed_33__53_,chained_data_delayed_33__52_,chained_data_delayed_33__51_,
  chained_data_delayed_33__50_,chained_data_delayed_33__49_,
  chained_data_delayed_33__48_,chained_data_delayed_33__47_,chained_data_delayed_33__46_,
  chained_data_delayed_33__45_,chained_data_delayed_33__44_,chained_data_delayed_33__43_,
  chained_data_delayed_33__42_,chained_data_delayed_33__41_,chained_data_delayed_33__40_,
  chained_data_delayed_33__39_,chained_data_delayed_33__38_,
  chained_data_delayed_33__37_,chained_data_delayed_33__36_,chained_data_delayed_33__35_,
  chained_data_delayed_33__34_,chained_data_delayed_33__33_,chained_data_delayed_33__32_,
  chained_data_delayed_33__31_,chained_data_delayed_33__30_,chained_data_delayed_33__29_,
  chained_data_delayed_33__28_,chained_data_delayed_33__27_,
  chained_data_delayed_33__26_,chained_data_delayed_33__25_,chained_data_delayed_33__24_,
  chained_data_delayed_33__23_,chained_data_delayed_33__22_,chained_data_delayed_33__21_,
  chained_data_delayed_33__20_,chained_data_delayed_33__19_,chained_data_delayed_33__18_,
  chained_data_delayed_33__17_,chained_data_delayed_33__16_,
  chained_data_delayed_33__15_,chained_data_delayed_33__14_,chained_data_delayed_33__13_,
  chained_data_delayed_33__12_,chained_data_delayed_33__11_,chained_data_delayed_33__10_,
  chained_data_delayed_33__9_,chained_data_delayed_33__8_,chained_data_delayed_33__7_,
  chained_data_delayed_33__6_,chained_data_delayed_33__5_,chained_data_delayed_33__4_,
  chained_data_delayed_33__3_,chained_data_delayed_33__2_,chained_data_delayed_33__1_,
  chained_data_delayed_33__0_,chained_data_delayed_48__63_,
  chained_data_delayed_48__62_,chained_data_delayed_48__61_,chained_data_delayed_48__60_,
  chained_data_delayed_48__59_,chained_data_delayed_48__58_,chained_data_delayed_48__57_,
  chained_data_delayed_48__56_,chained_data_delayed_48__55_,chained_data_delayed_48__54_,
  chained_data_delayed_48__53_,chained_data_delayed_48__52_,
  chained_data_delayed_48__51_,chained_data_delayed_48__50_,chained_data_delayed_48__49_,
  chained_data_delayed_48__48_,chained_data_delayed_48__47_,chained_data_delayed_48__46_,
  chained_data_delayed_48__45_,chained_data_delayed_48__44_,chained_data_delayed_48__43_,
  chained_data_delayed_48__42_,chained_data_delayed_48__41_,
  chained_data_delayed_48__40_,chained_data_delayed_48__39_,chained_data_delayed_48__38_,
  chained_data_delayed_48__37_,chained_data_delayed_48__36_,chained_data_delayed_48__35_,
  chained_data_delayed_48__34_,chained_data_delayed_48__33_,chained_data_delayed_48__32_,
  chained_data_delayed_48__31_,chained_data_delayed_48__30_,
  chained_data_delayed_48__29_,chained_data_delayed_48__28_,chained_data_delayed_48__27_,
  chained_data_delayed_48__26_,chained_data_delayed_48__25_,chained_data_delayed_48__24_,
  chained_data_delayed_48__23_,chained_data_delayed_48__22_,chained_data_delayed_48__21_,
  chained_data_delayed_48__20_,chained_data_delayed_48__19_,chained_data_delayed_48__18_,
  chained_data_delayed_48__17_,chained_data_delayed_48__16_,
  chained_data_delayed_48__15_,chained_data_delayed_48__14_,chained_data_delayed_48__13_,
  chained_data_delayed_48__12_,chained_data_delayed_48__11_,chained_data_delayed_48__10_,
  chained_data_delayed_48__9_,chained_data_delayed_48__8_,chained_data_delayed_48__7_,
  chained_data_delayed_48__6_,chained_data_delayed_48__5_,chained_data_delayed_48__4_,
  chained_data_delayed_48__3_,chained_data_delayed_48__2_,
  chained_data_delayed_48__1_,chained_data_delayed_48__0_,chained_data_delayed_47__63_,
  chained_data_delayed_47__62_,chained_data_delayed_47__61_,chained_data_delayed_47__60_,
  chained_data_delayed_47__59_,chained_data_delayed_47__58_,chained_data_delayed_47__57_,
  chained_data_delayed_47__56_,chained_data_delayed_47__55_,
  chained_data_delayed_47__54_,chained_data_delayed_47__53_,chained_data_delayed_47__52_,
  chained_data_delayed_47__51_,chained_data_delayed_47__50_,chained_data_delayed_47__49_,
  chained_data_delayed_47__48_,chained_data_delayed_47__47_,chained_data_delayed_47__46_,
  chained_data_delayed_47__45_,chained_data_delayed_47__44_,
  chained_data_delayed_47__43_,chained_data_delayed_47__42_,chained_data_delayed_47__41_,
  chained_data_delayed_47__40_,chained_data_delayed_47__39_,chained_data_delayed_47__38_,
  chained_data_delayed_47__37_,chained_data_delayed_47__36_,chained_data_delayed_47__35_,
  chained_data_delayed_47__34_,chained_data_delayed_47__33_,chained_data_delayed_47__32_,
  chained_data_delayed_47__31_,chained_data_delayed_47__30_,
  chained_data_delayed_47__29_,chained_data_delayed_47__28_,chained_data_delayed_47__27_,
  chained_data_delayed_47__26_,chained_data_delayed_47__25_,chained_data_delayed_47__24_,
  chained_data_delayed_47__23_,chained_data_delayed_47__22_,chained_data_delayed_47__21_,
  chained_data_delayed_47__20_,chained_data_delayed_47__19_,
  chained_data_delayed_47__18_,chained_data_delayed_47__17_,chained_data_delayed_47__16_,
  chained_data_delayed_47__15_,chained_data_delayed_47__14_,chained_data_delayed_47__13_,
  chained_data_delayed_47__12_,chained_data_delayed_47__11_,chained_data_delayed_47__10_,
  chained_data_delayed_47__9_,chained_data_delayed_47__8_,
  chained_data_delayed_47__7_,chained_data_delayed_47__6_,chained_data_delayed_47__5_,
  chained_data_delayed_47__4_,chained_data_delayed_47__3_,chained_data_delayed_47__2_,
  chained_data_delayed_47__1_,chained_data_delayed_47__0_,chained_data_delayed_46__63_,
  chained_data_delayed_46__62_,chained_data_delayed_46__61_,chained_data_delayed_46__60_,
  chained_data_delayed_46__59_,chained_data_delayed_46__58_,
  chained_data_delayed_46__57_,chained_data_delayed_46__56_,chained_data_delayed_46__55_,
  chained_data_delayed_46__54_,chained_data_delayed_46__53_,chained_data_delayed_46__52_,
  chained_data_delayed_46__51_,chained_data_delayed_46__50_,chained_data_delayed_46__49_,
  chained_data_delayed_46__48_,chained_data_delayed_46__47_,chained_data_delayed_46__46_,
  chained_data_delayed_46__45_,chained_data_delayed_46__44_,
  chained_data_delayed_46__43_,chained_data_delayed_46__42_,chained_data_delayed_46__41_,
  chained_data_delayed_46__40_,chained_data_delayed_46__39_,chained_data_delayed_46__38_,
  chained_data_delayed_46__37_,chained_data_delayed_46__36_,chained_data_delayed_46__35_,
  chained_data_delayed_46__34_,chained_data_delayed_46__33_,
  chained_data_delayed_46__32_,chained_data_delayed_46__31_,chained_data_delayed_46__30_,
  chained_data_delayed_46__29_,chained_data_delayed_46__28_,chained_data_delayed_46__27_,
  chained_data_delayed_46__26_,chained_data_delayed_46__25_,chained_data_delayed_46__24_,
  chained_data_delayed_46__23_,chained_data_delayed_46__22_,
  chained_data_delayed_46__21_,chained_data_delayed_46__20_,chained_data_delayed_46__19_,
  chained_data_delayed_46__18_,chained_data_delayed_46__17_,chained_data_delayed_46__16_,
  chained_data_delayed_46__15_,chained_data_delayed_46__14_,chained_data_delayed_46__13_,
  chained_data_delayed_46__12_,chained_data_delayed_46__11_,
  chained_data_delayed_46__10_,chained_data_delayed_46__9_,chained_data_delayed_46__8_,
  chained_data_delayed_46__7_,chained_data_delayed_46__6_,chained_data_delayed_46__5_,
  chained_data_delayed_46__4_,chained_data_delayed_46__3_,chained_data_delayed_46__2_,
  chained_data_delayed_46__1_,chained_data_delayed_46__0_,chained_data_delayed_45__63_,
  chained_data_delayed_45__62_,chained_data_delayed_45__61_,chained_data_delayed_45__60_,
  chained_data_delayed_45__59_,chained_data_delayed_45__58_,
  chained_data_delayed_45__57_,chained_data_delayed_45__56_,chained_data_delayed_45__55_,
  chained_data_delayed_45__54_,chained_data_delayed_45__53_,chained_data_delayed_45__52_,
  chained_data_delayed_45__51_,chained_data_delayed_45__50_,chained_data_delayed_45__49_,
  chained_data_delayed_45__48_,chained_data_delayed_45__47_,
  chained_data_delayed_45__46_,chained_data_delayed_45__45_,chained_data_delayed_45__44_,
  chained_data_delayed_45__43_,chained_data_delayed_45__42_,chained_data_delayed_45__41_,
  chained_data_delayed_45__40_,chained_data_delayed_45__39_,chained_data_delayed_45__38_,
  chained_data_delayed_45__37_,chained_data_delayed_45__36_,
  chained_data_delayed_45__35_,chained_data_delayed_45__34_,chained_data_delayed_45__33_,
  chained_data_delayed_45__32_,chained_data_delayed_45__31_,chained_data_delayed_45__30_,
  chained_data_delayed_45__29_,chained_data_delayed_45__28_,chained_data_delayed_45__27_,
  chained_data_delayed_45__26_,chained_data_delayed_45__25_,
  chained_data_delayed_45__24_,chained_data_delayed_45__23_,chained_data_delayed_45__22_,
  chained_data_delayed_45__21_,chained_data_delayed_45__20_,chained_data_delayed_45__19_,
  chained_data_delayed_45__18_,chained_data_delayed_45__17_,chained_data_delayed_45__16_,
  chained_data_delayed_45__15_,chained_data_delayed_45__14_,
  chained_data_delayed_45__13_,chained_data_delayed_45__12_,chained_data_delayed_45__11_,
  chained_data_delayed_45__10_,chained_data_delayed_45__9_,chained_data_delayed_45__8_,
  chained_data_delayed_45__7_,chained_data_delayed_45__6_,chained_data_delayed_45__5_,
  chained_data_delayed_45__4_,chained_data_delayed_45__3_,chained_data_delayed_45__2_,
  chained_data_delayed_45__1_,chained_data_delayed_45__0_,chained_data_delayed_44__63_,
  chained_data_delayed_44__62_,chained_data_delayed_44__61_,
  chained_data_delayed_44__60_,chained_data_delayed_44__59_,chained_data_delayed_44__58_,
  chained_data_delayed_44__57_,chained_data_delayed_44__56_,chained_data_delayed_44__55_,
  chained_data_delayed_44__54_,chained_data_delayed_44__53_,chained_data_delayed_44__52_,
  chained_data_delayed_44__51_,chained_data_delayed_44__50_,
  chained_data_delayed_44__49_,chained_data_delayed_44__48_,chained_data_delayed_44__47_,
  chained_data_delayed_44__46_,chained_data_delayed_44__45_,chained_data_delayed_44__44_,
  chained_data_delayed_44__43_,chained_data_delayed_44__42_,chained_data_delayed_44__41_,
  chained_data_delayed_44__40_,chained_data_delayed_44__39_,
  chained_data_delayed_44__38_,chained_data_delayed_44__37_,chained_data_delayed_44__36_,
  chained_data_delayed_44__35_,chained_data_delayed_44__34_,chained_data_delayed_44__33_,
  chained_data_delayed_44__32_,chained_data_delayed_44__31_,chained_data_delayed_44__30_,
  chained_data_delayed_44__29_,chained_data_delayed_44__28_,
  chained_data_delayed_44__27_,chained_data_delayed_44__26_,chained_data_delayed_44__25_,
  chained_data_delayed_44__24_,chained_data_delayed_44__23_,chained_data_delayed_44__22_,
  chained_data_delayed_44__21_,chained_data_delayed_44__20_,chained_data_delayed_44__19_,
  chained_data_delayed_44__18_,chained_data_delayed_44__17_,
  chained_data_delayed_44__16_,chained_data_delayed_44__15_,chained_data_delayed_44__14_,
  chained_data_delayed_44__13_,chained_data_delayed_44__12_,chained_data_delayed_44__11_,
  chained_data_delayed_44__10_,chained_data_delayed_44__9_,chained_data_delayed_44__8_,
  chained_data_delayed_44__7_,chained_data_delayed_44__6_,chained_data_delayed_44__5_,
  chained_data_delayed_44__4_,chained_data_delayed_44__3_,chained_data_delayed_44__2_,
  chained_data_delayed_44__1_,chained_data_delayed_44__0_,
  chained_data_delayed_43__63_,chained_data_delayed_43__62_,chained_data_delayed_43__61_,
  chained_data_delayed_43__60_,chained_data_delayed_43__59_,chained_data_delayed_43__58_,
  chained_data_delayed_43__57_,chained_data_delayed_43__56_,chained_data_delayed_43__55_,
  chained_data_delayed_43__54_,chained_data_delayed_43__53_,
  chained_data_delayed_43__52_,chained_data_delayed_43__51_,chained_data_delayed_43__50_,
  chained_data_delayed_43__49_,chained_data_delayed_43__48_,chained_data_delayed_43__47_,
  chained_data_delayed_43__46_,chained_data_delayed_43__45_,chained_data_delayed_43__44_,
  chained_data_delayed_43__43_,chained_data_delayed_43__42_,
  chained_data_delayed_43__41_,chained_data_delayed_43__40_,chained_data_delayed_43__39_,
  chained_data_delayed_43__38_,chained_data_delayed_43__37_,chained_data_delayed_43__36_,
  chained_data_delayed_43__35_,chained_data_delayed_43__34_,chained_data_delayed_43__33_,
  chained_data_delayed_43__32_,chained_data_delayed_43__31_,
  chained_data_delayed_43__30_,chained_data_delayed_43__29_,chained_data_delayed_43__28_,
  chained_data_delayed_43__27_,chained_data_delayed_43__26_,chained_data_delayed_43__25_,
  chained_data_delayed_43__24_,chained_data_delayed_43__23_,chained_data_delayed_43__22_,
  chained_data_delayed_43__21_,chained_data_delayed_43__20_,
  chained_data_delayed_43__19_,chained_data_delayed_43__18_,chained_data_delayed_43__17_,
  chained_data_delayed_43__16_,chained_data_delayed_43__15_,chained_data_delayed_43__14_,
  chained_data_delayed_43__13_,chained_data_delayed_43__12_,chained_data_delayed_43__11_,
  chained_data_delayed_43__10_,chained_data_delayed_43__9_,chained_data_delayed_43__8_,
  chained_data_delayed_43__7_,chained_data_delayed_43__6_,
  chained_data_delayed_43__5_,chained_data_delayed_43__4_,chained_data_delayed_43__3_,
  chained_data_delayed_43__2_,chained_data_delayed_43__1_,chained_data_delayed_43__0_,
  chained_data_delayed_42__63_,chained_data_delayed_42__62_,chained_data_delayed_42__61_,
  chained_data_delayed_42__60_,chained_data_delayed_42__59_,chained_data_delayed_42__58_,
  chained_data_delayed_42__57_,chained_data_delayed_42__56_,
  chained_data_delayed_42__55_,chained_data_delayed_42__54_,chained_data_delayed_42__53_,
  chained_data_delayed_42__52_,chained_data_delayed_42__51_,chained_data_delayed_42__50_,
  chained_data_delayed_42__49_,chained_data_delayed_42__48_,chained_data_delayed_42__47_,
  chained_data_delayed_42__46_,chained_data_delayed_42__45_,
  chained_data_delayed_42__44_,chained_data_delayed_42__43_,chained_data_delayed_42__42_,
  chained_data_delayed_42__41_,chained_data_delayed_42__40_,chained_data_delayed_42__39_,
  chained_data_delayed_42__38_,chained_data_delayed_42__37_,chained_data_delayed_42__36_,
  chained_data_delayed_42__35_,chained_data_delayed_42__34_,
  chained_data_delayed_42__33_,chained_data_delayed_42__32_,chained_data_delayed_42__31_,
  chained_data_delayed_42__30_,chained_data_delayed_42__29_,chained_data_delayed_42__28_,
  chained_data_delayed_42__27_,chained_data_delayed_42__26_,chained_data_delayed_42__25_,
  chained_data_delayed_42__24_,chained_data_delayed_42__23_,chained_data_delayed_42__22_,
  chained_data_delayed_42__21_,chained_data_delayed_42__20_,
  chained_data_delayed_42__19_,chained_data_delayed_42__18_,chained_data_delayed_42__17_,
  chained_data_delayed_42__16_,chained_data_delayed_42__15_,chained_data_delayed_42__14_,
  chained_data_delayed_42__13_,chained_data_delayed_42__12_,chained_data_delayed_42__11_,
  chained_data_delayed_42__10_,chained_data_delayed_42__9_,
  chained_data_delayed_42__8_,chained_data_delayed_42__7_,chained_data_delayed_42__6_,
  chained_data_delayed_42__5_,chained_data_delayed_42__4_,chained_data_delayed_42__3_,
  chained_data_delayed_42__2_,chained_data_delayed_42__1_,chained_data_delayed_42__0_,
  chained_data_delayed_41__63_,chained_data_delayed_41__62_,chained_data_delayed_41__61_,
  chained_data_delayed_41__60_,chained_data_delayed_41__59_,
  chained_data_delayed_41__58_,chained_data_delayed_41__57_,chained_data_delayed_41__56_,
  chained_data_delayed_41__55_,chained_data_delayed_41__54_,chained_data_delayed_41__53_,
  chained_data_delayed_41__52_,chained_data_delayed_41__51_,chained_data_delayed_41__50_,
  chained_data_delayed_41__49_,chained_data_delayed_41__48_,
  chained_data_delayed_41__47_,chained_data_delayed_41__46_,chained_data_delayed_41__45_,
  chained_data_delayed_41__44_,chained_data_delayed_41__43_,chained_data_delayed_41__42_,
  chained_data_delayed_41__41_,chained_data_delayed_41__40_,chained_data_delayed_41__39_,
  chained_data_delayed_41__38_,chained_data_delayed_41__37_,chained_data_delayed_41__36_,
  chained_data_delayed_41__35_,chained_data_delayed_41__34_,
  chained_data_delayed_41__33_,chained_data_delayed_41__32_,chained_data_delayed_41__31_,
  chained_data_delayed_41__30_,chained_data_delayed_41__29_,chained_data_delayed_41__28_,
  chained_data_delayed_41__27_,chained_data_delayed_41__26_,chained_data_delayed_41__25_,
  chained_data_delayed_41__24_,chained_data_delayed_41__23_,
  chained_data_delayed_41__22_,chained_data_delayed_41__21_,chained_data_delayed_41__20_,
  chained_data_delayed_41__19_,chained_data_delayed_41__18_,chained_data_delayed_41__17_,
  chained_data_delayed_41__16_,chained_data_delayed_41__15_,chained_data_delayed_41__14_,
  chained_data_delayed_41__13_,chained_data_delayed_41__12_,
  chained_data_delayed_41__11_,chained_data_delayed_41__10_,chained_data_delayed_41__9_,
  chained_data_delayed_41__8_,chained_data_delayed_41__7_,chained_data_delayed_41__6_,
  chained_data_delayed_41__5_,chained_data_delayed_41__4_,chained_data_delayed_41__3_,
  chained_data_delayed_41__2_,chained_data_delayed_41__1_,chained_data_delayed_41__0_,
  chained_data_delayed_56__63_,chained_data_delayed_56__62_,
  chained_data_delayed_56__61_,chained_data_delayed_56__60_,chained_data_delayed_56__59_,
  chained_data_delayed_56__58_,chained_data_delayed_56__57_,chained_data_delayed_56__56_,
  chained_data_delayed_56__55_,chained_data_delayed_56__54_,chained_data_delayed_56__53_,
  chained_data_delayed_56__52_,chained_data_delayed_56__51_,chained_data_delayed_56__50_,
  chained_data_delayed_56__49_,chained_data_delayed_56__48_,
  chained_data_delayed_56__47_,chained_data_delayed_56__46_,chained_data_delayed_56__45_,
  chained_data_delayed_56__44_,chained_data_delayed_56__43_,chained_data_delayed_56__42_,
  chained_data_delayed_56__41_,chained_data_delayed_56__40_,chained_data_delayed_56__39_,
  chained_data_delayed_56__38_,chained_data_delayed_56__37_,
  chained_data_delayed_56__36_,chained_data_delayed_56__35_,chained_data_delayed_56__34_,
  chained_data_delayed_56__33_,chained_data_delayed_56__32_,chained_data_delayed_56__31_,
  chained_data_delayed_56__30_,chained_data_delayed_56__29_,chained_data_delayed_56__28_,
  chained_data_delayed_56__27_,chained_data_delayed_56__26_,
  chained_data_delayed_56__25_,chained_data_delayed_56__24_,chained_data_delayed_56__23_,
  chained_data_delayed_56__22_,chained_data_delayed_56__21_,chained_data_delayed_56__20_,
  chained_data_delayed_56__19_,chained_data_delayed_56__18_,chained_data_delayed_56__17_,
  chained_data_delayed_56__16_,chained_data_delayed_56__15_,
  chained_data_delayed_56__14_,chained_data_delayed_56__13_,chained_data_delayed_56__12_,
  chained_data_delayed_56__11_,chained_data_delayed_56__10_,chained_data_delayed_56__9_,
  chained_data_delayed_56__8_,chained_data_delayed_56__7_,chained_data_delayed_56__6_,
  chained_data_delayed_56__5_,chained_data_delayed_56__4_,chained_data_delayed_56__3_,
  chained_data_delayed_56__2_,chained_data_delayed_56__1_,chained_data_delayed_56__0_,
  chained_data_delayed_55__63_,chained_data_delayed_55__62_,
  chained_data_delayed_55__61_,chained_data_delayed_55__60_,chained_data_delayed_55__59_,
  chained_data_delayed_55__58_,chained_data_delayed_55__57_,chained_data_delayed_55__56_,
  chained_data_delayed_55__55_,chained_data_delayed_55__54_,chained_data_delayed_55__53_,
  chained_data_delayed_55__52_,chained_data_delayed_55__51_,
  chained_data_delayed_55__50_,chained_data_delayed_55__49_,chained_data_delayed_55__48_,
  chained_data_delayed_55__47_,chained_data_delayed_55__46_,chained_data_delayed_55__45_,
  chained_data_delayed_55__44_,chained_data_delayed_55__43_,chained_data_delayed_55__42_,
  chained_data_delayed_55__41_,chained_data_delayed_55__40_,
  chained_data_delayed_55__39_,chained_data_delayed_55__38_,chained_data_delayed_55__37_,
  chained_data_delayed_55__36_,chained_data_delayed_55__35_,chained_data_delayed_55__34_,
  chained_data_delayed_55__33_,chained_data_delayed_55__32_,chained_data_delayed_55__31_,
  chained_data_delayed_55__30_,chained_data_delayed_55__29_,
  chained_data_delayed_55__28_,chained_data_delayed_55__27_,chained_data_delayed_55__26_,
  chained_data_delayed_55__25_,chained_data_delayed_55__24_,chained_data_delayed_55__23_,
  chained_data_delayed_55__22_,chained_data_delayed_55__21_,chained_data_delayed_55__20_,
  chained_data_delayed_55__19_,chained_data_delayed_55__18_,
  chained_data_delayed_55__17_,chained_data_delayed_55__16_,chained_data_delayed_55__15_,
  chained_data_delayed_55__14_,chained_data_delayed_55__13_,chained_data_delayed_55__12_,
  chained_data_delayed_55__11_,chained_data_delayed_55__10_,chained_data_delayed_55__9_,
  chained_data_delayed_55__8_,chained_data_delayed_55__7_,chained_data_delayed_55__6_,
  chained_data_delayed_55__5_,chained_data_delayed_55__4_,
  chained_data_delayed_55__3_,chained_data_delayed_55__2_,chained_data_delayed_55__1_,
  chained_data_delayed_55__0_,chained_data_delayed_54__63_,chained_data_delayed_54__62_,
  chained_data_delayed_54__61_,chained_data_delayed_54__60_,chained_data_delayed_54__59_,
  chained_data_delayed_54__58_,chained_data_delayed_54__57_,chained_data_delayed_54__56_,
  chained_data_delayed_54__55_,chained_data_delayed_54__54_,
  chained_data_delayed_54__53_,chained_data_delayed_54__52_,chained_data_delayed_54__51_,
  chained_data_delayed_54__50_,chained_data_delayed_54__49_,chained_data_delayed_54__48_,
  chained_data_delayed_54__47_,chained_data_delayed_54__46_,chained_data_delayed_54__45_,
  chained_data_delayed_54__44_,chained_data_delayed_54__43_,
  chained_data_delayed_54__42_,chained_data_delayed_54__41_,chained_data_delayed_54__40_,
  chained_data_delayed_54__39_,chained_data_delayed_54__38_,chained_data_delayed_54__37_,
  chained_data_delayed_54__36_,chained_data_delayed_54__35_,chained_data_delayed_54__34_,
  chained_data_delayed_54__33_,chained_data_delayed_54__32_,
  chained_data_delayed_54__31_,chained_data_delayed_54__30_,chained_data_delayed_54__29_,
  chained_data_delayed_54__28_,chained_data_delayed_54__27_,chained_data_delayed_54__26_,
  chained_data_delayed_54__25_,chained_data_delayed_54__24_,chained_data_delayed_54__23_,
  chained_data_delayed_54__22_,chained_data_delayed_54__21_,
  chained_data_delayed_54__20_,chained_data_delayed_54__19_,chained_data_delayed_54__18_,
  chained_data_delayed_54__17_,chained_data_delayed_54__16_,chained_data_delayed_54__15_,
  chained_data_delayed_54__14_,chained_data_delayed_54__13_,chained_data_delayed_54__12_,
  chained_data_delayed_54__11_,chained_data_delayed_54__10_,chained_data_delayed_54__9_,
  chained_data_delayed_54__8_,chained_data_delayed_54__7_,
  chained_data_delayed_54__6_,chained_data_delayed_54__5_,chained_data_delayed_54__4_,
  chained_data_delayed_54__3_,chained_data_delayed_54__2_,chained_data_delayed_54__1_,
  chained_data_delayed_54__0_,chained_data_delayed_53__63_,chained_data_delayed_53__62_,
  chained_data_delayed_53__61_,chained_data_delayed_53__60_,chained_data_delayed_53__59_,
  chained_data_delayed_53__58_,chained_data_delayed_53__57_,
  chained_data_delayed_53__56_,chained_data_delayed_53__55_,chained_data_delayed_53__54_,
  chained_data_delayed_53__53_,chained_data_delayed_53__52_,chained_data_delayed_53__51_,
  chained_data_delayed_53__50_,chained_data_delayed_53__49_,chained_data_delayed_53__48_,
  chained_data_delayed_53__47_,chained_data_delayed_53__46_,
  chained_data_delayed_53__45_,chained_data_delayed_53__44_,chained_data_delayed_53__43_,
  chained_data_delayed_53__42_,chained_data_delayed_53__41_,chained_data_delayed_53__40_,
  chained_data_delayed_53__39_,chained_data_delayed_53__38_,chained_data_delayed_53__37_,
  chained_data_delayed_53__36_,chained_data_delayed_53__35_,
  chained_data_delayed_53__34_,chained_data_delayed_53__33_,chained_data_delayed_53__32_,
  chained_data_delayed_53__31_,chained_data_delayed_53__30_,chained_data_delayed_53__29_,
  chained_data_delayed_53__28_,chained_data_delayed_53__27_,chained_data_delayed_53__26_,
  chained_data_delayed_53__25_,chained_data_delayed_53__24_,
  chained_data_delayed_53__23_,chained_data_delayed_53__22_,chained_data_delayed_53__21_,
  chained_data_delayed_53__20_,chained_data_delayed_53__19_,chained_data_delayed_53__18_,
  chained_data_delayed_53__17_,chained_data_delayed_53__16_,chained_data_delayed_53__15_,
  chained_data_delayed_53__14_,chained_data_delayed_53__13_,chained_data_delayed_53__12_,
  chained_data_delayed_53__11_,chained_data_delayed_53__10_,
  chained_data_delayed_53__9_,chained_data_delayed_53__8_,chained_data_delayed_53__7_,
  chained_data_delayed_53__6_,chained_data_delayed_53__5_,chained_data_delayed_53__4_,
  chained_data_delayed_53__3_,chained_data_delayed_53__2_,chained_data_delayed_53__1_,
  chained_data_delayed_53__0_,chained_data_delayed_52__63_,chained_data_delayed_52__62_,
  chained_data_delayed_52__61_,chained_data_delayed_52__60_,
  chained_data_delayed_52__59_,chained_data_delayed_52__58_,chained_data_delayed_52__57_,
  chained_data_delayed_52__56_,chained_data_delayed_52__55_,chained_data_delayed_52__54_,
  chained_data_delayed_52__53_,chained_data_delayed_52__52_,chained_data_delayed_52__51_,
  chained_data_delayed_52__50_,chained_data_delayed_52__49_,
  chained_data_delayed_52__48_,chained_data_delayed_52__47_,chained_data_delayed_52__46_,
  chained_data_delayed_52__45_,chained_data_delayed_52__44_,chained_data_delayed_52__43_,
  chained_data_delayed_52__42_,chained_data_delayed_52__41_,chained_data_delayed_52__40_,
  chained_data_delayed_52__39_,chained_data_delayed_52__38_,
  chained_data_delayed_52__37_,chained_data_delayed_52__36_,chained_data_delayed_52__35_,
  chained_data_delayed_52__34_,chained_data_delayed_52__33_,chained_data_delayed_52__32_,
  chained_data_delayed_52__31_,chained_data_delayed_52__30_,chained_data_delayed_52__29_,
  chained_data_delayed_52__28_,chained_data_delayed_52__27_,chained_data_delayed_52__26_,
  chained_data_delayed_52__25_,chained_data_delayed_52__24_,
  chained_data_delayed_52__23_,chained_data_delayed_52__22_,chained_data_delayed_52__21_,
  chained_data_delayed_52__20_,chained_data_delayed_52__19_,chained_data_delayed_52__18_,
  chained_data_delayed_52__17_,chained_data_delayed_52__16_,chained_data_delayed_52__15_,
  chained_data_delayed_52__14_,chained_data_delayed_52__13_,
  chained_data_delayed_52__12_,chained_data_delayed_52__11_,chained_data_delayed_52__10_,
  chained_data_delayed_52__9_,chained_data_delayed_52__8_,chained_data_delayed_52__7_,
  chained_data_delayed_52__6_,chained_data_delayed_52__5_,chained_data_delayed_52__4_,
  chained_data_delayed_52__3_,chained_data_delayed_52__2_,chained_data_delayed_52__1_,
  chained_data_delayed_52__0_,chained_data_delayed_51__63_,
  chained_data_delayed_51__62_,chained_data_delayed_51__61_,chained_data_delayed_51__60_,
  chained_data_delayed_51__59_,chained_data_delayed_51__58_,chained_data_delayed_51__57_,
  chained_data_delayed_51__56_,chained_data_delayed_51__55_,chained_data_delayed_51__54_,
  chained_data_delayed_51__53_,chained_data_delayed_51__52_,
  chained_data_delayed_51__51_,chained_data_delayed_51__50_,chained_data_delayed_51__49_,
  chained_data_delayed_51__48_,chained_data_delayed_51__47_,chained_data_delayed_51__46_,
  chained_data_delayed_51__45_,chained_data_delayed_51__44_,chained_data_delayed_51__43_,
  chained_data_delayed_51__42_,chained_data_delayed_51__41_,chained_data_delayed_51__40_,
  chained_data_delayed_51__39_,chained_data_delayed_51__38_,
  chained_data_delayed_51__37_,chained_data_delayed_51__36_,chained_data_delayed_51__35_,
  chained_data_delayed_51__34_,chained_data_delayed_51__33_,chained_data_delayed_51__32_,
  chained_data_delayed_51__31_,chained_data_delayed_51__30_,chained_data_delayed_51__29_,
  chained_data_delayed_51__28_,chained_data_delayed_51__27_,
  chained_data_delayed_51__26_,chained_data_delayed_51__25_,chained_data_delayed_51__24_,
  chained_data_delayed_51__23_,chained_data_delayed_51__22_,chained_data_delayed_51__21_,
  chained_data_delayed_51__20_,chained_data_delayed_51__19_,chained_data_delayed_51__18_,
  chained_data_delayed_51__17_,chained_data_delayed_51__16_,
  chained_data_delayed_51__15_,chained_data_delayed_51__14_,chained_data_delayed_51__13_,
  chained_data_delayed_51__12_,chained_data_delayed_51__11_,chained_data_delayed_51__10_,
  chained_data_delayed_51__9_,chained_data_delayed_51__8_,chained_data_delayed_51__7_,
  chained_data_delayed_51__6_,chained_data_delayed_51__5_,chained_data_delayed_51__4_,
  chained_data_delayed_51__3_,chained_data_delayed_51__2_,
  chained_data_delayed_51__1_,chained_data_delayed_51__0_,chained_data_delayed_50__63_,
  chained_data_delayed_50__62_,chained_data_delayed_50__61_,chained_data_delayed_50__60_,
  chained_data_delayed_50__59_,chained_data_delayed_50__58_,chained_data_delayed_50__57_,
  chained_data_delayed_50__56_,chained_data_delayed_50__55_,chained_data_delayed_50__54_,
  chained_data_delayed_50__53_,chained_data_delayed_50__52_,
  chained_data_delayed_50__51_,chained_data_delayed_50__50_,chained_data_delayed_50__49_,
  chained_data_delayed_50__48_,chained_data_delayed_50__47_,chained_data_delayed_50__46_,
  chained_data_delayed_50__45_,chained_data_delayed_50__44_,chained_data_delayed_50__43_,
  chained_data_delayed_50__42_,chained_data_delayed_50__41_,
  chained_data_delayed_50__40_,chained_data_delayed_50__39_,chained_data_delayed_50__38_,
  chained_data_delayed_50__37_,chained_data_delayed_50__36_,chained_data_delayed_50__35_,
  chained_data_delayed_50__34_,chained_data_delayed_50__33_,chained_data_delayed_50__32_,
  chained_data_delayed_50__31_,chained_data_delayed_50__30_,
  chained_data_delayed_50__29_,chained_data_delayed_50__28_,chained_data_delayed_50__27_,
  chained_data_delayed_50__26_,chained_data_delayed_50__25_,chained_data_delayed_50__24_,
  chained_data_delayed_50__23_,chained_data_delayed_50__22_,chained_data_delayed_50__21_,
  chained_data_delayed_50__20_,chained_data_delayed_50__19_,
  chained_data_delayed_50__18_,chained_data_delayed_50__17_,chained_data_delayed_50__16_,
  chained_data_delayed_50__15_,chained_data_delayed_50__14_,chained_data_delayed_50__13_,
  chained_data_delayed_50__12_,chained_data_delayed_50__11_,chained_data_delayed_50__10_,
  chained_data_delayed_50__9_,chained_data_delayed_50__8_,chained_data_delayed_50__7_,
  chained_data_delayed_50__6_,chained_data_delayed_50__5_,
  chained_data_delayed_50__4_,chained_data_delayed_50__3_,chained_data_delayed_50__2_,
  chained_data_delayed_50__1_,chained_data_delayed_50__0_,chained_data_delayed_49__63_,
  chained_data_delayed_49__62_,chained_data_delayed_49__61_,chained_data_delayed_49__60_,
  chained_data_delayed_49__59_,chained_data_delayed_49__58_,chained_data_delayed_49__57_,
  chained_data_delayed_49__56_,chained_data_delayed_49__55_,
  chained_data_delayed_49__54_,chained_data_delayed_49__53_,chained_data_delayed_49__52_,
  chained_data_delayed_49__51_,chained_data_delayed_49__50_,chained_data_delayed_49__49_,
  chained_data_delayed_49__48_,chained_data_delayed_49__47_,chained_data_delayed_49__46_,
  chained_data_delayed_49__45_,chained_data_delayed_49__44_,
  chained_data_delayed_49__43_,chained_data_delayed_49__42_,chained_data_delayed_49__41_,
  chained_data_delayed_49__40_,chained_data_delayed_49__39_,chained_data_delayed_49__38_,
  chained_data_delayed_49__37_,chained_data_delayed_49__36_,chained_data_delayed_49__35_,
  chained_data_delayed_49__34_,chained_data_delayed_49__33_,
  chained_data_delayed_49__32_,chained_data_delayed_49__31_,chained_data_delayed_49__30_,
  chained_data_delayed_49__29_,chained_data_delayed_49__28_,chained_data_delayed_49__27_,
  chained_data_delayed_49__26_,chained_data_delayed_49__25_,chained_data_delayed_49__24_,
  chained_data_delayed_49__23_,chained_data_delayed_49__22_,
  chained_data_delayed_49__21_,chained_data_delayed_49__20_,chained_data_delayed_49__19_,
  chained_data_delayed_49__18_,chained_data_delayed_49__17_,chained_data_delayed_49__16_,
  chained_data_delayed_49__15_,chained_data_delayed_49__14_,chained_data_delayed_49__13_,
  chained_data_delayed_49__12_,chained_data_delayed_49__11_,
  chained_data_delayed_49__10_,chained_data_delayed_49__9_,chained_data_delayed_49__8_,
  chained_data_delayed_49__7_,chained_data_delayed_49__6_,chained_data_delayed_49__5_,
  chained_data_delayed_49__4_,chained_data_delayed_49__3_,chained_data_delayed_49__2_,
  chained_data_delayed_49__1_,chained_data_delayed_49__0_;

  bsg_dff_width_p64
  chained_genblk1_1__ch_reg
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .data_o({ chained_data_delayed_1__63_, chained_data_delayed_1__62_, chained_data_delayed_1__61_, chained_data_delayed_1__60_, chained_data_delayed_1__59_, chained_data_delayed_1__58_, chained_data_delayed_1__57_, chained_data_delayed_1__56_, chained_data_delayed_1__55_, chained_data_delayed_1__54_, chained_data_delayed_1__53_, chained_data_delayed_1__52_, chained_data_delayed_1__51_, chained_data_delayed_1__50_, chained_data_delayed_1__49_, chained_data_delayed_1__48_, chained_data_delayed_1__47_, chained_data_delayed_1__46_, chained_data_delayed_1__45_, chained_data_delayed_1__44_, chained_data_delayed_1__43_, chained_data_delayed_1__42_, chained_data_delayed_1__41_, chained_data_delayed_1__40_, chained_data_delayed_1__39_, chained_data_delayed_1__38_, chained_data_delayed_1__37_, chained_data_delayed_1__36_, chained_data_delayed_1__35_, chained_data_delayed_1__34_, chained_data_delayed_1__33_, chained_data_delayed_1__32_, chained_data_delayed_1__31_, chained_data_delayed_1__30_, chained_data_delayed_1__29_, chained_data_delayed_1__28_, chained_data_delayed_1__27_, chained_data_delayed_1__26_, chained_data_delayed_1__25_, chained_data_delayed_1__24_, chained_data_delayed_1__23_, chained_data_delayed_1__22_, chained_data_delayed_1__21_, chained_data_delayed_1__20_, chained_data_delayed_1__19_, chained_data_delayed_1__18_, chained_data_delayed_1__17_, chained_data_delayed_1__16_, chained_data_delayed_1__15_, chained_data_delayed_1__14_, chained_data_delayed_1__13_, chained_data_delayed_1__12_, chained_data_delayed_1__11_, chained_data_delayed_1__10_, chained_data_delayed_1__9_, chained_data_delayed_1__8_, chained_data_delayed_1__7_, chained_data_delayed_1__6_, chained_data_delayed_1__5_, chained_data_delayed_1__4_, chained_data_delayed_1__3_, chained_data_delayed_1__2_, chained_data_delayed_1__1_, chained_data_delayed_1__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_2__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_1__63_, chained_data_delayed_1__62_, chained_data_delayed_1__61_, chained_data_delayed_1__60_, chained_data_delayed_1__59_, chained_data_delayed_1__58_, chained_data_delayed_1__57_, chained_data_delayed_1__56_, chained_data_delayed_1__55_, chained_data_delayed_1__54_, chained_data_delayed_1__53_, chained_data_delayed_1__52_, chained_data_delayed_1__51_, chained_data_delayed_1__50_, chained_data_delayed_1__49_, chained_data_delayed_1__48_, chained_data_delayed_1__47_, chained_data_delayed_1__46_, chained_data_delayed_1__45_, chained_data_delayed_1__44_, chained_data_delayed_1__43_, chained_data_delayed_1__42_, chained_data_delayed_1__41_, chained_data_delayed_1__40_, chained_data_delayed_1__39_, chained_data_delayed_1__38_, chained_data_delayed_1__37_, chained_data_delayed_1__36_, chained_data_delayed_1__35_, chained_data_delayed_1__34_, chained_data_delayed_1__33_, chained_data_delayed_1__32_, chained_data_delayed_1__31_, chained_data_delayed_1__30_, chained_data_delayed_1__29_, chained_data_delayed_1__28_, chained_data_delayed_1__27_, chained_data_delayed_1__26_, chained_data_delayed_1__25_, chained_data_delayed_1__24_, chained_data_delayed_1__23_, chained_data_delayed_1__22_, chained_data_delayed_1__21_, chained_data_delayed_1__20_, chained_data_delayed_1__19_, chained_data_delayed_1__18_, chained_data_delayed_1__17_, chained_data_delayed_1__16_, chained_data_delayed_1__15_, chained_data_delayed_1__14_, chained_data_delayed_1__13_, chained_data_delayed_1__12_, chained_data_delayed_1__11_, chained_data_delayed_1__10_, chained_data_delayed_1__9_, chained_data_delayed_1__8_, chained_data_delayed_1__7_, chained_data_delayed_1__6_, chained_data_delayed_1__5_, chained_data_delayed_1__4_, chained_data_delayed_1__3_, chained_data_delayed_1__2_, chained_data_delayed_1__1_, chained_data_delayed_1__0_ }),
    .data_o({ chained_data_delayed_2__63_, chained_data_delayed_2__62_, chained_data_delayed_2__61_, chained_data_delayed_2__60_, chained_data_delayed_2__59_, chained_data_delayed_2__58_, chained_data_delayed_2__57_, chained_data_delayed_2__56_, chained_data_delayed_2__55_, chained_data_delayed_2__54_, chained_data_delayed_2__53_, chained_data_delayed_2__52_, chained_data_delayed_2__51_, chained_data_delayed_2__50_, chained_data_delayed_2__49_, chained_data_delayed_2__48_, chained_data_delayed_2__47_, chained_data_delayed_2__46_, chained_data_delayed_2__45_, chained_data_delayed_2__44_, chained_data_delayed_2__43_, chained_data_delayed_2__42_, chained_data_delayed_2__41_, chained_data_delayed_2__40_, chained_data_delayed_2__39_, chained_data_delayed_2__38_, chained_data_delayed_2__37_, chained_data_delayed_2__36_, chained_data_delayed_2__35_, chained_data_delayed_2__34_, chained_data_delayed_2__33_, chained_data_delayed_2__32_, chained_data_delayed_2__31_, chained_data_delayed_2__30_, chained_data_delayed_2__29_, chained_data_delayed_2__28_, chained_data_delayed_2__27_, chained_data_delayed_2__26_, chained_data_delayed_2__25_, chained_data_delayed_2__24_, chained_data_delayed_2__23_, chained_data_delayed_2__22_, chained_data_delayed_2__21_, chained_data_delayed_2__20_, chained_data_delayed_2__19_, chained_data_delayed_2__18_, chained_data_delayed_2__17_, chained_data_delayed_2__16_, chained_data_delayed_2__15_, chained_data_delayed_2__14_, chained_data_delayed_2__13_, chained_data_delayed_2__12_, chained_data_delayed_2__11_, chained_data_delayed_2__10_, chained_data_delayed_2__9_, chained_data_delayed_2__8_, chained_data_delayed_2__7_, chained_data_delayed_2__6_, chained_data_delayed_2__5_, chained_data_delayed_2__4_, chained_data_delayed_2__3_, chained_data_delayed_2__2_, chained_data_delayed_2__1_, chained_data_delayed_2__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_3__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_2__63_, chained_data_delayed_2__62_, chained_data_delayed_2__61_, chained_data_delayed_2__60_, chained_data_delayed_2__59_, chained_data_delayed_2__58_, chained_data_delayed_2__57_, chained_data_delayed_2__56_, chained_data_delayed_2__55_, chained_data_delayed_2__54_, chained_data_delayed_2__53_, chained_data_delayed_2__52_, chained_data_delayed_2__51_, chained_data_delayed_2__50_, chained_data_delayed_2__49_, chained_data_delayed_2__48_, chained_data_delayed_2__47_, chained_data_delayed_2__46_, chained_data_delayed_2__45_, chained_data_delayed_2__44_, chained_data_delayed_2__43_, chained_data_delayed_2__42_, chained_data_delayed_2__41_, chained_data_delayed_2__40_, chained_data_delayed_2__39_, chained_data_delayed_2__38_, chained_data_delayed_2__37_, chained_data_delayed_2__36_, chained_data_delayed_2__35_, chained_data_delayed_2__34_, chained_data_delayed_2__33_, chained_data_delayed_2__32_, chained_data_delayed_2__31_, chained_data_delayed_2__30_, chained_data_delayed_2__29_, chained_data_delayed_2__28_, chained_data_delayed_2__27_, chained_data_delayed_2__26_, chained_data_delayed_2__25_, chained_data_delayed_2__24_, chained_data_delayed_2__23_, chained_data_delayed_2__22_, chained_data_delayed_2__21_, chained_data_delayed_2__20_, chained_data_delayed_2__19_, chained_data_delayed_2__18_, chained_data_delayed_2__17_, chained_data_delayed_2__16_, chained_data_delayed_2__15_, chained_data_delayed_2__14_, chained_data_delayed_2__13_, chained_data_delayed_2__12_, chained_data_delayed_2__11_, chained_data_delayed_2__10_, chained_data_delayed_2__9_, chained_data_delayed_2__8_, chained_data_delayed_2__7_, chained_data_delayed_2__6_, chained_data_delayed_2__5_, chained_data_delayed_2__4_, chained_data_delayed_2__3_, chained_data_delayed_2__2_, chained_data_delayed_2__1_, chained_data_delayed_2__0_ }),
    .data_o({ chained_data_delayed_3__63_, chained_data_delayed_3__62_, chained_data_delayed_3__61_, chained_data_delayed_3__60_, chained_data_delayed_3__59_, chained_data_delayed_3__58_, chained_data_delayed_3__57_, chained_data_delayed_3__56_, chained_data_delayed_3__55_, chained_data_delayed_3__54_, chained_data_delayed_3__53_, chained_data_delayed_3__52_, chained_data_delayed_3__51_, chained_data_delayed_3__50_, chained_data_delayed_3__49_, chained_data_delayed_3__48_, chained_data_delayed_3__47_, chained_data_delayed_3__46_, chained_data_delayed_3__45_, chained_data_delayed_3__44_, chained_data_delayed_3__43_, chained_data_delayed_3__42_, chained_data_delayed_3__41_, chained_data_delayed_3__40_, chained_data_delayed_3__39_, chained_data_delayed_3__38_, chained_data_delayed_3__37_, chained_data_delayed_3__36_, chained_data_delayed_3__35_, chained_data_delayed_3__34_, chained_data_delayed_3__33_, chained_data_delayed_3__32_, chained_data_delayed_3__31_, chained_data_delayed_3__30_, chained_data_delayed_3__29_, chained_data_delayed_3__28_, chained_data_delayed_3__27_, chained_data_delayed_3__26_, chained_data_delayed_3__25_, chained_data_delayed_3__24_, chained_data_delayed_3__23_, chained_data_delayed_3__22_, chained_data_delayed_3__21_, chained_data_delayed_3__20_, chained_data_delayed_3__19_, chained_data_delayed_3__18_, chained_data_delayed_3__17_, chained_data_delayed_3__16_, chained_data_delayed_3__15_, chained_data_delayed_3__14_, chained_data_delayed_3__13_, chained_data_delayed_3__12_, chained_data_delayed_3__11_, chained_data_delayed_3__10_, chained_data_delayed_3__9_, chained_data_delayed_3__8_, chained_data_delayed_3__7_, chained_data_delayed_3__6_, chained_data_delayed_3__5_, chained_data_delayed_3__4_, chained_data_delayed_3__3_, chained_data_delayed_3__2_, chained_data_delayed_3__1_, chained_data_delayed_3__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_4__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_3__63_, chained_data_delayed_3__62_, chained_data_delayed_3__61_, chained_data_delayed_3__60_, chained_data_delayed_3__59_, chained_data_delayed_3__58_, chained_data_delayed_3__57_, chained_data_delayed_3__56_, chained_data_delayed_3__55_, chained_data_delayed_3__54_, chained_data_delayed_3__53_, chained_data_delayed_3__52_, chained_data_delayed_3__51_, chained_data_delayed_3__50_, chained_data_delayed_3__49_, chained_data_delayed_3__48_, chained_data_delayed_3__47_, chained_data_delayed_3__46_, chained_data_delayed_3__45_, chained_data_delayed_3__44_, chained_data_delayed_3__43_, chained_data_delayed_3__42_, chained_data_delayed_3__41_, chained_data_delayed_3__40_, chained_data_delayed_3__39_, chained_data_delayed_3__38_, chained_data_delayed_3__37_, chained_data_delayed_3__36_, chained_data_delayed_3__35_, chained_data_delayed_3__34_, chained_data_delayed_3__33_, chained_data_delayed_3__32_, chained_data_delayed_3__31_, chained_data_delayed_3__30_, chained_data_delayed_3__29_, chained_data_delayed_3__28_, chained_data_delayed_3__27_, chained_data_delayed_3__26_, chained_data_delayed_3__25_, chained_data_delayed_3__24_, chained_data_delayed_3__23_, chained_data_delayed_3__22_, chained_data_delayed_3__21_, chained_data_delayed_3__20_, chained_data_delayed_3__19_, chained_data_delayed_3__18_, chained_data_delayed_3__17_, chained_data_delayed_3__16_, chained_data_delayed_3__15_, chained_data_delayed_3__14_, chained_data_delayed_3__13_, chained_data_delayed_3__12_, chained_data_delayed_3__11_, chained_data_delayed_3__10_, chained_data_delayed_3__9_, chained_data_delayed_3__8_, chained_data_delayed_3__7_, chained_data_delayed_3__6_, chained_data_delayed_3__5_, chained_data_delayed_3__4_, chained_data_delayed_3__3_, chained_data_delayed_3__2_, chained_data_delayed_3__1_, chained_data_delayed_3__0_ }),
    .data_o({ chained_data_delayed_4__63_, chained_data_delayed_4__62_, chained_data_delayed_4__61_, chained_data_delayed_4__60_, chained_data_delayed_4__59_, chained_data_delayed_4__58_, chained_data_delayed_4__57_, chained_data_delayed_4__56_, chained_data_delayed_4__55_, chained_data_delayed_4__54_, chained_data_delayed_4__53_, chained_data_delayed_4__52_, chained_data_delayed_4__51_, chained_data_delayed_4__50_, chained_data_delayed_4__49_, chained_data_delayed_4__48_, chained_data_delayed_4__47_, chained_data_delayed_4__46_, chained_data_delayed_4__45_, chained_data_delayed_4__44_, chained_data_delayed_4__43_, chained_data_delayed_4__42_, chained_data_delayed_4__41_, chained_data_delayed_4__40_, chained_data_delayed_4__39_, chained_data_delayed_4__38_, chained_data_delayed_4__37_, chained_data_delayed_4__36_, chained_data_delayed_4__35_, chained_data_delayed_4__34_, chained_data_delayed_4__33_, chained_data_delayed_4__32_, chained_data_delayed_4__31_, chained_data_delayed_4__30_, chained_data_delayed_4__29_, chained_data_delayed_4__28_, chained_data_delayed_4__27_, chained_data_delayed_4__26_, chained_data_delayed_4__25_, chained_data_delayed_4__24_, chained_data_delayed_4__23_, chained_data_delayed_4__22_, chained_data_delayed_4__21_, chained_data_delayed_4__20_, chained_data_delayed_4__19_, chained_data_delayed_4__18_, chained_data_delayed_4__17_, chained_data_delayed_4__16_, chained_data_delayed_4__15_, chained_data_delayed_4__14_, chained_data_delayed_4__13_, chained_data_delayed_4__12_, chained_data_delayed_4__11_, chained_data_delayed_4__10_, chained_data_delayed_4__9_, chained_data_delayed_4__8_, chained_data_delayed_4__7_, chained_data_delayed_4__6_, chained_data_delayed_4__5_, chained_data_delayed_4__4_, chained_data_delayed_4__3_, chained_data_delayed_4__2_, chained_data_delayed_4__1_, chained_data_delayed_4__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_5__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_4__63_, chained_data_delayed_4__62_, chained_data_delayed_4__61_, chained_data_delayed_4__60_, chained_data_delayed_4__59_, chained_data_delayed_4__58_, chained_data_delayed_4__57_, chained_data_delayed_4__56_, chained_data_delayed_4__55_, chained_data_delayed_4__54_, chained_data_delayed_4__53_, chained_data_delayed_4__52_, chained_data_delayed_4__51_, chained_data_delayed_4__50_, chained_data_delayed_4__49_, chained_data_delayed_4__48_, chained_data_delayed_4__47_, chained_data_delayed_4__46_, chained_data_delayed_4__45_, chained_data_delayed_4__44_, chained_data_delayed_4__43_, chained_data_delayed_4__42_, chained_data_delayed_4__41_, chained_data_delayed_4__40_, chained_data_delayed_4__39_, chained_data_delayed_4__38_, chained_data_delayed_4__37_, chained_data_delayed_4__36_, chained_data_delayed_4__35_, chained_data_delayed_4__34_, chained_data_delayed_4__33_, chained_data_delayed_4__32_, chained_data_delayed_4__31_, chained_data_delayed_4__30_, chained_data_delayed_4__29_, chained_data_delayed_4__28_, chained_data_delayed_4__27_, chained_data_delayed_4__26_, chained_data_delayed_4__25_, chained_data_delayed_4__24_, chained_data_delayed_4__23_, chained_data_delayed_4__22_, chained_data_delayed_4__21_, chained_data_delayed_4__20_, chained_data_delayed_4__19_, chained_data_delayed_4__18_, chained_data_delayed_4__17_, chained_data_delayed_4__16_, chained_data_delayed_4__15_, chained_data_delayed_4__14_, chained_data_delayed_4__13_, chained_data_delayed_4__12_, chained_data_delayed_4__11_, chained_data_delayed_4__10_, chained_data_delayed_4__9_, chained_data_delayed_4__8_, chained_data_delayed_4__7_, chained_data_delayed_4__6_, chained_data_delayed_4__5_, chained_data_delayed_4__4_, chained_data_delayed_4__3_, chained_data_delayed_4__2_, chained_data_delayed_4__1_, chained_data_delayed_4__0_ }),
    .data_o({ chained_data_delayed_5__63_, chained_data_delayed_5__62_, chained_data_delayed_5__61_, chained_data_delayed_5__60_, chained_data_delayed_5__59_, chained_data_delayed_5__58_, chained_data_delayed_5__57_, chained_data_delayed_5__56_, chained_data_delayed_5__55_, chained_data_delayed_5__54_, chained_data_delayed_5__53_, chained_data_delayed_5__52_, chained_data_delayed_5__51_, chained_data_delayed_5__50_, chained_data_delayed_5__49_, chained_data_delayed_5__48_, chained_data_delayed_5__47_, chained_data_delayed_5__46_, chained_data_delayed_5__45_, chained_data_delayed_5__44_, chained_data_delayed_5__43_, chained_data_delayed_5__42_, chained_data_delayed_5__41_, chained_data_delayed_5__40_, chained_data_delayed_5__39_, chained_data_delayed_5__38_, chained_data_delayed_5__37_, chained_data_delayed_5__36_, chained_data_delayed_5__35_, chained_data_delayed_5__34_, chained_data_delayed_5__33_, chained_data_delayed_5__32_, chained_data_delayed_5__31_, chained_data_delayed_5__30_, chained_data_delayed_5__29_, chained_data_delayed_5__28_, chained_data_delayed_5__27_, chained_data_delayed_5__26_, chained_data_delayed_5__25_, chained_data_delayed_5__24_, chained_data_delayed_5__23_, chained_data_delayed_5__22_, chained_data_delayed_5__21_, chained_data_delayed_5__20_, chained_data_delayed_5__19_, chained_data_delayed_5__18_, chained_data_delayed_5__17_, chained_data_delayed_5__16_, chained_data_delayed_5__15_, chained_data_delayed_5__14_, chained_data_delayed_5__13_, chained_data_delayed_5__12_, chained_data_delayed_5__11_, chained_data_delayed_5__10_, chained_data_delayed_5__9_, chained_data_delayed_5__8_, chained_data_delayed_5__7_, chained_data_delayed_5__6_, chained_data_delayed_5__5_, chained_data_delayed_5__4_, chained_data_delayed_5__3_, chained_data_delayed_5__2_, chained_data_delayed_5__1_, chained_data_delayed_5__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_6__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_5__63_, chained_data_delayed_5__62_, chained_data_delayed_5__61_, chained_data_delayed_5__60_, chained_data_delayed_5__59_, chained_data_delayed_5__58_, chained_data_delayed_5__57_, chained_data_delayed_5__56_, chained_data_delayed_5__55_, chained_data_delayed_5__54_, chained_data_delayed_5__53_, chained_data_delayed_5__52_, chained_data_delayed_5__51_, chained_data_delayed_5__50_, chained_data_delayed_5__49_, chained_data_delayed_5__48_, chained_data_delayed_5__47_, chained_data_delayed_5__46_, chained_data_delayed_5__45_, chained_data_delayed_5__44_, chained_data_delayed_5__43_, chained_data_delayed_5__42_, chained_data_delayed_5__41_, chained_data_delayed_5__40_, chained_data_delayed_5__39_, chained_data_delayed_5__38_, chained_data_delayed_5__37_, chained_data_delayed_5__36_, chained_data_delayed_5__35_, chained_data_delayed_5__34_, chained_data_delayed_5__33_, chained_data_delayed_5__32_, chained_data_delayed_5__31_, chained_data_delayed_5__30_, chained_data_delayed_5__29_, chained_data_delayed_5__28_, chained_data_delayed_5__27_, chained_data_delayed_5__26_, chained_data_delayed_5__25_, chained_data_delayed_5__24_, chained_data_delayed_5__23_, chained_data_delayed_5__22_, chained_data_delayed_5__21_, chained_data_delayed_5__20_, chained_data_delayed_5__19_, chained_data_delayed_5__18_, chained_data_delayed_5__17_, chained_data_delayed_5__16_, chained_data_delayed_5__15_, chained_data_delayed_5__14_, chained_data_delayed_5__13_, chained_data_delayed_5__12_, chained_data_delayed_5__11_, chained_data_delayed_5__10_, chained_data_delayed_5__9_, chained_data_delayed_5__8_, chained_data_delayed_5__7_, chained_data_delayed_5__6_, chained_data_delayed_5__5_, chained_data_delayed_5__4_, chained_data_delayed_5__3_, chained_data_delayed_5__2_, chained_data_delayed_5__1_, chained_data_delayed_5__0_ }),
    .data_o({ chained_data_delayed_6__63_, chained_data_delayed_6__62_, chained_data_delayed_6__61_, chained_data_delayed_6__60_, chained_data_delayed_6__59_, chained_data_delayed_6__58_, chained_data_delayed_6__57_, chained_data_delayed_6__56_, chained_data_delayed_6__55_, chained_data_delayed_6__54_, chained_data_delayed_6__53_, chained_data_delayed_6__52_, chained_data_delayed_6__51_, chained_data_delayed_6__50_, chained_data_delayed_6__49_, chained_data_delayed_6__48_, chained_data_delayed_6__47_, chained_data_delayed_6__46_, chained_data_delayed_6__45_, chained_data_delayed_6__44_, chained_data_delayed_6__43_, chained_data_delayed_6__42_, chained_data_delayed_6__41_, chained_data_delayed_6__40_, chained_data_delayed_6__39_, chained_data_delayed_6__38_, chained_data_delayed_6__37_, chained_data_delayed_6__36_, chained_data_delayed_6__35_, chained_data_delayed_6__34_, chained_data_delayed_6__33_, chained_data_delayed_6__32_, chained_data_delayed_6__31_, chained_data_delayed_6__30_, chained_data_delayed_6__29_, chained_data_delayed_6__28_, chained_data_delayed_6__27_, chained_data_delayed_6__26_, chained_data_delayed_6__25_, chained_data_delayed_6__24_, chained_data_delayed_6__23_, chained_data_delayed_6__22_, chained_data_delayed_6__21_, chained_data_delayed_6__20_, chained_data_delayed_6__19_, chained_data_delayed_6__18_, chained_data_delayed_6__17_, chained_data_delayed_6__16_, chained_data_delayed_6__15_, chained_data_delayed_6__14_, chained_data_delayed_6__13_, chained_data_delayed_6__12_, chained_data_delayed_6__11_, chained_data_delayed_6__10_, chained_data_delayed_6__9_, chained_data_delayed_6__8_, chained_data_delayed_6__7_, chained_data_delayed_6__6_, chained_data_delayed_6__5_, chained_data_delayed_6__4_, chained_data_delayed_6__3_, chained_data_delayed_6__2_, chained_data_delayed_6__1_, chained_data_delayed_6__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_7__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_6__63_, chained_data_delayed_6__62_, chained_data_delayed_6__61_, chained_data_delayed_6__60_, chained_data_delayed_6__59_, chained_data_delayed_6__58_, chained_data_delayed_6__57_, chained_data_delayed_6__56_, chained_data_delayed_6__55_, chained_data_delayed_6__54_, chained_data_delayed_6__53_, chained_data_delayed_6__52_, chained_data_delayed_6__51_, chained_data_delayed_6__50_, chained_data_delayed_6__49_, chained_data_delayed_6__48_, chained_data_delayed_6__47_, chained_data_delayed_6__46_, chained_data_delayed_6__45_, chained_data_delayed_6__44_, chained_data_delayed_6__43_, chained_data_delayed_6__42_, chained_data_delayed_6__41_, chained_data_delayed_6__40_, chained_data_delayed_6__39_, chained_data_delayed_6__38_, chained_data_delayed_6__37_, chained_data_delayed_6__36_, chained_data_delayed_6__35_, chained_data_delayed_6__34_, chained_data_delayed_6__33_, chained_data_delayed_6__32_, chained_data_delayed_6__31_, chained_data_delayed_6__30_, chained_data_delayed_6__29_, chained_data_delayed_6__28_, chained_data_delayed_6__27_, chained_data_delayed_6__26_, chained_data_delayed_6__25_, chained_data_delayed_6__24_, chained_data_delayed_6__23_, chained_data_delayed_6__22_, chained_data_delayed_6__21_, chained_data_delayed_6__20_, chained_data_delayed_6__19_, chained_data_delayed_6__18_, chained_data_delayed_6__17_, chained_data_delayed_6__16_, chained_data_delayed_6__15_, chained_data_delayed_6__14_, chained_data_delayed_6__13_, chained_data_delayed_6__12_, chained_data_delayed_6__11_, chained_data_delayed_6__10_, chained_data_delayed_6__9_, chained_data_delayed_6__8_, chained_data_delayed_6__7_, chained_data_delayed_6__6_, chained_data_delayed_6__5_, chained_data_delayed_6__4_, chained_data_delayed_6__3_, chained_data_delayed_6__2_, chained_data_delayed_6__1_, chained_data_delayed_6__0_ }),
    .data_o({ chained_data_delayed_7__63_, chained_data_delayed_7__62_, chained_data_delayed_7__61_, chained_data_delayed_7__60_, chained_data_delayed_7__59_, chained_data_delayed_7__58_, chained_data_delayed_7__57_, chained_data_delayed_7__56_, chained_data_delayed_7__55_, chained_data_delayed_7__54_, chained_data_delayed_7__53_, chained_data_delayed_7__52_, chained_data_delayed_7__51_, chained_data_delayed_7__50_, chained_data_delayed_7__49_, chained_data_delayed_7__48_, chained_data_delayed_7__47_, chained_data_delayed_7__46_, chained_data_delayed_7__45_, chained_data_delayed_7__44_, chained_data_delayed_7__43_, chained_data_delayed_7__42_, chained_data_delayed_7__41_, chained_data_delayed_7__40_, chained_data_delayed_7__39_, chained_data_delayed_7__38_, chained_data_delayed_7__37_, chained_data_delayed_7__36_, chained_data_delayed_7__35_, chained_data_delayed_7__34_, chained_data_delayed_7__33_, chained_data_delayed_7__32_, chained_data_delayed_7__31_, chained_data_delayed_7__30_, chained_data_delayed_7__29_, chained_data_delayed_7__28_, chained_data_delayed_7__27_, chained_data_delayed_7__26_, chained_data_delayed_7__25_, chained_data_delayed_7__24_, chained_data_delayed_7__23_, chained_data_delayed_7__22_, chained_data_delayed_7__21_, chained_data_delayed_7__20_, chained_data_delayed_7__19_, chained_data_delayed_7__18_, chained_data_delayed_7__17_, chained_data_delayed_7__16_, chained_data_delayed_7__15_, chained_data_delayed_7__14_, chained_data_delayed_7__13_, chained_data_delayed_7__12_, chained_data_delayed_7__11_, chained_data_delayed_7__10_, chained_data_delayed_7__9_, chained_data_delayed_7__8_, chained_data_delayed_7__7_, chained_data_delayed_7__6_, chained_data_delayed_7__5_, chained_data_delayed_7__4_, chained_data_delayed_7__3_, chained_data_delayed_7__2_, chained_data_delayed_7__1_, chained_data_delayed_7__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_8__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_7__63_, chained_data_delayed_7__62_, chained_data_delayed_7__61_, chained_data_delayed_7__60_, chained_data_delayed_7__59_, chained_data_delayed_7__58_, chained_data_delayed_7__57_, chained_data_delayed_7__56_, chained_data_delayed_7__55_, chained_data_delayed_7__54_, chained_data_delayed_7__53_, chained_data_delayed_7__52_, chained_data_delayed_7__51_, chained_data_delayed_7__50_, chained_data_delayed_7__49_, chained_data_delayed_7__48_, chained_data_delayed_7__47_, chained_data_delayed_7__46_, chained_data_delayed_7__45_, chained_data_delayed_7__44_, chained_data_delayed_7__43_, chained_data_delayed_7__42_, chained_data_delayed_7__41_, chained_data_delayed_7__40_, chained_data_delayed_7__39_, chained_data_delayed_7__38_, chained_data_delayed_7__37_, chained_data_delayed_7__36_, chained_data_delayed_7__35_, chained_data_delayed_7__34_, chained_data_delayed_7__33_, chained_data_delayed_7__32_, chained_data_delayed_7__31_, chained_data_delayed_7__30_, chained_data_delayed_7__29_, chained_data_delayed_7__28_, chained_data_delayed_7__27_, chained_data_delayed_7__26_, chained_data_delayed_7__25_, chained_data_delayed_7__24_, chained_data_delayed_7__23_, chained_data_delayed_7__22_, chained_data_delayed_7__21_, chained_data_delayed_7__20_, chained_data_delayed_7__19_, chained_data_delayed_7__18_, chained_data_delayed_7__17_, chained_data_delayed_7__16_, chained_data_delayed_7__15_, chained_data_delayed_7__14_, chained_data_delayed_7__13_, chained_data_delayed_7__12_, chained_data_delayed_7__11_, chained_data_delayed_7__10_, chained_data_delayed_7__9_, chained_data_delayed_7__8_, chained_data_delayed_7__7_, chained_data_delayed_7__6_, chained_data_delayed_7__5_, chained_data_delayed_7__4_, chained_data_delayed_7__3_, chained_data_delayed_7__2_, chained_data_delayed_7__1_, chained_data_delayed_7__0_ }),
    .data_o({ chained_data_delayed_8__63_, chained_data_delayed_8__62_, chained_data_delayed_8__61_, chained_data_delayed_8__60_, chained_data_delayed_8__59_, chained_data_delayed_8__58_, chained_data_delayed_8__57_, chained_data_delayed_8__56_, chained_data_delayed_8__55_, chained_data_delayed_8__54_, chained_data_delayed_8__53_, chained_data_delayed_8__52_, chained_data_delayed_8__51_, chained_data_delayed_8__50_, chained_data_delayed_8__49_, chained_data_delayed_8__48_, chained_data_delayed_8__47_, chained_data_delayed_8__46_, chained_data_delayed_8__45_, chained_data_delayed_8__44_, chained_data_delayed_8__43_, chained_data_delayed_8__42_, chained_data_delayed_8__41_, chained_data_delayed_8__40_, chained_data_delayed_8__39_, chained_data_delayed_8__38_, chained_data_delayed_8__37_, chained_data_delayed_8__36_, chained_data_delayed_8__35_, chained_data_delayed_8__34_, chained_data_delayed_8__33_, chained_data_delayed_8__32_, chained_data_delayed_8__31_, chained_data_delayed_8__30_, chained_data_delayed_8__29_, chained_data_delayed_8__28_, chained_data_delayed_8__27_, chained_data_delayed_8__26_, chained_data_delayed_8__25_, chained_data_delayed_8__24_, chained_data_delayed_8__23_, chained_data_delayed_8__22_, chained_data_delayed_8__21_, chained_data_delayed_8__20_, chained_data_delayed_8__19_, chained_data_delayed_8__18_, chained_data_delayed_8__17_, chained_data_delayed_8__16_, chained_data_delayed_8__15_, chained_data_delayed_8__14_, chained_data_delayed_8__13_, chained_data_delayed_8__12_, chained_data_delayed_8__11_, chained_data_delayed_8__10_, chained_data_delayed_8__9_, chained_data_delayed_8__8_, chained_data_delayed_8__7_, chained_data_delayed_8__6_, chained_data_delayed_8__5_, chained_data_delayed_8__4_, chained_data_delayed_8__3_, chained_data_delayed_8__2_, chained_data_delayed_8__1_, chained_data_delayed_8__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_9__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_8__63_, chained_data_delayed_8__62_, chained_data_delayed_8__61_, chained_data_delayed_8__60_, chained_data_delayed_8__59_, chained_data_delayed_8__58_, chained_data_delayed_8__57_, chained_data_delayed_8__56_, chained_data_delayed_8__55_, chained_data_delayed_8__54_, chained_data_delayed_8__53_, chained_data_delayed_8__52_, chained_data_delayed_8__51_, chained_data_delayed_8__50_, chained_data_delayed_8__49_, chained_data_delayed_8__48_, chained_data_delayed_8__47_, chained_data_delayed_8__46_, chained_data_delayed_8__45_, chained_data_delayed_8__44_, chained_data_delayed_8__43_, chained_data_delayed_8__42_, chained_data_delayed_8__41_, chained_data_delayed_8__40_, chained_data_delayed_8__39_, chained_data_delayed_8__38_, chained_data_delayed_8__37_, chained_data_delayed_8__36_, chained_data_delayed_8__35_, chained_data_delayed_8__34_, chained_data_delayed_8__33_, chained_data_delayed_8__32_, chained_data_delayed_8__31_, chained_data_delayed_8__30_, chained_data_delayed_8__29_, chained_data_delayed_8__28_, chained_data_delayed_8__27_, chained_data_delayed_8__26_, chained_data_delayed_8__25_, chained_data_delayed_8__24_, chained_data_delayed_8__23_, chained_data_delayed_8__22_, chained_data_delayed_8__21_, chained_data_delayed_8__20_, chained_data_delayed_8__19_, chained_data_delayed_8__18_, chained_data_delayed_8__17_, chained_data_delayed_8__16_, chained_data_delayed_8__15_, chained_data_delayed_8__14_, chained_data_delayed_8__13_, chained_data_delayed_8__12_, chained_data_delayed_8__11_, chained_data_delayed_8__10_, chained_data_delayed_8__9_, chained_data_delayed_8__8_, chained_data_delayed_8__7_, chained_data_delayed_8__6_, chained_data_delayed_8__5_, chained_data_delayed_8__4_, chained_data_delayed_8__3_, chained_data_delayed_8__2_, chained_data_delayed_8__1_, chained_data_delayed_8__0_ }),
    .data_o({ chained_data_delayed_9__63_, chained_data_delayed_9__62_, chained_data_delayed_9__61_, chained_data_delayed_9__60_, chained_data_delayed_9__59_, chained_data_delayed_9__58_, chained_data_delayed_9__57_, chained_data_delayed_9__56_, chained_data_delayed_9__55_, chained_data_delayed_9__54_, chained_data_delayed_9__53_, chained_data_delayed_9__52_, chained_data_delayed_9__51_, chained_data_delayed_9__50_, chained_data_delayed_9__49_, chained_data_delayed_9__48_, chained_data_delayed_9__47_, chained_data_delayed_9__46_, chained_data_delayed_9__45_, chained_data_delayed_9__44_, chained_data_delayed_9__43_, chained_data_delayed_9__42_, chained_data_delayed_9__41_, chained_data_delayed_9__40_, chained_data_delayed_9__39_, chained_data_delayed_9__38_, chained_data_delayed_9__37_, chained_data_delayed_9__36_, chained_data_delayed_9__35_, chained_data_delayed_9__34_, chained_data_delayed_9__33_, chained_data_delayed_9__32_, chained_data_delayed_9__31_, chained_data_delayed_9__30_, chained_data_delayed_9__29_, chained_data_delayed_9__28_, chained_data_delayed_9__27_, chained_data_delayed_9__26_, chained_data_delayed_9__25_, chained_data_delayed_9__24_, chained_data_delayed_9__23_, chained_data_delayed_9__22_, chained_data_delayed_9__21_, chained_data_delayed_9__20_, chained_data_delayed_9__19_, chained_data_delayed_9__18_, chained_data_delayed_9__17_, chained_data_delayed_9__16_, chained_data_delayed_9__15_, chained_data_delayed_9__14_, chained_data_delayed_9__13_, chained_data_delayed_9__12_, chained_data_delayed_9__11_, chained_data_delayed_9__10_, chained_data_delayed_9__9_, chained_data_delayed_9__8_, chained_data_delayed_9__7_, chained_data_delayed_9__6_, chained_data_delayed_9__5_, chained_data_delayed_9__4_, chained_data_delayed_9__3_, chained_data_delayed_9__2_, chained_data_delayed_9__1_, chained_data_delayed_9__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_10__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_9__63_, chained_data_delayed_9__62_, chained_data_delayed_9__61_, chained_data_delayed_9__60_, chained_data_delayed_9__59_, chained_data_delayed_9__58_, chained_data_delayed_9__57_, chained_data_delayed_9__56_, chained_data_delayed_9__55_, chained_data_delayed_9__54_, chained_data_delayed_9__53_, chained_data_delayed_9__52_, chained_data_delayed_9__51_, chained_data_delayed_9__50_, chained_data_delayed_9__49_, chained_data_delayed_9__48_, chained_data_delayed_9__47_, chained_data_delayed_9__46_, chained_data_delayed_9__45_, chained_data_delayed_9__44_, chained_data_delayed_9__43_, chained_data_delayed_9__42_, chained_data_delayed_9__41_, chained_data_delayed_9__40_, chained_data_delayed_9__39_, chained_data_delayed_9__38_, chained_data_delayed_9__37_, chained_data_delayed_9__36_, chained_data_delayed_9__35_, chained_data_delayed_9__34_, chained_data_delayed_9__33_, chained_data_delayed_9__32_, chained_data_delayed_9__31_, chained_data_delayed_9__30_, chained_data_delayed_9__29_, chained_data_delayed_9__28_, chained_data_delayed_9__27_, chained_data_delayed_9__26_, chained_data_delayed_9__25_, chained_data_delayed_9__24_, chained_data_delayed_9__23_, chained_data_delayed_9__22_, chained_data_delayed_9__21_, chained_data_delayed_9__20_, chained_data_delayed_9__19_, chained_data_delayed_9__18_, chained_data_delayed_9__17_, chained_data_delayed_9__16_, chained_data_delayed_9__15_, chained_data_delayed_9__14_, chained_data_delayed_9__13_, chained_data_delayed_9__12_, chained_data_delayed_9__11_, chained_data_delayed_9__10_, chained_data_delayed_9__9_, chained_data_delayed_9__8_, chained_data_delayed_9__7_, chained_data_delayed_9__6_, chained_data_delayed_9__5_, chained_data_delayed_9__4_, chained_data_delayed_9__3_, chained_data_delayed_9__2_, chained_data_delayed_9__1_, chained_data_delayed_9__0_ }),
    .data_o({ chained_data_delayed_10__63_, chained_data_delayed_10__62_, chained_data_delayed_10__61_, chained_data_delayed_10__60_, chained_data_delayed_10__59_, chained_data_delayed_10__58_, chained_data_delayed_10__57_, chained_data_delayed_10__56_, chained_data_delayed_10__55_, chained_data_delayed_10__54_, chained_data_delayed_10__53_, chained_data_delayed_10__52_, chained_data_delayed_10__51_, chained_data_delayed_10__50_, chained_data_delayed_10__49_, chained_data_delayed_10__48_, chained_data_delayed_10__47_, chained_data_delayed_10__46_, chained_data_delayed_10__45_, chained_data_delayed_10__44_, chained_data_delayed_10__43_, chained_data_delayed_10__42_, chained_data_delayed_10__41_, chained_data_delayed_10__40_, chained_data_delayed_10__39_, chained_data_delayed_10__38_, chained_data_delayed_10__37_, chained_data_delayed_10__36_, chained_data_delayed_10__35_, chained_data_delayed_10__34_, chained_data_delayed_10__33_, chained_data_delayed_10__32_, chained_data_delayed_10__31_, chained_data_delayed_10__30_, chained_data_delayed_10__29_, chained_data_delayed_10__28_, chained_data_delayed_10__27_, chained_data_delayed_10__26_, chained_data_delayed_10__25_, chained_data_delayed_10__24_, chained_data_delayed_10__23_, chained_data_delayed_10__22_, chained_data_delayed_10__21_, chained_data_delayed_10__20_, chained_data_delayed_10__19_, chained_data_delayed_10__18_, chained_data_delayed_10__17_, chained_data_delayed_10__16_, chained_data_delayed_10__15_, chained_data_delayed_10__14_, chained_data_delayed_10__13_, chained_data_delayed_10__12_, chained_data_delayed_10__11_, chained_data_delayed_10__10_, chained_data_delayed_10__9_, chained_data_delayed_10__8_, chained_data_delayed_10__7_, chained_data_delayed_10__6_, chained_data_delayed_10__5_, chained_data_delayed_10__4_, chained_data_delayed_10__3_, chained_data_delayed_10__2_, chained_data_delayed_10__1_, chained_data_delayed_10__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_11__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_10__63_, chained_data_delayed_10__62_, chained_data_delayed_10__61_, chained_data_delayed_10__60_, chained_data_delayed_10__59_, chained_data_delayed_10__58_, chained_data_delayed_10__57_, chained_data_delayed_10__56_, chained_data_delayed_10__55_, chained_data_delayed_10__54_, chained_data_delayed_10__53_, chained_data_delayed_10__52_, chained_data_delayed_10__51_, chained_data_delayed_10__50_, chained_data_delayed_10__49_, chained_data_delayed_10__48_, chained_data_delayed_10__47_, chained_data_delayed_10__46_, chained_data_delayed_10__45_, chained_data_delayed_10__44_, chained_data_delayed_10__43_, chained_data_delayed_10__42_, chained_data_delayed_10__41_, chained_data_delayed_10__40_, chained_data_delayed_10__39_, chained_data_delayed_10__38_, chained_data_delayed_10__37_, chained_data_delayed_10__36_, chained_data_delayed_10__35_, chained_data_delayed_10__34_, chained_data_delayed_10__33_, chained_data_delayed_10__32_, chained_data_delayed_10__31_, chained_data_delayed_10__30_, chained_data_delayed_10__29_, chained_data_delayed_10__28_, chained_data_delayed_10__27_, chained_data_delayed_10__26_, chained_data_delayed_10__25_, chained_data_delayed_10__24_, chained_data_delayed_10__23_, chained_data_delayed_10__22_, chained_data_delayed_10__21_, chained_data_delayed_10__20_, chained_data_delayed_10__19_, chained_data_delayed_10__18_, chained_data_delayed_10__17_, chained_data_delayed_10__16_, chained_data_delayed_10__15_, chained_data_delayed_10__14_, chained_data_delayed_10__13_, chained_data_delayed_10__12_, chained_data_delayed_10__11_, chained_data_delayed_10__10_, chained_data_delayed_10__9_, chained_data_delayed_10__8_, chained_data_delayed_10__7_, chained_data_delayed_10__6_, chained_data_delayed_10__5_, chained_data_delayed_10__4_, chained_data_delayed_10__3_, chained_data_delayed_10__2_, chained_data_delayed_10__1_, chained_data_delayed_10__0_ }),
    .data_o({ chained_data_delayed_11__63_, chained_data_delayed_11__62_, chained_data_delayed_11__61_, chained_data_delayed_11__60_, chained_data_delayed_11__59_, chained_data_delayed_11__58_, chained_data_delayed_11__57_, chained_data_delayed_11__56_, chained_data_delayed_11__55_, chained_data_delayed_11__54_, chained_data_delayed_11__53_, chained_data_delayed_11__52_, chained_data_delayed_11__51_, chained_data_delayed_11__50_, chained_data_delayed_11__49_, chained_data_delayed_11__48_, chained_data_delayed_11__47_, chained_data_delayed_11__46_, chained_data_delayed_11__45_, chained_data_delayed_11__44_, chained_data_delayed_11__43_, chained_data_delayed_11__42_, chained_data_delayed_11__41_, chained_data_delayed_11__40_, chained_data_delayed_11__39_, chained_data_delayed_11__38_, chained_data_delayed_11__37_, chained_data_delayed_11__36_, chained_data_delayed_11__35_, chained_data_delayed_11__34_, chained_data_delayed_11__33_, chained_data_delayed_11__32_, chained_data_delayed_11__31_, chained_data_delayed_11__30_, chained_data_delayed_11__29_, chained_data_delayed_11__28_, chained_data_delayed_11__27_, chained_data_delayed_11__26_, chained_data_delayed_11__25_, chained_data_delayed_11__24_, chained_data_delayed_11__23_, chained_data_delayed_11__22_, chained_data_delayed_11__21_, chained_data_delayed_11__20_, chained_data_delayed_11__19_, chained_data_delayed_11__18_, chained_data_delayed_11__17_, chained_data_delayed_11__16_, chained_data_delayed_11__15_, chained_data_delayed_11__14_, chained_data_delayed_11__13_, chained_data_delayed_11__12_, chained_data_delayed_11__11_, chained_data_delayed_11__10_, chained_data_delayed_11__9_, chained_data_delayed_11__8_, chained_data_delayed_11__7_, chained_data_delayed_11__6_, chained_data_delayed_11__5_, chained_data_delayed_11__4_, chained_data_delayed_11__3_, chained_data_delayed_11__2_, chained_data_delayed_11__1_, chained_data_delayed_11__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_12__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_11__63_, chained_data_delayed_11__62_, chained_data_delayed_11__61_, chained_data_delayed_11__60_, chained_data_delayed_11__59_, chained_data_delayed_11__58_, chained_data_delayed_11__57_, chained_data_delayed_11__56_, chained_data_delayed_11__55_, chained_data_delayed_11__54_, chained_data_delayed_11__53_, chained_data_delayed_11__52_, chained_data_delayed_11__51_, chained_data_delayed_11__50_, chained_data_delayed_11__49_, chained_data_delayed_11__48_, chained_data_delayed_11__47_, chained_data_delayed_11__46_, chained_data_delayed_11__45_, chained_data_delayed_11__44_, chained_data_delayed_11__43_, chained_data_delayed_11__42_, chained_data_delayed_11__41_, chained_data_delayed_11__40_, chained_data_delayed_11__39_, chained_data_delayed_11__38_, chained_data_delayed_11__37_, chained_data_delayed_11__36_, chained_data_delayed_11__35_, chained_data_delayed_11__34_, chained_data_delayed_11__33_, chained_data_delayed_11__32_, chained_data_delayed_11__31_, chained_data_delayed_11__30_, chained_data_delayed_11__29_, chained_data_delayed_11__28_, chained_data_delayed_11__27_, chained_data_delayed_11__26_, chained_data_delayed_11__25_, chained_data_delayed_11__24_, chained_data_delayed_11__23_, chained_data_delayed_11__22_, chained_data_delayed_11__21_, chained_data_delayed_11__20_, chained_data_delayed_11__19_, chained_data_delayed_11__18_, chained_data_delayed_11__17_, chained_data_delayed_11__16_, chained_data_delayed_11__15_, chained_data_delayed_11__14_, chained_data_delayed_11__13_, chained_data_delayed_11__12_, chained_data_delayed_11__11_, chained_data_delayed_11__10_, chained_data_delayed_11__9_, chained_data_delayed_11__8_, chained_data_delayed_11__7_, chained_data_delayed_11__6_, chained_data_delayed_11__5_, chained_data_delayed_11__4_, chained_data_delayed_11__3_, chained_data_delayed_11__2_, chained_data_delayed_11__1_, chained_data_delayed_11__0_ }),
    .data_o({ chained_data_delayed_12__63_, chained_data_delayed_12__62_, chained_data_delayed_12__61_, chained_data_delayed_12__60_, chained_data_delayed_12__59_, chained_data_delayed_12__58_, chained_data_delayed_12__57_, chained_data_delayed_12__56_, chained_data_delayed_12__55_, chained_data_delayed_12__54_, chained_data_delayed_12__53_, chained_data_delayed_12__52_, chained_data_delayed_12__51_, chained_data_delayed_12__50_, chained_data_delayed_12__49_, chained_data_delayed_12__48_, chained_data_delayed_12__47_, chained_data_delayed_12__46_, chained_data_delayed_12__45_, chained_data_delayed_12__44_, chained_data_delayed_12__43_, chained_data_delayed_12__42_, chained_data_delayed_12__41_, chained_data_delayed_12__40_, chained_data_delayed_12__39_, chained_data_delayed_12__38_, chained_data_delayed_12__37_, chained_data_delayed_12__36_, chained_data_delayed_12__35_, chained_data_delayed_12__34_, chained_data_delayed_12__33_, chained_data_delayed_12__32_, chained_data_delayed_12__31_, chained_data_delayed_12__30_, chained_data_delayed_12__29_, chained_data_delayed_12__28_, chained_data_delayed_12__27_, chained_data_delayed_12__26_, chained_data_delayed_12__25_, chained_data_delayed_12__24_, chained_data_delayed_12__23_, chained_data_delayed_12__22_, chained_data_delayed_12__21_, chained_data_delayed_12__20_, chained_data_delayed_12__19_, chained_data_delayed_12__18_, chained_data_delayed_12__17_, chained_data_delayed_12__16_, chained_data_delayed_12__15_, chained_data_delayed_12__14_, chained_data_delayed_12__13_, chained_data_delayed_12__12_, chained_data_delayed_12__11_, chained_data_delayed_12__10_, chained_data_delayed_12__9_, chained_data_delayed_12__8_, chained_data_delayed_12__7_, chained_data_delayed_12__6_, chained_data_delayed_12__5_, chained_data_delayed_12__4_, chained_data_delayed_12__3_, chained_data_delayed_12__2_, chained_data_delayed_12__1_, chained_data_delayed_12__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_13__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_12__63_, chained_data_delayed_12__62_, chained_data_delayed_12__61_, chained_data_delayed_12__60_, chained_data_delayed_12__59_, chained_data_delayed_12__58_, chained_data_delayed_12__57_, chained_data_delayed_12__56_, chained_data_delayed_12__55_, chained_data_delayed_12__54_, chained_data_delayed_12__53_, chained_data_delayed_12__52_, chained_data_delayed_12__51_, chained_data_delayed_12__50_, chained_data_delayed_12__49_, chained_data_delayed_12__48_, chained_data_delayed_12__47_, chained_data_delayed_12__46_, chained_data_delayed_12__45_, chained_data_delayed_12__44_, chained_data_delayed_12__43_, chained_data_delayed_12__42_, chained_data_delayed_12__41_, chained_data_delayed_12__40_, chained_data_delayed_12__39_, chained_data_delayed_12__38_, chained_data_delayed_12__37_, chained_data_delayed_12__36_, chained_data_delayed_12__35_, chained_data_delayed_12__34_, chained_data_delayed_12__33_, chained_data_delayed_12__32_, chained_data_delayed_12__31_, chained_data_delayed_12__30_, chained_data_delayed_12__29_, chained_data_delayed_12__28_, chained_data_delayed_12__27_, chained_data_delayed_12__26_, chained_data_delayed_12__25_, chained_data_delayed_12__24_, chained_data_delayed_12__23_, chained_data_delayed_12__22_, chained_data_delayed_12__21_, chained_data_delayed_12__20_, chained_data_delayed_12__19_, chained_data_delayed_12__18_, chained_data_delayed_12__17_, chained_data_delayed_12__16_, chained_data_delayed_12__15_, chained_data_delayed_12__14_, chained_data_delayed_12__13_, chained_data_delayed_12__12_, chained_data_delayed_12__11_, chained_data_delayed_12__10_, chained_data_delayed_12__9_, chained_data_delayed_12__8_, chained_data_delayed_12__7_, chained_data_delayed_12__6_, chained_data_delayed_12__5_, chained_data_delayed_12__4_, chained_data_delayed_12__3_, chained_data_delayed_12__2_, chained_data_delayed_12__1_, chained_data_delayed_12__0_ }),
    .data_o({ chained_data_delayed_13__63_, chained_data_delayed_13__62_, chained_data_delayed_13__61_, chained_data_delayed_13__60_, chained_data_delayed_13__59_, chained_data_delayed_13__58_, chained_data_delayed_13__57_, chained_data_delayed_13__56_, chained_data_delayed_13__55_, chained_data_delayed_13__54_, chained_data_delayed_13__53_, chained_data_delayed_13__52_, chained_data_delayed_13__51_, chained_data_delayed_13__50_, chained_data_delayed_13__49_, chained_data_delayed_13__48_, chained_data_delayed_13__47_, chained_data_delayed_13__46_, chained_data_delayed_13__45_, chained_data_delayed_13__44_, chained_data_delayed_13__43_, chained_data_delayed_13__42_, chained_data_delayed_13__41_, chained_data_delayed_13__40_, chained_data_delayed_13__39_, chained_data_delayed_13__38_, chained_data_delayed_13__37_, chained_data_delayed_13__36_, chained_data_delayed_13__35_, chained_data_delayed_13__34_, chained_data_delayed_13__33_, chained_data_delayed_13__32_, chained_data_delayed_13__31_, chained_data_delayed_13__30_, chained_data_delayed_13__29_, chained_data_delayed_13__28_, chained_data_delayed_13__27_, chained_data_delayed_13__26_, chained_data_delayed_13__25_, chained_data_delayed_13__24_, chained_data_delayed_13__23_, chained_data_delayed_13__22_, chained_data_delayed_13__21_, chained_data_delayed_13__20_, chained_data_delayed_13__19_, chained_data_delayed_13__18_, chained_data_delayed_13__17_, chained_data_delayed_13__16_, chained_data_delayed_13__15_, chained_data_delayed_13__14_, chained_data_delayed_13__13_, chained_data_delayed_13__12_, chained_data_delayed_13__11_, chained_data_delayed_13__10_, chained_data_delayed_13__9_, chained_data_delayed_13__8_, chained_data_delayed_13__7_, chained_data_delayed_13__6_, chained_data_delayed_13__5_, chained_data_delayed_13__4_, chained_data_delayed_13__3_, chained_data_delayed_13__2_, chained_data_delayed_13__1_, chained_data_delayed_13__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_14__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_13__63_, chained_data_delayed_13__62_, chained_data_delayed_13__61_, chained_data_delayed_13__60_, chained_data_delayed_13__59_, chained_data_delayed_13__58_, chained_data_delayed_13__57_, chained_data_delayed_13__56_, chained_data_delayed_13__55_, chained_data_delayed_13__54_, chained_data_delayed_13__53_, chained_data_delayed_13__52_, chained_data_delayed_13__51_, chained_data_delayed_13__50_, chained_data_delayed_13__49_, chained_data_delayed_13__48_, chained_data_delayed_13__47_, chained_data_delayed_13__46_, chained_data_delayed_13__45_, chained_data_delayed_13__44_, chained_data_delayed_13__43_, chained_data_delayed_13__42_, chained_data_delayed_13__41_, chained_data_delayed_13__40_, chained_data_delayed_13__39_, chained_data_delayed_13__38_, chained_data_delayed_13__37_, chained_data_delayed_13__36_, chained_data_delayed_13__35_, chained_data_delayed_13__34_, chained_data_delayed_13__33_, chained_data_delayed_13__32_, chained_data_delayed_13__31_, chained_data_delayed_13__30_, chained_data_delayed_13__29_, chained_data_delayed_13__28_, chained_data_delayed_13__27_, chained_data_delayed_13__26_, chained_data_delayed_13__25_, chained_data_delayed_13__24_, chained_data_delayed_13__23_, chained_data_delayed_13__22_, chained_data_delayed_13__21_, chained_data_delayed_13__20_, chained_data_delayed_13__19_, chained_data_delayed_13__18_, chained_data_delayed_13__17_, chained_data_delayed_13__16_, chained_data_delayed_13__15_, chained_data_delayed_13__14_, chained_data_delayed_13__13_, chained_data_delayed_13__12_, chained_data_delayed_13__11_, chained_data_delayed_13__10_, chained_data_delayed_13__9_, chained_data_delayed_13__8_, chained_data_delayed_13__7_, chained_data_delayed_13__6_, chained_data_delayed_13__5_, chained_data_delayed_13__4_, chained_data_delayed_13__3_, chained_data_delayed_13__2_, chained_data_delayed_13__1_, chained_data_delayed_13__0_ }),
    .data_o({ chained_data_delayed_14__63_, chained_data_delayed_14__62_, chained_data_delayed_14__61_, chained_data_delayed_14__60_, chained_data_delayed_14__59_, chained_data_delayed_14__58_, chained_data_delayed_14__57_, chained_data_delayed_14__56_, chained_data_delayed_14__55_, chained_data_delayed_14__54_, chained_data_delayed_14__53_, chained_data_delayed_14__52_, chained_data_delayed_14__51_, chained_data_delayed_14__50_, chained_data_delayed_14__49_, chained_data_delayed_14__48_, chained_data_delayed_14__47_, chained_data_delayed_14__46_, chained_data_delayed_14__45_, chained_data_delayed_14__44_, chained_data_delayed_14__43_, chained_data_delayed_14__42_, chained_data_delayed_14__41_, chained_data_delayed_14__40_, chained_data_delayed_14__39_, chained_data_delayed_14__38_, chained_data_delayed_14__37_, chained_data_delayed_14__36_, chained_data_delayed_14__35_, chained_data_delayed_14__34_, chained_data_delayed_14__33_, chained_data_delayed_14__32_, chained_data_delayed_14__31_, chained_data_delayed_14__30_, chained_data_delayed_14__29_, chained_data_delayed_14__28_, chained_data_delayed_14__27_, chained_data_delayed_14__26_, chained_data_delayed_14__25_, chained_data_delayed_14__24_, chained_data_delayed_14__23_, chained_data_delayed_14__22_, chained_data_delayed_14__21_, chained_data_delayed_14__20_, chained_data_delayed_14__19_, chained_data_delayed_14__18_, chained_data_delayed_14__17_, chained_data_delayed_14__16_, chained_data_delayed_14__15_, chained_data_delayed_14__14_, chained_data_delayed_14__13_, chained_data_delayed_14__12_, chained_data_delayed_14__11_, chained_data_delayed_14__10_, chained_data_delayed_14__9_, chained_data_delayed_14__8_, chained_data_delayed_14__7_, chained_data_delayed_14__6_, chained_data_delayed_14__5_, chained_data_delayed_14__4_, chained_data_delayed_14__3_, chained_data_delayed_14__2_, chained_data_delayed_14__1_, chained_data_delayed_14__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_15__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_14__63_, chained_data_delayed_14__62_, chained_data_delayed_14__61_, chained_data_delayed_14__60_, chained_data_delayed_14__59_, chained_data_delayed_14__58_, chained_data_delayed_14__57_, chained_data_delayed_14__56_, chained_data_delayed_14__55_, chained_data_delayed_14__54_, chained_data_delayed_14__53_, chained_data_delayed_14__52_, chained_data_delayed_14__51_, chained_data_delayed_14__50_, chained_data_delayed_14__49_, chained_data_delayed_14__48_, chained_data_delayed_14__47_, chained_data_delayed_14__46_, chained_data_delayed_14__45_, chained_data_delayed_14__44_, chained_data_delayed_14__43_, chained_data_delayed_14__42_, chained_data_delayed_14__41_, chained_data_delayed_14__40_, chained_data_delayed_14__39_, chained_data_delayed_14__38_, chained_data_delayed_14__37_, chained_data_delayed_14__36_, chained_data_delayed_14__35_, chained_data_delayed_14__34_, chained_data_delayed_14__33_, chained_data_delayed_14__32_, chained_data_delayed_14__31_, chained_data_delayed_14__30_, chained_data_delayed_14__29_, chained_data_delayed_14__28_, chained_data_delayed_14__27_, chained_data_delayed_14__26_, chained_data_delayed_14__25_, chained_data_delayed_14__24_, chained_data_delayed_14__23_, chained_data_delayed_14__22_, chained_data_delayed_14__21_, chained_data_delayed_14__20_, chained_data_delayed_14__19_, chained_data_delayed_14__18_, chained_data_delayed_14__17_, chained_data_delayed_14__16_, chained_data_delayed_14__15_, chained_data_delayed_14__14_, chained_data_delayed_14__13_, chained_data_delayed_14__12_, chained_data_delayed_14__11_, chained_data_delayed_14__10_, chained_data_delayed_14__9_, chained_data_delayed_14__8_, chained_data_delayed_14__7_, chained_data_delayed_14__6_, chained_data_delayed_14__5_, chained_data_delayed_14__4_, chained_data_delayed_14__3_, chained_data_delayed_14__2_, chained_data_delayed_14__1_, chained_data_delayed_14__0_ }),
    .data_o({ chained_data_delayed_15__63_, chained_data_delayed_15__62_, chained_data_delayed_15__61_, chained_data_delayed_15__60_, chained_data_delayed_15__59_, chained_data_delayed_15__58_, chained_data_delayed_15__57_, chained_data_delayed_15__56_, chained_data_delayed_15__55_, chained_data_delayed_15__54_, chained_data_delayed_15__53_, chained_data_delayed_15__52_, chained_data_delayed_15__51_, chained_data_delayed_15__50_, chained_data_delayed_15__49_, chained_data_delayed_15__48_, chained_data_delayed_15__47_, chained_data_delayed_15__46_, chained_data_delayed_15__45_, chained_data_delayed_15__44_, chained_data_delayed_15__43_, chained_data_delayed_15__42_, chained_data_delayed_15__41_, chained_data_delayed_15__40_, chained_data_delayed_15__39_, chained_data_delayed_15__38_, chained_data_delayed_15__37_, chained_data_delayed_15__36_, chained_data_delayed_15__35_, chained_data_delayed_15__34_, chained_data_delayed_15__33_, chained_data_delayed_15__32_, chained_data_delayed_15__31_, chained_data_delayed_15__30_, chained_data_delayed_15__29_, chained_data_delayed_15__28_, chained_data_delayed_15__27_, chained_data_delayed_15__26_, chained_data_delayed_15__25_, chained_data_delayed_15__24_, chained_data_delayed_15__23_, chained_data_delayed_15__22_, chained_data_delayed_15__21_, chained_data_delayed_15__20_, chained_data_delayed_15__19_, chained_data_delayed_15__18_, chained_data_delayed_15__17_, chained_data_delayed_15__16_, chained_data_delayed_15__15_, chained_data_delayed_15__14_, chained_data_delayed_15__13_, chained_data_delayed_15__12_, chained_data_delayed_15__11_, chained_data_delayed_15__10_, chained_data_delayed_15__9_, chained_data_delayed_15__8_, chained_data_delayed_15__7_, chained_data_delayed_15__6_, chained_data_delayed_15__5_, chained_data_delayed_15__4_, chained_data_delayed_15__3_, chained_data_delayed_15__2_, chained_data_delayed_15__1_, chained_data_delayed_15__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_16__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_15__63_, chained_data_delayed_15__62_, chained_data_delayed_15__61_, chained_data_delayed_15__60_, chained_data_delayed_15__59_, chained_data_delayed_15__58_, chained_data_delayed_15__57_, chained_data_delayed_15__56_, chained_data_delayed_15__55_, chained_data_delayed_15__54_, chained_data_delayed_15__53_, chained_data_delayed_15__52_, chained_data_delayed_15__51_, chained_data_delayed_15__50_, chained_data_delayed_15__49_, chained_data_delayed_15__48_, chained_data_delayed_15__47_, chained_data_delayed_15__46_, chained_data_delayed_15__45_, chained_data_delayed_15__44_, chained_data_delayed_15__43_, chained_data_delayed_15__42_, chained_data_delayed_15__41_, chained_data_delayed_15__40_, chained_data_delayed_15__39_, chained_data_delayed_15__38_, chained_data_delayed_15__37_, chained_data_delayed_15__36_, chained_data_delayed_15__35_, chained_data_delayed_15__34_, chained_data_delayed_15__33_, chained_data_delayed_15__32_, chained_data_delayed_15__31_, chained_data_delayed_15__30_, chained_data_delayed_15__29_, chained_data_delayed_15__28_, chained_data_delayed_15__27_, chained_data_delayed_15__26_, chained_data_delayed_15__25_, chained_data_delayed_15__24_, chained_data_delayed_15__23_, chained_data_delayed_15__22_, chained_data_delayed_15__21_, chained_data_delayed_15__20_, chained_data_delayed_15__19_, chained_data_delayed_15__18_, chained_data_delayed_15__17_, chained_data_delayed_15__16_, chained_data_delayed_15__15_, chained_data_delayed_15__14_, chained_data_delayed_15__13_, chained_data_delayed_15__12_, chained_data_delayed_15__11_, chained_data_delayed_15__10_, chained_data_delayed_15__9_, chained_data_delayed_15__8_, chained_data_delayed_15__7_, chained_data_delayed_15__6_, chained_data_delayed_15__5_, chained_data_delayed_15__4_, chained_data_delayed_15__3_, chained_data_delayed_15__2_, chained_data_delayed_15__1_, chained_data_delayed_15__0_ }),
    .data_o({ chained_data_delayed_16__63_, chained_data_delayed_16__62_, chained_data_delayed_16__61_, chained_data_delayed_16__60_, chained_data_delayed_16__59_, chained_data_delayed_16__58_, chained_data_delayed_16__57_, chained_data_delayed_16__56_, chained_data_delayed_16__55_, chained_data_delayed_16__54_, chained_data_delayed_16__53_, chained_data_delayed_16__52_, chained_data_delayed_16__51_, chained_data_delayed_16__50_, chained_data_delayed_16__49_, chained_data_delayed_16__48_, chained_data_delayed_16__47_, chained_data_delayed_16__46_, chained_data_delayed_16__45_, chained_data_delayed_16__44_, chained_data_delayed_16__43_, chained_data_delayed_16__42_, chained_data_delayed_16__41_, chained_data_delayed_16__40_, chained_data_delayed_16__39_, chained_data_delayed_16__38_, chained_data_delayed_16__37_, chained_data_delayed_16__36_, chained_data_delayed_16__35_, chained_data_delayed_16__34_, chained_data_delayed_16__33_, chained_data_delayed_16__32_, chained_data_delayed_16__31_, chained_data_delayed_16__30_, chained_data_delayed_16__29_, chained_data_delayed_16__28_, chained_data_delayed_16__27_, chained_data_delayed_16__26_, chained_data_delayed_16__25_, chained_data_delayed_16__24_, chained_data_delayed_16__23_, chained_data_delayed_16__22_, chained_data_delayed_16__21_, chained_data_delayed_16__20_, chained_data_delayed_16__19_, chained_data_delayed_16__18_, chained_data_delayed_16__17_, chained_data_delayed_16__16_, chained_data_delayed_16__15_, chained_data_delayed_16__14_, chained_data_delayed_16__13_, chained_data_delayed_16__12_, chained_data_delayed_16__11_, chained_data_delayed_16__10_, chained_data_delayed_16__9_, chained_data_delayed_16__8_, chained_data_delayed_16__7_, chained_data_delayed_16__6_, chained_data_delayed_16__5_, chained_data_delayed_16__4_, chained_data_delayed_16__3_, chained_data_delayed_16__2_, chained_data_delayed_16__1_, chained_data_delayed_16__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_17__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_16__63_, chained_data_delayed_16__62_, chained_data_delayed_16__61_, chained_data_delayed_16__60_, chained_data_delayed_16__59_, chained_data_delayed_16__58_, chained_data_delayed_16__57_, chained_data_delayed_16__56_, chained_data_delayed_16__55_, chained_data_delayed_16__54_, chained_data_delayed_16__53_, chained_data_delayed_16__52_, chained_data_delayed_16__51_, chained_data_delayed_16__50_, chained_data_delayed_16__49_, chained_data_delayed_16__48_, chained_data_delayed_16__47_, chained_data_delayed_16__46_, chained_data_delayed_16__45_, chained_data_delayed_16__44_, chained_data_delayed_16__43_, chained_data_delayed_16__42_, chained_data_delayed_16__41_, chained_data_delayed_16__40_, chained_data_delayed_16__39_, chained_data_delayed_16__38_, chained_data_delayed_16__37_, chained_data_delayed_16__36_, chained_data_delayed_16__35_, chained_data_delayed_16__34_, chained_data_delayed_16__33_, chained_data_delayed_16__32_, chained_data_delayed_16__31_, chained_data_delayed_16__30_, chained_data_delayed_16__29_, chained_data_delayed_16__28_, chained_data_delayed_16__27_, chained_data_delayed_16__26_, chained_data_delayed_16__25_, chained_data_delayed_16__24_, chained_data_delayed_16__23_, chained_data_delayed_16__22_, chained_data_delayed_16__21_, chained_data_delayed_16__20_, chained_data_delayed_16__19_, chained_data_delayed_16__18_, chained_data_delayed_16__17_, chained_data_delayed_16__16_, chained_data_delayed_16__15_, chained_data_delayed_16__14_, chained_data_delayed_16__13_, chained_data_delayed_16__12_, chained_data_delayed_16__11_, chained_data_delayed_16__10_, chained_data_delayed_16__9_, chained_data_delayed_16__8_, chained_data_delayed_16__7_, chained_data_delayed_16__6_, chained_data_delayed_16__5_, chained_data_delayed_16__4_, chained_data_delayed_16__3_, chained_data_delayed_16__2_, chained_data_delayed_16__1_, chained_data_delayed_16__0_ }),
    .data_o({ chained_data_delayed_17__63_, chained_data_delayed_17__62_, chained_data_delayed_17__61_, chained_data_delayed_17__60_, chained_data_delayed_17__59_, chained_data_delayed_17__58_, chained_data_delayed_17__57_, chained_data_delayed_17__56_, chained_data_delayed_17__55_, chained_data_delayed_17__54_, chained_data_delayed_17__53_, chained_data_delayed_17__52_, chained_data_delayed_17__51_, chained_data_delayed_17__50_, chained_data_delayed_17__49_, chained_data_delayed_17__48_, chained_data_delayed_17__47_, chained_data_delayed_17__46_, chained_data_delayed_17__45_, chained_data_delayed_17__44_, chained_data_delayed_17__43_, chained_data_delayed_17__42_, chained_data_delayed_17__41_, chained_data_delayed_17__40_, chained_data_delayed_17__39_, chained_data_delayed_17__38_, chained_data_delayed_17__37_, chained_data_delayed_17__36_, chained_data_delayed_17__35_, chained_data_delayed_17__34_, chained_data_delayed_17__33_, chained_data_delayed_17__32_, chained_data_delayed_17__31_, chained_data_delayed_17__30_, chained_data_delayed_17__29_, chained_data_delayed_17__28_, chained_data_delayed_17__27_, chained_data_delayed_17__26_, chained_data_delayed_17__25_, chained_data_delayed_17__24_, chained_data_delayed_17__23_, chained_data_delayed_17__22_, chained_data_delayed_17__21_, chained_data_delayed_17__20_, chained_data_delayed_17__19_, chained_data_delayed_17__18_, chained_data_delayed_17__17_, chained_data_delayed_17__16_, chained_data_delayed_17__15_, chained_data_delayed_17__14_, chained_data_delayed_17__13_, chained_data_delayed_17__12_, chained_data_delayed_17__11_, chained_data_delayed_17__10_, chained_data_delayed_17__9_, chained_data_delayed_17__8_, chained_data_delayed_17__7_, chained_data_delayed_17__6_, chained_data_delayed_17__5_, chained_data_delayed_17__4_, chained_data_delayed_17__3_, chained_data_delayed_17__2_, chained_data_delayed_17__1_, chained_data_delayed_17__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_18__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_17__63_, chained_data_delayed_17__62_, chained_data_delayed_17__61_, chained_data_delayed_17__60_, chained_data_delayed_17__59_, chained_data_delayed_17__58_, chained_data_delayed_17__57_, chained_data_delayed_17__56_, chained_data_delayed_17__55_, chained_data_delayed_17__54_, chained_data_delayed_17__53_, chained_data_delayed_17__52_, chained_data_delayed_17__51_, chained_data_delayed_17__50_, chained_data_delayed_17__49_, chained_data_delayed_17__48_, chained_data_delayed_17__47_, chained_data_delayed_17__46_, chained_data_delayed_17__45_, chained_data_delayed_17__44_, chained_data_delayed_17__43_, chained_data_delayed_17__42_, chained_data_delayed_17__41_, chained_data_delayed_17__40_, chained_data_delayed_17__39_, chained_data_delayed_17__38_, chained_data_delayed_17__37_, chained_data_delayed_17__36_, chained_data_delayed_17__35_, chained_data_delayed_17__34_, chained_data_delayed_17__33_, chained_data_delayed_17__32_, chained_data_delayed_17__31_, chained_data_delayed_17__30_, chained_data_delayed_17__29_, chained_data_delayed_17__28_, chained_data_delayed_17__27_, chained_data_delayed_17__26_, chained_data_delayed_17__25_, chained_data_delayed_17__24_, chained_data_delayed_17__23_, chained_data_delayed_17__22_, chained_data_delayed_17__21_, chained_data_delayed_17__20_, chained_data_delayed_17__19_, chained_data_delayed_17__18_, chained_data_delayed_17__17_, chained_data_delayed_17__16_, chained_data_delayed_17__15_, chained_data_delayed_17__14_, chained_data_delayed_17__13_, chained_data_delayed_17__12_, chained_data_delayed_17__11_, chained_data_delayed_17__10_, chained_data_delayed_17__9_, chained_data_delayed_17__8_, chained_data_delayed_17__7_, chained_data_delayed_17__6_, chained_data_delayed_17__5_, chained_data_delayed_17__4_, chained_data_delayed_17__3_, chained_data_delayed_17__2_, chained_data_delayed_17__1_, chained_data_delayed_17__0_ }),
    .data_o({ chained_data_delayed_18__63_, chained_data_delayed_18__62_, chained_data_delayed_18__61_, chained_data_delayed_18__60_, chained_data_delayed_18__59_, chained_data_delayed_18__58_, chained_data_delayed_18__57_, chained_data_delayed_18__56_, chained_data_delayed_18__55_, chained_data_delayed_18__54_, chained_data_delayed_18__53_, chained_data_delayed_18__52_, chained_data_delayed_18__51_, chained_data_delayed_18__50_, chained_data_delayed_18__49_, chained_data_delayed_18__48_, chained_data_delayed_18__47_, chained_data_delayed_18__46_, chained_data_delayed_18__45_, chained_data_delayed_18__44_, chained_data_delayed_18__43_, chained_data_delayed_18__42_, chained_data_delayed_18__41_, chained_data_delayed_18__40_, chained_data_delayed_18__39_, chained_data_delayed_18__38_, chained_data_delayed_18__37_, chained_data_delayed_18__36_, chained_data_delayed_18__35_, chained_data_delayed_18__34_, chained_data_delayed_18__33_, chained_data_delayed_18__32_, chained_data_delayed_18__31_, chained_data_delayed_18__30_, chained_data_delayed_18__29_, chained_data_delayed_18__28_, chained_data_delayed_18__27_, chained_data_delayed_18__26_, chained_data_delayed_18__25_, chained_data_delayed_18__24_, chained_data_delayed_18__23_, chained_data_delayed_18__22_, chained_data_delayed_18__21_, chained_data_delayed_18__20_, chained_data_delayed_18__19_, chained_data_delayed_18__18_, chained_data_delayed_18__17_, chained_data_delayed_18__16_, chained_data_delayed_18__15_, chained_data_delayed_18__14_, chained_data_delayed_18__13_, chained_data_delayed_18__12_, chained_data_delayed_18__11_, chained_data_delayed_18__10_, chained_data_delayed_18__9_, chained_data_delayed_18__8_, chained_data_delayed_18__7_, chained_data_delayed_18__6_, chained_data_delayed_18__5_, chained_data_delayed_18__4_, chained_data_delayed_18__3_, chained_data_delayed_18__2_, chained_data_delayed_18__1_, chained_data_delayed_18__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_19__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_18__63_, chained_data_delayed_18__62_, chained_data_delayed_18__61_, chained_data_delayed_18__60_, chained_data_delayed_18__59_, chained_data_delayed_18__58_, chained_data_delayed_18__57_, chained_data_delayed_18__56_, chained_data_delayed_18__55_, chained_data_delayed_18__54_, chained_data_delayed_18__53_, chained_data_delayed_18__52_, chained_data_delayed_18__51_, chained_data_delayed_18__50_, chained_data_delayed_18__49_, chained_data_delayed_18__48_, chained_data_delayed_18__47_, chained_data_delayed_18__46_, chained_data_delayed_18__45_, chained_data_delayed_18__44_, chained_data_delayed_18__43_, chained_data_delayed_18__42_, chained_data_delayed_18__41_, chained_data_delayed_18__40_, chained_data_delayed_18__39_, chained_data_delayed_18__38_, chained_data_delayed_18__37_, chained_data_delayed_18__36_, chained_data_delayed_18__35_, chained_data_delayed_18__34_, chained_data_delayed_18__33_, chained_data_delayed_18__32_, chained_data_delayed_18__31_, chained_data_delayed_18__30_, chained_data_delayed_18__29_, chained_data_delayed_18__28_, chained_data_delayed_18__27_, chained_data_delayed_18__26_, chained_data_delayed_18__25_, chained_data_delayed_18__24_, chained_data_delayed_18__23_, chained_data_delayed_18__22_, chained_data_delayed_18__21_, chained_data_delayed_18__20_, chained_data_delayed_18__19_, chained_data_delayed_18__18_, chained_data_delayed_18__17_, chained_data_delayed_18__16_, chained_data_delayed_18__15_, chained_data_delayed_18__14_, chained_data_delayed_18__13_, chained_data_delayed_18__12_, chained_data_delayed_18__11_, chained_data_delayed_18__10_, chained_data_delayed_18__9_, chained_data_delayed_18__8_, chained_data_delayed_18__7_, chained_data_delayed_18__6_, chained_data_delayed_18__5_, chained_data_delayed_18__4_, chained_data_delayed_18__3_, chained_data_delayed_18__2_, chained_data_delayed_18__1_, chained_data_delayed_18__0_ }),
    .data_o({ chained_data_delayed_19__63_, chained_data_delayed_19__62_, chained_data_delayed_19__61_, chained_data_delayed_19__60_, chained_data_delayed_19__59_, chained_data_delayed_19__58_, chained_data_delayed_19__57_, chained_data_delayed_19__56_, chained_data_delayed_19__55_, chained_data_delayed_19__54_, chained_data_delayed_19__53_, chained_data_delayed_19__52_, chained_data_delayed_19__51_, chained_data_delayed_19__50_, chained_data_delayed_19__49_, chained_data_delayed_19__48_, chained_data_delayed_19__47_, chained_data_delayed_19__46_, chained_data_delayed_19__45_, chained_data_delayed_19__44_, chained_data_delayed_19__43_, chained_data_delayed_19__42_, chained_data_delayed_19__41_, chained_data_delayed_19__40_, chained_data_delayed_19__39_, chained_data_delayed_19__38_, chained_data_delayed_19__37_, chained_data_delayed_19__36_, chained_data_delayed_19__35_, chained_data_delayed_19__34_, chained_data_delayed_19__33_, chained_data_delayed_19__32_, chained_data_delayed_19__31_, chained_data_delayed_19__30_, chained_data_delayed_19__29_, chained_data_delayed_19__28_, chained_data_delayed_19__27_, chained_data_delayed_19__26_, chained_data_delayed_19__25_, chained_data_delayed_19__24_, chained_data_delayed_19__23_, chained_data_delayed_19__22_, chained_data_delayed_19__21_, chained_data_delayed_19__20_, chained_data_delayed_19__19_, chained_data_delayed_19__18_, chained_data_delayed_19__17_, chained_data_delayed_19__16_, chained_data_delayed_19__15_, chained_data_delayed_19__14_, chained_data_delayed_19__13_, chained_data_delayed_19__12_, chained_data_delayed_19__11_, chained_data_delayed_19__10_, chained_data_delayed_19__9_, chained_data_delayed_19__8_, chained_data_delayed_19__7_, chained_data_delayed_19__6_, chained_data_delayed_19__5_, chained_data_delayed_19__4_, chained_data_delayed_19__3_, chained_data_delayed_19__2_, chained_data_delayed_19__1_, chained_data_delayed_19__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_20__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_19__63_, chained_data_delayed_19__62_, chained_data_delayed_19__61_, chained_data_delayed_19__60_, chained_data_delayed_19__59_, chained_data_delayed_19__58_, chained_data_delayed_19__57_, chained_data_delayed_19__56_, chained_data_delayed_19__55_, chained_data_delayed_19__54_, chained_data_delayed_19__53_, chained_data_delayed_19__52_, chained_data_delayed_19__51_, chained_data_delayed_19__50_, chained_data_delayed_19__49_, chained_data_delayed_19__48_, chained_data_delayed_19__47_, chained_data_delayed_19__46_, chained_data_delayed_19__45_, chained_data_delayed_19__44_, chained_data_delayed_19__43_, chained_data_delayed_19__42_, chained_data_delayed_19__41_, chained_data_delayed_19__40_, chained_data_delayed_19__39_, chained_data_delayed_19__38_, chained_data_delayed_19__37_, chained_data_delayed_19__36_, chained_data_delayed_19__35_, chained_data_delayed_19__34_, chained_data_delayed_19__33_, chained_data_delayed_19__32_, chained_data_delayed_19__31_, chained_data_delayed_19__30_, chained_data_delayed_19__29_, chained_data_delayed_19__28_, chained_data_delayed_19__27_, chained_data_delayed_19__26_, chained_data_delayed_19__25_, chained_data_delayed_19__24_, chained_data_delayed_19__23_, chained_data_delayed_19__22_, chained_data_delayed_19__21_, chained_data_delayed_19__20_, chained_data_delayed_19__19_, chained_data_delayed_19__18_, chained_data_delayed_19__17_, chained_data_delayed_19__16_, chained_data_delayed_19__15_, chained_data_delayed_19__14_, chained_data_delayed_19__13_, chained_data_delayed_19__12_, chained_data_delayed_19__11_, chained_data_delayed_19__10_, chained_data_delayed_19__9_, chained_data_delayed_19__8_, chained_data_delayed_19__7_, chained_data_delayed_19__6_, chained_data_delayed_19__5_, chained_data_delayed_19__4_, chained_data_delayed_19__3_, chained_data_delayed_19__2_, chained_data_delayed_19__1_, chained_data_delayed_19__0_ }),
    .data_o({ chained_data_delayed_20__63_, chained_data_delayed_20__62_, chained_data_delayed_20__61_, chained_data_delayed_20__60_, chained_data_delayed_20__59_, chained_data_delayed_20__58_, chained_data_delayed_20__57_, chained_data_delayed_20__56_, chained_data_delayed_20__55_, chained_data_delayed_20__54_, chained_data_delayed_20__53_, chained_data_delayed_20__52_, chained_data_delayed_20__51_, chained_data_delayed_20__50_, chained_data_delayed_20__49_, chained_data_delayed_20__48_, chained_data_delayed_20__47_, chained_data_delayed_20__46_, chained_data_delayed_20__45_, chained_data_delayed_20__44_, chained_data_delayed_20__43_, chained_data_delayed_20__42_, chained_data_delayed_20__41_, chained_data_delayed_20__40_, chained_data_delayed_20__39_, chained_data_delayed_20__38_, chained_data_delayed_20__37_, chained_data_delayed_20__36_, chained_data_delayed_20__35_, chained_data_delayed_20__34_, chained_data_delayed_20__33_, chained_data_delayed_20__32_, chained_data_delayed_20__31_, chained_data_delayed_20__30_, chained_data_delayed_20__29_, chained_data_delayed_20__28_, chained_data_delayed_20__27_, chained_data_delayed_20__26_, chained_data_delayed_20__25_, chained_data_delayed_20__24_, chained_data_delayed_20__23_, chained_data_delayed_20__22_, chained_data_delayed_20__21_, chained_data_delayed_20__20_, chained_data_delayed_20__19_, chained_data_delayed_20__18_, chained_data_delayed_20__17_, chained_data_delayed_20__16_, chained_data_delayed_20__15_, chained_data_delayed_20__14_, chained_data_delayed_20__13_, chained_data_delayed_20__12_, chained_data_delayed_20__11_, chained_data_delayed_20__10_, chained_data_delayed_20__9_, chained_data_delayed_20__8_, chained_data_delayed_20__7_, chained_data_delayed_20__6_, chained_data_delayed_20__5_, chained_data_delayed_20__4_, chained_data_delayed_20__3_, chained_data_delayed_20__2_, chained_data_delayed_20__1_, chained_data_delayed_20__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_21__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_20__63_, chained_data_delayed_20__62_, chained_data_delayed_20__61_, chained_data_delayed_20__60_, chained_data_delayed_20__59_, chained_data_delayed_20__58_, chained_data_delayed_20__57_, chained_data_delayed_20__56_, chained_data_delayed_20__55_, chained_data_delayed_20__54_, chained_data_delayed_20__53_, chained_data_delayed_20__52_, chained_data_delayed_20__51_, chained_data_delayed_20__50_, chained_data_delayed_20__49_, chained_data_delayed_20__48_, chained_data_delayed_20__47_, chained_data_delayed_20__46_, chained_data_delayed_20__45_, chained_data_delayed_20__44_, chained_data_delayed_20__43_, chained_data_delayed_20__42_, chained_data_delayed_20__41_, chained_data_delayed_20__40_, chained_data_delayed_20__39_, chained_data_delayed_20__38_, chained_data_delayed_20__37_, chained_data_delayed_20__36_, chained_data_delayed_20__35_, chained_data_delayed_20__34_, chained_data_delayed_20__33_, chained_data_delayed_20__32_, chained_data_delayed_20__31_, chained_data_delayed_20__30_, chained_data_delayed_20__29_, chained_data_delayed_20__28_, chained_data_delayed_20__27_, chained_data_delayed_20__26_, chained_data_delayed_20__25_, chained_data_delayed_20__24_, chained_data_delayed_20__23_, chained_data_delayed_20__22_, chained_data_delayed_20__21_, chained_data_delayed_20__20_, chained_data_delayed_20__19_, chained_data_delayed_20__18_, chained_data_delayed_20__17_, chained_data_delayed_20__16_, chained_data_delayed_20__15_, chained_data_delayed_20__14_, chained_data_delayed_20__13_, chained_data_delayed_20__12_, chained_data_delayed_20__11_, chained_data_delayed_20__10_, chained_data_delayed_20__9_, chained_data_delayed_20__8_, chained_data_delayed_20__7_, chained_data_delayed_20__6_, chained_data_delayed_20__5_, chained_data_delayed_20__4_, chained_data_delayed_20__3_, chained_data_delayed_20__2_, chained_data_delayed_20__1_, chained_data_delayed_20__0_ }),
    .data_o({ chained_data_delayed_21__63_, chained_data_delayed_21__62_, chained_data_delayed_21__61_, chained_data_delayed_21__60_, chained_data_delayed_21__59_, chained_data_delayed_21__58_, chained_data_delayed_21__57_, chained_data_delayed_21__56_, chained_data_delayed_21__55_, chained_data_delayed_21__54_, chained_data_delayed_21__53_, chained_data_delayed_21__52_, chained_data_delayed_21__51_, chained_data_delayed_21__50_, chained_data_delayed_21__49_, chained_data_delayed_21__48_, chained_data_delayed_21__47_, chained_data_delayed_21__46_, chained_data_delayed_21__45_, chained_data_delayed_21__44_, chained_data_delayed_21__43_, chained_data_delayed_21__42_, chained_data_delayed_21__41_, chained_data_delayed_21__40_, chained_data_delayed_21__39_, chained_data_delayed_21__38_, chained_data_delayed_21__37_, chained_data_delayed_21__36_, chained_data_delayed_21__35_, chained_data_delayed_21__34_, chained_data_delayed_21__33_, chained_data_delayed_21__32_, chained_data_delayed_21__31_, chained_data_delayed_21__30_, chained_data_delayed_21__29_, chained_data_delayed_21__28_, chained_data_delayed_21__27_, chained_data_delayed_21__26_, chained_data_delayed_21__25_, chained_data_delayed_21__24_, chained_data_delayed_21__23_, chained_data_delayed_21__22_, chained_data_delayed_21__21_, chained_data_delayed_21__20_, chained_data_delayed_21__19_, chained_data_delayed_21__18_, chained_data_delayed_21__17_, chained_data_delayed_21__16_, chained_data_delayed_21__15_, chained_data_delayed_21__14_, chained_data_delayed_21__13_, chained_data_delayed_21__12_, chained_data_delayed_21__11_, chained_data_delayed_21__10_, chained_data_delayed_21__9_, chained_data_delayed_21__8_, chained_data_delayed_21__7_, chained_data_delayed_21__6_, chained_data_delayed_21__5_, chained_data_delayed_21__4_, chained_data_delayed_21__3_, chained_data_delayed_21__2_, chained_data_delayed_21__1_, chained_data_delayed_21__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_22__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_21__63_, chained_data_delayed_21__62_, chained_data_delayed_21__61_, chained_data_delayed_21__60_, chained_data_delayed_21__59_, chained_data_delayed_21__58_, chained_data_delayed_21__57_, chained_data_delayed_21__56_, chained_data_delayed_21__55_, chained_data_delayed_21__54_, chained_data_delayed_21__53_, chained_data_delayed_21__52_, chained_data_delayed_21__51_, chained_data_delayed_21__50_, chained_data_delayed_21__49_, chained_data_delayed_21__48_, chained_data_delayed_21__47_, chained_data_delayed_21__46_, chained_data_delayed_21__45_, chained_data_delayed_21__44_, chained_data_delayed_21__43_, chained_data_delayed_21__42_, chained_data_delayed_21__41_, chained_data_delayed_21__40_, chained_data_delayed_21__39_, chained_data_delayed_21__38_, chained_data_delayed_21__37_, chained_data_delayed_21__36_, chained_data_delayed_21__35_, chained_data_delayed_21__34_, chained_data_delayed_21__33_, chained_data_delayed_21__32_, chained_data_delayed_21__31_, chained_data_delayed_21__30_, chained_data_delayed_21__29_, chained_data_delayed_21__28_, chained_data_delayed_21__27_, chained_data_delayed_21__26_, chained_data_delayed_21__25_, chained_data_delayed_21__24_, chained_data_delayed_21__23_, chained_data_delayed_21__22_, chained_data_delayed_21__21_, chained_data_delayed_21__20_, chained_data_delayed_21__19_, chained_data_delayed_21__18_, chained_data_delayed_21__17_, chained_data_delayed_21__16_, chained_data_delayed_21__15_, chained_data_delayed_21__14_, chained_data_delayed_21__13_, chained_data_delayed_21__12_, chained_data_delayed_21__11_, chained_data_delayed_21__10_, chained_data_delayed_21__9_, chained_data_delayed_21__8_, chained_data_delayed_21__7_, chained_data_delayed_21__6_, chained_data_delayed_21__5_, chained_data_delayed_21__4_, chained_data_delayed_21__3_, chained_data_delayed_21__2_, chained_data_delayed_21__1_, chained_data_delayed_21__0_ }),
    .data_o({ chained_data_delayed_22__63_, chained_data_delayed_22__62_, chained_data_delayed_22__61_, chained_data_delayed_22__60_, chained_data_delayed_22__59_, chained_data_delayed_22__58_, chained_data_delayed_22__57_, chained_data_delayed_22__56_, chained_data_delayed_22__55_, chained_data_delayed_22__54_, chained_data_delayed_22__53_, chained_data_delayed_22__52_, chained_data_delayed_22__51_, chained_data_delayed_22__50_, chained_data_delayed_22__49_, chained_data_delayed_22__48_, chained_data_delayed_22__47_, chained_data_delayed_22__46_, chained_data_delayed_22__45_, chained_data_delayed_22__44_, chained_data_delayed_22__43_, chained_data_delayed_22__42_, chained_data_delayed_22__41_, chained_data_delayed_22__40_, chained_data_delayed_22__39_, chained_data_delayed_22__38_, chained_data_delayed_22__37_, chained_data_delayed_22__36_, chained_data_delayed_22__35_, chained_data_delayed_22__34_, chained_data_delayed_22__33_, chained_data_delayed_22__32_, chained_data_delayed_22__31_, chained_data_delayed_22__30_, chained_data_delayed_22__29_, chained_data_delayed_22__28_, chained_data_delayed_22__27_, chained_data_delayed_22__26_, chained_data_delayed_22__25_, chained_data_delayed_22__24_, chained_data_delayed_22__23_, chained_data_delayed_22__22_, chained_data_delayed_22__21_, chained_data_delayed_22__20_, chained_data_delayed_22__19_, chained_data_delayed_22__18_, chained_data_delayed_22__17_, chained_data_delayed_22__16_, chained_data_delayed_22__15_, chained_data_delayed_22__14_, chained_data_delayed_22__13_, chained_data_delayed_22__12_, chained_data_delayed_22__11_, chained_data_delayed_22__10_, chained_data_delayed_22__9_, chained_data_delayed_22__8_, chained_data_delayed_22__7_, chained_data_delayed_22__6_, chained_data_delayed_22__5_, chained_data_delayed_22__4_, chained_data_delayed_22__3_, chained_data_delayed_22__2_, chained_data_delayed_22__1_, chained_data_delayed_22__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_23__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_22__63_, chained_data_delayed_22__62_, chained_data_delayed_22__61_, chained_data_delayed_22__60_, chained_data_delayed_22__59_, chained_data_delayed_22__58_, chained_data_delayed_22__57_, chained_data_delayed_22__56_, chained_data_delayed_22__55_, chained_data_delayed_22__54_, chained_data_delayed_22__53_, chained_data_delayed_22__52_, chained_data_delayed_22__51_, chained_data_delayed_22__50_, chained_data_delayed_22__49_, chained_data_delayed_22__48_, chained_data_delayed_22__47_, chained_data_delayed_22__46_, chained_data_delayed_22__45_, chained_data_delayed_22__44_, chained_data_delayed_22__43_, chained_data_delayed_22__42_, chained_data_delayed_22__41_, chained_data_delayed_22__40_, chained_data_delayed_22__39_, chained_data_delayed_22__38_, chained_data_delayed_22__37_, chained_data_delayed_22__36_, chained_data_delayed_22__35_, chained_data_delayed_22__34_, chained_data_delayed_22__33_, chained_data_delayed_22__32_, chained_data_delayed_22__31_, chained_data_delayed_22__30_, chained_data_delayed_22__29_, chained_data_delayed_22__28_, chained_data_delayed_22__27_, chained_data_delayed_22__26_, chained_data_delayed_22__25_, chained_data_delayed_22__24_, chained_data_delayed_22__23_, chained_data_delayed_22__22_, chained_data_delayed_22__21_, chained_data_delayed_22__20_, chained_data_delayed_22__19_, chained_data_delayed_22__18_, chained_data_delayed_22__17_, chained_data_delayed_22__16_, chained_data_delayed_22__15_, chained_data_delayed_22__14_, chained_data_delayed_22__13_, chained_data_delayed_22__12_, chained_data_delayed_22__11_, chained_data_delayed_22__10_, chained_data_delayed_22__9_, chained_data_delayed_22__8_, chained_data_delayed_22__7_, chained_data_delayed_22__6_, chained_data_delayed_22__5_, chained_data_delayed_22__4_, chained_data_delayed_22__3_, chained_data_delayed_22__2_, chained_data_delayed_22__1_, chained_data_delayed_22__0_ }),
    .data_o({ chained_data_delayed_23__63_, chained_data_delayed_23__62_, chained_data_delayed_23__61_, chained_data_delayed_23__60_, chained_data_delayed_23__59_, chained_data_delayed_23__58_, chained_data_delayed_23__57_, chained_data_delayed_23__56_, chained_data_delayed_23__55_, chained_data_delayed_23__54_, chained_data_delayed_23__53_, chained_data_delayed_23__52_, chained_data_delayed_23__51_, chained_data_delayed_23__50_, chained_data_delayed_23__49_, chained_data_delayed_23__48_, chained_data_delayed_23__47_, chained_data_delayed_23__46_, chained_data_delayed_23__45_, chained_data_delayed_23__44_, chained_data_delayed_23__43_, chained_data_delayed_23__42_, chained_data_delayed_23__41_, chained_data_delayed_23__40_, chained_data_delayed_23__39_, chained_data_delayed_23__38_, chained_data_delayed_23__37_, chained_data_delayed_23__36_, chained_data_delayed_23__35_, chained_data_delayed_23__34_, chained_data_delayed_23__33_, chained_data_delayed_23__32_, chained_data_delayed_23__31_, chained_data_delayed_23__30_, chained_data_delayed_23__29_, chained_data_delayed_23__28_, chained_data_delayed_23__27_, chained_data_delayed_23__26_, chained_data_delayed_23__25_, chained_data_delayed_23__24_, chained_data_delayed_23__23_, chained_data_delayed_23__22_, chained_data_delayed_23__21_, chained_data_delayed_23__20_, chained_data_delayed_23__19_, chained_data_delayed_23__18_, chained_data_delayed_23__17_, chained_data_delayed_23__16_, chained_data_delayed_23__15_, chained_data_delayed_23__14_, chained_data_delayed_23__13_, chained_data_delayed_23__12_, chained_data_delayed_23__11_, chained_data_delayed_23__10_, chained_data_delayed_23__9_, chained_data_delayed_23__8_, chained_data_delayed_23__7_, chained_data_delayed_23__6_, chained_data_delayed_23__5_, chained_data_delayed_23__4_, chained_data_delayed_23__3_, chained_data_delayed_23__2_, chained_data_delayed_23__1_, chained_data_delayed_23__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_24__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_23__63_, chained_data_delayed_23__62_, chained_data_delayed_23__61_, chained_data_delayed_23__60_, chained_data_delayed_23__59_, chained_data_delayed_23__58_, chained_data_delayed_23__57_, chained_data_delayed_23__56_, chained_data_delayed_23__55_, chained_data_delayed_23__54_, chained_data_delayed_23__53_, chained_data_delayed_23__52_, chained_data_delayed_23__51_, chained_data_delayed_23__50_, chained_data_delayed_23__49_, chained_data_delayed_23__48_, chained_data_delayed_23__47_, chained_data_delayed_23__46_, chained_data_delayed_23__45_, chained_data_delayed_23__44_, chained_data_delayed_23__43_, chained_data_delayed_23__42_, chained_data_delayed_23__41_, chained_data_delayed_23__40_, chained_data_delayed_23__39_, chained_data_delayed_23__38_, chained_data_delayed_23__37_, chained_data_delayed_23__36_, chained_data_delayed_23__35_, chained_data_delayed_23__34_, chained_data_delayed_23__33_, chained_data_delayed_23__32_, chained_data_delayed_23__31_, chained_data_delayed_23__30_, chained_data_delayed_23__29_, chained_data_delayed_23__28_, chained_data_delayed_23__27_, chained_data_delayed_23__26_, chained_data_delayed_23__25_, chained_data_delayed_23__24_, chained_data_delayed_23__23_, chained_data_delayed_23__22_, chained_data_delayed_23__21_, chained_data_delayed_23__20_, chained_data_delayed_23__19_, chained_data_delayed_23__18_, chained_data_delayed_23__17_, chained_data_delayed_23__16_, chained_data_delayed_23__15_, chained_data_delayed_23__14_, chained_data_delayed_23__13_, chained_data_delayed_23__12_, chained_data_delayed_23__11_, chained_data_delayed_23__10_, chained_data_delayed_23__9_, chained_data_delayed_23__8_, chained_data_delayed_23__7_, chained_data_delayed_23__6_, chained_data_delayed_23__5_, chained_data_delayed_23__4_, chained_data_delayed_23__3_, chained_data_delayed_23__2_, chained_data_delayed_23__1_, chained_data_delayed_23__0_ }),
    .data_o({ chained_data_delayed_24__63_, chained_data_delayed_24__62_, chained_data_delayed_24__61_, chained_data_delayed_24__60_, chained_data_delayed_24__59_, chained_data_delayed_24__58_, chained_data_delayed_24__57_, chained_data_delayed_24__56_, chained_data_delayed_24__55_, chained_data_delayed_24__54_, chained_data_delayed_24__53_, chained_data_delayed_24__52_, chained_data_delayed_24__51_, chained_data_delayed_24__50_, chained_data_delayed_24__49_, chained_data_delayed_24__48_, chained_data_delayed_24__47_, chained_data_delayed_24__46_, chained_data_delayed_24__45_, chained_data_delayed_24__44_, chained_data_delayed_24__43_, chained_data_delayed_24__42_, chained_data_delayed_24__41_, chained_data_delayed_24__40_, chained_data_delayed_24__39_, chained_data_delayed_24__38_, chained_data_delayed_24__37_, chained_data_delayed_24__36_, chained_data_delayed_24__35_, chained_data_delayed_24__34_, chained_data_delayed_24__33_, chained_data_delayed_24__32_, chained_data_delayed_24__31_, chained_data_delayed_24__30_, chained_data_delayed_24__29_, chained_data_delayed_24__28_, chained_data_delayed_24__27_, chained_data_delayed_24__26_, chained_data_delayed_24__25_, chained_data_delayed_24__24_, chained_data_delayed_24__23_, chained_data_delayed_24__22_, chained_data_delayed_24__21_, chained_data_delayed_24__20_, chained_data_delayed_24__19_, chained_data_delayed_24__18_, chained_data_delayed_24__17_, chained_data_delayed_24__16_, chained_data_delayed_24__15_, chained_data_delayed_24__14_, chained_data_delayed_24__13_, chained_data_delayed_24__12_, chained_data_delayed_24__11_, chained_data_delayed_24__10_, chained_data_delayed_24__9_, chained_data_delayed_24__8_, chained_data_delayed_24__7_, chained_data_delayed_24__6_, chained_data_delayed_24__5_, chained_data_delayed_24__4_, chained_data_delayed_24__3_, chained_data_delayed_24__2_, chained_data_delayed_24__1_, chained_data_delayed_24__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_25__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_24__63_, chained_data_delayed_24__62_, chained_data_delayed_24__61_, chained_data_delayed_24__60_, chained_data_delayed_24__59_, chained_data_delayed_24__58_, chained_data_delayed_24__57_, chained_data_delayed_24__56_, chained_data_delayed_24__55_, chained_data_delayed_24__54_, chained_data_delayed_24__53_, chained_data_delayed_24__52_, chained_data_delayed_24__51_, chained_data_delayed_24__50_, chained_data_delayed_24__49_, chained_data_delayed_24__48_, chained_data_delayed_24__47_, chained_data_delayed_24__46_, chained_data_delayed_24__45_, chained_data_delayed_24__44_, chained_data_delayed_24__43_, chained_data_delayed_24__42_, chained_data_delayed_24__41_, chained_data_delayed_24__40_, chained_data_delayed_24__39_, chained_data_delayed_24__38_, chained_data_delayed_24__37_, chained_data_delayed_24__36_, chained_data_delayed_24__35_, chained_data_delayed_24__34_, chained_data_delayed_24__33_, chained_data_delayed_24__32_, chained_data_delayed_24__31_, chained_data_delayed_24__30_, chained_data_delayed_24__29_, chained_data_delayed_24__28_, chained_data_delayed_24__27_, chained_data_delayed_24__26_, chained_data_delayed_24__25_, chained_data_delayed_24__24_, chained_data_delayed_24__23_, chained_data_delayed_24__22_, chained_data_delayed_24__21_, chained_data_delayed_24__20_, chained_data_delayed_24__19_, chained_data_delayed_24__18_, chained_data_delayed_24__17_, chained_data_delayed_24__16_, chained_data_delayed_24__15_, chained_data_delayed_24__14_, chained_data_delayed_24__13_, chained_data_delayed_24__12_, chained_data_delayed_24__11_, chained_data_delayed_24__10_, chained_data_delayed_24__9_, chained_data_delayed_24__8_, chained_data_delayed_24__7_, chained_data_delayed_24__6_, chained_data_delayed_24__5_, chained_data_delayed_24__4_, chained_data_delayed_24__3_, chained_data_delayed_24__2_, chained_data_delayed_24__1_, chained_data_delayed_24__0_ }),
    .data_o({ chained_data_delayed_25__63_, chained_data_delayed_25__62_, chained_data_delayed_25__61_, chained_data_delayed_25__60_, chained_data_delayed_25__59_, chained_data_delayed_25__58_, chained_data_delayed_25__57_, chained_data_delayed_25__56_, chained_data_delayed_25__55_, chained_data_delayed_25__54_, chained_data_delayed_25__53_, chained_data_delayed_25__52_, chained_data_delayed_25__51_, chained_data_delayed_25__50_, chained_data_delayed_25__49_, chained_data_delayed_25__48_, chained_data_delayed_25__47_, chained_data_delayed_25__46_, chained_data_delayed_25__45_, chained_data_delayed_25__44_, chained_data_delayed_25__43_, chained_data_delayed_25__42_, chained_data_delayed_25__41_, chained_data_delayed_25__40_, chained_data_delayed_25__39_, chained_data_delayed_25__38_, chained_data_delayed_25__37_, chained_data_delayed_25__36_, chained_data_delayed_25__35_, chained_data_delayed_25__34_, chained_data_delayed_25__33_, chained_data_delayed_25__32_, chained_data_delayed_25__31_, chained_data_delayed_25__30_, chained_data_delayed_25__29_, chained_data_delayed_25__28_, chained_data_delayed_25__27_, chained_data_delayed_25__26_, chained_data_delayed_25__25_, chained_data_delayed_25__24_, chained_data_delayed_25__23_, chained_data_delayed_25__22_, chained_data_delayed_25__21_, chained_data_delayed_25__20_, chained_data_delayed_25__19_, chained_data_delayed_25__18_, chained_data_delayed_25__17_, chained_data_delayed_25__16_, chained_data_delayed_25__15_, chained_data_delayed_25__14_, chained_data_delayed_25__13_, chained_data_delayed_25__12_, chained_data_delayed_25__11_, chained_data_delayed_25__10_, chained_data_delayed_25__9_, chained_data_delayed_25__8_, chained_data_delayed_25__7_, chained_data_delayed_25__6_, chained_data_delayed_25__5_, chained_data_delayed_25__4_, chained_data_delayed_25__3_, chained_data_delayed_25__2_, chained_data_delayed_25__1_, chained_data_delayed_25__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_26__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_25__63_, chained_data_delayed_25__62_, chained_data_delayed_25__61_, chained_data_delayed_25__60_, chained_data_delayed_25__59_, chained_data_delayed_25__58_, chained_data_delayed_25__57_, chained_data_delayed_25__56_, chained_data_delayed_25__55_, chained_data_delayed_25__54_, chained_data_delayed_25__53_, chained_data_delayed_25__52_, chained_data_delayed_25__51_, chained_data_delayed_25__50_, chained_data_delayed_25__49_, chained_data_delayed_25__48_, chained_data_delayed_25__47_, chained_data_delayed_25__46_, chained_data_delayed_25__45_, chained_data_delayed_25__44_, chained_data_delayed_25__43_, chained_data_delayed_25__42_, chained_data_delayed_25__41_, chained_data_delayed_25__40_, chained_data_delayed_25__39_, chained_data_delayed_25__38_, chained_data_delayed_25__37_, chained_data_delayed_25__36_, chained_data_delayed_25__35_, chained_data_delayed_25__34_, chained_data_delayed_25__33_, chained_data_delayed_25__32_, chained_data_delayed_25__31_, chained_data_delayed_25__30_, chained_data_delayed_25__29_, chained_data_delayed_25__28_, chained_data_delayed_25__27_, chained_data_delayed_25__26_, chained_data_delayed_25__25_, chained_data_delayed_25__24_, chained_data_delayed_25__23_, chained_data_delayed_25__22_, chained_data_delayed_25__21_, chained_data_delayed_25__20_, chained_data_delayed_25__19_, chained_data_delayed_25__18_, chained_data_delayed_25__17_, chained_data_delayed_25__16_, chained_data_delayed_25__15_, chained_data_delayed_25__14_, chained_data_delayed_25__13_, chained_data_delayed_25__12_, chained_data_delayed_25__11_, chained_data_delayed_25__10_, chained_data_delayed_25__9_, chained_data_delayed_25__8_, chained_data_delayed_25__7_, chained_data_delayed_25__6_, chained_data_delayed_25__5_, chained_data_delayed_25__4_, chained_data_delayed_25__3_, chained_data_delayed_25__2_, chained_data_delayed_25__1_, chained_data_delayed_25__0_ }),
    .data_o({ chained_data_delayed_26__63_, chained_data_delayed_26__62_, chained_data_delayed_26__61_, chained_data_delayed_26__60_, chained_data_delayed_26__59_, chained_data_delayed_26__58_, chained_data_delayed_26__57_, chained_data_delayed_26__56_, chained_data_delayed_26__55_, chained_data_delayed_26__54_, chained_data_delayed_26__53_, chained_data_delayed_26__52_, chained_data_delayed_26__51_, chained_data_delayed_26__50_, chained_data_delayed_26__49_, chained_data_delayed_26__48_, chained_data_delayed_26__47_, chained_data_delayed_26__46_, chained_data_delayed_26__45_, chained_data_delayed_26__44_, chained_data_delayed_26__43_, chained_data_delayed_26__42_, chained_data_delayed_26__41_, chained_data_delayed_26__40_, chained_data_delayed_26__39_, chained_data_delayed_26__38_, chained_data_delayed_26__37_, chained_data_delayed_26__36_, chained_data_delayed_26__35_, chained_data_delayed_26__34_, chained_data_delayed_26__33_, chained_data_delayed_26__32_, chained_data_delayed_26__31_, chained_data_delayed_26__30_, chained_data_delayed_26__29_, chained_data_delayed_26__28_, chained_data_delayed_26__27_, chained_data_delayed_26__26_, chained_data_delayed_26__25_, chained_data_delayed_26__24_, chained_data_delayed_26__23_, chained_data_delayed_26__22_, chained_data_delayed_26__21_, chained_data_delayed_26__20_, chained_data_delayed_26__19_, chained_data_delayed_26__18_, chained_data_delayed_26__17_, chained_data_delayed_26__16_, chained_data_delayed_26__15_, chained_data_delayed_26__14_, chained_data_delayed_26__13_, chained_data_delayed_26__12_, chained_data_delayed_26__11_, chained_data_delayed_26__10_, chained_data_delayed_26__9_, chained_data_delayed_26__8_, chained_data_delayed_26__7_, chained_data_delayed_26__6_, chained_data_delayed_26__5_, chained_data_delayed_26__4_, chained_data_delayed_26__3_, chained_data_delayed_26__2_, chained_data_delayed_26__1_, chained_data_delayed_26__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_27__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_26__63_, chained_data_delayed_26__62_, chained_data_delayed_26__61_, chained_data_delayed_26__60_, chained_data_delayed_26__59_, chained_data_delayed_26__58_, chained_data_delayed_26__57_, chained_data_delayed_26__56_, chained_data_delayed_26__55_, chained_data_delayed_26__54_, chained_data_delayed_26__53_, chained_data_delayed_26__52_, chained_data_delayed_26__51_, chained_data_delayed_26__50_, chained_data_delayed_26__49_, chained_data_delayed_26__48_, chained_data_delayed_26__47_, chained_data_delayed_26__46_, chained_data_delayed_26__45_, chained_data_delayed_26__44_, chained_data_delayed_26__43_, chained_data_delayed_26__42_, chained_data_delayed_26__41_, chained_data_delayed_26__40_, chained_data_delayed_26__39_, chained_data_delayed_26__38_, chained_data_delayed_26__37_, chained_data_delayed_26__36_, chained_data_delayed_26__35_, chained_data_delayed_26__34_, chained_data_delayed_26__33_, chained_data_delayed_26__32_, chained_data_delayed_26__31_, chained_data_delayed_26__30_, chained_data_delayed_26__29_, chained_data_delayed_26__28_, chained_data_delayed_26__27_, chained_data_delayed_26__26_, chained_data_delayed_26__25_, chained_data_delayed_26__24_, chained_data_delayed_26__23_, chained_data_delayed_26__22_, chained_data_delayed_26__21_, chained_data_delayed_26__20_, chained_data_delayed_26__19_, chained_data_delayed_26__18_, chained_data_delayed_26__17_, chained_data_delayed_26__16_, chained_data_delayed_26__15_, chained_data_delayed_26__14_, chained_data_delayed_26__13_, chained_data_delayed_26__12_, chained_data_delayed_26__11_, chained_data_delayed_26__10_, chained_data_delayed_26__9_, chained_data_delayed_26__8_, chained_data_delayed_26__7_, chained_data_delayed_26__6_, chained_data_delayed_26__5_, chained_data_delayed_26__4_, chained_data_delayed_26__3_, chained_data_delayed_26__2_, chained_data_delayed_26__1_, chained_data_delayed_26__0_ }),
    .data_o({ chained_data_delayed_27__63_, chained_data_delayed_27__62_, chained_data_delayed_27__61_, chained_data_delayed_27__60_, chained_data_delayed_27__59_, chained_data_delayed_27__58_, chained_data_delayed_27__57_, chained_data_delayed_27__56_, chained_data_delayed_27__55_, chained_data_delayed_27__54_, chained_data_delayed_27__53_, chained_data_delayed_27__52_, chained_data_delayed_27__51_, chained_data_delayed_27__50_, chained_data_delayed_27__49_, chained_data_delayed_27__48_, chained_data_delayed_27__47_, chained_data_delayed_27__46_, chained_data_delayed_27__45_, chained_data_delayed_27__44_, chained_data_delayed_27__43_, chained_data_delayed_27__42_, chained_data_delayed_27__41_, chained_data_delayed_27__40_, chained_data_delayed_27__39_, chained_data_delayed_27__38_, chained_data_delayed_27__37_, chained_data_delayed_27__36_, chained_data_delayed_27__35_, chained_data_delayed_27__34_, chained_data_delayed_27__33_, chained_data_delayed_27__32_, chained_data_delayed_27__31_, chained_data_delayed_27__30_, chained_data_delayed_27__29_, chained_data_delayed_27__28_, chained_data_delayed_27__27_, chained_data_delayed_27__26_, chained_data_delayed_27__25_, chained_data_delayed_27__24_, chained_data_delayed_27__23_, chained_data_delayed_27__22_, chained_data_delayed_27__21_, chained_data_delayed_27__20_, chained_data_delayed_27__19_, chained_data_delayed_27__18_, chained_data_delayed_27__17_, chained_data_delayed_27__16_, chained_data_delayed_27__15_, chained_data_delayed_27__14_, chained_data_delayed_27__13_, chained_data_delayed_27__12_, chained_data_delayed_27__11_, chained_data_delayed_27__10_, chained_data_delayed_27__9_, chained_data_delayed_27__8_, chained_data_delayed_27__7_, chained_data_delayed_27__6_, chained_data_delayed_27__5_, chained_data_delayed_27__4_, chained_data_delayed_27__3_, chained_data_delayed_27__2_, chained_data_delayed_27__1_, chained_data_delayed_27__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_28__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_27__63_, chained_data_delayed_27__62_, chained_data_delayed_27__61_, chained_data_delayed_27__60_, chained_data_delayed_27__59_, chained_data_delayed_27__58_, chained_data_delayed_27__57_, chained_data_delayed_27__56_, chained_data_delayed_27__55_, chained_data_delayed_27__54_, chained_data_delayed_27__53_, chained_data_delayed_27__52_, chained_data_delayed_27__51_, chained_data_delayed_27__50_, chained_data_delayed_27__49_, chained_data_delayed_27__48_, chained_data_delayed_27__47_, chained_data_delayed_27__46_, chained_data_delayed_27__45_, chained_data_delayed_27__44_, chained_data_delayed_27__43_, chained_data_delayed_27__42_, chained_data_delayed_27__41_, chained_data_delayed_27__40_, chained_data_delayed_27__39_, chained_data_delayed_27__38_, chained_data_delayed_27__37_, chained_data_delayed_27__36_, chained_data_delayed_27__35_, chained_data_delayed_27__34_, chained_data_delayed_27__33_, chained_data_delayed_27__32_, chained_data_delayed_27__31_, chained_data_delayed_27__30_, chained_data_delayed_27__29_, chained_data_delayed_27__28_, chained_data_delayed_27__27_, chained_data_delayed_27__26_, chained_data_delayed_27__25_, chained_data_delayed_27__24_, chained_data_delayed_27__23_, chained_data_delayed_27__22_, chained_data_delayed_27__21_, chained_data_delayed_27__20_, chained_data_delayed_27__19_, chained_data_delayed_27__18_, chained_data_delayed_27__17_, chained_data_delayed_27__16_, chained_data_delayed_27__15_, chained_data_delayed_27__14_, chained_data_delayed_27__13_, chained_data_delayed_27__12_, chained_data_delayed_27__11_, chained_data_delayed_27__10_, chained_data_delayed_27__9_, chained_data_delayed_27__8_, chained_data_delayed_27__7_, chained_data_delayed_27__6_, chained_data_delayed_27__5_, chained_data_delayed_27__4_, chained_data_delayed_27__3_, chained_data_delayed_27__2_, chained_data_delayed_27__1_, chained_data_delayed_27__0_ }),
    .data_o({ chained_data_delayed_28__63_, chained_data_delayed_28__62_, chained_data_delayed_28__61_, chained_data_delayed_28__60_, chained_data_delayed_28__59_, chained_data_delayed_28__58_, chained_data_delayed_28__57_, chained_data_delayed_28__56_, chained_data_delayed_28__55_, chained_data_delayed_28__54_, chained_data_delayed_28__53_, chained_data_delayed_28__52_, chained_data_delayed_28__51_, chained_data_delayed_28__50_, chained_data_delayed_28__49_, chained_data_delayed_28__48_, chained_data_delayed_28__47_, chained_data_delayed_28__46_, chained_data_delayed_28__45_, chained_data_delayed_28__44_, chained_data_delayed_28__43_, chained_data_delayed_28__42_, chained_data_delayed_28__41_, chained_data_delayed_28__40_, chained_data_delayed_28__39_, chained_data_delayed_28__38_, chained_data_delayed_28__37_, chained_data_delayed_28__36_, chained_data_delayed_28__35_, chained_data_delayed_28__34_, chained_data_delayed_28__33_, chained_data_delayed_28__32_, chained_data_delayed_28__31_, chained_data_delayed_28__30_, chained_data_delayed_28__29_, chained_data_delayed_28__28_, chained_data_delayed_28__27_, chained_data_delayed_28__26_, chained_data_delayed_28__25_, chained_data_delayed_28__24_, chained_data_delayed_28__23_, chained_data_delayed_28__22_, chained_data_delayed_28__21_, chained_data_delayed_28__20_, chained_data_delayed_28__19_, chained_data_delayed_28__18_, chained_data_delayed_28__17_, chained_data_delayed_28__16_, chained_data_delayed_28__15_, chained_data_delayed_28__14_, chained_data_delayed_28__13_, chained_data_delayed_28__12_, chained_data_delayed_28__11_, chained_data_delayed_28__10_, chained_data_delayed_28__9_, chained_data_delayed_28__8_, chained_data_delayed_28__7_, chained_data_delayed_28__6_, chained_data_delayed_28__5_, chained_data_delayed_28__4_, chained_data_delayed_28__3_, chained_data_delayed_28__2_, chained_data_delayed_28__1_, chained_data_delayed_28__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_29__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_28__63_, chained_data_delayed_28__62_, chained_data_delayed_28__61_, chained_data_delayed_28__60_, chained_data_delayed_28__59_, chained_data_delayed_28__58_, chained_data_delayed_28__57_, chained_data_delayed_28__56_, chained_data_delayed_28__55_, chained_data_delayed_28__54_, chained_data_delayed_28__53_, chained_data_delayed_28__52_, chained_data_delayed_28__51_, chained_data_delayed_28__50_, chained_data_delayed_28__49_, chained_data_delayed_28__48_, chained_data_delayed_28__47_, chained_data_delayed_28__46_, chained_data_delayed_28__45_, chained_data_delayed_28__44_, chained_data_delayed_28__43_, chained_data_delayed_28__42_, chained_data_delayed_28__41_, chained_data_delayed_28__40_, chained_data_delayed_28__39_, chained_data_delayed_28__38_, chained_data_delayed_28__37_, chained_data_delayed_28__36_, chained_data_delayed_28__35_, chained_data_delayed_28__34_, chained_data_delayed_28__33_, chained_data_delayed_28__32_, chained_data_delayed_28__31_, chained_data_delayed_28__30_, chained_data_delayed_28__29_, chained_data_delayed_28__28_, chained_data_delayed_28__27_, chained_data_delayed_28__26_, chained_data_delayed_28__25_, chained_data_delayed_28__24_, chained_data_delayed_28__23_, chained_data_delayed_28__22_, chained_data_delayed_28__21_, chained_data_delayed_28__20_, chained_data_delayed_28__19_, chained_data_delayed_28__18_, chained_data_delayed_28__17_, chained_data_delayed_28__16_, chained_data_delayed_28__15_, chained_data_delayed_28__14_, chained_data_delayed_28__13_, chained_data_delayed_28__12_, chained_data_delayed_28__11_, chained_data_delayed_28__10_, chained_data_delayed_28__9_, chained_data_delayed_28__8_, chained_data_delayed_28__7_, chained_data_delayed_28__6_, chained_data_delayed_28__5_, chained_data_delayed_28__4_, chained_data_delayed_28__3_, chained_data_delayed_28__2_, chained_data_delayed_28__1_, chained_data_delayed_28__0_ }),
    .data_o({ chained_data_delayed_29__63_, chained_data_delayed_29__62_, chained_data_delayed_29__61_, chained_data_delayed_29__60_, chained_data_delayed_29__59_, chained_data_delayed_29__58_, chained_data_delayed_29__57_, chained_data_delayed_29__56_, chained_data_delayed_29__55_, chained_data_delayed_29__54_, chained_data_delayed_29__53_, chained_data_delayed_29__52_, chained_data_delayed_29__51_, chained_data_delayed_29__50_, chained_data_delayed_29__49_, chained_data_delayed_29__48_, chained_data_delayed_29__47_, chained_data_delayed_29__46_, chained_data_delayed_29__45_, chained_data_delayed_29__44_, chained_data_delayed_29__43_, chained_data_delayed_29__42_, chained_data_delayed_29__41_, chained_data_delayed_29__40_, chained_data_delayed_29__39_, chained_data_delayed_29__38_, chained_data_delayed_29__37_, chained_data_delayed_29__36_, chained_data_delayed_29__35_, chained_data_delayed_29__34_, chained_data_delayed_29__33_, chained_data_delayed_29__32_, chained_data_delayed_29__31_, chained_data_delayed_29__30_, chained_data_delayed_29__29_, chained_data_delayed_29__28_, chained_data_delayed_29__27_, chained_data_delayed_29__26_, chained_data_delayed_29__25_, chained_data_delayed_29__24_, chained_data_delayed_29__23_, chained_data_delayed_29__22_, chained_data_delayed_29__21_, chained_data_delayed_29__20_, chained_data_delayed_29__19_, chained_data_delayed_29__18_, chained_data_delayed_29__17_, chained_data_delayed_29__16_, chained_data_delayed_29__15_, chained_data_delayed_29__14_, chained_data_delayed_29__13_, chained_data_delayed_29__12_, chained_data_delayed_29__11_, chained_data_delayed_29__10_, chained_data_delayed_29__9_, chained_data_delayed_29__8_, chained_data_delayed_29__7_, chained_data_delayed_29__6_, chained_data_delayed_29__5_, chained_data_delayed_29__4_, chained_data_delayed_29__3_, chained_data_delayed_29__2_, chained_data_delayed_29__1_, chained_data_delayed_29__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_30__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_29__63_, chained_data_delayed_29__62_, chained_data_delayed_29__61_, chained_data_delayed_29__60_, chained_data_delayed_29__59_, chained_data_delayed_29__58_, chained_data_delayed_29__57_, chained_data_delayed_29__56_, chained_data_delayed_29__55_, chained_data_delayed_29__54_, chained_data_delayed_29__53_, chained_data_delayed_29__52_, chained_data_delayed_29__51_, chained_data_delayed_29__50_, chained_data_delayed_29__49_, chained_data_delayed_29__48_, chained_data_delayed_29__47_, chained_data_delayed_29__46_, chained_data_delayed_29__45_, chained_data_delayed_29__44_, chained_data_delayed_29__43_, chained_data_delayed_29__42_, chained_data_delayed_29__41_, chained_data_delayed_29__40_, chained_data_delayed_29__39_, chained_data_delayed_29__38_, chained_data_delayed_29__37_, chained_data_delayed_29__36_, chained_data_delayed_29__35_, chained_data_delayed_29__34_, chained_data_delayed_29__33_, chained_data_delayed_29__32_, chained_data_delayed_29__31_, chained_data_delayed_29__30_, chained_data_delayed_29__29_, chained_data_delayed_29__28_, chained_data_delayed_29__27_, chained_data_delayed_29__26_, chained_data_delayed_29__25_, chained_data_delayed_29__24_, chained_data_delayed_29__23_, chained_data_delayed_29__22_, chained_data_delayed_29__21_, chained_data_delayed_29__20_, chained_data_delayed_29__19_, chained_data_delayed_29__18_, chained_data_delayed_29__17_, chained_data_delayed_29__16_, chained_data_delayed_29__15_, chained_data_delayed_29__14_, chained_data_delayed_29__13_, chained_data_delayed_29__12_, chained_data_delayed_29__11_, chained_data_delayed_29__10_, chained_data_delayed_29__9_, chained_data_delayed_29__8_, chained_data_delayed_29__7_, chained_data_delayed_29__6_, chained_data_delayed_29__5_, chained_data_delayed_29__4_, chained_data_delayed_29__3_, chained_data_delayed_29__2_, chained_data_delayed_29__1_, chained_data_delayed_29__0_ }),
    .data_o({ chained_data_delayed_30__63_, chained_data_delayed_30__62_, chained_data_delayed_30__61_, chained_data_delayed_30__60_, chained_data_delayed_30__59_, chained_data_delayed_30__58_, chained_data_delayed_30__57_, chained_data_delayed_30__56_, chained_data_delayed_30__55_, chained_data_delayed_30__54_, chained_data_delayed_30__53_, chained_data_delayed_30__52_, chained_data_delayed_30__51_, chained_data_delayed_30__50_, chained_data_delayed_30__49_, chained_data_delayed_30__48_, chained_data_delayed_30__47_, chained_data_delayed_30__46_, chained_data_delayed_30__45_, chained_data_delayed_30__44_, chained_data_delayed_30__43_, chained_data_delayed_30__42_, chained_data_delayed_30__41_, chained_data_delayed_30__40_, chained_data_delayed_30__39_, chained_data_delayed_30__38_, chained_data_delayed_30__37_, chained_data_delayed_30__36_, chained_data_delayed_30__35_, chained_data_delayed_30__34_, chained_data_delayed_30__33_, chained_data_delayed_30__32_, chained_data_delayed_30__31_, chained_data_delayed_30__30_, chained_data_delayed_30__29_, chained_data_delayed_30__28_, chained_data_delayed_30__27_, chained_data_delayed_30__26_, chained_data_delayed_30__25_, chained_data_delayed_30__24_, chained_data_delayed_30__23_, chained_data_delayed_30__22_, chained_data_delayed_30__21_, chained_data_delayed_30__20_, chained_data_delayed_30__19_, chained_data_delayed_30__18_, chained_data_delayed_30__17_, chained_data_delayed_30__16_, chained_data_delayed_30__15_, chained_data_delayed_30__14_, chained_data_delayed_30__13_, chained_data_delayed_30__12_, chained_data_delayed_30__11_, chained_data_delayed_30__10_, chained_data_delayed_30__9_, chained_data_delayed_30__8_, chained_data_delayed_30__7_, chained_data_delayed_30__6_, chained_data_delayed_30__5_, chained_data_delayed_30__4_, chained_data_delayed_30__3_, chained_data_delayed_30__2_, chained_data_delayed_30__1_, chained_data_delayed_30__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_31__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_30__63_, chained_data_delayed_30__62_, chained_data_delayed_30__61_, chained_data_delayed_30__60_, chained_data_delayed_30__59_, chained_data_delayed_30__58_, chained_data_delayed_30__57_, chained_data_delayed_30__56_, chained_data_delayed_30__55_, chained_data_delayed_30__54_, chained_data_delayed_30__53_, chained_data_delayed_30__52_, chained_data_delayed_30__51_, chained_data_delayed_30__50_, chained_data_delayed_30__49_, chained_data_delayed_30__48_, chained_data_delayed_30__47_, chained_data_delayed_30__46_, chained_data_delayed_30__45_, chained_data_delayed_30__44_, chained_data_delayed_30__43_, chained_data_delayed_30__42_, chained_data_delayed_30__41_, chained_data_delayed_30__40_, chained_data_delayed_30__39_, chained_data_delayed_30__38_, chained_data_delayed_30__37_, chained_data_delayed_30__36_, chained_data_delayed_30__35_, chained_data_delayed_30__34_, chained_data_delayed_30__33_, chained_data_delayed_30__32_, chained_data_delayed_30__31_, chained_data_delayed_30__30_, chained_data_delayed_30__29_, chained_data_delayed_30__28_, chained_data_delayed_30__27_, chained_data_delayed_30__26_, chained_data_delayed_30__25_, chained_data_delayed_30__24_, chained_data_delayed_30__23_, chained_data_delayed_30__22_, chained_data_delayed_30__21_, chained_data_delayed_30__20_, chained_data_delayed_30__19_, chained_data_delayed_30__18_, chained_data_delayed_30__17_, chained_data_delayed_30__16_, chained_data_delayed_30__15_, chained_data_delayed_30__14_, chained_data_delayed_30__13_, chained_data_delayed_30__12_, chained_data_delayed_30__11_, chained_data_delayed_30__10_, chained_data_delayed_30__9_, chained_data_delayed_30__8_, chained_data_delayed_30__7_, chained_data_delayed_30__6_, chained_data_delayed_30__5_, chained_data_delayed_30__4_, chained_data_delayed_30__3_, chained_data_delayed_30__2_, chained_data_delayed_30__1_, chained_data_delayed_30__0_ }),
    .data_o({ chained_data_delayed_31__63_, chained_data_delayed_31__62_, chained_data_delayed_31__61_, chained_data_delayed_31__60_, chained_data_delayed_31__59_, chained_data_delayed_31__58_, chained_data_delayed_31__57_, chained_data_delayed_31__56_, chained_data_delayed_31__55_, chained_data_delayed_31__54_, chained_data_delayed_31__53_, chained_data_delayed_31__52_, chained_data_delayed_31__51_, chained_data_delayed_31__50_, chained_data_delayed_31__49_, chained_data_delayed_31__48_, chained_data_delayed_31__47_, chained_data_delayed_31__46_, chained_data_delayed_31__45_, chained_data_delayed_31__44_, chained_data_delayed_31__43_, chained_data_delayed_31__42_, chained_data_delayed_31__41_, chained_data_delayed_31__40_, chained_data_delayed_31__39_, chained_data_delayed_31__38_, chained_data_delayed_31__37_, chained_data_delayed_31__36_, chained_data_delayed_31__35_, chained_data_delayed_31__34_, chained_data_delayed_31__33_, chained_data_delayed_31__32_, chained_data_delayed_31__31_, chained_data_delayed_31__30_, chained_data_delayed_31__29_, chained_data_delayed_31__28_, chained_data_delayed_31__27_, chained_data_delayed_31__26_, chained_data_delayed_31__25_, chained_data_delayed_31__24_, chained_data_delayed_31__23_, chained_data_delayed_31__22_, chained_data_delayed_31__21_, chained_data_delayed_31__20_, chained_data_delayed_31__19_, chained_data_delayed_31__18_, chained_data_delayed_31__17_, chained_data_delayed_31__16_, chained_data_delayed_31__15_, chained_data_delayed_31__14_, chained_data_delayed_31__13_, chained_data_delayed_31__12_, chained_data_delayed_31__11_, chained_data_delayed_31__10_, chained_data_delayed_31__9_, chained_data_delayed_31__8_, chained_data_delayed_31__7_, chained_data_delayed_31__6_, chained_data_delayed_31__5_, chained_data_delayed_31__4_, chained_data_delayed_31__3_, chained_data_delayed_31__2_, chained_data_delayed_31__1_, chained_data_delayed_31__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_32__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_31__63_, chained_data_delayed_31__62_, chained_data_delayed_31__61_, chained_data_delayed_31__60_, chained_data_delayed_31__59_, chained_data_delayed_31__58_, chained_data_delayed_31__57_, chained_data_delayed_31__56_, chained_data_delayed_31__55_, chained_data_delayed_31__54_, chained_data_delayed_31__53_, chained_data_delayed_31__52_, chained_data_delayed_31__51_, chained_data_delayed_31__50_, chained_data_delayed_31__49_, chained_data_delayed_31__48_, chained_data_delayed_31__47_, chained_data_delayed_31__46_, chained_data_delayed_31__45_, chained_data_delayed_31__44_, chained_data_delayed_31__43_, chained_data_delayed_31__42_, chained_data_delayed_31__41_, chained_data_delayed_31__40_, chained_data_delayed_31__39_, chained_data_delayed_31__38_, chained_data_delayed_31__37_, chained_data_delayed_31__36_, chained_data_delayed_31__35_, chained_data_delayed_31__34_, chained_data_delayed_31__33_, chained_data_delayed_31__32_, chained_data_delayed_31__31_, chained_data_delayed_31__30_, chained_data_delayed_31__29_, chained_data_delayed_31__28_, chained_data_delayed_31__27_, chained_data_delayed_31__26_, chained_data_delayed_31__25_, chained_data_delayed_31__24_, chained_data_delayed_31__23_, chained_data_delayed_31__22_, chained_data_delayed_31__21_, chained_data_delayed_31__20_, chained_data_delayed_31__19_, chained_data_delayed_31__18_, chained_data_delayed_31__17_, chained_data_delayed_31__16_, chained_data_delayed_31__15_, chained_data_delayed_31__14_, chained_data_delayed_31__13_, chained_data_delayed_31__12_, chained_data_delayed_31__11_, chained_data_delayed_31__10_, chained_data_delayed_31__9_, chained_data_delayed_31__8_, chained_data_delayed_31__7_, chained_data_delayed_31__6_, chained_data_delayed_31__5_, chained_data_delayed_31__4_, chained_data_delayed_31__3_, chained_data_delayed_31__2_, chained_data_delayed_31__1_, chained_data_delayed_31__0_ }),
    .data_o({ chained_data_delayed_32__63_, chained_data_delayed_32__62_, chained_data_delayed_32__61_, chained_data_delayed_32__60_, chained_data_delayed_32__59_, chained_data_delayed_32__58_, chained_data_delayed_32__57_, chained_data_delayed_32__56_, chained_data_delayed_32__55_, chained_data_delayed_32__54_, chained_data_delayed_32__53_, chained_data_delayed_32__52_, chained_data_delayed_32__51_, chained_data_delayed_32__50_, chained_data_delayed_32__49_, chained_data_delayed_32__48_, chained_data_delayed_32__47_, chained_data_delayed_32__46_, chained_data_delayed_32__45_, chained_data_delayed_32__44_, chained_data_delayed_32__43_, chained_data_delayed_32__42_, chained_data_delayed_32__41_, chained_data_delayed_32__40_, chained_data_delayed_32__39_, chained_data_delayed_32__38_, chained_data_delayed_32__37_, chained_data_delayed_32__36_, chained_data_delayed_32__35_, chained_data_delayed_32__34_, chained_data_delayed_32__33_, chained_data_delayed_32__32_, chained_data_delayed_32__31_, chained_data_delayed_32__30_, chained_data_delayed_32__29_, chained_data_delayed_32__28_, chained_data_delayed_32__27_, chained_data_delayed_32__26_, chained_data_delayed_32__25_, chained_data_delayed_32__24_, chained_data_delayed_32__23_, chained_data_delayed_32__22_, chained_data_delayed_32__21_, chained_data_delayed_32__20_, chained_data_delayed_32__19_, chained_data_delayed_32__18_, chained_data_delayed_32__17_, chained_data_delayed_32__16_, chained_data_delayed_32__15_, chained_data_delayed_32__14_, chained_data_delayed_32__13_, chained_data_delayed_32__12_, chained_data_delayed_32__11_, chained_data_delayed_32__10_, chained_data_delayed_32__9_, chained_data_delayed_32__8_, chained_data_delayed_32__7_, chained_data_delayed_32__6_, chained_data_delayed_32__5_, chained_data_delayed_32__4_, chained_data_delayed_32__3_, chained_data_delayed_32__2_, chained_data_delayed_32__1_, chained_data_delayed_32__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_33__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_32__63_, chained_data_delayed_32__62_, chained_data_delayed_32__61_, chained_data_delayed_32__60_, chained_data_delayed_32__59_, chained_data_delayed_32__58_, chained_data_delayed_32__57_, chained_data_delayed_32__56_, chained_data_delayed_32__55_, chained_data_delayed_32__54_, chained_data_delayed_32__53_, chained_data_delayed_32__52_, chained_data_delayed_32__51_, chained_data_delayed_32__50_, chained_data_delayed_32__49_, chained_data_delayed_32__48_, chained_data_delayed_32__47_, chained_data_delayed_32__46_, chained_data_delayed_32__45_, chained_data_delayed_32__44_, chained_data_delayed_32__43_, chained_data_delayed_32__42_, chained_data_delayed_32__41_, chained_data_delayed_32__40_, chained_data_delayed_32__39_, chained_data_delayed_32__38_, chained_data_delayed_32__37_, chained_data_delayed_32__36_, chained_data_delayed_32__35_, chained_data_delayed_32__34_, chained_data_delayed_32__33_, chained_data_delayed_32__32_, chained_data_delayed_32__31_, chained_data_delayed_32__30_, chained_data_delayed_32__29_, chained_data_delayed_32__28_, chained_data_delayed_32__27_, chained_data_delayed_32__26_, chained_data_delayed_32__25_, chained_data_delayed_32__24_, chained_data_delayed_32__23_, chained_data_delayed_32__22_, chained_data_delayed_32__21_, chained_data_delayed_32__20_, chained_data_delayed_32__19_, chained_data_delayed_32__18_, chained_data_delayed_32__17_, chained_data_delayed_32__16_, chained_data_delayed_32__15_, chained_data_delayed_32__14_, chained_data_delayed_32__13_, chained_data_delayed_32__12_, chained_data_delayed_32__11_, chained_data_delayed_32__10_, chained_data_delayed_32__9_, chained_data_delayed_32__8_, chained_data_delayed_32__7_, chained_data_delayed_32__6_, chained_data_delayed_32__5_, chained_data_delayed_32__4_, chained_data_delayed_32__3_, chained_data_delayed_32__2_, chained_data_delayed_32__1_, chained_data_delayed_32__0_ }),
    .data_o({ chained_data_delayed_33__63_, chained_data_delayed_33__62_, chained_data_delayed_33__61_, chained_data_delayed_33__60_, chained_data_delayed_33__59_, chained_data_delayed_33__58_, chained_data_delayed_33__57_, chained_data_delayed_33__56_, chained_data_delayed_33__55_, chained_data_delayed_33__54_, chained_data_delayed_33__53_, chained_data_delayed_33__52_, chained_data_delayed_33__51_, chained_data_delayed_33__50_, chained_data_delayed_33__49_, chained_data_delayed_33__48_, chained_data_delayed_33__47_, chained_data_delayed_33__46_, chained_data_delayed_33__45_, chained_data_delayed_33__44_, chained_data_delayed_33__43_, chained_data_delayed_33__42_, chained_data_delayed_33__41_, chained_data_delayed_33__40_, chained_data_delayed_33__39_, chained_data_delayed_33__38_, chained_data_delayed_33__37_, chained_data_delayed_33__36_, chained_data_delayed_33__35_, chained_data_delayed_33__34_, chained_data_delayed_33__33_, chained_data_delayed_33__32_, chained_data_delayed_33__31_, chained_data_delayed_33__30_, chained_data_delayed_33__29_, chained_data_delayed_33__28_, chained_data_delayed_33__27_, chained_data_delayed_33__26_, chained_data_delayed_33__25_, chained_data_delayed_33__24_, chained_data_delayed_33__23_, chained_data_delayed_33__22_, chained_data_delayed_33__21_, chained_data_delayed_33__20_, chained_data_delayed_33__19_, chained_data_delayed_33__18_, chained_data_delayed_33__17_, chained_data_delayed_33__16_, chained_data_delayed_33__15_, chained_data_delayed_33__14_, chained_data_delayed_33__13_, chained_data_delayed_33__12_, chained_data_delayed_33__11_, chained_data_delayed_33__10_, chained_data_delayed_33__9_, chained_data_delayed_33__8_, chained_data_delayed_33__7_, chained_data_delayed_33__6_, chained_data_delayed_33__5_, chained_data_delayed_33__4_, chained_data_delayed_33__3_, chained_data_delayed_33__2_, chained_data_delayed_33__1_, chained_data_delayed_33__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_34__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_33__63_, chained_data_delayed_33__62_, chained_data_delayed_33__61_, chained_data_delayed_33__60_, chained_data_delayed_33__59_, chained_data_delayed_33__58_, chained_data_delayed_33__57_, chained_data_delayed_33__56_, chained_data_delayed_33__55_, chained_data_delayed_33__54_, chained_data_delayed_33__53_, chained_data_delayed_33__52_, chained_data_delayed_33__51_, chained_data_delayed_33__50_, chained_data_delayed_33__49_, chained_data_delayed_33__48_, chained_data_delayed_33__47_, chained_data_delayed_33__46_, chained_data_delayed_33__45_, chained_data_delayed_33__44_, chained_data_delayed_33__43_, chained_data_delayed_33__42_, chained_data_delayed_33__41_, chained_data_delayed_33__40_, chained_data_delayed_33__39_, chained_data_delayed_33__38_, chained_data_delayed_33__37_, chained_data_delayed_33__36_, chained_data_delayed_33__35_, chained_data_delayed_33__34_, chained_data_delayed_33__33_, chained_data_delayed_33__32_, chained_data_delayed_33__31_, chained_data_delayed_33__30_, chained_data_delayed_33__29_, chained_data_delayed_33__28_, chained_data_delayed_33__27_, chained_data_delayed_33__26_, chained_data_delayed_33__25_, chained_data_delayed_33__24_, chained_data_delayed_33__23_, chained_data_delayed_33__22_, chained_data_delayed_33__21_, chained_data_delayed_33__20_, chained_data_delayed_33__19_, chained_data_delayed_33__18_, chained_data_delayed_33__17_, chained_data_delayed_33__16_, chained_data_delayed_33__15_, chained_data_delayed_33__14_, chained_data_delayed_33__13_, chained_data_delayed_33__12_, chained_data_delayed_33__11_, chained_data_delayed_33__10_, chained_data_delayed_33__9_, chained_data_delayed_33__8_, chained_data_delayed_33__7_, chained_data_delayed_33__6_, chained_data_delayed_33__5_, chained_data_delayed_33__4_, chained_data_delayed_33__3_, chained_data_delayed_33__2_, chained_data_delayed_33__1_, chained_data_delayed_33__0_ }),
    .data_o({ chained_data_delayed_34__63_, chained_data_delayed_34__62_, chained_data_delayed_34__61_, chained_data_delayed_34__60_, chained_data_delayed_34__59_, chained_data_delayed_34__58_, chained_data_delayed_34__57_, chained_data_delayed_34__56_, chained_data_delayed_34__55_, chained_data_delayed_34__54_, chained_data_delayed_34__53_, chained_data_delayed_34__52_, chained_data_delayed_34__51_, chained_data_delayed_34__50_, chained_data_delayed_34__49_, chained_data_delayed_34__48_, chained_data_delayed_34__47_, chained_data_delayed_34__46_, chained_data_delayed_34__45_, chained_data_delayed_34__44_, chained_data_delayed_34__43_, chained_data_delayed_34__42_, chained_data_delayed_34__41_, chained_data_delayed_34__40_, chained_data_delayed_34__39_, chained_data_delayed_34__38_, chained_data_delayed_34__37_, chained_data_delayed_34__36_, chained_data_delayed_34__35_, chained_data_delayed_34__34_, chained_data_delayed_34__33_, chained_data_delayed_34__32_, chained_data_delayed_34__31_, chained_data_delayed_34__30_, chained_data_delayed_34__29_, chained_data_delayed_34__28_, chained_data_delayed_34__27_, chained_data_delayed_34__26_, chained_data_delayed_34__25_, chained_data_delayed_34__24_, chained_data_delayed_34__23_, chained_data_delayed_34__22_, chained_data_delayed_34__21_, chained_data_delayed_34__20_, chained_data_delayed_34__19_, chained_data_delayed_34__18_, chained_data_delayed_34__17_, chained_data_delayed_34__16_, chained_data_delayed_34__15_, chained_data_delayed_34__14_, chained_data_delayed_34__13_, chained_data_delayed_34__12_, chained_data_delayed_34__11_, chained_data_delayed_34__10_, chained_data_delayed_34__9_, chained_data_delayed_34__8_, chained_data_delayed_34__7_, chained_data_delayed_34__6_, chained_data_delayed_34__5_, chained_data_delayed_34__4_, chained_data_delayed_34__3_, chained_data_delayed_34__2_, chained_data_delayed_34__1_, chained_data_delayed_34__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_35__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_34__63_, chained_data_delayed_34__62_, chained_data_delayed_34__61_, chained_data_delayed_34__60_, chained_data_delayed_34__59_, chained_data_delayed_34__58_, chained_data_delayed_34__57_, chained_data_delayed_34__56_, chained_data_delayed_34__55_, chained_data_delayed_34__54_, chained_data_delayed_34__53_, chained_data_delayed_34__52_, chained_data_delayed_34__51_, chained_data_delayed_34__50_, chained_data_delayed_34__49_, chained_data_delayed_34__48_, chained_data_delayed_34__47_, chained_data_delayed_34__46_, chained_data_delayed_34__45_, chained_data_delayed_34__44_, chained_data_delayed_34__43_, chained_data_delayed_34__42_, chained_data_delayed_34__41_, chained_data_delayed_34__40_, chained_data_delayed_34__39_, chained_data_delayed_34__38_, chained_data_delayed_34__37_, chained_data_delayed_34__36_, chained_data_delayed_34__35_, chained_data_delayed_34__34_, chained_data_delayed_34__33_, chained_data_delayed_34__32_, chained_data_delayed_34__31_, chained_data_delayed_34__30_, chained_data_delayed_34__29_, chained_data_delayed_34__28_, chained_data_delayed_34__27_, chained_data_delayed_34__26_, chained_data_delayed_34__25_, chained_data_delayed_34__24_, chained_data_delayed_34__23_, chained_data_delayed_34__22_, chained_data_delayed_34__21_, chained_data_delayed_34__20_, chained_data_delayed_34__19_, chained_data_delayed_34__18_, chained_data_delayed_34__17_, chained_data_delayed_34__16_, chained_data_delayed_34__15_, chained_data_delayed_34__14_, chained_data_delayed_34__13_, chained_data_delayed_34__12_, chained_data_delayed_34__11_, chained_data_delayed_34__10_, chained_data_delayed_34__9_, chained_data_delayed_34__8_, chained_data_delayed_34__7_, chained_data_delayed_34__6_, chained_data_delayed_34__5_, chained_data_delayed_34__4_, chained_data_delayed_34__3_, chained_data_delayed_34__2_, chained_data_delayed_34__1_, chained_data_delayed_34__0_ }),
    .data_o({ chained_data_delayed_35__63_, chained_data_delayed_35__62_, chained_data_delayed_35__61_, chained_data_delayed_35__60_, chained_data_delayed_35__59_, chained_data_delayed_35__58_, chained_data_delayed_35__57_, chained_data_delayed_35__56_, chained_data_delayed_35__55_, chained_data_delayed_35__54_, chained_data_delayed_35__53_, chained_data_delayed_35__52_, chained_data_delayed_35__51_, chained_data_delayed_35__50_, chained_data_delayed_35__49_, chained_data_delayed_35__48_, chained_data_delayed_35__47_, chained_data_delayed_35__46_, chained_data_delayed_35__45_, chained_data_delayed_35__44_, chained_data_delayed_35__43_, chained_data_delayed_35__42_, chained_data_delayed_35__41_, chained_data_delayed_35__40_, chained_data_delayed_35__39_, chained_data_delayed_35__38_, chained_data_delayed_35__37_, chained_data_delayed_35__36_, chained_data_delayed_35__35_, chained_data_delayed_35__34_, chained_data_delayed_35__33_, chained_data_delayed_35__32_, chained_data_delayed_35__31_, chained_data_delayed_35__30_, chained_data_delayed_35__29_, chained_data_delayed_35__28_, chained_data_delayed_35__27_, chained_data_delayed_35__26_, chained_data_delayed_35__25_, chained_data_delayed_35__24_, chained_data_delayed_35__23_, chained_data_delayed_35__22_, chained_data_delayed_35__21_, chained_data_delayed_35__20_, chained_data_delayed_35__19_, chained_data_delayed_35__18_, chained_data_delayed_35__17_, chained_data_delayed_35__16_, chained_data_delayed_35__15_, chained_data_delayed_35__14_, chained_data_delayed_35__13_, chained_data_delayed_35__12_, chained_data_delayed_35__11_, chained_data_delayed_35__10_, chained_data_delayed_35__9_, chained_data_delayed_35__8_, chained_data_delayed_35__7_, chained_data_delayed_35__6_, chained_data_delayed_35__5_, chained_data_delayed_35__4_, chained_data_delayed_35__3_, chained_data_delayed_35__2_, chained_data_delayed_35__1_, chained_data_delayed_35__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_36__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_35__63_, chained_data_delayed_35__62_, chained_data_delayed_35__61_, chained_data_delayed_35__60_, chained_data_delayed_35__59_, chained_data_delayed_35__58_, chained_data_delayed_35__57_, chained_data_delayed_35__56_, chained_data_delayed_35__55_, chained_data_delayed_35__54_, chained_data_delayed_35__53_, chained_data_delayed_35__52_, chained_data_delayed_35__51_, chained_data_delayed_35__50_, chained_data_delayed_35__49_, chained_data_delayed_35__48_, chained_data_delayed_35__47_, chained_data_delayed_35__46_, chained_data_delayed_35__45_, chained_data_delayed_35__44_, chained_data_delayed_35__43_, chained_data_delayed_35__42_, chained_data_delayed_35__41_, chained_data_delayed_35__40_, chained_data_delayed_35__39_, chained_data_delayed_35__38_, chained_data_delayed_35__37_, chained_data_delayed_35__36_, chained_data_delayed_35__35_, chained_data_delayed_35__34_, chained_data_delayed_35__33_, chained_data_delayed_35__32_, chained_data_delayed_35__31_, chained_data_delayed_35__30_, chained_data_delayed_35__29_, chained_data_delayed_35__28_, chained_data_delayed_35__27_, chained_data_delayed_35__26_, chained_data_delayed_35__25_, chained_data_delayed_35__24_, chained_data_delayed_35__23_, chained_data_delayed_35__22_, chained_data_delayed_35__21_, chained_data_delayed_35__20_, chained_data_delayed_35__19_, chained_data_delayed_35__18_, chained_data_delayed_35__17_, chained_data_delayed_35__16_, chained_data_delayed_35__15_, chained_data_delayed_35__14_, chained_data_delayed_35__13_, chained_data_delayed_35__12_, chained_data_delayed_35__11_, chained_data_delayed_35__10_, chained_data_delayed_35__9_, chained_data_delayed_35__8_, chained_data_delayed_35__7_, chained_data_delayed_35__6_, chained_data_delayed_35__5_, chained_data_delayed_35__4_, chained_data_delayed_35__3_, chained_data_delayed_35__2_, chained_data_delayed_35__1_, chained_data_delayed_35__0_ }),
    .data_o({ chained_data_delayed_36__63_, chained_data_delayed_36__62_, chained_data_delayed_36__61_, chained_data_delayed_36__60_, chained_data_delayed_36__59_, chained_data_delayed_36__58_, chained_data_delayed_36__57_, chained_data_delayed_36__56_, chained_data_delayed_36__55_, chained_data_delayed_36__54_, chained_data_delayed_36__53_, chained_data_delayed_36__52_, chained_data_delayed_36__51_, chained_data_delayed_36__50_, chained_data_delayed_36__49_, chained_data_delayed_36__48_, chained_data_delayed_36__47_, chained_data_delayed_36__46_, chained_data_delayed_36__45_, chained_data_delayed_36__44_, chained_data_delayed_36__43_, chained_data_delayed_36__42_, chained_data_delayed_36__41_, chained_data_delayed_36__40_, chained_data_delayed_36__39_, chained_data_delayed_36__38_, chained_data_delayed_36__37_, chained_data_delayed_36__36_, chained_data_delayed_36__35_, chained_data_delayed_36__34_, chained_data_delayed_36__33_, chained_data_delayed_36__32_, chained_data_delayed_36__31_, chained_data_delayed_36__30_, chained_data_delayed_36__29_, chained_data_delayed_36__28_, chained_data_delayed_36__27_, chained_data_delayed_36__26_, chained_data_delayed_36__25_, chained_data_delayed_36__24_, chained_data_delayed_36__23_, chained_data_delayed_36__22_, chained_data_delayed_36__21_, chained_data_delayed_36__20_, chained_data_delayed_36__19_, chained_data_delayed_36__18_, chained_data_delayed_36__17_, chained_data_delayed_36__16_, chained_data_delayed_36__15_, chained_data_delayed_36__14_, chained_data_delayed_36__13_, chained_data_delayed_36__12_, chained_data_delayed_36__11_, chained_data_delayed_36__10_, chained_data_delayed_36__9_, chained_data_delayed_36__8_, chained_data_delayed_36__7_, chained_data_delayed_36__6_, chained_data_delayed_36__5_, chained_data_delayed_36__4_, chained_data_delayed_36__3_, chained_data_delayed_36__2_, chained_data_delayed_36__1_, chained_data_delayed_36__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_37__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_36__63_, chained_data_delayed_36__62_, chained_data_delayed_36__61_, chained_data_delayed_36__60_, chained_data_delayed_36__59_, chained_data_delayed_36__58_, chained_data_delayed_36__57_, chained_data_delayed_36__56_, chained_data_delayed_36__55_, chained_data_delayed_36__54_, chained_data_delayed_36__53_, chained_data_delayed_36__52_, chained_data_delayed_36__51_, chained_data_delayed_36__50_, chained_data_delayed_36__49_, chained_data_delayed_36__48_, chained_data_delayed_36__47_, chained_data_delayed_36__46_, chained_data_delayed_36__45_, chained_data_delayed_36__44_, chained_data_delayed_36__43_, chained_data_delayed_36__42_, chained_data_delayed_36__41_, chained_data_delayed_36__40_, chained_data_delayed_36__39_, chained_data_delayed_36__38_, chained_data_delayed_36__37_, chained_data_delayed_36__36_, chained_data_delayed_36__35_, chained_data_delayed_36__34_, chained_data_delayed_36__33_, chained_data_delayed_36__32_, chained_data_delayed_36__31_, chained_data_delayed_36__30_, chained_data_delayed_36__29_, chained_data_delayed_36__28_, chained_data_delayed_36__27_, chained_data_delayed_36__26_, chained_data_delayed_36__25_, chained_data_delayed_36__24_, chained_data_delayed_36__23_, chained_data_delayed_36__22_, chained_data_delayed_36__21_, chained_data_delayed_36__20_, chained_data_delayed_36__19_, chained_data_delayed_36__18_, chained_data_delayed_36__17_, chained_data_delayed_36__16_, chained_data_delayed_36__15_, chained_data_delayed_36__14_, chained_data_delayed_36__13_, chained_data_delayed_36__12_, chained_data_delayed_36__11_, chained_data_delayed_36__10_, chained_data_delayed_36__9_, chained_data_delayed_36__8_, chained_data_delayed_36__7_, chained_data_delayed_36__6_, chained_data_delayed_36__5_, chained_data_delayed_36__4_, chained_data_delayed_36__3_, chained_data_delayed_36__2_, chained_data_delayed_36__1_, chained_data_delayed_36__0_ }),
    .data_o({ chained_data_delayed_37__63_, chained_data_delayed_37__62_, chained_data_delayed_37__61_, chained_data_delayed_37__60_, chained_data_delayed_37__59_, chained_data_delayed_37__58_, chained_data_delayed_37__57_, chained_data_delayed_37__56_, chained_data_delayed_37__55_, chained_data_delayed_37__54_, chained_data_delayed_37__53_, chained_data_delayed_37__52_, chained_data_delayed_37__51_, chained_data_delayed_37__50_, chained_data_delayed_37__49_, chained_data_delayed_37__48_, chained_data_delayed_37__47_, chained_data_delayed_37__46_, chained_data_delayed_37__45_, chained_data_delayed_37__44_, chained_data_delayed_37__43_, chained_data_delayed_37__42_, chained_data_delayed_37__41_, chained_data_delayed_37__40_, chained_data_delayed_37__39_, chained_data_delayed_37__38_, chained_data_delayed_37__37_, chained_data_delayed_37__36_, chained_data_delayed_37__35_, chained_data_delayed_37__34_, chained_data_delayed_37__33_, chained_data_delayed_37__32_, chained_data_delayed_37__31_, chained_data_delayed_37__30_, chained_data_delayed_37__29_, chained_data_delayed_37__28_, chained_data_delayed_37__27_, chained_data_delayed_37__26_, chained_data_delayed_37__25_, chained_data_delayed_37__24_, chained_data_delayed_37__23_, chained_data_delayed_37__22_, chained_data_delayed_37__21_, chained_data_delayed_37__20_, chained_data_delayed_37__19_, chained_data_delayed_37__18_, chained_data_delayed_37__17_, chained_data_delayed_37__16_, chained_data_delayed_37__15_, chained_data_delayed_37__14_, chained_data_delayed_37__13_, chained_data_delayed_37__12_, chained_data_delayed_37__11_, chained_data_delayed_37__10_, chained_data_delayed_37__9_, chained_data_delayed_37__8_, chained_data_delayed_37__7_, chained_data_delayed_37__6_, chained_data_delayed_37__5_, chained_data_delayed_37__4_, chained_data_delayed_37__3_, chained_data_delayed_37__2_, chained_data_delayed_37__1_, chained_data_delayed_37__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_38__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_37__63_, chained_data_delayed_37__62_, chained_data_delayed_37__61_, chained_data_delayed_37__60_, chained_data_delayed_37__59_, chained_data_delayed_37__58_, chained_data_delayed_37__57_, chained_data_delayed_37__56_, chained_data_delayed_37__55_, chained_data_delayed_37__54_, chained_data_delayed_37__53_, chained_data_delayed_37__52_, chained_data_delayed_37__51_, chained_data_delayed_37__50_, chained_data_delayed_37__49_, chained_data_delayed_37__48_, chained_data_delayed_37__47_, chained_data_delayed_37__46_, chained_data_delayed_37__45_, chained_data_delayed_37__44_, chained_data_delayed_37__43_, chained_data_delayed_37__42_, chained_data_delayed_37__41_, chained_data_delayed_37__40_, chained_data_delayed_37__39_, chained_data_delayed_37__38_, chained_data_delayed_37__37_, chained_data_delayed_37__36_, chained_data_delayed_37__35_, chained_data_delayed_37__34_, chained_data_delayed_37__33_, chained_data_delayed_37__32_, chained_data_delayed_37__31_, chained_data_delayed_37__30_, chained_data_delayed_37__29_, chained_data_delayed_37__28_, chained_data_delayed_37__27_, chained_data_delayed_37__26_, chained_data_delayed_37__25_, chained_data_delayed_37__24_, chained_data_delayed_37__23_, chained_data_delayed_37__22_, chained_data_delayed_37__21_, chained_data_delayed_37__20_, chained_data_delayed_37__19_, chained_data_delayed_37__18_, chained_data_delayed_37__17_, chained_data_delayed_37__16_, chained_data_delayed_37__15_, chained_data_delayed_37__14_, chained_data_delayed_37__13_, chained_data_delayed_37__12_, chained_data_delayed_37__11_, chained_data_delayed_37__10_, chained_data_delayed_37__9_, chained_data_delayed_37__8_, chained_data_delayed_37__7_, chained_data_delayed_37__6_, chained_data_delayed_37__5_, chained_data_delayed_37__4_, chained_data_delayed_37__3_, chained_data_delayed_37__2_, chained_data_delayed_37__1_, chained_data_delayed_37__0_ }),
    .data_o({ chained_data_delayed_38__63_, chained_data_delayed_38__62_, chained_data_delayed_38__61_, chained_data_delayed_38__60_, chained_data_delayed_38__59_, chained_data_delayed_38__58_, chained_data_delayed_38__57_, chained_data_delayed_38__56_, chained_data_delayed_38__55_, chained_data_delayed_38__54_, chained_data_delayed_38__53_, chained_data_delayed_38__52_, chained_data_delayed_38__51_, chained_data_delayed_38__50_, chained_data_delayed_38__49_, chained_data_delayed_38__48_, chained_data_delayed_38__47_, chained_data_delayed_38__46_, chained_data_delayed_38__45_, chained_data_delayed_38__44_, chained_data_delayed_38__43_, chained_data_delayed_38__42_, chained_data_delayed_38__41_, chained_data_delayed_38__40_, chained_data_delayed_38__39_, chained_data_delayed_38__38_, chained_data_delayed_38__37_, chained_data_delayed_38__36_, chained_data_delayed_38__35_, chained_data_delayed_38__34_, chained_data_delayed_38__33_, chained_data_delayed_38__32_, chained_data_delayed_38__31_, chained_data_delayed_38__30_, chained_data_delayed_38__29_, chained_data_delayed_38__28_, chained_data_delayed_38__27_, chained_data_delayed_38__26_, chained_data_delayed_38__25_, chained_data_delayed_38__24_, chained_data_delayed_38__23_, chained_data_delayed_38__22_, chained_data_delayed_38__21_, chained_data_delayed_38__20_, chained_data_delayed_38__19_, chained_data_delayed_38__18_, chained_data_delayed_38__17_, chained_data_delayed_38__16_, chained_data_delayed_38__15_, chained_data_delayed_38__14_, chained_data_delayed_38__13_, chained_data_delayed_38__12_, chained_data_delayed_38__11_, chained_data_delayed_38__10_, chained_data_delayed_38__9_, chained_data_delayed_38__8_, chained_data_delayed_38__7_, chained_data_delayed_38__6_, chained_data_delayed_38__5_, chained_data_delayed_38__4_, chained_data_delayed_38__3_, chained_data_delayed_38__2_, chained_data_delayed_38__1_, chained_data_delayed_38__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_39__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_38__63_, chained_data_delayed_38__62_, chained_data_delayed_38__61_, chained_data_delayed_38__60_, chained_data_delayed_38__59_, chained_data_delayed_38__58_, chained_data_delayed_38__57_, chained_data_delayed_38__56_, chained_data_delayed_38__55_, chained_data_delayed_38__54_, chained_data_delayed_38__53_, chained_data_delayed_38__52_, chained_data_delayed_38__51_, chained_data_delayed_38__50_, chained_data_delayed_38__49_, chained_data_delayed_38__48_, chained_data_delayed_38__47_, chained_data_delayed_38__46_, chained_data_delayed_38__45_, chained_data_delayed_38__44_, chained_data_delayed_38__43_, chained_data_delayed_38__42_, chained_data_delayed_38__41_, chained_data_delayed_38__40_, chained_data_delayed_38__39_, chained_data_delayed_38__38_, chained_data_delayed_38__37_, chained_data_delayed_38__36_, chained_data_delayed_38__35_, chained_data_delayed_38__34_, chained_data_delayed_38__33_, chained_data_delayed_38__32_, chained_data_delayed_38__31_, chained_data_delayed_38__30_, chained_data_delayed_38__29_, chained_data_delayed_38__28_, chained_data_delayed_38__27_, chained_data_delayed_38__26_, chained_data_delayed_38__25_, chained_data_delayed_38__24_, chained_data_delayed_38__23_, chained_data_delayed_38__22_, chained_data_delayed_38__21_, chained_data_delayed_38__20_, chained_data_delayed_38__19_, chained_data_delayed_38__18_, chained_data_delayed_38__17_, chained_data_delayed_38__16_, chained_data_delayed_38__15_, chained_data_delayed_38__14_, chained_data_delayed_38__13_, chained_data_delayed_38__12_, chained_data_delayed_38__11_, chained_data_delayed_38__10_, chained_data_delayed_38__9_, chained_data_delayed_38__8_, chained_data_delayed_38__7_, chained_data_delayed_38__6_, chained_data_delayed_38__5_, chained_data_delayed_38__4_, chained_data_delayed_38__3_, chained_data_delayed_38__2_, chained_data_delayed_38__1_, chained_data_delayed_38__0_ }),
    .data_o({ chained_data_delayed_39__63_, chained_data_delayed_39__62_, chained_data_delayed_39__61_, chained_data_delayed_39__60_, chained_data_delayed_39__59_, chained_data_delayed_39__58_, chained_data_delayed_39__57_, chained_data_delayed_39__56_, chained_data_delayed_39__55_, chained_data_delayed_39__54_, chained_data_delayed_39__53_, chained_data_delayed_39__52_, chained_data_delayed_39__51_, chained_data_delayed_39__50_, chained_data_delayed_39__49_, chained_data_delayed_39__48_, chained_data_delayed_39__47_, chained_data_delayed_39__46_, chained_data_delayed_39__45_, chained_data_delayed_39__44_, chained_data_delayed_39__43_, chained_data_delayed_39__42_, chained_data_delayed_39__41_, chained_data_delayed_39__40_, chained_data_delayed_39__39_, chained_data_delayed_39__38_, chained_data_delayed_39__37_, chained_data_delayed_39__36_, chained_data_delayed_39__35_, chained_data_delayed_39__34_, chained_data_delayed_39__33_, chained_data_delayed_39__32_, chained_data_delayed_39__31_, chained_data_delayed_39__30_, chained_data_delayed_39__29_, chained_data_delayed_39__28_, chained_data_delayed_39__27_, chained_data_delayed_39__26_, chained_data_delayed_39__25_, chained_data_delayed_39__24_, chained_data_delayed_39__23_, chained_data_delayed_39__22_, chained_data_delayed_39__21_, chained_data_delayed_39__20_, chained_data_delayed_39__19_, chained_data_delayed_39__18_, chained_data_delayed_39__17_, chained_data_delayed_39__16_, chained_data_delayed_39__15_, chained_data_delayed_39__14_, chained_data_delayed_39__13_, chained_data_delayed_39__12_, chained_data_delayed_39__11_, chained_data_delayed_39__10_, chained_data_delayed_39__9_, chained_data_delayed_39__8_, chained_data_delayed_39__7_, chained_data_delayed_39__6_, chained_data_delayed_39__5_, chained_data_delayed_39__4_, chained_data_delayed_39__3_, chained_data_delayed_39__2_, chained_data_delayed_39__1_, chained_data_delayed_39__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_40__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_39__63_, chained_data_delayed_39__62_, chained_data_delayed_39__61_, chained_data_delayed_39__60_, chained_data_delayed_39__59_, chained_data_delayed_39__58_, chained_data_delayed_39__57_, chained_data_delayed_39__56_, chained_data_delayed_39__55_, chained_data_delayed_39__54_, chained_data_delayed_39__53_, chained_data_delayed_39__52_, chained_data_delayed_39__51_, chained_data_delayed_39__50_, chained_data_delayed_39__49_, chained_data_delayed_39__48_, chained_data_delayed_39__47_, chained_data_delayed_39__46_, chained_data_delayed_39__45_, chained_data_delayed_39__44_, chained_data_delayed_39__43_, chained_data_delayed_39__42_, chained_data_delayed_39__41_, chained_data_delayed_39__40_, chained_data_delayed_39__39_, chained_data_delayed_39__38_, chained_data_delayed_39__37_, chained_data_delayed_39__36_, chained_data_delayed_39__35_, chained_data_delayed_39__34_, chained_data_delayed_39__33_, chained_data_delayed_39__32_, chained_data_delayed_39__31_, chained_data_delayed_39__30_, chained_data_delayed_39__29_, chained_data_delayed_39__28_, chained_data_delayed_39__27_, chained_data_delayed_39__26_, chained_data_delayed_39__25_, chained_data_delayed_39__24_, chained_data_delayed_39__23_, chained_data_delayed_39__22_, chained_data_delayed_39__21_, chained_data_delayed_39__20_, chained_data_delayed_39__19_, chained_data_delayed_39__18_, chained_data_delayed_39__17_, chained_data_delayed_39__16_, chained_data_delayed_39__15_, chained_data_delayed_39__14_, chained_data_delayed_39__13_, chained_data_delayed_39__12_, chained_data_delayed_39__11_, chained_data_delayed_39__10_, chained_data_delayed_39__9_, chained_data_delayed_39__8_, chained_data_delayed_39__7_, chained_data_delayed_39__6_, chained_data_delayed_39__5_, chained_data_delayed_39__4_, chained_data_delayed_39__3_, chained_data_delayed_39__2_, chained_data_delayed_39__1_, chained_data_delayed_39__0_ }),
    .data_o({ chained_data_delayed_40__63_, chained_data_delayed_40__62_, chained_data_delayed_40__61_, chained_data_delayed_40__60_, chained_data_delayed_40__59_, chained_data_delayed_40__58_, chained_data_delayed_40__57_, chained_data_delayed_40__56_, chained_data_delayed_40__55_, chained_data_delayed_40__54_, chained_data_delayed_40__53_, chained_data_delayed_40__52_, chained_data_delayed_40__51_, chained_data_delayed_40__50_, chained_data_delayed_40__49_, chained_data_delayed_40__48_, chained_data_delayed_40__47_, chained_data_delayed_40__46_, chained_data_delayed_40__45_, chained_data_delayed_40__44_, chained_data_delayed_40__43_, chained_data_delayed_40__42_, chained_data_delayed_40__41_, chained_data_delayed_40__40_, chained_data_delayed_40__39_, chained_data_delayed_40__38_, chained_data_delayed_40__37_, chained_data_delayed_40__36_, chained_data_delayed_40__35_, chained_data_delayed_40__34_, chained_data_delayed_40__33_, chained_data_delayed_40__32_, chained_data_delayed_40__31_, chained_data_delayed_40__30_, chained_data_delayed_40__29_, chained_data_delayed_40__28_, chained_data_delayed_40__27_, chained_data_delayed_40__26_, chained_data_delayed_40__25_, chained_data_delayed_40__24_, chained_data_delayed_40__23_, chained_data_delayed_40__22_, chained_data_delayed_40__21_, chained_data_delayed_40__20_, chained_data_delayed_40__19_, chained_data_delayed_40__18_, chained_data_delayed_40__17_, chained_data_delayed_40__16_, chained_data_delayed_40__15_, chained_data_delayed_40__14_, chained_data_delayed_40__13_, chained_data_delayed_40__12_, chained_data_delayed_40__11_, chained_data_delayed_40__10_, chained_data_delayed_40__9_, chained_data_delayed_40__8_, chained_data_delayed_40__7_, chained_data_delayed_40__6_, chained_data_delayed_40__5_, chained_data_delayed_40__4_, chained_data_delayed_40__3_, chained_data_delayed_40__2_, chained_data_delayed_40__1_, chained_data_delayed_40__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_41__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_40__63_, chained_data_delayed_40__62_, chained_data_delayed_40__61_, chained_data_delayed_40__60_, chained_data_delayed_40__59_, chained_data_delayed_40__58_, chained_data_delayed_40__57_, chained_data_delayed_40__56_, chained_data_delayed_40__55_, chained_data_delayed_40__54_, chained_data_delayed_40__53_, chained_data_delayed_40__52_, chained_data_delayed_40__51_, chained_data_delayed_40__50_, chained_data_delayed_40__49_, chained_data_delayed_40__48_, chained_data_delayed_40__47_, chained_data_delayed_40__46_, chained_data_delayed_40__45_, chained_data_delayed_40__44_, chained_data_delayed_40__43_, chained_data_delayed_40__42_, chained_data_delayed_40__41_, chained_data_delayed_40__40_, chained_data_delayed_40__39_, chained_data_delayed_40__38_, chained_data_delayed_40__37_, chained_data_delayed_40__36_, chained_data_delayed_40__35_, chained_data_delayed_40__34_, chained_data_delayed_40__33_, chained_data_delayed_40__32_, chained_data_delayed_40__31_, chained_data_delayed_40__30_, chained_data_delayed_40__29_, chained_data_delayed_40__28_, chained_data_delayed_40__27_, chained_data_delayed_40__26_, chained_data_delayed_40__25_, chained_data_delayed_40__24_, chained_data_delayed_40__23_, chained_data_delayed_40__22_, chained_data_delayed_40__21_, chained_data_delayed_40__20_, chained_data_delayed_40__19_, chained_data_delayed_40__18_, chained_data_delayed_40__17_, chained_data_delayed_40__16_, chained_data_delayed_40__15_, chained_data_delayed_40__14_, chained_data_delayed_40__13_, chained_data_delayed_40__12_, chained_data_delayed_40__11_, chained_data_delayed_40__10_, chained_data_delayed_40__9_, chained_data_delayed_40__8_, chained_data_delayed_40__7_, chained_data_delayed_40__6_, chained_data_delayed_40__5_, chained_data_delayed_40__4_, chained_data_delayed_40__3_, chained_data_delayed_40__2_, chained_data_delayed_40__1_, chained_data_delayed_40__0_ }),
    .data_o({ chained_data_delayed_41__63_, chained_data_delayed_41__62_, chained_data_delayed_41__61_, chained_data_delayed_41__60_, chained_data_delayed_41__59_, chained_data_delayed_41__58_, chained_data_delayed_41__57_, chained_data_delayed_41__56_, chained_data_delayed_41__55_, chained_data_delayed_41__54_, chained_data_delayed_41__53_, chained_data_delayed_41__52_, chained_data_delayed_41__51_, chained_data_delayed_41__50_, chained_data_delayed_41__49_, chained_data_delayed_41__48_, chained_data_delayed_41__47_, chained_data_delayed_41__46_, chained_data_delayed_41__45_, chained_data_delayed_41__44_, chained_data_delayed_41__43_, chained_data_delayed_41__42_, chained_data_delayed_41__41_, chained_data_delayed_41__40_, chained_data_delayed_41__39_, chained_data_delayed_41__38_, chained_data_delayed_41__37_, chained_data_delayed_41__36_, chained_data_delayed_41__35_, chained_data_delayed_41__34_, chained_data_delayed_41__33_, chained_data_delayed_41__32_, chained_data_delayed_41__31_, chained_data_delayed_41__30_, chained_data_delayed_41__29_, chained_data_delayed_41__28_, chained_data_delayed_41__27_, chained_data_delayed_41__26_, chained_data_delayed_41__25_, chained_data_delayed_41__24_, chained_data_delayed_41__23_, chained_data_delayed_41__22_, chained_data_delayed_41__21_, chained_data_delayed_41__20_, chained_data_delayed_41__19_, chained_data_delayed_41__18_, chained_data_delayed_41__17_, chained_data_delayed_41__16_, chained_data_delayed_41__15_, chained_data_delayed_41__14_, chained_data_delayed_41__13_, chained_data_delayed_41__12_, chained_data_delayed_41__11_, chained_data_delayed_41__10_, chained_data_delayed_41__9_, chained_data_delayed_41__8_, chained_data_delayed_41__7_, chained_data_delayed_41__6_, chained_data_delayed_41__5_, chained_data_delayed_41__4_, chained_data_delayed_41__3_, chained_data_delayed_41__2_, chained_data_delayed_41__1_, chained_data_delayed_41__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_42__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_41__63_, chained_data_delayed_41__62_, chained_data_delayed_41__61_, chained_data_delayed_41__60_, chained_data_delayed_41__59_, chained_data_delayed_41__58_, chained_data_delayed_41__57_, chained_data_delayed_41__56_, chained_data_delayed_41__55_, chained_data_delayed_41__54_, chained_data_delayed_41__53_, chained_data_delayed_41__52_, chained_data_delayed_41__51_, chained_data_delayed_41__50_, chained_data_delayed_41__49_, chained_data_delayed_41__48_, chained_data_delayed_41__47_, chained_data_delayed_41__46_, chained_data_delayed_41__45_, chained_data_delayed_41__44_, chained_data_delayed_41__43_, chained_data_delayed_41__42_, chained_data_delayed_41__41_, chained_data_delayed_41__40_, chained_data_delayed_41__39_, chained_data_delayed_41__38_, chained_data_delayed_41__37_, chained_data_delayed_41__36_, chained_data_delayed_41__35_, chained_data_delayed_41__34_, chained_data_delayed_41__33_, chained_data_delayed_41__32_, chained_data_delayed_41__31_, chained_data_delayed_41__30_, chained_data_delayed_41__29_, chained_data_delayed_41__28_, chained_data_delayed_41__27_, chained_data_delayed_41__26_, chained_data_delayed_41__25_, chained_data_delayed_41__24_, chained_data_delayed_41__23_, chained_data_delayed_41__22_, chained_data_delayed_41__21_, chained_data_delayed_41__20_, chained_data_delayed_41__19_, chained_data_delayed_41__18_, chained_data_delayed_41__17_, chained_data_delayed_41__16_, chained_data_delayed_41__15_, chained_data_delayed_41__14_, chained_data_delayed_41__13_, chained_data_delayed_41__12_, chained_data_delayed_41__11_, chained_data_delayed_41__10_, chained_data_delayed_41__9_, chained_data_delayed_41__8_, chained_data_delayed_41__7_, chained_data_delayed_41__6_, chained_data_delayed_41__5_, chained_data_delayed_41__4_, chained_data_delayed_41__3_, chained_data_delayed_41__2_, chained_data_delayed_41__1_, chained_data_delayed_41__0_ }),
    .data_o({ chained_data_delayed_42__63_, chained_data_delayed_42__62_, chained_data_delayed_42__61_, chained_data_delayed_42__60_, chained_data_delayed_42__59_, chained_data_delayed_42__58_, chained_data_delayed_42__57_, chained_data_delayed_42__56_, chained_data_delayed_42__55_, chained_data_delayed_42__54_, chained_data_delayed_42__53_, chained_data_delayed_42__52_, chained_data_delayed_42__51_, chained_data_delayed_42__50_, chained_data_delayed_42__49_, chained_data_delayed_42__48_, chained_data_delayed_42__47_, chained_data_delayed_42__46_, chained_data_delayed_42__45_, chained_data_delayed_42__44_, chained_data_delayed_42__43_, chained_data_delayed_42__42_, chained_data_delayed_42__41_, chained_data_delayed_42__40_, chained_data_delayed_42__39_, chained_data_delayed_42__38_, chained_data_delayed_42__37_, chained_data_delayed_42__36_, chained_data_delayed_42__35_, chained_data_delayed_42__34_, chained_data_delayed_42__33_, chained_data_delayed_42__32_, chained_data_delayed_42__31_, chained_data_delayed_42__30_, chained_data_delayed_42__29_, chained_data_delayed_42__28_, chained_data_delayed_42__27_, chained_data_delayed_42__26_, chained_data_delayed_42__25_, chained_data_delayed_42__24_, chained_data_delayed_42__23_, chained_data_delayed_42__22_, chained_data_delayed_42__21_, chained_data_delayed_42__20_, chained_data_delayed_42__19_, chained_data_delayed_42__18_, chained_data_delayed_42__17_, chained_data_delayed_42__16_, chained_data_delayed_42__15_, chained_data_delayed_42__14_, chained_data_delayed_42__13_, chained_data_delayed_42__12_, chained_data_delayed_42__11_, chained_data_delayed_42__10_, chained_data_delayed_42__9_, chained_data_delayed_42__8_, chained_data_delayed_42__7_, chained_data_delayed_42__6_, chained_data_delayed_42__5_, chained_data_delayed_42__4_, chained_data_delayed_42__3_, chained_data_delayed_42__2_, chained_data_delayed_42__1_, chained_data_delayed_42__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_43__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_42__63_, chained_data_delayed_42__62_, chained_data_delayed_42__61_, chained_data_delayed_42__60_, chained_data_delayed_42__59_, chained_data_delayed_42__58_, chained_data_delayed_42__57_, chained_data_delayed_42__56_, chained_data_delayed_42__55_, chained_data_delayed_42__54_, chained_data_delayed_42__53_, chained_data_delayed_42__52_, chained_data_delayed_42__51_, chained_data_delayed_42__50_, chained_data_delayed_42__49_, chained_data_delayed_42__48_, chained_data_delayed_42__47_, chained_data_delayed_42__46_, chained_data_delayed_42__45_, chained_data_delayed_42__44_, chained_data_delayed_42__43_, chained_data_delayed_42__42_, chained_data_delayed_42__41_, chained_data_delayed_42__40_, chained_data_delayed_42__39_, chained_data_delayed_42__38_, chained_data_delayed_42__37_, chained_data_delayed_42__36_, chained_data_delayed_42__35_, chained_data_delayed_42__34_, chained_data_delayed_42__33_, chained_data_delayed_42__32_, chained_data_delayed_42__31_, chained_data_delayed_42__30_, chained_data_delayed_42__29_, chained_data_delayed_42__28_, chained_data_delayed_42__27_, chained_data_delayed_42__26_, chained_data_delayed_42__25_, chained_data_delayed_42__24_, chained_data_delayed_42__23_, chained_data_delayed_42__22_, chained_data_delayed_42__21_, chained_data_delayed_42__20_, chained_data_delayed_42__19_, chained_data_delayed_42__18_, chained_data_delayed_42__17_, chained_data_delayed_42__16_, chained_data_delayed_42__15_, chained_data_delayed_42__14_, chained_data_delayed_42__13_, chained_data_delayed_42__12_, chained_data_delayed_42__11_, chained_data_delayed_42__10_, chained_data_delayed_42__9_, chained_data_delayed_42__8_, chained_data_delayed_42__7_, chained_data_delayed_42__6_, chained_data_delayed_42__5_, chained_data_delayed_42__4_, chained_data_delayed_42__3_, chained_data_delayed_42__2_, chained_data_delayed_42__1_, chained_data_delayed_42__0_ }),
    .data_o({ chained_data_delayed_43__63_, chained_data_delayed_43__62_, chained_data_delayed_43__61_, chained_data_delayed_43__60_, chained_data_delayed_43__59_, chained_data_delayed_43__58_, chained_data_delayed_43__57_, chained_data_delayed_43__56_, chained_data_delayed_43__55_, chained_data_delayed_43__54_, chained_data_delayed_43__53_, chained_data_delayed_43__52_, chained_data_delayed_43__51_, chained_data_delayed_43__50_, chained_data_delayed_43__49_, chained_data_delayed_43__48_, chained_data_delayed_43__47_, chained_data_delayed_43__46_, chained_data_delayed_43__45_, chained_data_delayed_43__44_, chained_data_delayed_43__43_, chained_data_delayed_43__42_, chained_data_delayed_43__41_, chained_data_delayed_43__40_, chained_data_delayed_43__39_, chained_data_delayed_43__38_, chained_data_delayed_43__37_, chained_data_delayed_43__36_, chained_data_delayed_43__35_, chained_data_delayed_43__34_, chained_data_delayed_43__33_, chained_data_delayed_43__32_, chained_data_delayed_43__31_, chained_data_delayed_43__30_, chained_data_delayed_43__29_, chained_data_delayed_43__28_, chained_data_delayed_43__27_, chained_data_delayed_43__26_, chained_data_delayed_43__25_, chained_data_delayed_43__24_, chained_data_delayed_43__23_, chained_data_delayed_43__22_, chained_data_delayed_43__21_, chained_data_delayed_43__20_, chained_data_delayed_43__19_, chained_data_delayed_43__18_, chained_data_delayed_43__17_, chained_data_delayed_43__16_, chained_data_delayed_43__15_, chained_data_delayed_43__14_, chained_data_delayed_43__13_, chained_data_delayed_43__12_, chained_data_delayed_43__11_, chained_data_delayed_43__10_, chained_data_delayed_43__9_, chained_data_delayed_43__8_, chained_data_delayed_43__7_, chained_data_delayed_43__6_, chained_data_delayed_43__5_, chained_data_delayed_43__4_, chained_data_delayed_43__3_, chained_data_delayed_43__2_, chained_data_delayed_43__1_, chained_data_delayed_43__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_44__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_43__63_, chained_data_delayed_43__62_, chained_data_delayed_43__61_, chained_data_delayed_43__60_, chained_data_delayed_43__59_, chained_data_delayed_43__58_, chained_data_delayed_43__57_, chained_data_delayed_43__56_, chained_data_delayed_43__55_, chained_data_delayed_43__54_, chained_data_delayed_43__53_, chained_data_delayed_43__52_, chained_data_delayed_43__51_, chained_data_delayed_43__50_, chained_data_delayed_43__49_, chained_data_delayed_43__48_, chained_data_delayed_43__47_, chained_data_delayed_43__46_, chained_data_delayed_43__45_, chained_data_delayed_43__44_, chained_data_delayed_43__43_, chained_data_delayed_43__42_, chained_data_delayed_43__41_, chained_data_delayed_43__40_, chained_data_delayed_43__39_, chained_data_delayed_43__38_, chained_data_delayed_43__37_, chained_data_delayed_43__36_, chained_data_delayed_43__35_, chained_data_delayed_43__34_, chained_data_delayed_43__33_, chained_data_delayed_43__32_, chained_data_delayed_43__31_, chained_data_delayed_43__30_, chained_data_delayed_43__29_, chained_data_delayed_43__28_, chained_data_delayed_43__27_, chained_data_delayed_43__26_, chained_data_delayed_43__25_, chained_data_delayed_43__24_, chained_data_delayed_43__23_, chained_data_delayed_43__22_, chained_data_delayed_43__21_, chained_data_delayed_43__20_, chained_data_delayed_43__19_, chained_data_delayed_43__18_, chained_data_delayed_43__17_, chained_data_delayed_43__16_, chained_data_delayed_43__15_, chained_data_delayed_43__14_, chained_data_delayed_43__13_, chained_data_delayed_43__12_, chained_data_delayed_43__11_, chained_data_delayed_43__10_, chained_data_delayed_43__9_, chained_data_delayed_43__8_, chained_data_delayed_43__7_, chained_data_delayed_43__6_, chained_data_delayed_43__5_, chained_data_delayed_43__4_, chained_data_delayed_43__3_, chained_data_delayed_43__2_, chained_data_delayed_43__1_, chained_data_delayed_43__0_ }),
    .data_o({ chained_data_delayed_44__63_, chained_data_delayed_44__62_, chained_data_delayed_44__61_, chained_data_delayed_44__60_, chained_data_delayed_44__59_, chained_data_delayed_44__58_, chained_data_delayed_44__57_, chained_data_delayed_44__56_, chained_data_delayed_44__55_, chained_data_delayed_44__54_, chained_data_delayed_44__53_, chained_data_delayed_44__52_, chained_data_delayed_44__51_, chained_data_delayed_44__50_, chained_data_delayed_44__49_, chained_data_delayed_44__48_, chained_data_delayed_44__47_, chained_data_delayed_44__46_, chained_data_delayed_44__45_, chained_data_delayed_44__44_, chained_data_delayed_44__43_, chained_data_delayed_44__42_, chained_data_delayed_44__41_, chained_data_delayed_44__40_, chained_data_delayed_44__39_, chained_data_delayed_44__38_, chained_data_delayed_44__37_, chained_data_delayed_44__36_, chained_data_delayed_44__35_, chained_data_delayed_44__34_, chained_data_delayed_44__33_, chained_data_delayed_44__32_, chained_data_delayed_44__31_, chained_data_delayed_44__30_, chained_data_delayed_44__29_, chained_data_delayed_44__28_, chained_data_delayed_44__27_, chained_data_delayed_44__26_, chained_data_delayed_44__25_, chained_data_delayed_44__24_, chained_data_delayed_44__23_, chained_data_delayed_44__22_, chained_data_delayed_44__21_, chained_data_delayed_44__20_, chained_data_delayed_44__19_, chained_data_delayed_44__18_, chained_data_delayed_44__17_, chained_data_delayed_44__16_, chained_data_delayed_44__15_, chained_data_delayed_44__14_, chained_data_delayed_44__13_, chained_data_delayed_44__12_, chained_data_delayed_44__11_, chained_data_delayed_44__10_, chained_data_delayed_44__9_, chained_data_delayed_44__8_, chained_data_delayed_44__7_, chained_data_delayed_44__6_, chained_data_delayed_44__5_, chained_data_delayed_44__4_, chained_data_delayed_44__3_, chained_data_delayed_44__2_, chained_data_delayed_44__1_, chained_data_delayed_44__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_45__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_44__63_, chained_data_delayed_44__62_, chained_data_delayed_44__61_, chained_data_delayed_44__60_, chained_data_delayed_44__59_, chained_data_delayed_44__58_, chained_data_delayed_44__57_, chained_data_delayed_44__56_, chained_data_delayed_44__55_, chained_data_delayed_44__54_, chained_data_delayed_44__53_, chained_data_delayed_44__52_, chained_data_delayed_44__51_, chained_data_delayed_44__50_, chained_data_delayed_44__49_, chained_data_delayed_44__48_, chained_data_delayed_44__47_, chained_data_delayed_44__46_, chained_data_delayed_44__45_, chained_data_delayed_44__44_, chained_data_delayed_44__43_, chained_data_delayed_44__42_, chained_data_delayed_44__41_, chained_data_delayed_44__40_, chained_data_delayed_44__39_, chained_data_delayed_44__38_, chained_data_delayed_44__37_, chained_data_delayed_44__36_, chained_data_delayed_44__35_, chained_data_delayed_44__34_, chained_data_delayed_44__33_, chained_data_delayed_44__32_, chained_data_delayed_44__31_, chained_data_delayed_44__30_, chained_data_delayed_44__29_, chained_data_delayed_44__28_, chained_data_delayed_44__27_, chained_data_delayed_44__26_, chained_data_delayed_44__25_, chained_data_delayed_44__24_, chained_data_delayed_44__23_, chained_data_delayed_44__22_, chained_data_delayed_44__21_, chained_data_delayed_44__20_, chained_data_delayed_44__19_, chained_data_delayed_44__18_, chained_data_delayed_44__17_, chained_data_delayed_44__16_, chained_data_delayed_44__15_, chained_data_delayed_44__14_, chained_data_delayed_44__13_, chained_data_delayed_44__12_, chained_data_delayed_44__11_, chained_data_delayed_44__10_, chained_data_delayed_44__9_, chained_data_delayed_44__8_, chained_data_delayed_44__7_, chained_data_delayed_44__6_, chained_data_delayed_44__5_, chained_data_delayed_44__4_, chained_data_delayed_44__3_, chained_data_delayed_44__2_, chained_data_delayed_44__1_, chained_data_delayed_44__0_ }),
    .data_o({ chained_data_delayed_45__63_, chained_data_delayed_45__62_, chained_data_delayed_45__61_, chained_data_delayed_45__60_, chained_data_delayed_45__59_, chained_data_delayed_45__58_, chained_data_delayed_45__57_, chained_data_delayed_45__56_, chained_data_delayed_45__55_, chained_data_delayed_45__54_, chained_data_delayed_45__53_, chained_data_delayed_45__52_, chained_data_delayed_45__51_, chained_data_delayed_45__50_, chained_data_delayed_45__49_, chained_data_delayed_45__48_, chained_data_delayed_45__47_, chained_data_delayed_45__46_, chained_data_delayed_45__45_, chained_data_delayed_45__44_, chained_data_delayed_45__43_, chained_data_delayed_45__42_, chained_data_delayed_45__41_, chained_data_delayed_45__40_, chained_data_delayed_45__39_, chained_data_delayed_45__38_, chained_data_delayed_45__37_, chained_data_delayed_45__36_, chained_data_delayed_45__35_, chained_data_delayed_45__34_, chained_data_delayed_45__33_, chained_data_delayed_45__32_, chained_data_delayed_45__31_, chained_data_delayed_45__30_, chained_data_delayed_45__29_, chained_data_delayed_45__28_, chained_data_delayed_45__27_, chained_data_delayed_45__26_, chained_data_delayed_45__25_, chained_data_delayed_45__24_, chained_data_delayed_45__23_, chained_data_delayed_45__22_, chained_data_delayed_45__21_, chained_data_delayed_45__20_, chained_data_delayed_45__19_, chained_data_delayed_45__18_, chained_data_delayed_45__17_, chained_data_delayed_45__16_, chained_data_delayed_45__15_, chained_data_delayed_45__14_, chained_data_delayed_45__13_, chained_data_delayed_45__12_, chained_data_delayed_45__11_, chained_data_delayed_45__10_, chained_data_delayed_45__9_, chained_data_delayed_45__8_, chained_data_delayed_45__7_, chained_data_delayed_45__6_, chained_data_delayed_45__5_, chained_data_delayed_45__4_, chained_data_delayed_45__3_, chained_data_delayed_45__2_, chained_data_delayed_45__1_, chained_data_delayed_45__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_46__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_45__63_, chained_data_delayed_45__62_, chained_data_delayed_45__61_, chained_data_delayed_45__60_, chained_data_delayed_45__59_, chained_data_delayed_45__58_, chained_data_delayed_45__57_, chained_data_delayed_45__56_, chained_data_delayed_45__55_, chained_data_delayed_45__54_, chained_data_delayed_45__53_, chained_data_delayed_45__52_, chained_data_delayed_45__51_, chained_data_delayed_45__50_, chained_data_delayed_45__49_, chained_data_delayed_45__48_, chained_data_delayed_45__47_, chained_data_delayed_45__46_, chained_data_delayed_45__45_, chained_data_delayed_45__44_, chained_data_delayed_45__43_, chained_data_delayed_45__42_, chained_data_delayed_45__41_, chained_data_delayed_45__40_, chained_data_delayed_45__39_, chained_data_delayed_45__38_, chained_data_delayed_45__37_, chained_data_delayed_45__36_, chained_data_delayed_45__35_, chained_data_delayed_45__34_, chained_data_delayed_45__33_, chained_data_delayed_45__32_, chained_data_delayed_45__31_, chained_data_delayed_45__30_, chained_data_delayed_45__29_, chained_data_delayed_45__28_, chained_data_delayed_45__27_, chained_data_delayed_45__26_, chained_data_delayed_45__25_, chained_data_delayed_45__24_, chained_data_delayed_45__23_, chained_data_delayed_45__22_, chained_data_delayed_45__21_, chained_data_delayed_45__20_, chained_data_delayed_45__19_, chained_data_delayed_45__18_, chained_data_delayed_45__17_, chained_data_delayed_45__16_, chained_data_delayed_45__15_, chained_data_delayed_45__14_, chained_data_delayed_45__13_, chained_data_delayed_45__12_, chained_data_delayed_45__11_, chained_data_delayed_45__10_, chained_data_delayed_45__9_, chained_data_delayed_45__8_, chained_data_delayed_45__7_, chained_data_delayed_45__6_, chained_data_delayed_45__5_, chained_data_delayed_45__4_, chained_data_delayed_45__3_, chained_data_delayed_45__2_, chained_data_delayed_45__1_, chained_data_delayed_45__0_ }),
    .data_o({ chained_data_delayed_46__63_, chained_data_delayed_46__62_, chained_data_delayed_46__61_, chained_data_delayed_46__60_, chained_data_delayed_46__59_, chained_data_delayed_46__58_, chained_data_delayed_46__57_, chained_data_delayed_46__56_, chained_data_delayed_46__55_, chained_data_delayed_46__54_, chained_data_delayed_46__53_, chained_data_delayed_46__52_, chained_data_delayed_46__51_, chained_data_delayed_46__50_, chained_data_delayed_46__49_, chained_data_delayed_46__48_, chained_data_delayed_46__47_, chained_data_delayed_46__46_, chained_data_delayed_46__45_, chained_data_delayed_46__44_, chained_data_delayed_46__43_, chained_data_delayed_46__42_, chained_data_delayed_46__41_, chained_data_delayed_46__40_, chained_data_delayed_46__39_, chained_data_delayed_46__38_, chained_data_delayed_46__37_, chained_data_delayed_46__36_, chained_data_delayed_46__35_, chained_data_delayed_46__34_, chained_data_delayed_46__33_, chained_data_delayed_46__32_, chained_data_delayed_46__31_, chained_data_delayed_46__30_, chained_data_delayed_46__29_, chained_data_delayed_46__28_, chained_data_delayed_46__27_, chained_data_delayed_46__26_, chained_data_delayed_46__25_, chained_data_delayed_46__24_, chained_data_delayed_46__23_, chained_data_delayed_46__22_, chained_data_delayed_46__21_, chained_data_delayed_46__20_, chained_data_delayed_46__19_, chained_data_delayed_46__18_, chained_data_delayed_46__17_, chained_data_delayed_46__16_, chained_data_delayed_46__15_, chained_data_delayed_46__14_, chained_data_delayed_46__13_, chained_data_delayed_46__12_, chained_data_delayed_46__11_, chained_data_delayed_46__10_, chained_data_delayed_46__9_, chained_data_delayed_46__8_, chained_data_delayed_46__7_, chained_data_delayed_46__6_, chained_data_delayed_46__5_, chained_data_delayed_46__4_, chained_data_delayed_46__3_, chained_data_delayed_46__2_, chained_data_delayed_46__1_, chained_data_delayed_46__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_47__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_46__63_, chained_data_delayed_46__62_, chained_data_delayed_46__61_, chained_data_delayed_46__60_, chained_data_delayed_46__59_, chained_data_delayed_46__58_, chained_data_delayed_46__57_, chained_data_delayed_46__56_, chained_data_delayed_46__55_, chained_data_delayed_46__54_, chained_data_delayed_46__53_, chained_data_delayed_46__52_, chained_data_delayed_46__51_, chained_data_delayed_46__50_, chained_data_delayed_46__49_, chained_data_delayed_46__48_, chained_data_delayed_46__47_, chained_data_delayed_46__46_, chained_data_delayed_46__45_, chained_data_delayed_46__44_, chained_data_delayed_46__43_, chained_data_delayed_46__42_, chained_data_delayed_46__41_, chained_data_delayed_46__40_, chained_data_delayed_46__39_, chained_data_delayed_46__38_, chained_data_delayed_46__37_, chained_data_delayed_46__36_, chained_data_delayed_46__35_, chained_data_delayed_46__34_, chained_data_delayed_46__33_, chained_data_delayed_46__32_, chained_data_delayed_46__31_, chained_data_delayed_46__30_, chained_data_delayed_46__29_, chained_data_delayed_46__28_, chained_data_delayed_46__27_, chained_data_delayed_46__26_, chained_data_delayed_46__25_, chained_data_delayed_46__24_, chained_data_delayed_46__23_, chained_data_delayed_46__22_, chained_data_delayed_46__21_, chained_data_delayed_46__20_, chained_data_delayed_46__19_, chained_data_delayed_46__18_, chained_data_delayed_46__17_, chained_data_delayed_46__16_, chained_data_delayed_46__15_, chained_data_delayed_46__14_, chained_data_delayed_46__13_, chained_data_delayed_46__12_, chained_data_delayed_46__11_, chained_data_delayed_46__10_, chained_data_delayed_46__9_, chained_data_delayed_46__8_, chained_data_delayed_46__7_, chained_data_delayed_46__6_, chained_data_delayed_46__5_, chained_data_delayed_46__4_, chained_data_delayed_46__3_, chained_data_delayed_46__2_, chained_data_delayed_46__1_, chained_data_delayed_46__0_ }),
    .data_o({ chained_data_delayed_47__63_, chained_data_delayed_47__62_, chained_data_delayed_47__61_, chained_data_delayed_47__60_, chained_data_delayed_47__59_, chained_data_delayed_47__58_, chained_data_delayed_47__57_, chained_data_delayed_47__56_, chained_data_delayed_47__55_, chained_data_delayed_47__54_, chained_data_delayed_47__53_, chained_data_delayed_47__52_, chained_data_delayed_47__51_, chained_data_delayed_47__50_, chained_data_delayed_47__49_, chained_data_delayed_47__48_, chained_data_delayed_47__47_, chained_data_delayed_47__46_, chained_data_delayed_47__45_, chained_data_delayed_47__44_, chained_data_delayed_47__43_, chained_data_delayed_47__42_, chained_data_delayed_47__41_, chained_data_delayed_47__40_, chained_data_delayed_47__39_, chained_data_delayed_47__38_, chained_data_delayed_47__37_, chained_data_delayed_47__36_, chained_data_delayed_47__35_, chained_data_delayed_47__34_, chained_data_delayed_47__33_, chained_data_delayed_47__32_, chained_data_delayed_47__31_, chained_data_delayed_47__30_, chained_data_delayed_47__29_, chained_data_delayed_47__28_, chained_data_delayed_47__27_, chained_data_delayed_47__26_, chained_data_delayed_47__25_, chained_data_delayed_47__24_, chained_data_delayed_47__23_, chained_data_delayed_47__22_, chained_data_delayed_47__21_, chained_data_delayed_47__20_, chained_data_delayed_47__19_, chained_data_delayed_47__18_, chained_data_delayed_47__17_, chained_data_delayed_47__16_, chained_data_delayed_47__15_, chained_data_delayed_47__14_, chained_data_delayed_47__13_, chained_data_delayed_47__12_, chained_data_delayed_47__11_, chained_data_delayed_47__10_, chained_data_delayed_47__9_, chained_data_delayed_47__8_, chained_data_delayed_47__7_, chained_data_delayed_47__6_, chained_data_delayed_47__5_, chained_data_delayed_47__4_, chained_data_delayed_47__3_, chained_data_delayed_47__2_, chained_data_delayed_47__1_, chained_data_delayed_47__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_48__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_47__63_, chained_data_delayed_47__62_, chained_data_delayed_47__61_, chained_data_delayed_47__60_, chained_data_delayed_47__59_, chained_data_delayed_47__58_, chained_data_delayed_47__57_, chained_data_delayed_47__56_, chained_data_delayed_47__55_, chained_data_delayed_47__54_, chained_data_delayed_47__53_, chained_data_delayed_47__52_, chained_data_delayed_47__51_, chained_data_delayed_47__50_, chained_data_delayed_47__49_, chained_data_delayed_47__48_, chained_data_delayed_47__47_, chained_data_delayed_47__46_, chained_data_delayed_47__45_, chained_data_delayed_47__44_, chained_data_delayed_47__43_, chained_data_delayed_47__42_, chained_data_delayed_47__41_, chained_data_delayed_47__40_, chained_data_delayed_47__39_, chained_data_delayed_47__38_, chained_data_delayed_47__37_, chained_data_delayed_47__36_, chained_data_delayed_47__35_, chained_data_delayed_47__34_, chained_data_delayed_47__33_, chained_data_delayed_47__32_, chained_data_delayed_47__31_, chained_data_delayed_47__30_, chained_data_delayed_47__29_, chained_data_delayed_47__28_, chained_data_delayed_47__27_, chained_data_delayed_47__26_, chained_data_delayed_47__25_, chained_data_delayed_47__24_, chained_data_delayed_47__23_, chained_data_delayed_47__22_, chained_data_delayed_47__21_, chained_data_delayed_47__20_, chained_data_delayed_47__19_, chained_data_delayed_47__18_, chained_data_delayed_47__17_, chained_data_delayed_47__16_, chained_data_delayed_47__15_, chained_data_delayed_47__14_, chained_data_delayed_47__13_, chained_data_delayed_47__12_, chained_data_delayed_47__11_, chained_data_delayed_47__10_, chained_data_delayed_47__9_, chained_data_delayed_47__8_, chained_data_delayed_47__7_, chained_data_delayed_47__6_, chained_data_delayed_47__5_, chained_data_delayed_47__4_, chained_data_delayed_47__3_, chained_data_delayed_47__2_, chained_data_delayed_47__1_, chained_data_delayed_47__0_ }),
    .data_o({ chained_data_delayed_48__63_, chained_data_delayed_48__62_, chained_data_delayed_48__61_, chained_data_delayed_48__60_, chained_data_delayed_48__59_, chained_data_delayed_48__58_, chained_data_delayed_48__57_, chained_data_delayed_48__56_, chained_data_delayed_48__55_, chained_data_delayed_48__54_, chained_data_delayed_48__53_, chained_data_delayed_48__52_, chained_data_delayed_48__51_, chained_data_delayed_48__50_, chained_data_delayed_48__49_, chained_data_delayed_48__48_, chained_data_delayed_48__47_, chained_data_delayed_48__46_, chained_data_delayed_48__45_, chained_data_delayed_48__44_, chained_data_delayed_48__43_, chained_data_delayed_48__42_, chained_data_delayed_48__41_, chained_data_delayed_48__40_, chained_data_delayed_48__39_, chained_data_delayed_48__38_, chained_data_delayed_48__37_, chained_data_delayed_48__36_, chained_data_delayed_48__35_, chained_data_delayed_48__34_, chained_data_delayed_48__33_, chained_data_delayed_48__32_, chained_data_delayed_48__31_, chained_data_delayed_48__30_, chained_data_delayed_48__29_, chained_data_delayed_48__28_, chained_data_delayed_48__27_, chained_data_delayed_48__26_, chained_data_delayed_48__25_, chained_data_delayed_48__24_, chained_data_delayed_48__23_, chained_data_delayed_48__22_, chained_data_delayed_48__21_, chained_data_delayed_48__20_, chained_data_delayed_48__19_, chained_data_delayed_48__18_, chained_data_delayed_48__17_, chained_data_delayed_48__16_, chained_data_delayed_48__15_, chained_data_delayed_48__14_, chained_data_delayed_48__13_, chained_data_delayed_48__12_, chained_data_delayed_48__11_, chained_data_delayed_48__10_, chained_data_delayed_48__9_, chained_data_delayed_48__8_, chained_data_delayed_48__7_, chained_data_delayed_48__6_, chained_data_delayed_48__5_, chained_data_delayed_48__4_, chained_data_delayed_48__3_, chained_data_delayed_48__2_, chained_data_delayed_48__1_, chained_data_delayed_48__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_49__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_48__63_, chained_data_delayed_48__62_, chained_data_delayed_48__61_, chained_data_delayed_48__60_, chained_data_delayed_48__59_, chained_data_delayed_48__58_, chained_data_delayed_48__57_, chained_data_delayed_48__56_, chained_data_delayed_48__55_, chained_data_delayed_48__54_, chained_data_delayed_48__53_, chained_data_delayed_48__52_, chained_data_delayed_48__51_, chained_data_delayed_48__50_, chained_data_delayed_48__49_, chained_data_delayed_48__48_, chained_data_delayed_48__47_, chained_data_delayed_48__46_, chained_data_delayed_48__45_, chained_data_delayed_48__44_, chained_data_delayed_48__43_, chained_data_delayed_48__42_, chained_data_delayed_48__41_, chained_data_delayed_48__40_, chained_data_delayed_48__39_, chained_data_delayed_48__38_, chained_data_delayed_48__37_, chained_data_delayed_48__36_, chained_data_delayed_48__35_, chained_data_delayed_48__34_, chained_data_delayed_48__33_, chained_data_delayed_48__32_, chained_data_delayed_48__31_, chained_data_delayed_48__30_, chained_data_delayed_48__29_, chained_data_delayed_48__28_, chained_data_delayed_48__27_, chained_data_delayed_48__26_, chained_data_delayed_48__25_, chained_data_delayed_48__24_, chained_data_delayed_48__23_, chained_data_delayed_48__22_, chained_data_delayed_48__21_, chained_data_delayed_48__20_, chained_data_delayed_48__19_, chained_data_delayed_48__18_, chained_data_delayed_48__17_, chained_data_delayed_48__16_, chained_data_delayed_48__15_, chained_data_delayed_48__14_, chained_data_delayed_48__13_, chained_data_delayed_48__12_, chained_data_delayed_48__11_, chained_data_delayed_48__10_, chained_data_delayed_48__9_, chained_data_delayed_48__8_, chained_data_delayed_48__7_, chained_data_delayed_48__6_, chained_data_delayed_48__5_, chained_data_delayed_48__4_, chained_data_delayed_48__3_, chained_data_delayed_48__2_, chained_data_delayed_48__1_, chained_data_delayed_48__0_ }),
    .data_o({ chained_data_delayed_49__63_, chained_data_delayed_49__62_, chained_data_delayed_49__61_, chained_data_delayed_49__60_, chained_data_delayed_49__59_, chained_data_delayed_49__58_, chained_data_delayed_49__57_, chained_data_delayed_49__56_, chained_data_delayed_49__55_, chained_data_delayed_49__54_, chained_data_delayed_49__53_, chained_data_delayed_49__52_, chained_data_delayed_49__51_, chained_data_delayed_49__50_, chained_data_delayed_49__49_, chained_data_delayed_49__48_, chained_data_delayed_49__47_, chained_data_delayed_49__46_, chained_data_delayed_49__45_, chained_data_delayed_49__44_, chained_data_delayed_49__43_, chained_data_delayed_49__42_, chained_data_delayed_49__41_, chained_data_delayed_49__40_, chained_data_delayed_49__39_, chained_data_delayed_49__38_, chained_data_delayed_49__37_, chained_data_delayed_49__36_, chained_data_delayed_49__35_, chained_data_delayed_49__34_, chained_data_delayed_49__33_, chained_data_delayed_49__32_, chained_data_delayed_49__31_, chained_data_delayed_49__30_, chained_data_delayed_49__29_, chained_data_delayed_49__28_, chained_data_delayed_49__27_, chained_data_delayed_49__26_, chained_data_delayed_49__25_, chained_data_delayed_49__24_, chained_data_delayed_49__23_, chained_data_delayed_49__22_, chained_data_delayed_49__21_, chained_data_delayed_49__20_, chained_data_delayed_49__19_, chained_data_delayed_49__18_, chained_data_delayed_49__17_, chained_data_delayed_49__16_, chained_data_delayed_49__15_, chained_data_delayed_49__14_, chained_data_delayed_49__13_, chained_data_delayed_49__12_, chained_data_delayed_49__11_, chained_data_delayed_49__10_, chained_data_delayed_49__9_, chained_data_delayed_49__8_, chained_data_delayed_49__7_, chained_data_delayed_49__6_, chained_data_delayed_49__5_, chained_data_delayed_49__4_, chained_data_delayed_49__3_, chained_data_delayed_49__2_, chained_data_delayed_49__1_, chained_data_delayed_49__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_50__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_49__63_, chained_data_delayed_49__62_, chained_data_delayed_49__61_, chained_data_delayed_49__60_, chained_data_delayed_49__59_, chained_data_delayed_49__58_, chained_data_delayed_49__57_, chained_data_delayed_49__56_, chained_data_delayed_49__55_, chained_data_delayed_49__54_, chained_data_delayed_49__53_, chained_data_delayed_49__52_, chained_data_delayed_49__51_, chained_data_delayed_49__50_, chained_data_delayed_49__49_, chained_data_delayed_49__48_, chained_data_delayed_49__47_, chained_data_delayed_49__46_, chained_data_delayed_49__45_, chained_data_delayed_49__44_, chained_data_delayed_49__43_, chained_data_delayed_49__42_, chained_data_delayed_49__41_, chained_data_delayed_49__40_, chained_data_delayed_49__39_, chained_data_delayed_49__38_, chained_data_delayed_49__37_, chained_data_delayed_49__36_, chained_data_delayed_49__35_, chained_data_delayed_49__34_, chained_data_delayed_49__33_, chained_data_delayed_49__32_, chained_data_delayed_49__31_, chained_data_delayed_49__30_, chained_data_delayed_49__29_, chained_data_delayed_49__28_, chained_data_delayed_49__27_, chained_data_delayed_49__26_, chained_data_delayed_49__25_, chained_data_delayed_49__24_, chained_data_delayed_49__23_, chained_data_delayed_49__22_, chained_data_delayed_49__21_, chained_data_delayed_49__20_, chained_data_delayed_49__19_, chained_data_delayed_49__18_, chained_data_delayed_49__17_, chained_data_delayed_49__16_, chained_data_delayed_49__15_, chained_data_delayed_49__14_, chained_data_delayed_49__13_, chained_data_delayed_49__12_, chained_data_delayed_49__11_, chained_data_delayed_49__10_, chained_data_delayed_49__9_, chained_data_delayed_49__8_, chained_data_delayed_49__7_, chained_data_delayed_49__6_, chained_data_delayed_49__5_, chained_data_delayed_49__4_, chained_data_delayed_49__3_, chained_data_delayed_49__2_, chained_data_delayed_49__1_, chained_data_delayed_49__0_ }),
    .data_o({ chained_data_delayed_50__63_, chained_data_delayed_50__62_, chained_data_delayed_50__61_, chained_data_delayed_50__60_, chained_data_delayed_50__59_, chained_data_delayed_50__58_, chained_data_delayed_50__57_, chained_data_delayed_50__56_, chained_data_delayed_50__55_, chained_data_delayed_50__54_, chained_data_delayed_50__53_, chained_data_delayed_50__52_, chained_data_delayed_50__51_, chained_data_delayed_50__50_, chained_data_delayed_50__49_, chained_data_delayed_50__48_, chained_data_delayed_50__47_, chained_data_delayed_50__46_, chained_data_delayed_50__45_, chained_data_delayed_50__44_, chained_data_delayed_50__43_, chained_data_delayed_50__42_, chained_data_delayed_50__41_, chained_data_delayed_50__40_, chained_data_delayed_50__39_, chained_data_delayed_50__38_, chained_data_delayed_50__37_, chained_data_delayed_50__36_, chained_data_delayed_50__35_, chained_data_delayed_50__34_, chained_data_delayed_50__33_, chained_data_delayed_50__32_, chained_data_delayed_50__31_, chained_data_delayed_50__30_, chained_data_delayed_50__29_, chained_data_delayed_50__28_, chained_data_delayed_50__27_, chained_data_delayed_50__26_, chained_data_delayed_50__25_, chained_data_delayed_50__24_, chained_data_delayed_50__23_, chained_data_delayed_50__22_, chained_data_delayed_50__21_, chained_data_delayed_50__20_, chained_data_delayed_50__19_, chained_data_delayed_50__18_, chained_data_delayed_50__17_, chained_data_delayed_50__16_, chained_data_delayed_50__15_, chained_data_delayed_50__14_, chained_data_delayed_50__13_, chained_data_delayed_50__12_, chained_data_delayed_50__11_, chained_data_delayed_50__10_, chained_data_delayed_50__9_, chained_data_delayed_50__8_, chained_data_delayed_50__7_, chained_data_delayed_50__6_, chained_data_delayed_50__5_, chained_data_delayed_50__4_, chained_data_delayed_50__3_, chained_data_delayed_50__2_, chained_data_delayed_50__1_, chained_data_delayed_50__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_51__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_50__63_, chained_data_delayed_50__62_, chained_data_delayed_50__61_, chained_data_delayed_50__60_, chained_data_delayed_50__59_, chained_data_delayed_50__58_, chained_data_delayed_50__57_, chained_data_delayed_50__56_, chained_data_delayed_50__55_, chained_data_delayed_50__54_, chained_data_delayed_50__53_, chained_data_delayed_50__52_, chained_data_delayed_50__51_, chained_data_delayed_50__50_, chained_data_delayed_50__49_, chained_data_delayed_50__48_, chained_data_delayed_50__47_, chained_data_delayed_50__46_, chained_data_delayed_50__45_, chained_data_delayed_50__44_, chained_data_delayed_50__43_, chained_data_delayed_50__42_, chained_data_delayed_50__41_, chained_data_delayed_50__40_, chained_data_delayed_50__39_, chained_data_delayed_50__38_, chained_data_delayed_50__37_, chained_data_delayed_50__36_, chained_data_delayed_50__35_, chained_data_delayed_50__34_, chained_data_delayed_50__33_, chained_data_delayed_50__32_, chained_data_delayed_50__31_, chained_data_delayed_50__30_, chained_data_delayed_50__29_, chained_data_delayed_50__28_, chained_data_delayed_50__27_, chained_data_delayed_50__26_, chained_data_delayed_50__25_, chained_data_delayed_50__24_, chained_data_delayed_50__23_, chained_data_delayed_50__22_, chained_data_delayed_50__21_, chained_data_delayed_50__20_, chained_data_delayed_50__19_, chained_data_delayed_50__18_, chained_data_delayed_50__17_, chained_data_delayed_50__16_, chained_data_delayed_50__15_, chained_data_delayed_50__14_, chained_data_delayed_50__13_, chained_data_delayed_50__12_, chained_data_delayed_50__11_, chained_data_delayed_50__10_, chained_data_delayed_50__9_, chained_data_delayed_50__8_, chained_data_delayed_50__7_, chained_data_delayed_50__6_, chained_data_delayed_50__5_, chained_data_delayed_50__4_, chained_data_delayed_50__3_, chained_data_delayed_50__2_, chained_data_delayed_50__1_, chained_data_delayed_50__0_ }),
    .data_o({ chained_data_delayed_51__63_, chained_data_delayed_51__62_, chained_data_delayed_51__61_, chained_data_delayed_51__60_, chained_data_delayed_51__59_, chained_data_delayed_51__58_, chained_data_delayed_51__57_, chained_data_delayed_51__56_, chained_data_delayed_51__55_, chained_data_delayed_51__54_, chained_data_delayed_51__53_, chained_data_delayed_51__52_, chained_data_delayed_51__51_, chained_data_delayed_51__50_, chained_data_delayed_51__49_, chained_data_delayed_51__48_, chained_data_delayed_51__47_, chained_data_delayed_51__46_, chained_data_delayed_51__45_, chained_data_delayed_51__44_, chained_data_delayed_51__43_, chained_data_delayed_51__42_, chained_data_delayed_51__41_, chained_data_delayed_51__40_, chained_data_delayed_51__39_, chained_data_delayed_51__38_, chained_data_delayed_51__37_, chained_data_delayed_51__36_, chained_data_delayed_51__35_, chained_data_delayed_51__34_, chained_data_delayed_51__33_, chained_data_delayed_51__32_, chained_data_delayed_51__31_, chained_data_delayed_51__30_, chained_data_delayed_51__29_, chained_data_delayed_51__28_, chained_data_delayed_51__27_, chained_data_delayed_51__26_, chained_data_delayed_51__25_, chained_data_delayed_51__24_, chained_data_delayed_51__23_, chained_data_delayed_51__22_, chained_data_delayed_51__21_, chained_data_delayed_51__20_, chained_data_delayed_51__19_, chained_data_delayed_51__18_, chained_data_delayed_51__17_, chained_data_delayed_51__16_, chained_data_delayed_51__15_, chained_data_delayed_51__14_, chained_data_delayed_51__13_, chained_data_delayed_51__12_, chained_data_delayed_51__11_, chained_data_delayed_51__10_, chained_data_delayed_51__9_, chained_data_delayed_51__8_, chained_data_delayed_51__7_, chained_data_delayed_51__6_, chained_data_delayed_51__5_, chained_data_delayed_51__4_, chained_data_delayed_51__3_, chained_data_delayed_51__2_, chained_data_delayed_51__1_, chained_data_delayed_51__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_52__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_51__63_, chained_data_delayed_51__62_, chained_data_delayed_51__61_, chained_data_delayed_51__60_, chained_data_delayed_51__59_, chained_data_delayed_51__58_, chained_data_delayed_51__57_, chained_data_delayed_51__56_, chained_data_delayed_51__55_, chained_data_delayed_51__54_, chained_data_delayed_51__53_, chained_data_delayed_51__52_, chained_data_delayed_51__51_, chained_data_delayed_51__50_, chained_data_delayed_51__49_, chained_data_delayed_51__48_, chained_data_delayed_51__47_, chained_data_delayed_51__46_, chained_data_delayed_51__45_, chained_data_delayed_51__44_, chained_data_delayed_51__43_, chained_data_delayed_51__42_, chained_data_delayed_51__41_, chained_data_delayed_51__40_, chained_data_delayed_51__39_, chained_data_delayed_51__38_, chained_data_delayed_51__37_, chained_data_delayed_51__36_, chained_data_delayed_51__35_, chained_data_delayed_51__34_, chained_data_delayed_51__33_, chained_data_delayed_51__32_, chained_data_delayed_51__31_, chained_data_delayed_51__30_, chained_data_delayed_51__29_, chained_data_delayed_51__28_, chained_data_delayed_51__27_, chained_data_delayed_51__26_, chained_data_delayed_51__25_, chained_data_delayed_51__24_, chained_data_delayed_51__23_, chained_data_delayed_51__22_, chained_data_delayed_51__21_, chained_data_delayed_51__20_, chained_data_delayed_51__19_, chained_data_delayed_51__18_, chained_data_delayed_51__17_, chained_data_delayed_51__16_, chained_data_delayed_51__15_, chained_data_delayed_51__14_, chained_data_delayed_51__13_, chained_data_delayed_51__12_, chained_data_delayed_51__11_, chained_data_delayed_51__10_, chained_data_delayed_51__9_, chained_data_delayed_51__8_, chained_data_delayed_51__7_, chained_data_delayed_51__6_, chained_data_delayed_51__5_, chained_data_delayed_51__4_, chained_data_delayed_51__3_, chained_data_delayed_51__2_, chained_data_delayed_51__1_, chained_data_delayed_51__0_ }),
    .data_o({ chained_data_delayed_52__63_, chained_data_delayed_52__62_, chained_data_delayed_52__61_, chained_data_delayed_52__60_, chained_data_delayed_52__59_, chained_data_delayed_52__58_, chained_data_delayed_52__57_, chained_data_delayed_52__56_, chained_data_delayed_52__55_, chained_data_delayed_52__54_, chained_data_delayed_52__53_, chained_data_delayed_52__52_, chained_data_delayed_52__51_, chained_data_delayed_52__50_, chained_data_delayed_52__49_, chained_data_delayed_52__48_, chained_data_delayed_52__47_, chained_data_delayed_52__46_, chained_data_delayed_52__45_, chained_data_delayed_52__44_, chained_data_delayed_52__43_, chained_data_delayed_52__42_, chained_data_delayed_52__41_, chained_data_delayed_52__40_, chained_data_delayed_52__39_, chained_data_delayed_52__38_, chained_data_delayed_52__37_, chained_data_delayed_52__36_, chained_data_delayed_52__35_, chained_data_delayed_52__34_, chained_data_delayed_52__33_, chained_data_delayed_52__32_, chained_data_delayed_52__31_, chained_data_delayed_52__30_, chained_data_delayed_52__29_, chained_data_delayed_52__28_, chained_data_delayed_52__27_, chained_data_delayed_52__26_, chained_data_delayed_52__25_, chained_data_delayed_52__24_, chained_data_delayed_52__23_, chained_data_delayed_52__22_, chained_data_delayed_52__21_, chained_data_delayed_52__20_, chained_data_delayed_52__19_, chained_data_delayed_52__18_, chained_data_delayed_52__17_, chained_data_delayed_52__16_, chained_data_delayed_52__15_, chained_data_delayed_52__14_, chained_data_delayed_52__13_, chained_data_delayed_52__12_, chained_data_delayed_52__11_, chained_data_delayed_52__10_, chained_data_delayed_52__9_, chained_data_delayed_52__8_, chained_data_delayed_52__7_, chained_data_delayed_52__6_, chained_data_delayed_52__5_, chained_data_delayed_52__4_, chained_data_delayed_52__3_, chained_data_delayed_52__2_, chained_data_delayed_52__1_, chained_data_delayed_52__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_53__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_52__63_, chained_data_delayed_52__62_, chained_data_delayed_52__61_, chained_data_delayed_52__60_, chained_data_delayed_52__59_, chained_data_delayed_52__58_, chained_data_delayed_52__57_, chained_data_delayed_52__56_, chained_data_delayed_52__55_, chained_data_delayed_52__54_, chained_data_delayed_52__53_, chained_data_delayed_52__52_, chained_data_delayed_52__51_, chained_data_delayed_52__50_, chained_data_delayed_52__49_, chained_data_delayed_52__48_, chained_data_delayed_52__47_, chained_data_delayed_52__46_, chained_data_delayed_52__45_, chained_data_delayed_52__44_, chained_data_delayed_52__43_, chained_data_delayed_52__42_, chained_data_delayed_52__41_, chained_data_delayed_52__40_, chained_data_delayed_52__39_, chained_data_delayed_52__38_, chained_data_delayed_52__37_, chained_data_delayed_52__36_, chained_data_delayed_52__35_, chained_data_delayed_52__34_, chained_data_delayed_52__33_, chained_data_delayed_52__32_, chained_data_delayed_52__31_, chained_data_delayed_52__30_, chained_data_delayed_52__29_, chained_data_delayed_52__28_, chained_data_delayed_52__27_, chained_data_delayed_52__26_, chained_data_delayed_52__25_, chained_data_delayed_52__24_, chained_data_delayed_52__23_, chained_data_delayed_52__22_, chained_data_delayed_52__21_, chained_data_delayed_52__20_, chained_data_delayed_52__19_, chained_data_delayed_52__18_, chained_data_delayed_52__17_, chained_data_delayed_52__16_, chained_data_delayed_52__15_, chained_data_delayed_52__14_, chained_data_delayed_52__13_, chained_data_delayed_52__12_, chained_data_delayed_52__11_, chained_data_delayed_52__10_, chained_data_delayed_52__9_, chained_data_delayed_52__8_, chained_data_delayed_52__7_, chained_data_delayed_52__6_, chained_data_delayed_52__5_, chained_data_delayed_52__4_, chained_data_delayed_52__3_, chained_data_delayed_52__2_, chained_data_delayed_52__1_, chained_data_delayed_52__0_ }),
    .data_o({ chained_data_delayed_53__63_, chained_data_delayed_53__62_, chained_data_delayed_53__61_, chained_data_delayed_53__60_, chained_data_delayed_53__59_, chained_data_delayed_53__58_, chained_data_delayed_53__57_, chained_data_delayed_53__56_, chained_data_delayed_53__55_, chained_data_delayed_53__54_, chained_data_delayed_53__53_, chained_data_delayed_53__52_, chained_data_delayed_53__51_, chained_data_delayed_53__50_, chained_data_delayed_53__49_, chained_data_delayed_53__48_, chained_data_delayed_53__47_, chained_data_delayed_53__46_, chained_data_delayed_53__45_, chained_data_delayed_53__44_, chained_data_delayed_53__43_, chained_data_delayed_53__42_, chained_data_delayed_53__41_, chained_data_delayed_53__40_, chained_data_delayed_53__39_, chained_data_delayed_53__38_, chained_data_delayed_53__37_, chained_data_delayed_53__36_, chained_data_delayed_53__35_, chained_data_delayed_53__34_, chained_data_delayed_53__33_, chained_data_delayed_53__32_, chained_data_delayed_53__31_, chained_data_delayed_53__30_, chained_data_delayed_53__29_, chained_data_delayed_53__28_, chained_data_delayed_53__27_, chained_data_delayed_53__26_, chained_data_delayed_53__25_, chained_data_delayed_53__24_, chained_data_delayed_53__23_, chained_data_delayed_53__22_, chained_data_delayed_53__21_, chained_data_delayed_53__20_, chained_data_delayed_53__19_, chained_data_delayed_53__18_, chained_data_delayed_53__17_, chained_data_delayed_53__16_, chained_data_delayed_53__15_, chained_data_delayed_53__14_, chained_data_delayed_53__13_, chained_data_delayed_53__12_, chained_data_delayed_53__11_, chained_data_delayed_53__10_, chained_data_delayed_53__9_, chained_data_delayed_53__8_, chained_data_delayed_53__7_, chained_data_delayed_53__6_, chained_data_delayed_53__5_, chained_data_delayed_53__4_, chained_data_delayed_53__3_, chained_data_delayed_53__2_, chained_data_delayed_53__1_, chained_data_delayed_53__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_54__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_53__63_, chained_data_delayed_53__62_, chained_data_delayed_53__61_, chained_data_delayed_53__60_, chained_data_delayed_53__59_, chained_data_delayed_53__58_, chained_data_delayed_53__57_, chained_data_delayed_53__56_, chained_data_delayed_53__55_, chained_data_delayed_53__54_, chained_data_delayed_53__53_, chained_data_delayed_53__52_, chained_data_delayed_53__51_, chained_data_delayed_53__50_, chained_data_delayed_53__49_, chained_data_delayed_53__48_, chained_data_delayed_53__47_, chained_data_delayed_53__46_, chained_data_delayed_53__45_, chained_data_delayed_53__44_, chained_data_delayed_53__43_, chained_data_delayed_53__42_, chained_data_delayed_53__41_, chained_data_delayed_53__40_, chained_data_delayed_53__39_, chained_data_delayed_53__38_, chained_data_delayed_53__37_, chained_data_delayed_53__36_, chained_data_delayed_53__35_, chained_data_delayed_53__34_, chained_data_delayed_53__33_, chained_data_delayed_53__32_, chained_data_delayed_53__31_, chained_data_delayed_53__30_, chained_data_delayed_53__29_, chained_data_delayed_53__28_, chained_data_delayed_53__27_, chained_data_delayed_53__26_, chained_data_delayed_53__25_, chained_data_delayed_53__24_, chained_data_delayed_53__23_, chained_data_delayed_53__22_, chained_data_delayed_53__21_, chained_data_delayed_53__20_, chained_data_delayed_53__19_, chained_data_delayed_53__18_, chained_data_delayed_53__17_, chained_data_delayed_53__16_, chained_data_delayed_53__15_, chained_data_delayed_53__14_, chained_data_delayed_53__13_, chained_data_delayed_53__12_, chained_data_delayed_53__11_, chained_data_delayed_53__10_, chained_data_delayed_53__9_, chained_data_delayed_53__8_, chained_data_delayed_53__7_, chained_data_delayed_53__6_, chained_data_delayed_53__5_, chained_data_delayed_53__4_, chained_data_delayed_53__3_, chained_data_delayed_53__2_, chained_data_delayed_53__1_, chained_data_delayed_53__0_ }),
    .data_o({ chained_data_delayed_54__63_, chained_data_delayed_54__62_, chained_data_delayed_54__61_, chained_data_delayed_54__60_, chained_data_delayed_54__59_, chained_data_delayed_54__58_, chained_data_delayed_54__57_, chained_data_delayed_54__56_, chained_data_delayed_54__55_, chained_data_delayed_54__54_, chained_data_delayed_54__53_, chained_data_delayed_54__52_, chained_data_delayed_54__51_, chained_data_delayed_54__50_, chained_data_delayed_54__49_, chained_data_delayed_54__48_, chained_data_delayed_54__47_, chained_data_delayed_54__46_, chained_data_delayed_54__45_, chained_data_delayed_54__44_, chained_data_delayed_54__43_, chained_data_delayed_54__42_, chained_data_delayed_54__41_, chained_data_delayed_54__40_, chained_data_delayed_54__39_, chained_data_delayed_54__38_, chained_data_delayed_54__37_, chained_data_delayed_54__36_, chained_data_delayed_54__35_, chained_data_delayed_54__34_, chained_data_delayed_54__33_, chained_data_delayed_54__32_, chained_data_delayed_54__31_, chained_data_delayed_54__30_, chained_data_delayed_54__29_, chained_data_delayed_54__28_, chained_data_delayed_54__27_, chained_data_delayed_54__26_, chained_data_delayed_54__25_, chained_data_delayed_54__24_, chained_data_delayed_54__23_, chained_data_delayed_54__22_, chained_data_delayed_54__21_, chained_data_delayed_54__20_, chained_data_delayed_54__19_, chained_data_delayed_54__18_, chained_data_delayed_54__17_, chained_data_delayed_54__16_, chained_data_delayed_54__15_, chained_data_delayed_54__14_, chained_data_delayed_54__13_, chained_data_delayed_54__12_, chained_data_delayed_54__11_, chained_data_delayed_54__10_, chained_data_delayed_54__9_, chained_data_delayed_54__8_, chained_data_delayed_54__7_, chained_data_delayed_54__6_, chained_data_delayed_54__5_, chained_data_delayed_54__4_, chained_data_delayed_54__3_, chained_data_delayed_54__2_, chained_data_delayed_54__1_, chained_data_delayed_54__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_55__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_54__63_, chained_data_delayed_54__62_, chained_data_delayed_54__61_, chained_data_delayed_54__60_, chained_data_delayed_54__59_, chained_data_delayed_54__58_, chained_data_delayed_54__57_, chained_data_delayed_54__56_, chained_data_delayed_54__55_, chained_data_delayed_54__54_, chained_data_delayed_54__53_, chained_data_delayed_54__52_, chained_data_delayed_54__51_, chained_data_delayed_54__50_, chained_data_delayed_54__49_, chained_data_delayed_54__48_, chained_data_delayed_54__47_, chained_data_delayed_54__46_, chained_data_delayed_54__45_, chained_data_delayed_54__44_, chained_data_delayed_54__43_, chained_data_delayed_54__42_, chained_data_delayed_54__41_, chained_data_delayed_54__40_, chained_data_delayed_54__39_, chained_data_delayed_54__38_, chained_data_delayed_54__37_, chained_data_delayed_54__36_, chained_data_delayed_54__35_, chained_data_delayed_54__34_, chained_data_delayed_54__33_, chained_data_delayed_54__32_, chained_data_delayed_54__31_, chained_data_delayed_54__30_, chained_data_delayed_54__29_, chained_data_delayed_54__28_, chained_data_delayed_54__27_, chained_data_delayed_54__26_, chained_data_delayed_54__25_, chained_data_delayed_54__24_, chained_data_delayed_54__23_, chained_data_delayed_54__22_, chained_data_delayed_54__21_, chained_data_delayed_54__20_, chained_data_delayed_54__19_, chained_data_delayed_54__18_, chained_data_delayed_54__17_, chained_data_delayed_54__16_, chained_data_delayed_54__15_, chained_data_delayed_54__14_, chained_data_delayed_54__13_, chained_data_delayed_54__12_, chained_data_delayed_54__11_, chained_data_delayed_54__10_, chained_data_delayed_54__9_, chained_data_delayed_54__8_, chained_data_delayed_54__7_, chained_data_delayed_54__6_, chained_data_delayed_54__5_, chained_data_delayed_54__4_, chained_data_delayed_54__3_, chained_data_delayed_54__2_, chained_data_delayed_54__1_, chained_data_delayed_54__0_ }),
    .data_o({ chained_data_delayed_55__63_, chained_data_delayed_55__62_, chained_data_delayed_55__61_, chained_data_delayed_55__60_, chained_data_delayed_55__59_, chained_data_delayed_55__58_, chained_data_delayed_55__57_, chained_data_delayed_55__56_, chained_data_delayed_55__55_, chained_data_delayed_55__54_, chained_data_delayed_55__53_, chained_data_delayed_55__52_, chained_data_delayed_55__51_, chained_data_delayed_55__50_, chained_data_delayed_55__49_, chained_data_delayed_55__48_, chained_data_delayed_55__47_, chained_data_delayed_55__46_, chained_data_delayed_55__45_, chained_data_delayed_55__44_, chained_data_delayed_55__43_, chained_data_delayed_55__42_, chained_data_delayed_55__41_, chained_data_delayed_55__40_, chained_data_delayed_55__39_, chained_data_delayed_55__38_, chained_data_delayed_55__37_, chained_data_delayed_55__36_, chained_data_delayed_55__35_, chained_data_delayed_55__34_, chained_data_delayed_55__33_, chained_data_delayed_55__32_, chained_data_delayed_55__31_, chained_data_delayed_55__30_, chained_data_delayed_55__29_, chained_data_delayed_55__28_, chained_data_delayed_55__27_, chained_data_delayed_55__26_, chained_data_delayed_55__25_, chained_data_delayed_55__24_, chained_data_delayed_55__23_, chained_data_delayed_55__22_, chained_data_delayed_55__21_, chained_data_delayed_55__20_, chained_data_delayed_55__19_, chained_data_delayed_55__18_, chained_data_delayed_55__17_, chained_data_delayed_55__16_, chained_data_delayed_55__15_, chained_data_delayed_55__14_, chained_data_delayed_55__13_, chained_data_delayed_55__12_, chained_data_delayed_55__11_, chained_data_delayed_55__10_, chained_data_delayed_55__9_, chained_data_delayed_55__8_, chained_data_delayed_55__7_, chained_data_delayed_55__6_, chained_data_delayed_55__5_, chained_data_delayed_55__4_, chained_data_delayed_55__3_, chained_data_delayed_55__2_, chained_data_delayed_55__1_, chained_data_delayed_55__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_56__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_55__63_, chained_data_delayed_55__62_, chained_data_delayed_55__61_, chained_data_delayed_55__60_, chained_data_delayed_55__59_, chained_data_delayed_55__58_, chained_data_delayed_55__57_, chained_data_delayed_55__56_, chained_data_delayed_55__55_, chained_data_delayed_55__54_, chained_data_delayed_55__53_, chained_data_delayed_55__52_, chained_data_delayed_55__51_, chained_data_delayed_55__50_, chained_data_delayed_55__49_, chained_data_delayed_55__48_, chained_data_delayed_55__47_, chained_data_delayed_55__46_, chained_data_delayed_55__45_, chained_data_delayed_55__44_, chained_data_delayed_55__43_, chained_data_delayed_55__42_, chained_data_delayed_55__41_, chained_data_delayed_55__40_, chained_data_delayed_55__39_, chained_data_delayed_55__38_, chained_data_delayed_55__37_, chained_data_delayed_55__36_, chained_data_delayed_55__35_, chained_data_delayed_55__34_, chained_data_delayed_55__33_, chained_data_delayed_55__32_, chained_data_delayed_55__31_, chained_data_delayed_55__30_, chained_data_delayed_55__29_, chained_data_delayed_55__28_, chained_data_delayed_55__27_, chained_data_delayed_55__26_, chained_data_delayed_55__25_, chained_data_delayed_55__24_, chained_data_delayed_55__23_, chained_data_delayed_55__22_, chained_data_delayed_55__21_, chained_data_delayed_55__20_, chained_data_delayed_55__19_, chained_data_delayed_55__18_, chained_data_delayed_55__17_, chained_data_delayed_55__16_, chained_data_delayed_55__15_, chained_data_delayed_55__14_, chained_data_delayed_55__13_, chained_data_delayed_55__12_, chained_data_delayed_55__11_, chained_data_delayed_55__10_, chained_data_delayed_55__9_, chained_data_delayed_55__8_, chained_data_delayed_55__7_, chained_data_delayed_55__6_, chained_data_delayed_55__5_, chained_data_delayed_55__4_, chained_data_delayed_55__3_, chained_data_delayed_55__2_, chained_data_delayed_55__1_, chained_data_delayed_55__0_ }),
    .data_o({ chained_data_delayed_56__63_, chained_data_delayed_56__62_, chained_data_delayed_56__61_, chained_data_delayed_56__60_, chained_data_delayed_56__59_, chained_data_delayed_56__58_, chained_data_delayed_56__57_, chained_data_delayed_56__56_, chained_data_delayed_56__55_, chained_data_delayed_56__54_, chained_data_delayed_56__53_, chained_data_delayed_56__52_, chained_data_delayed_56__51_, chained_data_delayed_56__50_, chained_data_delayed_56__49_, chained_data_delayed_56__48_, chained_data_delayed_56__47_, chained_data_delayed_56__46_, chained_data_delayed_56__45_, chained_data_delayed_56__44_, chained_data_delayed_56__43_, chained_data_delayed_56__42_, chained_data_delayed_56__41_, chained_data_delayed_56__40_, chained_data_delayed_56__39_, chained_data_delayed_56__38_, chained_data_delayed_56__37_, chained_data_delayed_56__36_, chained_data_delayed_56__35_, chained_data_delayed_56__34_, chained_data_delayed_56__33_, chained_data_delayed_56__32_, chained_data_delayed_56__31_, chained_data_delayed_56__30_, chained_data_delayed_56__29_, chained_data_delayed_56__28_, chained_data_delayed_56__27_, chained_data_delayed_56__26_, chained_data_delayed_56__25_, chained_data_delayed_56__24_, chained_data_delayed_56__23_, chained_data_delayed_56__22_, chained_data_delayed_56__21_, chained_data_delayed_56__20_, chained_data_delayed_56__19_, chained_data_delayed_56__18_, chained_data_delayed_56__17_, chained_data_delayed_56__16_, chained_data_delayed_56__15_, chained_data_delayed_56__14_, chained_data_delayed_56__13_, chained_data_delayed_56__12_, chained_data_delayed_56__11_, chained_data_delayed_56__10_, chained_data_delayed_56__9_, chained_data_delayed_56__8_, chained_data_delayed_56__7_, chained_data_delayed_56__6_, chained_data_delayed_56__5_, chained_data_delayed_56__4_, chained_data_delayed_56__3_, chained_data_delayed_56__2_, chained_data_delayed_56__1_, chained_data_delayed_56__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_57__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_56__63_, chained_data_delayed_56__62_, chained_data_delayed_56__61_, chained_data_delayed_56__60_, chained_data_delayed_56__59_, chained_data_delayed_56__58_, chained_data_delayed_56__57_, chained_data_delayed_56__56_, chained_data_delayed_56__55_, chained_data_delayed_56__54_, chained_data_delayed_56__53_, chained_data_delayed_56__52_, chained_data_delayed_56__51_, chained_data_delayed_56__50_, chained_data_delayed_56__49_, chained_data_delayed_56__48_, chained_data_delayed_56__47_, chained_data_delayed_56__46_, chained_data_delayed_56__45_, chained_data_delayed_56__44_, chained_data_delayed_56__43_, chained_data_delayed_56__42_, chained_data_delayed_56__41_, chained_data_delayed_56__40_, chained_data_delayed_56__39_, chained_data_delayed_56__38_, chained_data_delayed_56__37_, chained_data_delayed_56__36_, chained_data_delayed_56__35_, chained_data_delayed_56__34_, chained_data_delayed_56__33_, chained_data_delayed_56__32_, chained_data_delayed_56__31_, chained_data_delayed_56__30_, chained_data_delayed_56__29_, chained_data_delayed_56__28_, chained_data_delayed_56__27_, chained_data_delayed_56__26_, chained_data_delayed_56__25_, chained_data_delayed_56__24_, chained_data_delayed_56__23_, chained_data_delayed_56__22_, chained_data_delayed_56__21_, chained_data_delayed_56__20_, chained_data_delayed_56__19_, chained_data_delayed_56__18_, chained_data_delayed_56__17_, chained_data_delayed_56__16_, chained_data_delayed_56__15_, chained_data_delayed_56__14_, chained_data_delayed_56__13_, chained_data_delayed_56__12_, chained_data_delayed_56__11_, chained_data_delayed_56__10_, chained_data_delayed_56__9_, chained_data_delayed_56__8_, chained_data_delayed_56__7_, chained_data_delayed_56__6_, chained_data_delayed_56__5_, chained_data_delayed_56__4_, chained_data_delayed_56__3_, chained_data_delayed_56__2_, chained_data_delayed_56__1_, chained_data_delayed_56__0_ }),
    .data_o({ chained_data_delayed_57__63_, chained_data_delayed_57__62_, chained_data_delayed_57__61_, chained_data_delayed_57__60_, chained_data_delayed_57__59_, chained_data_delayed_57__58_, chained_data_delayed_57__57_, chained_data_delayed_57__56_, chained_data_delayed_57__55_, chained_data_delayed_57__54_, chained_data_delayed_57__53_, chained_data_delayed_57__52_, chained_data_delayed_57__51_, chained_data_delayed_57__50_, chained_data_delayed_57__49_, chained_data_delayed_57__48_, chained_data_delayed_57__47_, chained_data_delayed_57__46_, chained_data_delayed_57__45_, chained_data_delayed_57__44_, chained_data_delayed_57__43_, chained_data_delayed_57__42_, chained_data_delayed_57__41_, chained_data_delayed_57__40_, chained_data_delayed_57__39_, chained_data_delayed_57__38_, chained_data_delayed_57__37_, chained_data_delayed_57__36_, chained_data_delayed_57__35_, chained_data_delayed_57__34_, chained_data_delayed_57__33_, chained_data_delayed_57__32_, chained_data_delayed_57__31_, chained_data_delayed_57__30_, chained_data_delayed_57__29_, chained_data_delayed_57__28_, chained_data_delayed_57__27_, chained_data_delayed_57__26_, chained_data_delayed_57__25_, chained_data_delayed_57__24_, chained_data_delayed_57__23_, chained_data_delayed_57__22_, chained_data_delayed_57__21_, chained_data_delayed_57__20_, chained_data_delayed_57__19_, chained_data_delayed_57__18_, chained_data_delayed_57__17_, chained_data_delayed_57__16_, chained_data_delayed_57__15_, chained_data_delayed_57__14_, chained_data_delayed_57__13_, chained_data_delayed_57__12_, chained_data_delayed_57__11_, chained_data_delayed_57__10_, chained_data_delayed_57__9_, chained_data_delayed_57__8_, chained_data_delayed_57__7_, chained_data_delayed_57__6_, chained_data_delayed_57__5_, chained_data_delayed_57__4_, chained_data_delayed_57__3_, chained_data_delayed_57__2_, chained_data_delayed_57__1_, chained_data_delayed_57__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_58__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_57__63_, chained_data_delayed_57__62_, chained_data_delayed_57__61_, chained_data_delayed_57__60_, chained_data_delayed_57__59_, chained_data_delayed_57__58_, chained_data_delayed_57__57_, chained_data_delayed_57__56_, chained_data_delayed_57__55_, chained_data_delayed_57__54_, chained_data_delayed_57__53_, chained_data_delayed_57__52_, chained_data_delayed_57__51_, chained_data_delayed_57__50_, chained_data_delayed_57__49_, chained_data_delayed_57__48_, chained_data_delayed_57__47_, chained_data_delayed_57__46_, chained_data_delayed_57__45_, chained_data_delayed_57__44_, chained_data_delayed_57__43_, chained_data_delayed_57__42_, chained_data_delayed_57__41_, chained_data_delayed_57__40_, chained_data_delayed_57__39_, chained_data_delayed_57__38_, chained_data_delayed_57__37_, chained_data_delayed_57__36_, chained_data_delayed_57__35_, chained_data_delayed_57__34_, chained_data_delayed_57__33_, chained_data_delayed_57__32_, chained_data_delayed_57__31_, chained_data_delayed_57__30_, chained_data_delayed_57__29_, chained_data_delayed_57__28_, chained_data_delayed_57__27_, chained_data_delayed_57__26_, chained_data_delayed_57__25_, chained_data_delayed_57__24_, chained_data_delayed_57__23_, chained_data_delayed_57__22_, chained_data_delayed_57__21_, chained_data_delayed_57__20_, chained_data_delayed_57__19_, chained_data_delayed_57__18_, chained_data_delayed_57__17_, chained_data_delayed_57__16_, chained_data_delayed_57__15_, chained_data_delayed_57__14_, chained_data_delayed_57__13_, chained_data_delayed_57__12_, chained_data_delayed_57__11_, chained_data_delayed_57__10_, chained_data_delayed_57__9_, chained_data_delayed_57__8_, chained_data_delayed_57__7_, chained_data_delayed_57__6_, chained_data_delayed_57__5_, chained_data_delayed_57__4_, chained_data_delayed_57__3_, chained_data_delayed_57__2_, chained_data_delayed_57__1_, chained_data_delayed_57__0_ }),
    .data_o({ chained_data_delayed_58__63_, chained_data_delayed_58__62_, chained_data_delayed_58__61_, chained_data_delayed_58__60_, chained_data_delayed_58__59_, chained_data_delayed_58__58_, chained_data_delayed_58__57_, chained_data_delayed_58__56_, chained_data_delayed_58__55_, chained_data_delayed_58__54_, chained_data_delayed_58__53_, chained_data_delayed_58__52_, chained_data_delayed_58__51_, chained_data_delayed_58__50_, chained_data_delayed_58__49_, chained_data_delayed_58__48_, chained_data_delayed_58__47_, chained_data_delayed_58__46_, chained_data_delayed_58__45_, chained_data_delayed_58__44_, chained_data_delayed_58__43_, chained_data_delayed_58__42_, chained_data_delayed_58__41_, chained_data_delayed_58__40_, chained_data_delayed_58__39_, chained_data_delayed_58__38_, chained_data_delayed_58__37_, chained_data_delayed_58__36_, chained_data_delayed_58__35_, chained_data_delayed_58__34_, chained_data_delayed_58__33_, chained_data_delayed_58__32_, chained_data_delayed_58__31_, chained_data_delayed_58__30_, chained_data_delayed_58__29_, chained_data_delayed_58__28_, chained_data_delayed_58__27_, chained_data_delayed_58__26_, chained_data_delayed_58__25_, chained_data_delayed_58__24_, chained_data_delayed_58__23_, chained_data_delayed_58__22_, chained_data_delayed_58__21_, chained_data_delayed_58__20_, chained_data_delayed_58__19_, chained_data_delayed_58__18_, chained_data_delayed_58__17_, chained_data_delayed_58__16_, chained_data_delayed_58__15_, chained_data_delayed_58__14_, chained_data_delayed_58__13_, chained_data_delayed_58__12_, chained_data_delayed_58__11_, chained_data_delayed_58__10_, chained_data_delayed_58__9_, chained_data_delayed_58__8_, chained_data_delayed_58__7_, chained_data_delayed_58__6_, chained_data_delayed_58__5_, chained_data_delayed_58__4_, chained_data_delayed_58__3_, chained_data_delayed_58__2_, chained_data_delayed_58__1_, chained_data_delayed_58__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_59__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_58__63_, chained_data_delayed_58__62_, chained_data_delayed_58__61_, chained_data_delayed_58__60_, chained_data_delayed_58__59_, chained_data_delayed_58__58_, chained_data_delayed_58__57_, chained_data_delayed_58__56_, chained_data_delayed_58__55_, chained_data_delayed_58__54_, chained_data_delayed_58__53_, chained_data_delayed_58__52_, chained_data_delayed_58__51_, chained_data_delayed_58__50_, chained_data_delayed_58__49_, chained_data_delayed_58__48_, chained_data_delayed_58__47_, chained_data_delayed_58__46_, chained_data_delayed_58__45_, chained_data_delayed_58__44_, chained_data_delayed_58__43_, chained_data_delayed_58__42_, chained_data_delayed_58__41_, chained_data_delayed_58__40_, chained_data_delayed_58__39_, chained_data_delayed_58__38_, chained_data_delayed_58__37_, chained_data_delayed_58__36_, chained_data_delayed_58__35_, chained_data_delayed_58__34_, chained_data_delayed_58__33_, chained_data_delayed_58__32_, chained_data_delayed_58__31_, chained_data_delayed_58__30_, chained_data_delayed_58__29_, chained_data_delayed_58__28_, chained_data_delayed_58__27_, chained_data_delayed_58__26_, chained_data_delayed_58__25_, chained_data_delayed_58__24_, chained_data_delayed_58__23_, chained_data_delayed_58__22_, chained_data_delayed_58__21_, chained_data_delayed_58__20_, chained_data_delayed_58__19_, chained_data_delayed_58__18_, chained_data_delayed_58__17_, chained_data_delayed_58__16_, chained_data_delayed_58__15_, chained_data_delayed_58__14_, chained_data_delayed_58__13_, chained_data_delayed_58__12_, chained_data_delayed_58__11_, chained_data_delayed_58__10_, chained_data_delayed_58__9_, chained_data_delayed_58__8_, chained_data_delayed_58__7_, chained_data_delayed_58__6_, chained_data_delayed_58__5_, chained_data_delayed_58__4_, chained_data_delayed_58__3_, chained_data_delayed_58__2_, chained_data_delayed_58__1_, chained_data_delayed_58__0_ }),
    .data_o({ chained_data_delayed_59__63_, chained_data_delayed_59__62_, chained_data_delayed_59__61_, chained_data_delayed_59__60_, chained_data_delayed_59__59_, chained_data_delayed_59__58_, chained_data_delayed_59__57_, chained_data_delayed_59__56_, chained_data_delayed_59__55_, chained_data_delayed_59__54_, chained_data_delayed_59__53_, chained_data_delayed_59__52_, chained_data_delayed_59__51_, chained_data_delayed_59__50_, chained_data_delayed_59__49_, chained_data_delayed_59__48_, chained_data_delayed_59__47_, chained_data_delayed_59__46_, chained_data_delayed_59__45_, chained_data_delayed_59__44_, chained_data_delayed_59__43_, chained_data_delayed_59__42_, chained_data_delayed_59__41_, chained_data_delayed_59__40_, chained_data_delayed_59__39_, chained_data_delayed_59__38_, chained_data_delayed_59__37_, chained_data_delayed_59__36_, chained_data_delayed_59__35_, chained_data_delayed_59__34_, chained_data_delayed_59__33_, chained_data_delayed_59__32_, chained_data_delayed_59__31_, chained_data_delayed_59__30_, chained_data_delayed_59__29_, chained_data_delayed_59__28_, chained_data_delayed_59__27_, chained_data_delayed_59__26_, chained_data_delayed_59__25_, chained_data_delayed_59__24_, chained_data_delayed_59__23_, chained_data_delayed_59__22_, chained_data_delayed_59__21_, chained_data_delayed_59__20_, chained_data_delayed_59__19_, chained_data_delayed_59__18_, chained_data_delayed_59__17_, chained_data_delayed_59__16_, chained_data_delayed_59__15_, chained_data_delayed_59__14_, chained_data_delayed_59__13_, chained_data_delayed_59__12_, chained_data_delayed_59__11_, chained_data_delayed_59__10_, chained_data_delayed_59__9_, chained_data_delayed_59__8_, chained_data_delayed_59__7_, chained_data_delayed_59__6_, chained_data_delayed_59__5_, chained_data_delayed_59__4_, chained_data_delayed_59__3_, chained_data_delayed_59__2_, chained_data_delayed_59__1_, chained_data_delayed_59__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_60__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_59__63_, chained_data_delayed_59__62_, chained_data_delayed_59__61_, chained_data_delayed_59__60_, chained_data_delayed_59__59_, chained_data_delayed_59__58_, chained_data_delayed_59__57_, chained_data_delayed_59__56_, chained_data_delayed_59__55_, chained_data_delayed_59__54_, chained_data_delayed_59__53_, chained_data_delayed_59__52_, chained_data_delayed_59__51_, chained_data_delayed_59__50_, chained_data_delayed_59__49_, chained_data_delayed_59__48_, chained_data_delayed_59__47_, chained_data_delayed_59__46_, chained_data_delayed_59__45_, chained_data_delayed_59__44_, chained_data_delayed_59__43_, chained_data_delayed_59__42_, chained_data_delayed_59__41_, chained_data_delayed_59__40_, chained_data_delayed_59__39_, chained_data_delayed_59__38_, chained_data_delayed_59__37_, chained_data_delayed_59__36_, chained_data_delayed_59__35_, chained_data_delayed_59__34_, chained_data_delayed_59__33_, chained_data_delayed_59__32_, chained_data_delayed_59__31_, chained_data_delayed_59__30_, chained_data_delayed_59__29_, chained_data_delayed_59__28_, chained_data_delayed_59__27_, chained_data_delayed_59__26_, chained_data_delayed_59__25_, chained_data_delayed_59__24_, chained_data_delayed_59__23_, chained_data_delayed_59__22_, chained_data_delayed_59__21_, chained_data_delayed_59__20_, chained_data_delayed_59__19_, chained_data_delayed_59__18_, chained_data_delayed_59__17_, chained_data_delayed_59__16_, chained_data_delayed_59__15_, chained_data_delayed_59__14_, chained_data_delayed_59__13_, chained_data_delayed_59__12_, chained_data_delayed_59__11_, chained_data_delayed_59__10_, chained_data_delayed_59__9_, chained_data_delayed_59__8_, chained_data_delayed_59__7_, chained_data_delayed_59__6_, chained_data_delayed_59__5_, chained_data_delayed_59__4_, chained_data_delayed_59__3_, chained_data_delayed_59__2_, chained_data_delayed_59__1_, chained_data_delayed_59__0_ }),
    .data_o({ chained_data_delayed_60__63_, chained_data_delayed_60__62_, chained_data_delayed_60__61_, chained_data_delayed_60__60_, chained_data_delayed_60__59_, chained_data_delayed_60__58_, chained_data_delayed_60__57_, chained_data_delayed_60__56_, chained_data_delayed_60__55_, chained_data_delayed_60__54_, chained_data_delayed_60__53_, chained_data_delayed_60__52_, chained_data_delayed_60__51_, chained_data_delayed_60__50_, chained_data_delayed_60__49_, chained_data_delayed_60__48_, chained_data_delayed_60__47_, chained_data_delayed_60__46_, chained_data_delayed_60__45_, chained_data_delayed_60__44_, chained_data_delayed_60__43_, chained_data_delayed_60__42_, chained_data_delayed_60__41_, chained_data_delayed_60__40_, chained_data_delayed_60__39_, chained_data_delayed_60__38_, chained_data_delayed_60__37_, chained_data_delayed_60__36_, chained_data_delayed_60__35_, chained_data_delayed_60__34_, chained_data_delayed_60__33_, chained_data_delayed_60__32_, chained_data_delayed_60__31_, chained_data_delayed_60__30_, chained_data_delayed_60__29_, chained_data_delayed_60__28_, chained_data_delayed_60__27_, chained_data_delayed_60__26_, chained_data_delayed_60__25_, chained_data_delayed_60__24_, chained_data_delayed_60__23_, chained_data_delayed_60__22_, chained_data_delayed_60__21_, chained_data_delayed_60__20_, chained_data_delayed_60__19_, chained_data_delayed_60__18_, chained_data_delayed_60__17_, chained_data_delayed_60__16_, chained_data_delayed_60__15_, chained_data_delayed_60__14_, chained_data_delayed_60__13_, chained_data_delayed_60__12_, chained_data_delayed_60__11_, chained_data_delayed_60__10_, chained_data_delayed_60__9_, chained_data_delayed_60__8_, chained_data_delayed_60__7_, chained_data_delayed_60__6_, chained_data_delayed_60__5_, chained_data_delayed_60__4_, chained_data_delayed_60__3_, chained_data_delayed_60__2_, chained_data_delayed_60__1_, chained_data_delayed_60__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_61__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_60__63_, chained_data_delayed_60__62_, chained_data_delayed_60__61_, chained_data_delayed_60__60_, chained_data_delayed_60__59_, chained_data_delayed_60__58_, chained_data_delayed_60__57_, chained_data_delayed_60__56_, chained_data_delayed_60__55_, chained_data_delayed_60__54_, chained_data_delayed_60__53_, chained_data_delayed_60__52_, chained_data_delayed_60__51_, chained_data_delayed_60__50_, chained_data_delayed_60__49_, chained_data_delayed_60__48_, chained_data_delayed_60__47_, chained_data_delayed_60__46_, chained_data_delayed_60__45_, chained_data_delayed_60__44_, chained_data_delayed_60__43_, chained_data_delayed_60__42_, chained_data_delayed_60__41_, chained_data_delayed_60__40_, chained_data_delayed_60__39_, chained_data_delayed_60__38_, chained_data_delayed_60__37_, chained_data_delayed_60__36_, chained_data_delayed_60__35_, chained_data_delayed_60__34_, chained_data_delayed_60__33_, chained_data_delayed_60__32_, chained_data_delayed_60__31_, chained_data_delayed_60__30_, chained_data_delayed_60__29_, chained_data_delayed_60__28_, chained_data_delayed_60__27_, chained_data_delayed_60__26_, chained_data_delayed_60__25_, chained_data_delayed_60__24_, chained_data_delayed_60__23_, chained_data_delayed_60__22_, chained_data_delayed_60__21_, chained_data_delayed_60__20_, chained_data_delayed_60__19_, chained_data_delayed_60__18_, chained_data_delayed_60__17_, chained_data_delayed_60__16_, chained_data_delayed_60__15_, chained_data_delayed_60__14_, chained_data_delayed_60__13_, chained_data_delayed_60__12_, chained_data_delayed_60__11_, chained_data_delayed_60__10_, chained_data_delayed_60__9_, chained_data_delayed_60__8_, chained_data_delayed_60__7_, chained_data_delayed_60__6_, chained_data_delayed_60__5_, chained_data_delayed_60__4_, chained_data_delayed_60__3_, chained_data_delayed_60__2_, chained_data_delayed_60__1_, chained_data_delayed_60__0_ }),
    .data_o({ chained_data_delayed_61__63_, chained_data_delayed_61__62_, chained_data_delayed_61__61_, chained_data_delayed_61__60_, chained_data_delayed_61__59_, chained_data_delayed_61__58_, chained_data_delayed_61__57_, chained_data_delayed_61__56_, chained_data_delayed_61__55_, chained_data_delayed_61__54_, chained_data_delayed_61__53_, chained_data_delayed_61__52_, chained_data_delayed_61__51_, chained_data_delayed_61__50_, chained_data_delayed_61__49_, chained_data_delayed_61__48_, chained_data_delayed_61__47_, chained_data_delayed_61__46_, chained_data_delayed_61__45_, chained_data_delayed_61__44_, chained_data_delayed_61__43_, chained_data_delayed_61__42_, chained_data_delayed_61__41_, chained_data_delayed_61__40_, chained_data_delayed_61__39_, chained_data_delayed_61__38_, chained_data_delayed_61__37_, chained_data_delayed_61__36_, chained_data_delayed_61__35_, chained_data_delayed_61__34_, chained_data_delayed_61__33_, chained_data_delayed_61__32_, chained_data_delayed_61__31_, chained_data_delayed_61__30_, chained_data_delayed_61__29_, chained_data_delayed_61__28_, chained_data_delayed_61__27_, chained_data_delayed_61__26_, chained_data_delayed_61__25_, chained_data_delayed_61__24_, chained_data_delayed_61__23_, chained_data_delayed_61__22_, chained_data_delayed_61__21_, chained_data_delayed_61__20_, chained_data_delayed_61__19_, chained_data_delayed_61__18_, chained_data_delayed_61__17_, chained_data_delayed_61__16_, chained_data_delayed_61__15_, chained_data_delayed_61__14_, chained_data_delayed_61__13_, chained_data_delayed_61__12_, chained_data_delayed_61__11_, chained_data_delayed_61__10_, chained_data_delayed_61__9_, chained_data_delayed_61__8_, chained_data_delayed_61__7_, chained_data_delayed_61__6_, chained_data_delayed_61__5_, chained_data_delayed_61__4_, chained_data_delayed_61__3_, chained_data_delayed_61__2_, chained_data_delayed_61__1_, chained_data_delayed_61__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_62__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_61__63_, chained_data_delayed_61__62_, chained_data_delayed_61__61_, chained_data_delayed_61__60_, chained_data_delayed_61__59_, chained_data_delayed_61__58_, chained_data_delayed_61__57_, chained_data_delayed_61__56_, chained_data_delayed_61__55_, chained_data_delayed_61__54_, chained_data_delayed_61__53_, chained_data_delayed_61__52_, chained_data_delayed_61__51_, chained_data_delayed_61__50_, chained_data_delayed_61__49_, chained_data_delayed_61__48_, chained_data_delayed_61__47_, chained_data_delayed_61__46_, chained_data_delayed_61__45_, chained_data_delayed_61__44_, chained_data_delayed_61__43_, chained_data_delayed_61__42_, chained_data_delayed_61__41_, chained_data_delayed_61__40_, chained_data_delayed_61__39_, chained_data_delayed_61__38_, chained_data_delayed_61__37_, chained_data_delayed_61__36_, chained_data_delayed_61__35_, chained_data_delayed_61__34_, chained_data_delayed_61__33_, chained_data_delayed_61__32_, chained_data_delayed_61__31_, chained_data_delayed_61__30_, chained_data_delayed_61__29_, chained_data_delayed_61__28_, chained_data_delayed_61__27_, chained_data_delayed_61__26_, chained_data_delayed_61__25_, chained_data_delayed_61__24_, chained_data_delayed_61__23_, chained_data_delayed_61__22_, chained_data_delayed_61__21_, chained_data_delayed_61__20_, chained_data_delayed_61__19_, chained_data_delayed_61__18_, chained_data_delayed_61__17_, chained_data_delayed_61__16_, chained_data_delayed_61__15_, chained_data_delayed_61__14_, chained_data_delayed_61__13_, chained_data_delayed_61__12_, chained_data_delayed_61__11_, chained_data_delayed_61__10_, chained_data_delayed_61__9_, chained_data_delayed_61__8_, chained_data_delayed_61__7_, chained_data_delayed_61__6_, chained_data_delayed_61__5_, chained_data_delayed_61__4_, chained_data_delayed_61__3_, chained_data_delayed_61__2_, chained_data_delayed_61__1_, chained_data_delayed_61__0_ }),
    .data_o({ chained_data_delayed_62__63_, chained_data_delayed_62__62_, chained_data_delayed_62__61_, chained_data_delayed_62__60_, chained_data_delayed_62__59_, chained_data_delayed_62__58_, chained_data_delayed_62__57_, chained_data_delayed_62__56_, chained_data_delayed_62__55_, chained_data_delayed_62__54_, chained_data_delayed_62__53_, chained_data_delayed_62__52_, chained_data_delayed_62__51_, chained_data_delayed_62__50_, chained_data_delayed_62__49_, chained_data_delayed_62__48_, chained_data_delayed_62__47_, chained_data_delayed_62__46_, chained_data_delayed_62__45_, chained_data_delayed_62__44_, chained_data_delayed_62__43_, chained_data_delayed_62__42_, chained_data_delayed_62__41_, chained_data_delayed_62__40_, chained_data_delayed_62__39_, chained_data_delayed_62__38_, chained_data_delayed_62__37_, chained_data_delayed_62__36_, chained_data_delayed_62__35_, chained_data_delayed_62__34_, chained_data_delayed_62__33_, chained_data_delayed_62__32_, chained_data_delayed_62__31_, chained_data_delayed_62__30_, chained_data_delayed_62__29_, chained_data_delayed_62__28_, chained_data_delayed_62__27_, chained_data_delayed_62__26_, chained_data_delayed_62__25_, chained_data_delayed_62__24_, chained_data_delayed_62__23_, chained_data_delayed_62__22_, chained_data_delayed_62__21_, chained_data_delayed_62__20_, chained_data_delayed_62__19_, chained_data_delayed_62__18_, chained_data_delayed_62__17_, chained_data_delayed_62__16_, chained_data_delayed_62__15_, chained_data_delayed_62__14_, chained_data_delayed_62__13_, chained_data_delayed_62__12_, chained_data_delayed_62__11_, chained_data_delayed_62__10_, chained_data_delayed_62__9_, chained_data_delayed_62__8_, chained_data_delayed_62__7_, chained_data_delayed_62__6_, chained_data_delayed_62__5_, chained_data_delayed_62__4_, chained_data_delayed_62__3_, chained_data_delayed_62__2_, chained_data_delayed_62__1_, chained_data_delayed_62__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_63__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_62__63_, chained_data_delayed_62__62_, chained_data_delayed_62__61_, chained_data_delayed_62__60_, chained_data_delayed_62__59_, chained_data_delayed_62__58_, chained_data_delayed_62__57_, chained_data_delayed_62__56_, chained_data_delayed_62__55_, chained_data_delayed_62__54_, chained_data_delayed_62__53_, chained_data_delayed_62__52_, chained_data_delayed_62__51_, chained_data_delayed_62__50_, chained_data_delayed_62__49_, chained_data_delayed_62__48_, chained_data_delayed_62__47_, chained_data_delayed_62__46_, chained_data_delayed_62__45_, chained_data_delayed_62__44_, chained_data_delayed_62__43_, chained_data_delayed_62__42_, chained_data_delayed_62__41_, chained_data_delayed_62__40_, chained_data_delayed_62__39_, chained_data_delayed_62__38_, chained_data_delayed_62__37_, chained_data_delayed_62__36_, chained_data_delayed_62__35_, chained_data_delayed_62__34_, chained_data_delayed_62__33_, chained_data_delayed_62__32_, chained_data_delayed_62__31_, chained_data_delayed_62__30_, chained_data_delayed_62__29_, chained_data_delayed_62__28_, chained_data_delayed_62__27_, chained_data_delayed_62__26_, chained_data_delayed_62__25_, chained_data_delayed_62__24_, chained_data_delayed_62__23_, chained_data_delayed_62__22_, chained_data_delayed_62__21_, chained_data_delayed_62__20_, chained_data_delayed_62__19_, chained_data_delayed_62__18_, chained_data_delayed_62__17_, chained_data_delayed_62__16_, chained_data_delayed_62__15_, chained_data_delayed_62__14_, chained_data_delayed_62__13_, chained_data_delayed_62__12_, chained_data_delayed_62__11_, chained_data_delayed_62__10_, chained_data_delayed_62__9_, chained_data_delayed_62__8_, chained_data_delayed_62__7_, chained_data_delayed_62__6_, chained_data_delayed_62__5_, chained_data_delayed_62__4_, chained_data_delayed_62__3_, chained_data_delayed_62__2_, chained_data_delayed_62__1_, chained_data_delayed_62__0_ }),
    .data_o({ chained_data_delayed_63__63_, chained_data_delayed_63__62_, chained_data_delayed_63__61_, chained_data_delayed_63__60_, chained_data_delayed_63__59_, chained_data_delayed_63__58_, chained_data_delayed_63__57_, chained_data_delayed_63__56_, chained_data_delayed_63__55_, chained_data_delayed_63__54_, chained_data_delayed_63__53_, chained_data_delayed_63__52_, chained_data_delayed_63__51_, chained_data_delayed_63__50_, chained_data_delayed_63__49_, chained_data_delayed_63__48_, chained_data_delayed_63__47_, chained_data_delayed_63__46_, chained_data_delayed_63__45_, chained_data_delayed_63__44_, chained_data_delayed_63__43_, chained_data_delayed_63__42_, chained_data_delayed_63__41_, chained_data_delayed_63__40_, chained_data_delayed_63__39_, chained_data_delayed_63__38_, chained_data_delayed_63__37_, chained_data_delayed_63__36_, chained_data_delayed_63__35_, chained_data_delayed_63__34_, chained_data_delayed_63__33_, chained_data_delayed_63__32_, chained_data_delayed_63__31_, chained_data_delayed_63__30_, chained_data_delayed_63__29_, chained_data_delayed_63__28_, chained_data_delayed_63__27_, chained_data_delayed_63__26_, chained_data_delayed_63__25_, chained_data_delayed_63__24_, chained_data_delayed_63__23_, chained_data_delayed_63__22_, chained_data_delayed_63__21_, chained_data_delayed_63__20_, chained_data_delayed_63__19_, chained_data_delayed_63__18_, chained_data_delayed_63__17_, chained_data_delayed_63__16_, chained_data_delayed_63__15_, chained_data_delayed_63__14_, chained_data_delayed_63__13_, chained_data_delayed_63__12_, chained_data_delayed_63__11_, chained_data_delayed_63__10_, chained_data_delayed_63__9_, chained_data_delayed_63__8_, chained_data_delayed_63__7_, chained_data_delayed_63__6_, chained_data_delayed_63__5_, chained_data_delayed_63__4_, chained_data_delayed_63__3_, chained_data_delayed_63__2_, chained_data_delayed_63__1_, chained_data_delayed_63__0_ })
  );


  bsg_dff_width_p64
  chained_genblk1_64__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_63__63_, chained_data_delayed_63__62_, chained_data_delayed_63__61_, chained_data_delayed_63__60_, chained_data_delayed_63__59_, chained_data_delayed_63__58_, chained_data_delayed_63__57_, chained_data_delayed_63__56_, chained_data_delayed_63__55_, chained_data_delayed_63__54_, chained_data_delayed_63__53_, chained_data_delayed_63__52_, chained_data_delayed_63__51_, chained_data_delayed_63__50_, chained_data_delayed_63__49_, chained_data_delayed_63__48_, chained_data_delayed_63__47_, chained_data_delayed_63__46_, chained_data_delayed_63__45_, chained_data_delayed_63__44_, chained_data_delayed_63__43_, chained_data_delayed_63__42_, chained_data_delayed_63__41_, chained_data_delayed_63__40_, chained_data_delayed_63__39_, chained_data_delayed_63__38_, chained_data_delayed_63__37_, chained_data_delayed_63__36_, chained_data_delayed_63__35_, chained_data_delayed_63__34_, chained_data_delayed_63__33_, chained_data_delayed_63__32_, chained_data_delayed_63__31_, chained_data_delayed_63__30_, chained_data_delayed_63__29_, chained_data_delayed_63__28_, chained_data_delayed_63__27_, chained_data_delayed_63__26_, chained_data_delayed_63__25_, chained_data_delayed_63__24_, chained_data_delayed_63__23_, chained_data_delayed_63__22_, chained_data_delayed_63__21_, chained_data_delayed_63__20_, chained_data_delayed_63__19_, chained_data_delayed_63__18_, chained_data_delayed_63__17_, chained_data_delayed_63__16_, chained_data_delayed_63__15_, chained_data_delayed_63__14_, chained_data_delayed_63__13_, chained_data_delayed_63__12_, chained_data_delayed_63__11_, chained_data_delayed_63__10_, chained_data_delayed_63__9_, chained_data_delayed_63__8_, chained_data_delayed_63__7_, chained_data_delayed_63__6_, chained_data_delayed_63__5_, chained_data_delayed_63__4_, chained_data_delayed_63__3_, chained_data_delayed_63__2_, chained_data_delayed_63__1_, chained_data_delayed_63__0_ }),
    .data_o(data_o)
  );


endmodule

