

module top
(
  i,
  o
);

  input [63999:0] i;
  output [63999:0] o;

  bsg_flatten_2D_array
  wrapper
  (
    .i(i),
    .o(o)
  );


endmodule



module bsg_flatten_2D_array
(
  i,
  o
);

  input [63999:0] i;
  output [63999:0] o;
  wire [63999:0] o;
  assign o[63999] = i[63999];
  assign o[63998] = i[63998];
  assign o[63997] = i[63997];
  assign o[63996] = i[63996];
  assign o[63995] = i[63995];
  assign o[63994] = i[63994];
  assign o[63993] = i[63993];
  assign o[63992] = i[63992];
  assign o[63991] = i[63991];
  assign o[63990] = i[63990];
  assign o[63989] = i[63989];
  assign o[63988] = i[63988];
  assign o[63987] = i[63987];
  assign o[63986] = i[63986];
  assign o[63985] = i[63985];
  assign o[63984] = i[63984];
  assign o[63983] = i[63983];
  assign o[63982] = i[63982];
  assign o[63981] = i[63981];
  assign o[63980] = i[63980];
  assign o[63979] = i[63979];
  assign o[63978] = i[63978];
  assign o[63977] = i[63977];
  assign o[63976] = i[63976];
  assign o[63975] = i[63975];
  assign o[63974] = i[63974];
  assign o[63973] = i[63973];
  assign o[63972] = i[63972];
  assign o[63971] = i[63971];
  assign o[63970] = i[63970];
  assign o[63969] = i[63969];
  assign o[63968] = i[63968];
  assign o[63967] = i[63967];
  assign o[63966] = i[63966];
  assign o[63965] = i[63965];
  assign o[63964] = i[63964];
  assign o[63963] = i[63963];
  assign o[63962] = i[63962];
  assign o[63961] = i[63961];
  assign o[63960] = i[63960];
  assign o[63959] = i[63959];
  assign o[63958] = i[63958];
  assign o[63957] = i[63957];
  assign o[63956] = i[63956];
  assign o[63955] = i[63955];
  assign o[63954] = i[63954];
  assign o[63953] = i[63953];
  assign o[63952] = i[63952];
  assign o[63951] = i[63951];
  assign o[63950] = i[63950];
  assign o[63949] = i[63949];
  assign o[63948] = i[63948];
  assign o[63947] = i[63947];
  assign o[63946] = i[63946];
  assign o[63945] = i[63945];
  assign o[63944] = i[63944];
  assign o[63943] = i[63943];
  assign o[63942] = i[63942];
  assign o[63941] = i[63941];
  assign o[63940] = i[63940];
  assign o[63939] = i[63939];
  assign o[63938] = i[63938];
  assign o[63937] = i[63937];
  assign o[63936] = i[63936];
  assign o[63935] = i[63935];
  assign o[63934] = i[63934];
  assign o[63933] = i[63933];
  assign o[63932] = i[63932];
  assign o[63931] = i[63931];
  assign o[63930] = i[63930];
  assign o[63929] = i[63929];
  assign o[63928] = i[63928];
  assign o[63927] = i[63927];
  assign o[63926] = i[63926];
  assign o[63925] = i[63925];
  assign o[63924] = i[63924];
  assign o[63923] = i[63923];
  assign o[63922] = i[63922];
  assign o[63921] = i[63921];
  assign o[63920] = i[63920];
  assign o[63919] = i[63919];
  assign o[63918] = i[63918];
  assign o[63917] = i[63917];
  assign o[63916] = i[63916];
  assign o[63915] = i[63915];
  assign o[63914] = i[63914];
  assign o[63913] = i[63913];
  assign o[63912] = i[63912];
  assign o[63911] = i[63911];
  assign o[63910] = i[63910];
  assign o[63909] = i[63909];
  assign o[63908] = i[63908];
  assign o[63907] = i[63907];
  assign o[63906] = i[63906];
  assign o[63905] = i[63905];
  assign o[63904] = i[63904];
  assign o[63903] = i[63903];
  assign o[63902] = i[63902];
  assign o[63901] = i[63901];
  assign o[63900] = i[63900];
  assign o[63899] = i[63899];
  assign o[63898] = i[63898];
  assign o[63897] = i[63897];
  assign o[63896] = i[63896];
  assign o[63895] = i[63895];
  assign o[63894] = i[63894];
  assign o[63893] = i[63893];
  assign o[63892] = i[63892];
  assign o[63891] = i[63891];
  assign o[63890] = i[63890];
  assign o[63889] = i[63889];
  assign o[63888] = i[63888];
  assign o[63887] = i[63887];
  assign o[63886] = i[63886];
  assign o[63885] = i[63885];
  assign o[63884] = i[63884];
  assign o[63883] = i[63883];
  assign o[63882] = i[63882];
  assign o[63881] = i[63881];
  assign o[63880] = i[63880];
  assign o[63879] = i[63879];
  assign o[63878] = i[63878];
  assign o[63877] = i[63877];
  assign o[63876] = i[63876];
  assign o[63875] = i[63875];
  assign o[63874] = i[63874];
  assign o[63873] = i[63873];
  assign o[63872] = i[63872];
  assign o[63871] = i[63871];
  assign o[63870] = i[63870];
  assign o[63869] = i[63869];
  assign o[63868] = i[63868];
  assign o[63867] = i[63867];
  assign o[63866] = i[63866];
  assign o[63865] = i[63865];
  assign o[63864] = i[63864];
  assign o[63863] = i[63863];
  assign o[63862] = i[63862];
  assign o[63861] = i[63861];
  assign o[63860] = i[63860];
  assign o[63859] = i[63859];
  assign o[63858] = i[63858];
  assign o[63857] = i[63857];
  assign o[63856] = i[63856];
  assign o[63855] = i[63855];
  assign o[63854] = i[63854];
  assign o[63853] = i[63853];
  assign o[63852] = i[63852];
  assign o[63851] = i[63851];
  assign o[63850] = i[63850];
  assign o[63849] = i[63849];
  assign o[63848] = i[63848];
  assign o[63847] = i[63847];
  assign o[63846] = i[63846];
  assign o[63845] = i[63845];
  assign o[63844] = i[63844];
  assign o[63843] = i[63843];
  assign o[63842] = i[63842];
  assign o[63841] = i[63841];
  assign o[63840] = i[63840];
  assign o[63839] = i[63839];
  assign o[63838] = i[63838];
  assign o[63837] = i[63837];
  assign o[63836] = i[63836];
  assign o[63835] = i[63835];
  assign o[63834] = i[63834];
  assign o[63833] = i[63833];
  assign o[63832] = i[63832];
  assign o[63831] = i[63831];
  assign o[63830] = i[63830];
  assign o[63829] = i[63829];
  assign o[63828] = i[63828];
  assign o[63827] = i[63827];
  assign o[63826] = i[63826];
  assign o[63825] = i[63825];
  assign o[63824] = i[63824];
  assign o[63823] = i[63823];
  assign o[63822] = i[63822];
  assign o[63821] = i[63821];
  assign o[63820] = i[63820];
  assign o[63819] = i[63819];
  assign o[63818] = i[63818];
  assign o[63817] = i[63817];
  assign o[63816] = i[63816];
  assign o[63815] = i[63815];
  assign o[63814] = i[63814];
  assign o[63813] = i[63813];
  assign o[63812] = i[63812];
  assign o[63811] = i[63811];
  assign o[63810] = i[63810];
  assign o[63809] = i[63809];
  assign o[63808] = i[63808];
  assign o[63807] = i[63807];
  assign o[63806] = i[63806];
  assign o[63805] = i[63805];
  assign o[63804] = i[63804];
  assign o[63803] = i[63803];
  assign o[63802] = i[63802];
  assign o[63801] = i[63801];
  assign o[63800] = i[63800];
  assign o[63799] = i[63799];
  assign o[63798] = i[63798];
  assign o[63797] = i[63797];
  assign o[63796] = i[63796];
  assign o[63795] = i[63795];
  assign o[63794] = i[63794];
  assign o[63793] = i[63793];
  assign o[63792] = i[63792];
  assign o[63791] = i[63791];
  assign o[63790] = i[63790];
  assign o[63789] = i[63789];
  assign o[63788] = i[63788];
  assign o[63787] = i[63787];
  assign o[63786] = i[63786];
  assign o[63785] = i[63785];
  assign o[63784] = i[63784];
  assign o[63783] = i[63783];
  assign o[63782] = i[63782];
  assign o[63781] = i[63781];
  assign o[63780] = i[63780];
  assign o[63779] = i[63779];
  assign o[63778] = i[63778];
  assign o[63777] = i[63777];
  assign o[63776] = i[63776];
  assign o[63775] = i[63775];
  assign o[63774] = i[63774];
  assign o[63773] = i[63773];
  assign o[63772] = i[63772];
  assign o[63771] = i[63771];
  assign o[63770] = i[63770];
  assign o[63769] = i[63769];
  assign o[63768] = i[63768];
  assign o[63767] = i[63767];
  assign o[63766] = i[63766];
  assign o[63765] = i[63765];
  assign o[63764] = i[63764];
  assign o[63763] = i[63763];
  assign o[63762] = i[63762];
  assign o[63761] = i[63761];
  assign o[63760] = i[63760];
  assign o[63759] = i[63759];
  assign o[63758] = i[63758];
  assign o[63757] = i[63757];
  assign o[63756] = i[63756];
  assign o[63755] = i[63755];
  assign o[63754] = i[63754];
  assign o[63753] = i[63753];
  assign o[63752] = i[63752];
  assign o[63751] = i[63751];
  assign o[63750] = i[63750];
  assign o[63749] = i[63749];
  assign o[63748] = i[63748];
  assign o[63747] = i[63747];
  assign o[63746] = i[63746];
  assign o[63745] = i[63745];
  assign o[63744] = i[63744];
  assign o[63743] = i[63743];
  assign o[63742] = i[63742];
  assign o[63741] = i[63741];
  assign o[63740] = i[63740];
  assign o[63739] = i[63739];
  assign o[63738] = i[63738];
  assign o[63737] = i[63737];
  assign o[63736] = i[63736];
  assign o[63735] = i[63735];
  assign o[63734] = i[63734];
  assign o[63733] = i[63733];
  assign o[63732] = i[63732];
  assign o[63731] = i[63731];
  assign o[63730] = i[63730];
  assign o[63729] = i[63729];
  assign o[63728] = i[63728];
  assign o[63727] = i[63727];
  assign o[63726] = i[63726];
  assign o[63725] = i[63725];
  assign o[63724] = i[63724];
  assign o[63723] = i[63723];
  assign o[63722] = i[63722];
  assign o[63721] = i[63721];
  assign o[63720] = i[63720];
  assign o[63719] = i[63719];
  assign o[63718] = i[63718];
  assign o[63717] = i[63717];
  assign o[63716] = i[63716];
  assign o[63715] = i[63715];
  assign o[63714] = i[63714];
  assign o[63713] = i[63713];
  assign o[63712] = i[63712];
  assign o[63711] = i[63711];
  assign o[63710] = i[63710];
  assign o[63709] = i[63709];
  assign o[63708] = i[63708];
  assign o[63707] = i[63707];
  assign o[63706] = i[63706];
  assign o[63705] = i[63705];
  assign o[63704] = i[63704];
  assign o[63703] = i[63703];
  assign o[63702] = i[63702];
  assign o[63701] = i[63701];
  assign o[63700] = i[63700];
  assign o[63699] = i[63699];
  assign o[63698] = i[63698];
  assign o[63697] = i[63697];
  assign o[63696] = i[63696];
  assign o[63695] = i[63695];
  assign o[63694] = i[63694];
  assign o[63693] = i[63693];
  assign o[63692] = i[63692];
  assign o[63691] = i[63691];
  assign o[63690] = i[63690];
  assign o[63689] = i[63689];
  assign o[63688] = i[63688];
  assign o[63687] = i[63687];
  assign o[63686] = i[63686];
  assign o[63685] = i[63685];
  assign o[63684] = i[63684];
  assign o[63683] = i[63683];
  assign o[63682] = i[63682];
  assign o[63681] = i[63681];
  assign o[63680] = i[63680];
  assign o[63679] = i[63679];
  assign o[63678] = i[63678];
  assign o[63677] = i[63677];
  assign o[63676] = i[63676];
  assign o[63675] = i[63675];
  assign o[63674] = i[63674];
  assign o[63673] = i[63673];
  assign o[63672] = i[63672];
  assign o[63671] = i[63671];
  assign o[63670] = i[63670];
  assign o[63669] = i[63669];
  assign o[63668] = i[63668];
  assign o[63667] = i[63667];
  assign o[63666] = i[63666];
  assign o[63665] = i[63665];
  assign o[63664] = i[63664];
  assign o[63663] = i[63663];
  assign o[63662] = i[63662];
  assign o[63661] = i[63661];
  assign o[63660] = i[63660];
  assign o[63659] = i[63659];
  assign o[63658] = i[63658];
  assign o[63657] = i[63657];
  assign o[63656] = i[63656];
  assign o[63655] = i[63655];
  assign o[63654] = i[63654];
  assign o[63653] = i[63653];
  assign o[63652] = i[63652];
  assign o[63651] = i[63651];
  assign o[63650] = i[63650];
  assign o[63649] = i[63649];
  assign o[63648] = i[63648];
  assign o[63647] = i[63647];
  assign o[63646] = i[63646];
  assign o[63645] = i[63645];
  assign o[63644] = i[63644];
  assign o[63643] = i[63643];
  assign o[63642] = i[63642];
  assign o[63641] = i[63641];
  assign o[63640] = i[63640];
  assign o[63639] = i[63639];
  assign o[63638] = i[63638];
  assign o[63637] = i[63637];
  assign o[63636] = i[63636];
  assign o[63635] = i[63635];
  assign o[63634] = i[63634];
  assign o[63633] = i[63633];
  assign o[63632] = i[63632];
  assign o[63631] = i[63631];
  assign o[63630] = i[63630];
  assign o[63629] = i[63629];
  assign o[63628] = i[63628];
  assign o[63627] = i[63627];
  assign o[63626] = i[63626];
  assign o[63625] = i[63625];
  assign o[63624] = i[63624];
  assign o[63623] = i[63623];
  assign o[63622] = i[63622];
  assign o[63621] = i[63621];
  assign o[63620] = i[63620];
  assign o[63619] = i[63619];
  assign o[63618] = i[63618];
  assign o[63617] = i[63617];
  assign o[63616] = i[63616];
  assign o[63615] = i[63615];
  assign o[63614] = i[63614];
  assign o[63613] = i[63613];
  assign o[63612] = i[63612];
  assign o[63611] = i[63611];
  assign o[63610] = i[63610];
  assign o[63609] = i[63609];
  assign o[63608] = i[63608];
  assign o[63607] = i[63607];
  assign o[63606] = i[63606];
  assign o[63605] = i[63605];
  assign o[63604] = i[63604];
  assign o[63603] = i[63603];
  assign o[63602] = i[63602];
  assign o[63601] = i[63601];
  assign o[63600] = i[63600];
  assign o[63599] = i[63599];
  assign o[63598] = i[63598];
  assign o[63597] = i[63597];
  assign o[63596] = i[63596];
  assign o[63595] = i[63595];
  assign o[63594] = i[63594];
  assign o[63593] = i[63593];
  assign o[63592] = i[63592];
  assign o[63591] = i[63591];
  assign o[63590] = i[63590];
  assign o[63589] = i[63589];
  assign o[63588] = i[63588];
  assign o[63587] = i[63587];
  assign o[63586] = i[63586];
  assign o[63585] = i[63585];
  assign o[63584] = i[63584];
  assign o[63583] = i[63583];
  assign o[63582] = i[63582];
  assign o[63581] = i[63581];
  assign o[63580] = i[63580];
  assign o[63579] = i[63579];
  assign o[63578] = i[63578];
  assign o[63577] = i[63577];
  assign o[63576] = i[63576];
  assign o[63575] = i[63575];
  assign o[63574] = i[63574];
  assign o[63573] = i[63573];
  assign o[63572] = i[63572];
  assign o[63571] = i[63571];
  assign o[63570] = i[63570];
  assign o[63569] = i[63569];
  assign o[63568] = i[63568];
  assign o[63567] = i[63567];
  assign o[63566] = i[63566];
  assign o[63565] = i[63565];
  assign o[63564] = i[63564];
  assign o[63563] = i[63563];
  assign o[63562] = i[63562];
  assign o[63561] = i[63561];
  assign o[63560] = i[63560];
  assign o[63559] = i[63559];
  assign o[63558] = i[63558];
  assign o[63557] = i[63557];
  assign o[63556] = i[63556];
  assign o[63555] = i[63555];
  assign o[63554] = i[63554];
  assign o[63553] = i[63553];
  assign o[63552] = i[63552];
  assign o[63551] = i[63551];
  assign o[63550] = i[63550];
  assign o[63549] = i[63549];
  assign o[63548] = i[63548];
  assign o[63547] = i[63547];
  assign o[63546] = i[63546];
  assign o[63545] = i[63545];
  assign o[63544] = i[63544];
  assign o[63543] = i[63543];
  assign o[63542] = i[63542];
  assign o[63541] = i[63541];
  assign o[63540] = i[63540];
  assign o[63539] = i[63539];
  assign o[63538] = i[63538];
  assign o[63537] = i[63537];
  assign o[63536] = i[63536];
  assign o[63535] = i[63535];
  assign o[63534] = i[63534];
  assign o[63533] = i[63533];
  assign o[63532] = i[63532];
  assign o[63531] = i[63531];
  assign o[63530] = i[63530];
  assign o[63529] = i[63529];
  assign o[63528] = i[63528];
  assign o[63527] = i[63527];
  assign o[63526] = i[63526];
  assign o[63525] = i[63525];
  assign o[63524] = i[63524];
  assign o[63523] = i[63523];
  assign o[63522] = i[63522];
  assign o[63521] = i[63521];
  assign o[63520] = i[63520];
  assign o[63519] = i[63519];
  assign o[63518] = i[63518];
  assign o[63517] = i[63517];
  assign o[63516] = i[63516];
  assign o[63515] = i[63515];
  assign o[63514] = i[63514];
  assign o[63513] = i[63513];
  assign o[63512] = i[63512];
  assign o[63511] = i[63511];
  assign o[63510] = i[63510];
  assign o[63509] = i[63509];
  assign o[63508] = i[63508];
  assign o[63507] = i[63507];
  assign o[63506] = i[63506];
  assign o[63505] = i[63505];
  assign o[63504] = i[63504];
  assign o[63503] = i[63503];
  assign o[63502] = i[63502];
  assign o[63501] = i[63501];
  assign o[63500] = i[63500];
  assign o[63499] = i[63499];
  assign o[63498] = i[63498];
  assign o[63497] = i[63497];
  assign o[63496] = i[63496];
  assign o[63495] = i[63495];
  assign o[63494] = i[63494];
  assign o[63493] = i[63493];
  assign o[63492] = i[63492];
  assign o[63491] = i[63491];
  assign o[63490] = i[63490];
  assign o[63489] = i[63489];
  assign o[63488] = i[63488];
  assign o[63487] = i[63487];
  assign o[63486] = i[63486];
  assign o[63485] = i[63485];
  assign o[63484] = i[63484];
  assign o[63483] = i[63483];
  assign o[63482] = i[63482];
  assign o[63481] = i[63481];
  assign o[63480] = i[63480];
  assign o[63479] = i[63479];
  assign o[63478] = i[63478];
  assign o[63477] = i[63477];
  assign o[63476] = i[63476];
  assign o[63475] = i[63475];
  assign o[63474] = i[63474];
  assign o[63473] = i[63473];
  assign o[63472] = i[63472];
  assign o[63471] = i[63471];
  assign o[63470] = i[63470];
  assign o[63469] = i[63469];
  assign o[63468] = i[63468];
  assign o[63467] = i[63467];
  assign o[63466] = i[63466];
  assign o[63465] = i[63465];
  assign o[63464] = i[63464];
  assign o[63463] = i[63463];
  assign o[63462] = i[63462];
  assign o[63461] = i[63461];
  assign o[63460] = i[63460];
  assign o[63459] = i[63459];
  assign o[63458] = i[63458];
  assign o[63457] = i[63457];
  assign o[63456] = i[63456];
  assign o[63455] = i[63455];
  assign o[63454] = i[63454];
  assign o[63453] = i[63453];
  assign o[63452] = i[63452];
  assign o[63451] = i[63451];
  assign o[63450] = i[63450];
  assign o[63449] = i[63449];
  assign o[63448] = i[63448];
  assign o[63447] = i[63447];
  assign o[63446] = i[63446];
  assign o[63445] = i[63445];
  assign o[63444] = i[63444];
  assign o[63443] = i[63443];
  assign o[63442] = i[63442];
  assign o[63441] = i[63441];
  assign o[63440] = i[63440];
  assign o[63439] = i[63439];
  assign o[63438] = i[63438];
  assign o[63437] = i[63437];
  assign o[63436] = i[63436];
  assign o[63435] = i[63435];
  assign o[63434] = i[63434];
  assign o[63433] = i[63433];
  assign o[63432] = i[63432];
  assign o[63431] = i[63431];
  assign o[63430] = i[63430];
  assign o[63429] = i[63429];
  assign o[63428] = i[63428];
  assign o[63427] = i[63427];
  assign o[63426] = i[63426];
  assign o[63425] = i[63425];
  assign o[63424] = i[63424];
  assign o[63423] = i[63423];
  assign o[63422] = i[63422];
  assign o[63421] = i[63421];
  assign o[63420] = i[63420];
  assign o[63419] = i[63419];
  assign o[63418] = i[63418];
  assign o[63417] = i[63417];
  assign o[63416] = i[63416];
  assign o[63415] = i[63415];
  assign o[63414] = i[63414];
  assign o[63413] = i[63413];
  assign o[63412] = i[63412];
  assign o[63411] = i[63411];
  assign o[63410] = i[63410];
  assign o[63409] = i[63409];
  assign o[63408] = i[63408];
  assign o[63407] = i[63407];
  assign o[63406] = i[63406];
  assign o[63405] = i[63405];
  assign o[63404] = i[63404];
  assign o[63403] = i[63403];
  assign o[63402] = i[63402];
  assign o[63401] = i[63401];
  assign o[63400] = i[63400];
  assign o[63399] = i[63399];
  assign o[63398] = i[63398];
  assign o[63397] = i[63397];
  assign o[63396] = i[63396];
  assign o[63395] = i[63395];
  assign o[63394] = i[63394];
  assign o[63393] = i[63393];
  assign o[63392] = i[63392];
  assign o[63391] = i[63391];
  assign o[63390] = i[63390];
  assign o[63389] = i[63389];
  assign o[63388] = i[63388];
  assign o[63387] = i[63387];
  assign o[63386] = i[63386];
  assign o[63385] = i[63385];
  assign o[63384] = i[63384];
  assign o[63383] = i[63383];
  assign o[63382] = i[63382];
  assign o[63381] = i[63381];
  assign o[63380] = i[63380];
  assign o[63379] = i[63379];
  assign o[63378] = i[63378];
  assign o[63377] = i[63377];
  assign o[63376] = i[63376];
  assign o[63375] = i[63375];
  assign o[63374] = i[63374];
  assign o[63373] = i[63373];
  assign o[63372] = i[63372];
  assign o[63371] = i[63371];
  assign o[63370] = i[63370];
  assign o[63369] = i[63369];
  assign o[63368] = i[63368];
  assign o[63367] = i[63367];
  assign o[63366] = i[63366];
  assign o[63365] = i[63365];
  assign o[63364] = i[63364];
  assign o[63363] = i[63363];
  assign o[63362] = i[63362];
  assign o[63361] = i[63361];
  assign o[63360] = i[63360];
  assign o[63359] = i[63359];
  assign o[63358] = i[63358];
  assign o[63357] = i[63357];
  assign o[63356] = i[63356];
  assign o[63355] = i[63355];
  assign o[63354] = i[63354];
  assign o[63353] = i[63353];
  assign o[63352] = i[63352];
  assign o[63351] = i[63351];
  assign o[63350] = i[63350];
  assign o[63349] = i[63349];
  assign o[63348] = i[63348];
  assign o[63347] = i[63347];
  assign o[63346] = i[63346];
  assign o[63345] = i[63345];
  assign o[63344] = i[63344];
  assign o[63343] = i[63343];
  assign o[63342] = i[63342];
  assign o[63341] = i[63341];
  assign o[63340] = i[63340];
  assign o[63339] = i[63339];
  assign o[63338] = i[63338];
  assign o[63337] = i[63337];
  assign o[63336] = i[63336];
  assign o[63335] = i[63335];
  assign o[63334] = i[63334];
  assign o[63333] = i[63333];
  assign o[63332] = i[63332];
  assign o[63331] = i[63331];
  assign o[63330] = i[63330];
  assign o[63329] = i[63329];
  assign o[63328] = i[63328];
  assign o[63327] = i[63327];
  assign o[63326] = i[63326];
  assign o[63325] = i[63325];
  assign o[63324] = i[63324];
  assign o[63323] = i[63323];
  assign o[63322] = i[63322];
  assign o[63321] = i[63321];
  assign o[63320] = i[63320];
  assign o[63319] = i[63319];
  assign o[63318] = i[63318];
  assign o[63317] = i[63317];
  assign o[63316] = i[63316];
  assign o[63315] = i[63315];
  assign o[63314] = i[63314];
  assign o[63313] = i[63313];
  assign o[63312] = i[63312];
  assign o[63311] = i[63311];
  assign o[63310] = i[63310];
  assign o[63309] = i[63309];
  assign o[63308] = i[63308];
  assign o[63307] = i[63307];
  assign o[63306] = i[63306];
  assign o[63305] = i[63305];
  assign o[63304] = i[63304];
  assign o[63303] = i[63303];
  assign o[63302] = i[63302];
  assign o[63301] = i[63301];
  assign o[63300] = i[63300];
  assign o[63299] = i[63299];
  assign o[63298] = i[63298];
  assign o[63297] = i[63297];
  assign o[63296] = i[63296];
  assign o[63295] = i[63295];
  assign o[63294] = i[63294];
  assign o[63293] = i[63293];
  assign o[63292] = i[63292];
  assign o[63291] = i[63291];
  assign o[63290] = i[63290];
  assign o[63289] = i[63289];
  assign o[63288] = i[63288];
  assign o[63287] = i[63287];
  assign o[63286] = i[63286];
  assign o[63285] = i[63285];
  assign o[63284] = i[63284];
  assign o[63283] = i[63283];
  assign o[63282] = i[63282];
  assign o[63281] = i[63281];
  assign o[63280] = i[63280];
  assign o[63279] = i[63279];
  assign o[63278] = i[63278];
  assign o[63277] = i[63277];
  assign o[63276] = i[63276];
  assign o[63275] = i[63275];
  assign o[63274] = i[63274];
  assign o[63273] = i[63273];
  assign o[63272] = i[63272];
  assign o[63271] = i[63271];
  assign o[63270] = i[63270];
  assign o[63269] = i[63269];
  assign o[63268] = i[63268];
  assign o[63267] = i[63267];
  assign o[63266] = i[63266];
  assign o[63265] = i[63265];
  assign o[63264] = i[63264];
  assign o[63263] = i[63263];
  assign o[63262] = i[63262];
  assign o[63261] = i[63261];
  assign o[63260] = i[63260];
  assign o[63259] = i[63259];
  assign o[63258] = i[63258];
  assign o[63257] = i[63257];
  assign o[63256] = i[63256];
  assign o[63255] = i[63255];
  assign o[63254] = i[63254];
  assign o[63253] = i[63253];
  assign o[63252] = i[63252];
  assign o[63251] = i[63251];
  assign o[63250] = i[63250];
  assign o[63249] = i[63249];
  assign o[63248] = i[63248];
  assign o[63247] = i[63247];
  assign o[63246] = i[63246];
  assign o[63245] = i[63245];
  assign o[63244] = i[63244];
  assign o[63243] = i[63243];
  assign o[63242] = i[63242];
  assign o[63241] = i[63241];
  assign o[63240] = i[63240];
  assign o[63239] = i[63239];
  assign o[63238] = i[63238];
  assign o[63237] = i[63237];
  assign o[63236] = i[63236];
  assign o[63235] = i[63235];
  assign o[63234] = i[63234];
  assign o[63233] = i[63233];
  assign o[63232] = i[63232];
  assign o[63231] = i[63231];
  assign o[63230] = i[63230];
  assign o[63229] = i[63229];
  assign o[63228] = i[63228];
  assign o[63227] = i[63227];
  assign o[63226] = i[63226];
  assign o[63225] = i[63225];
  assign o[63224] = i[63224];
  assign o[63223] = i[63223];
  assign o[63222] = i[63222];
  assign o[63221] = i[63221];
  assign o[63220] = i[63220];
  assign o[63219] = i[63219];
  assign o[63218] = i[63218];
  assign o[63217] = i[63217];
  assign o[63216] = i[63216];
  assign o[63215] = i[63215];
  assign o[63214] = i[63214];
  assign o[63213] = i[63213];
  assign o[63212] = i[63212];
  assign o[63211] = i[63211];
  assign o[63210] = i[63210];
  assign o[63209] = i[63209];
  assign o[63208] = i[63208];
  assign o[63207] = i[63207];
  assign o[63206] = i[63206];
  assign o[63205] = i[63205];
  assign o[63204] = i[63204];
  assign o[63203] = i[63203];
  assign o[63202] = i[63202];
  assign o[63201] = i[63201];
  assign o[63200] = i[63200];
  assign o[63199] = i[63199];
  assign o[63198] = i[63198];
  assign o[63197] = i[63197];
  assign o[63196] = i[63196];
  assign o[63195] = i[63195];
  assign o[63194] = i[63194];
  assign o[63193] = i[63193];
  assign o[63192] = i[63192];
  assign o[63191] = i[63191];
  assign o[63190] = i[63190];
  assign o[63189] = i[63189];
  assign o[63188] = i[63188];
  assign o[63187] = i[63187];
  assign o[63186] = i[63186];
  assign o[63185] = i[63185];
  assign o[63184] = i[63184];
  assign o[63183] = i[63183];
  assign o[63182] = i[63182];
  assign o[63181] = i[63181];
  assign o[63180] = i[63180];
  assign o[63179] = i[63179];
  assign o[63178] = i[63178];
  assign o[63177] = i[63177];
  assign o[63176] = i[63176];
  assign o[63175] = i[63175];
  assign o[63174] = i[63174];
  assign o[63173] = i[63173];
  assign o[63172] = i[63172];
  assign o[63171] = i[63171];
  assign o[63170] = i[63170];
  assign o[63169] = i[63169];
  assign o[63168] = i[63168];
  assign o[63167] = i[63167];
  assign o[63166] = i[63166];
  assign o[63165] = i[63165];
  assign o[63164] = i[63164];
  assign o[63163] = i[63163];
  assign o[63162] = i[63162];
  assign o[63161] = i[63161];
  assign o[63160] = i[63160];
  assign o[63159] = i[63159];
  assign o[63158] = i[63158];
  assign o[63157] = i[63157];
  assign o[63156] = i[63156];
  assign o[63155] = i[63155];
  assign o[63154] = i[63154];
  assign o[63153] = i[63153];
  assign o[63152] = i[63152];
  assign o[63151] = i[63151];
  assign o[63150] = i[63150];
  assign o[63149] = i[63149];
  assign o[63148] = i[63148];
  assign o[63147] = i[63147];
  assign o[63146] = i[63146];
  assign o[63145] = i[63145];
  assign o[63144] = i[63144];
  assign o[63143] = i[63143];
  assign o[63142] = i[63142];
  assign o[63141] = i[63141];
  assign o[63140] = i[63140];
  assign o[63139] = i[63139];
  assign o[63138] = i[63138];
  assign o[63137] = i[63137];
  assign o[63136] = i[63136];
  assign o[63135] = i[63135];
  assign o[63134] = i[63134];
  assign o[63133] = i[63133];
  assign o[63132] = i[63132];
  assign o[63131] = i[63131];
  assign o[63130] = i[63130];
  assign o[63129] = i[63129];
  assign o[63128] = i[63128];
  assign o[63127] = i[63127];
  assign o[63126] = i[63126];
  assign o[63125] = i[63125];
  assign o[63124] = i[63124];
  assign o[63123] = i[63123];
  assign o[63122] = i[63122];
  assign o[63121] = i[63121];
  assign o[63120] = i[63120];
  assign o[63119] = i[63119];
  assign o[63118] = i[63118];
  assign o[63117] = i[63117];
  assign o[63116] = i[63116];
  assign o[63115] = i[63115];
  assign o[63114] = i[63114];
  assign o[63113] = i[63113];
  assign o[63112] = i[63112];
  assign o[63111] = i[63111];
  assign o[63110] = i[63110];
  assign o[63109] = i[63109];
  assign o[63108] = i[63108];
  assign o[63107] = i[63107];
  assign o[63106] = i[63106];
  assign o[63105] = i[63105];
  assign o[63104] = i[63104];
  assign o[63103] = i[63103];
  assign o[63102] = i[63102];
  assign o[63101] = i[63101];
  assign o[63100] = i[63100];
  assign o[63099] = i[63099];
  assign o[63098] = i[63098];
  assign o[63097] = i[63097];
  assign o[63096] = i[63096];
  assign o[63095] = i[63095];
  assign o[63094] = i[63094];
  assign o[63093] = i[63093];
  assign o[63092] = i[63092];
  assign o[63091] = i[63091];
  assign o[63090] = i[63090];
  assign o[63089] = i[63089];
  assign o[63088] = i[63088];
  assign o[63087] = i[63087];
  assign o[63086] = i[63086];
  assign o[63085] = i[63085];
  assign o[63084] = i[63084];
  assign o[63083] = i[63083];
  assign o[63082] = i[63082];
  assign o[63081] = i[63081];
  assign o[63080] = i[63080];
  assign o[63079] = i[63079];
  assign o[63078] = i[63078];
  assign o[63077] = i[63077];
  assign o[63076] = i[63076];
  assign o[63075] = i[63075];
  assign o[63074] = i[63074];
  assign o[63073] = i[63073];
  assign o[63072] = i[63072];
  assign o[63071] = i[63071];
  assign o[63070] = i[63070];
  assign o[63069] = i[63069];
  assign o[63068] = i[63068];
  assign o[63067] = i[63067];
  assign o[63066] = i[63066];
  assign o[63065] = i[63065];
  assign o[63064] = i[63064];
  assign o[63063] = i[63063];
  assign o[63062] = i[63062];
  assign o[63061] = i[63061];
  assign o[63060] = i[63060];
  assign o[63059] = i[63059];
  assign o[63058] = i[63058];
  assign o[63057] = i[63057];
  assign o[63056] = i[63056];
  assign o[63055] = i[63055];
  assign o[63054] = i[63054];
  assign o[63053] = i[63053];
  assign o[63052] = i[63052];
  assign o[63051] = i[63051];
  assign o[63050] = i[63050];
  assign o[63049] = i[63049];
  assign o[63048] = i[63048];
  assign o[63047] = i[63047];
  assign o[63046] = i[63046];
  assign o[63045] = i[63045];
  assign o[63044] = i[63044];
  assign o[63043] = i[63043];
  assign o[63042] = i[63042];
  assign o[63041] = i[63041];
  assign o[63040] = i[63040];
  assign o[63039] = i[63039];
  assign o[63038] = i[63038];
  assign o[63037] = i[63037];
  assign o[63036] = i[63036];
  assign o[63035] = i[63035];
  assign o[63034] = i[63034];
  assign o[63033] = i[63033];
  assign o[63032] = i[63032];
  assign o[63031] = i[63031];
  assign o[63030] = i[63030];
  assign o[63029] = i[63029];
  assign o[63028] = i[63028];
  assign o[63027] = i[63027];
  assign o[63026] = i[63026];
  assign o[63025] = i[63025];
  assign o[63024] = i[63024];
  assign o[63023] = i[63023];
  assign o[63022] = i[63022];
  assign o[63021] = i[63021];
  assign o[63020] = i[63020];
  assign o[63019] = i[63019];
  assign o[63018] = i[63018];
  assign o[63017] = i[63017];
  assign o[63016] = i[63016];
  assign o[63015] = i[63015];
  assign o[63014] = i[63014];
  assign o[63013] = i[63013];
  assign o[63012] = i[63012];
  assign o[63011] = i[63011];
  assign o[63010] = i[63010];
  assign o[63009] = i[63009];
  assign o[63008] = i[63008];
  assign o[63007] = i[63007];
  assign o[63006] = i[63006];
  assign o[63005] = i[63005];
  assign o[63004] = i[63004];
  assign o[63003] = i[63003];
  assign o[63002] = i[63002];
  assign o[63001] = i[63001];
  assign o[63000] = i[63000];
  assign o[62999] = i[62999];
  assign o[62998] = i[62998];
  assign o[62997] = i[62997];
  assign o[62996] = i[62996];
  assign o[62995] = i[62995];
  assign o[62994] = i[62994];
  assign o[62993] = i[62993];
  assign o[62992] = i[62992];
  assign o[62991] = i[62991];
  assign o[62990] = i[62990];
  assign o[62989] = i[62989];
  assign o[62988] = i[62988];
  assign o[62987] = i[62987];
  assign o[62986] = i[62986];
  assign o[62985] = i[62985];
  assign o[62984] = i[62984];
  assign o[62983] = i[62983];
  assign o[62982] = i[62982];
  assign o[62981] = i[62981];
  assign o[62980] = i[62980];
  assign o[62979] = i[62979];
  assign o[62978] = i[62978];
  assign o[62977] = i[62977];
  assign o[62976] = i[62976];
  assign o[62975] = i[62975];
  assign o[62974] = i[62974];
  assign o[62973] = i[62973];
  assign o[62972] = i[62972];
  assign o[62971] = i[62971];
  assign o[62970] = i[62970];
  assign o[62969] = i[62969];
  assign o[62968] = i[62968];
  assign o[62967] = i[62967];
  assign o[62966] = i[62966];
  assign o[62965] = i[62965];
  assign o[62964] = i[62964];
  assign o[62963] = i[62963];
  assign o[62962] = i[62962];
  assign o[62961] = i[62961];
  assign o[62960] = i[62960];
  assign o[62959] = i[62959];
  assign o[62958] = i[62958];
  assign o[62957] = i[62957];
  assign o[62956] = i[62956];
  assign o[62955] = i[62955];
  assign o[62954] = i[62954];
  assign o[62953] = i[62953];
  assign o[62952] = i[62952];
  assign o[62951] = i[62951];
  assign o[62950] = i[62950];
  assign o[62949] = i[62949];
  assign o[62948] = i[62948];
  assign o[62947] = i[62947];
  assign o[62946] = i[62946];
  assign o[62945] = i[62945];
  assign o[62944] = i[62944];
  assign o[62943] = i[62943];
  assign o[62942] = i[62942];
  assign o[62941] = i[62941];
  assign o[62940] = i[62940];
  assign o[62939] = i[62939];
  assign o[62938] = i[62938];
  assign o[62937] = i[62937];
  assign o[62936] = i[62936];
  assign o[62935] = i[62935];
  assign o[62934] = i[62934];
  assign o[62933] = i[62933];
  assign o[62932] = i[62932];
  assign o[62931] = i[62931];
  assign o[62930] = i[62930];
  assign o[62929] = i[62929];
  assign o[62928] = i[62928];
  assign o[62927] = i[62927];
  assign o[62926] = i[62926];
  assign o[62925] = i[62925];
  assign o[62924] = i[62924];
  assign o[62923] = i[62923];
  assign o[62922] = i[62922];
  assign o[62921] = i[62921];
  assign o[62920] = i[62920];
  assign o[62919] = i[62919];
  assign o[62918] = i[62918];
  assign o[62917] = i[62917];
  assign o[62916] = i[62916];
  assign o[62915] = i[62915];
  assign o[62914] = i[62914];
  assign o[62913] = i[62913];
  assign o[62912] = i[62912];
  assign o[62911] = i[62911];
  assign o[62910] = i[62910];
  assign o[62909] = i[62909];
  assign o[62908] = i[62908];
  assign o[62907] = i[62907];
  assign o[62906] = i[62906];
  assign o[62905] = i[62905];
  assign o[62904] = i[62904];
  assign o[62903] = i[62903];
  assign o[62902] = i[62902];
  assign o[62901] = i[62901];
  assign o[62900] = i[62900];
  assign o[62899] = i[62899];
  assign o[62898] = i[62898];
  assign o[62897] = i[62897];
  assign o[62896] = i[62896];
  assign o[62895] = i[62895];
  assign o[62894] = i[62894];
  assign o[62893] = i[62893];
  assign o[62892] = i[62892];
  assign o[62891] = i[62891];
  assign o[62890] = i[62890];
  assign o[62889] = i[62889];
  assign o[62888] = i[62888];
  assign o[62887] = i[62887];
  assign o[62886] = i[62886];
  assign o[62885] = i[62885];
  assign o[62884] = i[62884];
  assign o[62883] = i[62883];
  assign o[62882] = i[62882];
  assign o[62881] = i[62881];
  assign o[62880] = i[62880];
  assign o[62879] = i[62879];
  assign o[62878] = i[62878];
  assign o[62877] = i[62877];
  assign o[62876] = i[62876];
  assign o[62875] = i[62875];
  assign o[62874] = i[62874];
  assign o[62873] = i[62873];
  assign o[62872] = i[62872];
  assign o[62871] = i[62871];
  assign o[62870] = i[62870];
  assign o[62869] = i[62869];
  assign o[62868] = i[62868];
  assign o[62867] = i[62867];
  assign o[62866] = i[62866];
  assign o[62865] = i[62865];
  assign o[62864] = i[62864];
  assign o[62863] = i[62863];
  assign o[62862] = i[62862];
  assign o[62861] = i[62861];
  assign o[62860] = i[62860];
  assign o[62859] = i[62859];
  assign o[62858] = i[62858];
  assign o[62857] = i[62857];
  assign o[62856] = i[62856];
  assign o[62855] = i[62855];
  assign o[62854] = i[62854];
  assign o[62853] = i[62853];
  assign o[62852] = i[62852];
  assign o[62851] = i[62851];
  assign o[62850] = i[62850];
  assign o[62849] = i[62849];
  assign o[62848] = i[62848];
  assign o[62847] = i[62847];
  assign o[62846] = i[62846];
  assign o[62845] = i[62845];
  assign o[62844] = i[62844];
  assign o[62843] = i[62843];
  assign o[62842] = i[62842];
  assign o[62841] = i[62841];
  assign o[62840] = i[62840];
  assign o[62839] = i[62839];
  assign o[62838] = i[62838];
  assign o[62837] = i[62837];
  assign o[62836] = i[62836];
  assign o[62835] = i[62835];
  assign o[62834] = i[62834];
  assign o[62833] = i[62833];
  assign o[62832] = i[62832];
  assign o[62831] = i[62831];
  assign o[62830] = i[62830];
  assign o[62829] = i[62829];
  assign o[62828] = i[62828];
  assign o[62827] = i[62827];
  assign o[62826] = i[62826];
  assign o[62825] = i[62825];
  assign o[62824] = i[62824];
  assign o[62823] = i[62823];
  assign o[62822] = i[62822];
  assign o[62821] = i[62821];
  assign o[62820] = i[62820];
  assign o[62819] = i[62819];
  assign o[62818] = i[62818];
  assign o[62817] = i[62817];
  assign o[62816] = i[62816];
  assign o[62815] = i[62815];
  assign o[62814] = i[62814];
  assign o[62813] = i[62813];
  assign o[62812] = i[62812];
  assign o[62811] = i[62811];
  assign o[62810] = i[62810];
  assign o[62809] = i[62809];
  assign o[62808] = i[62808];
  assign o[62807] = i[62807];
  assign o[62806] = i[62806];
  assign o[62805] = i[62805];
  assign o[62804] = i[62804];
  assign o[62803] = i[62803];
  assign o[62802] = i[62802];
  assign o[62801] = i[62801];
  assign o[62800] = i[62800];
  assign o[62799] = i[62799];
  assign o[62798] = i[62798];
  assign o[62797] = i[62797];
  assign o[62796] = i[62796];
  assign o[62795] = i[62795];
  assign o[62794] = i[62794];
  assign o[62793] = i[62793];
  assign o[62792] = i[62792];
  assign o[62791] = i[62791];
  assign o[62790] = i[62790];
  assign o[62789] = i[62789];
  assign o[62788] = i[62788];
  assign o[62787] = i[62787];
  assign o[62786] = i[62786];
  assign o[62785] = i[62785];
  assign o[62784] = i[62784];
  assign o[62783] = i[62783];
  assign o[62782] = i[62782];
  assign o[62781] = i[62781];
  assign o[62780] = i[62780];
  assign o[62779] = i[62779];
  assign o[62778] = i[62778];
  assign o[62777] = i[62777];
  assign o[62776] = i[62776];
  assign o[62775] = i[62775];
  assign o[62774] = i[62774];
  assign o[62773] = i[62773];
  assign o[62772] = i[62772];
  assign o[62771] = i[62771];
  assign o[62770] = i[62770];
  assign o[62769] = i[62769];
  assign o[62768] = i[62768];
  assign o[62767] = i[62767];
  assign o[62766] = i[62766];
  assign o[62765] = i[62765];
  assign o[62764] = i[62764];
  assign o[62763] = i[62763];
  assign o[62762] = i[62762];
  assign o[62761] = i[62761];
  assign o[62760] = i[62760];
  assign o[62759] = i[62759];
  assign o[62758] = i[62758];
  assign o[62757] = i[62757];
  assign o[62756] = i[62756];
  assign o[62755] = i[62755];
  assign o[62754] = i[62754];
  assign o[62753] = i[62753];
  assign o[62752] = i[62752];
  assign o[62751] = i[62751];
  assign o[62750] = i[62750];
  assign o[62749] = i[62749];
  assign o[62748] = i[62748];
  assign o[62747] = i[62747];
  assign o[62746] = i[62746];
  assign o[62745] = i[62745];
  assign o[62744] = i[62744];
  assign o[62743] = i[62743];
  assign o[62742] = i[62742];
  assign o[62741] = i[62741];
  assign o[62740] = i[62740];
  assign o[62739] = i[62739];
  assign o[62738] = i[62738];
  assign o[62737] = i[62737];
  assign o[62736] = i[62736];
  assign o[62735] = i[62735];
  assign o[62734] = i[62734];
  assign o[62733] = i[62733];
  assign o[62732] = i[62732];
  assign o[62731] = i[62731];
  assign o[62730] = i[62730];
  assign o[62729] = i[62729];
  assign o[62728] = i[62728];
  assign o[62727] = i[62727];
  assign o[62726] = i[62726];
  assign o[62725] = i[62725];
  assign o[62724] = i[62724];
  assign o[62723] = i[62723];
  assign o[62722] = i[62722];
  assign o[62721] = i[62721];
  assign o[62720] = i[62720];
  assign o[62719] = i[62719];
  assign o[62718] = i[62718];
  assign o[62717] = i[62717];
  assign o[62716] = i[62716];
  assign o[62715] = i[62715];
  assign o[62714] = i[62714];
  assign o[62713] = i[62713];
  assign o[62712] = i[62712];
  assign o[62711] = i[62711];
  assign o[62710] = i[62710];
  assign o[62709] = i[62709];
  assign o[62708] = i[62708];
  assign o[62707] = i[62707];
  assign o[62706] = i[62706];
  assign o[62705] = i[62705];
  assign o[62704] = i[62704];
  assign o[62703] = i[62703];
  assign o[62702] = i[62702];
  assign o[62701] = i[62701];
  assign o[62700] = i[62700];
  assign o[62699] = i[62699];
  assign o[62698] = i[62698];
  assign o[62697] = i[62697];
  assign o[62696] = i[62696];
  assign o[62695] = i[62695];
  assign o[62694] = i[62694];
  assign o[62693] = i[62693];
  assign o[62692] = i[62692];
  assign o[62691] = i[62691];
  assign o[62690] = i[62690];
  assign o[62689] = i[62689];
  assign o[62688] = i[62688];
  assign o[62687] = i[62687];
  assign o[62686] = i[62686];
  assign o[62685] = i[62685];
  assign o[62684] = i[62684];
  assign o[62683] = i[62683];
  assign o[62682] = i[62682];
  assign o[62681] = i[62681];
  assign o[62680] = i[62680];
  assign o[62679] = i[62679];
  assign o[62678] = i[62678];
  assign o[62677] = i[62677];
  assign o[62676] = i[62676];
  assign o[62675] = i[62675];
  assign o[62674] = i[62674];
  assign o[62673] = i[62673];
  assign o[62672] = i[62672];
  assign o[62671] = i[62671];
  assign o[62670] = i[62670];
  assign o[62669] = i[62669];
  assign o[62668] = i[62668];
  assign o[62667] = i[62667];
  assign o[62666] = i[62666];
  assign o[62665] = i[62665];
  assign o[62664] = i[62664];
  assign o[62663] = i[62663];
  assign o[62662] = i[62662];
  assign o[62661] = i[62661];
  assign o[62660] = i[62660];
  assign o[62659] = i[62659];
  assign o[62658] = i[62658];
  assign o[62657] = i[62657];
  assign o[62656] = i[62656];
  assign o[62655] = i[62655];
  assign o[62654] = i[62654];
  assign o[62653] = i[62653];
  assign o[62652] = i[62652];
  assign o[62651] = i[62651];
  assign o[62650] = i[62650];
  assign o[62649] = i[62649];
  assign o[62648] = i[62648];
  assign o[62647] = i[62647];
  assign o[62646] = i[62646];
  assign o[62645] = i[62645];
  assign o[62644] = i[62644];
  assign o[62643] = i[62643];
  assign o[62642] = i[62642];
  assign o[62641] = i[62641];
  assign o[62640] = i[62640];
  assign o[62639] = i[62639];
  assign o[62638] = i[62638];
  assign o[62637] = i[62637];
  assign o[62636] = i[62636];
  assign o[62635] = i[62635];
  assign o[62634] = i[62634];
  assign o[62633] = i[62633];
  assign o[62632] = i[62632];
  assign o[62631] = i[62631];
  assign o[62630] = i[62630];
  assign o[62629] = i[62629];
  assign o[62628] = i[62628];
  assign o[62627] = i[62627];
  assign o[62626] = i[62626];
  assign o[62625] = i[62625];
  assign o[62624] = i[62624];
  assign o[62623] = i[62623];
  assign o[62622] = i[62622];
  assign o[62621] = i[62621];
  assign o[62620] = i[62620];
  assign o[62619] = i[62619];
  assign o[62618] = i[62618];
  assign o[62617] = i[62617];
  assign o[62616] = i[62616];
  assign o[62615] = i[62615];
  assign o[62614] = i[62614];
  assign o[62613] = i[62613];
  assign o[62612] = i[62612];
  assign o[62611] = i[62611];
  assign o[62610] = i[62610];
  assign o[62609] = i[62609];
  assign o[62608] = i[62608];
  assign o[62607] = i[62607];
  assign o[62606] = i[62606];
  assign o[62605] = i[62605];
  assign o[62604] = i[62604];
  assign o[62603] = i[62603];
  assign o[62602] = i[62602];
  assign o[62601] = i[62601];
  assign o[62600] = i[62600];
  assign o[62599] = i[62599];
  assign o[62598] = i[62598];
  assign o[62597] = i[62597];
  assign o[62596] = i[62596];
  assign o[62595] = i[62595];
  assign o[62594] = i[62594];
  assign o[62593] = i[62593];
  assign o[62592] = i[62592];
  assign o[62591] = i[62591];
  assign o[62590] = i[62590];
  assign o[62589] = i[62589];
  assign o[62588] = i[62588];
  assign o[62587] = i[62587];
  assign o[62586] = i[62586];
  assign o[62585] = i[62585];
  assign o[62584] = i[62584];
  assign o[62583] = i[62583];
  assign o[62582] = i[62582];
  assign o[62581] = i[62581];
  assign o[62580] = i[62580];
  assign o[62579] = i[62579];
  assign o[62578] = i[62578];
  assign o[62577] = i[62577];
  assign o[62576] = i[62576];
  assign o[62575] = i[62575];
  assign o[62574] = i[62574];
  assign o[62573] = i[62573];
  assign o[62572] = i[62572];
  assign o[62571] = i[62571];
  assign o[62570] = i[62570];
  assign o[62569] = i[62569];
  assign o[62568] = i[62568];
  assign o[62567] = i[62567];
  assign o[62566] = i[62566];
  assign o[62565] = i[62565];
  assign o[62564] = i[62564];
  assign o[62563] = i[62563];
  assign o[62562] = i[62562];
  assign o[62561] = i[62561];
  assign o[62560] = i[62560];
  assign o[62559] = i[62559];
  assign o[62558] = i[62558];
  assign o[62557] = i[62557];
  assign o[62556] = i[62556];
  assign o[62555] = i[62555];
  assign o[62554] = i[62554];
  assign o[62553] = i[62553];
  assign o[62552] = i[62552];
  assign o[62551] = i[62551];
  assign o[62550] = i[62550];
  assign o[62549] = i[62549];
  assign o[62548] = i[62548];
  assign o[62547] = i[62547];
  assign o[62546] = i[62546];
  assign o[62545] = i[62545];
  assign o[62544] = i[62544];
  assign o[62543] = i[62543];
  assign o[62542] = i[62542];
  assign o[62541] = i[62541];
  assign o[62540] = i[62540];
  assign o[62539] = i[62539];
  assign o[62538] = i[62538];
  assign o[62537] = i[62537];
  assign o[62536] = i[62536];
  assign o[62535] = i[62535];
  assign o[62534] = i[62534];
  assign o[62533] = i[62533];
  assign o[62532] = i[62532];
  assign o[62531] = i[62531];
  assign o[62530] = i[62530];
  assign o[62529] = i[62529];
  assign o[62528] = i[62528];
  assign o[62527] = i[62527];
  assign o[62526] = i[62526];
  assign o[62525] = i[62525];
  assign o[62524] = i[62524];
  assign o[62523] = i[62523];
  assign o[62522] = i[62522];
  assign o[62521] = i[62521];
  assign o[62520] = i[62520];
  assign o[62519] = i[62519];
  assign o[62518] = i[62518];
  assign o[62517] = i[62517];
  assign o[62516] = i[62516];
  assign o[62515] = i[62515];
  assign o[62514] = i[62514];
  assign o[62513] = i[62513];
  assign o[62512] = i[62512];
  assign o[62511] = i[62511];
  assign o[62510] = i[62510];
  assign o[62509] = i[62509];
  assign o[62508] = i[62508];
  assign o[62507] = i[62507];
  assign o[62506] = i[62506];
  assign o[62505] = i[62505];
  assign o[62504] = i[62504];
  assign o[62503] = i[62503];
  assign o[62502] = i[62502];
  assign o[62501] = i[62501];
  assign o[62500] = i[62500];
  assign o[62499] = i[62499];
  assign o[62498] = i[62498];
  assign o[62497] = i[62497];
  assign o[62496] = i[62496];
  assign o[62495] = i[62495];
  assign o[62494] = i[62494];
  assign o[62493] = i[62493];
  assign o[62492] = i[62492];
  assign o[62491] = i[62491];
  assign o[62490] = i[62490];
  assign o[62489] = i[62489];
  assign o[62488] = i[62488];
  assign o[62487] = i[62487];
  assign o[62486] = i[62486];
  assign o[62485] = i[62485];
  assign o[62484] = i[62484];
  assign o[62483] = i[62483];
  assign o[62482] = i[62482];
  assign o[62481] = i[62481];
  assign o[62480] = i[62480];
  assign o[62479] = i[62479];
  assign o[62478] = i[62478];
  assign o[62477] = i[62477];
  assign o[62476] = i[62476];
  assign o[62475] = i[62475];
  assign o[62474] = i[62474];
  assign o[62473] = i[62473];
  assign o[62472] = i[62472];
  assign o[62471] = i[62471];
  assign o[62470] = i[62470];
  assign o[62469] = i[62469];
  assign o[62468] = i[62468];
  assign o[62467] = i[62467];
  assign o[62466] = i[62466];
  assign o[62465] = i[62465];
  assign o[62464] = i[62464];
  assign o[62463] = i[62463];
  assign o[62462] = i[62462];
  assign o[62461] = i[62461];
  assign o[62460] = i[62460];
  assign o[62459] = i[62459];
  assign o[62458] = i[62458];
  assign o[62457] = i[62457];
  assign o[62456] = i[62456];
  assign o[62455] = i[62455];
  assign o[62454] = i[62454];
  assign o[62453] = i[62453];
  assign o[62452] = i[62452];
  assign o[62451] = i[62451];
  assign o[62450] = i[62450];
  assign o[62449] = i[62449];
  assign o[62448] = i[62448];
  assign o[62447] = i[62447];
  assign o[62446] = i[62446];
  assign o[62445] = i[62445];
  assign o[62444] = i[62444];
  assign o[62443] = i[62443];
  assign o[62442] = i[62442];
  assign o[62441] = i[62441];
  assign o[62440] = i[62440];
  assign o[62439] = i[62439];
  assign o[62438] = i[62438];
  assign o[62437] = i[62437];
  assign o[62436] = i[62436];
  assign o[62435] = i[62435];
  assign o[62434] = i[62434];
  assign o[62433] = i[62433];
  assign o[62432] = i[62432];
  assign o[62431] = i[62431];
  assign o[62430] = i[62430];
  assign o[62429] = i[62429];
  assign o[62428] = i[62428];
  assign o[62427] = i[62427];
  assign o[62426] = i[62426];
  assign o[62425] = i[62425];
  assign o[62424] = i[62424];
  assign o[62423] = i[62423];
  assign o[62422] = i[62422];
  assign o[62421] = i[62421];
  assign o[62420] = i[62420];
  assign o[62419] = i[62419];
  assign o[62418] = i[62418];
  assign o[62417] = i[62417];
  assign o[62416] = i[62416];
  assign o[62415] = i[62415];
  assign o[62414] = i[62414];
  assign o[62413] = i[62413];
  assign o[62412] = i[62412];
  assign o[62411] = i[62411];
  assign o[62410] = i[62410];
  assign o[62409] = i[62409];
  assign o[62408] = i[62408];
  assign o[62407] = i[62407];
  assign o[62406] = i[62406];
  assign o[62405] = i[62405];
  assign o[62404] = i[62404];
  assign o[62403] = i[62403];
  assign o[62402] = i[62402];
  assign o[62401] = i[62401];
  assign o[62400] = i[62400];
  assign o[62399] = i[62399];
  assign o[62398] = i[62398];
  assign o[62397] = i[62397];
  assign o[62396] = i[62396];
  assign o[62395] = i[62395];
  assign o[62394] = i[62394];
  assign o[62393] = i[62393];
  assign o[62392] = i[62392];
  assign o[62391] = i[62391];
  assign o[62390] = i[62390];
  assign o[62389] = i[62389];
  assign o[62388] = i[62388];
  assign o[62387] = i[62387];
  assign o[62386] = i[62386];
  assign o[62385] = i[62385];
  assign o[62384] = i[62384];
  assign o[62383] = i[62383];
  assign o[62382] = i[62382];
  assign o[62381] = i[62381];
  assign o[62380] = i[62380];
  assign o[62379] = i[62379];
  assign o[62378] = i[62378];
  assign o[62377] = i[62377];
  assign o[62376] = i[62376];
  assign o[62375] = i[62375];
  assign o[62374] = i[62374];
  assign o[62373] = i[62373];
  assign o[62372] = i[62372];
  assign o[62371] = i[62371];
  assign o[62370] = i[62370];
  assign o[62369] = i[62369];
  assign o[62368] = i[62368];
  assign o[62367] = i[62367];
  assign o[62366] = i[62366];
  assign o[62365] = i[62365];
  assign o[62364] = i[62364];
  assign o[62363] = i[62363];
  assign o[62362] = i[62362];
  assign o[62361] = i[62361];
  assign o[62360] = i[62360];
  assign o[62359] = i[62359];
  assign o[62358] = i[62358];
  assign o[62357] = i[62357];
  assign o[62356] = i[62356];
  assign o[62355] = i[62355];
  assign o[62354] = i[62354];
  assign o[62353] = i[62353];
  assign o[62352] = i[62352];
  assign o[62351] = i[62351];
  assign o[62350] = i[62350];
  assign o[62349] = i[62349];
  assign o[62348] = i[62348];
  assign o[62347] = i[62347];
  assign o[62346] = i[62346];
  assign o[62345] = i[62345];
  assign o[62344] = i[62344];
  assign o[62343] = i[62343];
  assign o[62342] = i[62342];
  assign o[62341] = i[62341];
  assign o[62340] = i[62340];
  assign o[62339] = i[62339];
  assign o[62338] = i[62338];
  assign o[62337] = i[62337];
  assign o[62336] = i[62336];
  assign o[62335] = i[62335];
  assign o[62334] = i[62334];
  assign o[62333] = i[62333];
  assign o[62332] = i[62332];
  assign o[62331] = i[62331];
  assign o[62330] = i[62330];
  assign o[62329] = i[62329];
  assign o[62328] = i[62328];
  assign o[62327] = i[62327];
  assign o[62326] = i[62326];
  assign o[62325] = i[62325];
  assign o[62324] = i[62324];
  assign o[62323] = i[62323];
  assign o[62322] = i[62322];
  assign o[62321] = i[62321];
  assign o[62320] = i[62320];
  assign o[62319] = i[62319];
  assign o[62318] = i[62318];
  assign o[62317] = i[62317];
  assign o[62316] = i[62316];
  assign o[62315] = i[62315];
  assign o[62314] = i[62314];
  assign o[62313] = i[62313];
  assign o[62312] = i[62312];
  assign o[62311] = i[62311];
  assign o[62310] = i[62310];
  assign o[62309] = i[62309];
  assign o[62308] = i[62308];
  assign o[62307] = i[62307];
  assign o[62306] = i[62306];
  assign o[62305] = i[62305];
  assign o[62304] = i[62304];
  assign o[62303] = i[62303];
  assign o[62302] = i[62302];
  assign o[62301] = i[62301];
  assign o[62300] = i[62300];
  assign o[62299] = i[62299];
  assign o[62298] = i[62298];
  assign o[62297] = i[62297];
  assign o[62296] = i[62296];
  assign o[62295] = i[62295];
  assign o[62294] = i[62294];
  assign o[62293] = i[62293];
  assign o[62292] = i[62292];
  assign o[62291] = i[62291];
  assign o[62290] = i[62290];
  assign o[62289] = i[62289];
  assign o[62288] = i[62288];
  assign o[62287] = i[62287];
  assign o[62286] = i[62286];
  assign o[62285] = i[62285];
  assign o[62284] = i[62284];
  assign o[62283] = i[62283];
  assign o[62282] = i[62282];
  assign o[62281] = i[62281];
  assign o[62280] = i[62280];
  assign o[62279] = i[62279];
  assign o[62278] = i[62278];
  assign o[62277] = i[62277];
  assign o[62276] = i[62276];
  assign o[62275] = i[62275];
  assign o[62274] = i[62274];
  assign o[62273] = i[62273];
  assign o[62272] = i[62272];
  assign o[62271] = i[62271];
  assign o[62270] = i[62270];
  assign o[62269] = i[62269];
  assign o[62268] = i[62268];
  assign o[62267] = i[62267];
  assign o[62266] = i[62266];
  assign o[62265] = i[62265];
  assign o[62264] = i[62264];
  assign o[62263] = i[62263];
  assign o[62262] = i[62262];
  assign o[62261] = i[62261];
  assign o[62260] = i[62260];
  assign o[62259] = i[62259];
  assign o[62258] = i[62258];
  assign o[62257] = i[62257];
  assign o[62256] = i[62256];
  assign o[62255] = i[62255];
  assign o[62254] = i[62254];
  assign o[62253] = i[62253];
  assign o[62252] = i[62252];
  assign o[62251] = i[62251];
  assign o[62250] = i[62250];
  assign o[62249] = i[62249];
  assign o[62248] = i[62248];
  assign o[62247] = i[62247];
  assign o[62246] = i[62246];
  assign o[62245] = i[62245];
  assign o[62244] = i[62244];
  assign o[62243] = i[62243];
  assign o[62242] = i[62242];
  assign o[62241] = i[62241];
  assign o[62240] = i[62240];
  assign o[62239] = i[62239];
  assign o[62238] = i[62238];
  assign o[62237] = i[62237];
  assign o[62236] = i[62236];
  assign o[62235] = i[62235];
  assign o[62234] = i[62234];
  assign o[62233] = i[62233];
  assign o[62232] = i[62232];
  assign o[62231] = i[62231];
  assign o[62230] = i[62230];
  assign o[62229] = i[62229];
  assign o[62228] = i[62228];
  assign o[62227] = i[62227];
  assign o[62226] = i[62226];
  assign o[62225] = i[62225];
  assign o[62224] = i[62224];
  assign o[62223] = i[62223];
  assign o[62222] = i[62222];
  assign o[62221] = i[62221];
  assign o[62220] = i[62220];
  assign o[62219] = i[62219];
  assign o[62218] = i[62218];
  assign o[62217] = i[62217];
  assign o[62216] = i[62216];
  assign o[62215] = i[62215];
  assign o[62214] = i[62214];
  assign o[62213] = i[62213];
  assign o[62212] = i[62212];
  assign o[62211] = i[62211];
  assign o[62210] = i[62210];
  assign o[62209] = i[62209];
  assign o[62208] = i[62208];
  assign o[62207] = i[62207];
  assign o[62206] = i[62206];
  assign o[62205] = i[62205];
  assign o[62204] = i[62204];
  assign o[62203] = i[62203];
  assign o[62202] = i[62202];
  assign o[62201] = i[62201];
  assign o[62200] = i[62200];
  assign o[62199] = i[62199];
  assign o[62198] = i[62198];
  assign o[62197] = i[62197];
  assign o[62196] = i[62196];
  assign o[62195] = i[62195];
  assign o[62194] = i[62194];
  assign o[62193] = i[62193];
  assign o[62192] = i[62192];
  assign o[62191] = i[62191];
  assign o[62190] = i[62190];
  assign o[62189] = i[62189];
  assign o[62188] = i[62188];
  assign o[62187] = i[62187];
  assign o[62186] = i[62186];
  assign o[62185] = i[62185];
  assign o[62184] = i[62184];
  assign o[62183] = i[62183];
  assign o[62182] = i[62182];
  assign o[62181] = i[62181];
  assign o[62180] = i[62180];
  assign o[62179] = i[62179];
  assign o[62178] = i[62178];
  assign o[62177] = i[62177];
  assign o[62176] = i[62176];
  assign o[62175] = i[62175];
  assign o[62174] = i[62174];
  assign o[62173] = i[62173];
  assign o[62172] = i[62172];
  assign o[62171] = i[62171];
  assign o[62170] = i[62170];
  assign o[62169] = i[62169];
  assign o[62168] = i[62168];
  assign o[62167] = i[62167];
  assign o[62166] = i[62166];
  assign o[62165] = i[62165];
  assign o[62164] = i[62164];
  assign o[62163] = i[62163];
  assign o[62162] = i[62162];
  assign o[62161] = i[62161];
  assign o[62160] = i[62160];
  assign o[62159] = i[62159];
  assign o[62158] = i[62158];
  assign o[62157] = i[62157];
  assign o[62156] = i[62156];
  assign o[62155] = i[62155];
  assign o[62154] = i[62154];
  assign o[62153] = i[62153];
  assign o[62152] = i[62152];
  assign o[62151] = i[62151];
  assign o[62150] = i[62150];
  assign o[62149] = i[62149];
  assign o[62148] = i[62148];
  assign o[62147] = i[62147];
  assign o[62146] = i[62146];
  assign o[62145] = i[62145];
  assign o[62144] = i[62144];
  assign o[62143] = i[62143];
  assign o[62142] = i[62142];
  assign o[62141] = i[62141];
  assign o[62140] = i[62140];
  assign o[62139] = i[62139];
  assign o[62138] = i[62138];
  assign o[62137] = i[62137];
  assign o[62136] = i[62136];
  assign o[62135] = i[62135];
  assign o[62134] = i[62134];
  assign o[62133] = i[62133];
  assign o[62132] = i[62132];
  assign o[62131] = i[62131];
  assign o[62130] = i[62130];
  assign o[62129] = i[62129];
  assign o[62128] = i[62128];
  assign o[62127] = i[62127];
  assign o[62126] = i[62126];
  assign o[62125] = i[62125];
  assign o[62124] = i[62124];
  assign o[62123] = i[62123];
  assign o[62122] = i[62122];
  assign o[62121] = i[62121];
  assign o[62120] = i[62120];
  assign o[62119] = i[62119];
  assign o[62118] = i[62118];
  assign o[62117] = i[62117];
  assign o[62116] = i[62116];
  assign o[62115] = i[62115];
  assign o[62114] = i[62114];
  assign o[62113] = i[62113];
  assign o[62112] = i[62112];
  assign o[62111] = i[62111];
  assign o[62110] = i[62110];
  assign o[62109] = i[62109];
  assign o[62108] = i[62108];
  assign o[62107] = i[62107];
  assign o[62106] = i[62106];
  assign o[62105] = i[62105];
  assign o[62104] = i[62104];
  assign o[62103] = i[62103];
  assign o[62102] = i[62102];
  assign o[62101] = i[62101];
  assign o[62100] = i[62100];
  assign o[62099] = i[62099];
  assign o[62098] = i[62098];
  assign o[62097] = i[62097];
  assign o[62096] = i[62096];
  assign o[62095] = i[62095];
  assign o[62094] = i[62094];
  assign o[62093] = i[62093];
  assign o[62092] = i[62092];
  assign o[62091] = i[62091];
  assign o[62090] = i[62090];
  assign o[62089] = i[62089];
  assign o[62088] = i[62088];
  assign o[62087] = i[62087];
  assign o[62086] = i[62086];
  assign o[62085] = i[62085];
  assign o[62084] = i[62084];
  assign o[62083] = i[62083];
  assign o[62082] = i[62082];
  assign o[62081] = i[62081];
  assign o[62080] = i[62080];
  assign o[62079] = i[62079];
  assign o[62078] = i[62078];
  assign o[62077] = i[62077];
  assign o[62076] = i[62076];
  assign o[62075] = i[62075];
  assign o[62074] = i[62074];
  assign o[62073] = i[62073];
  assign o[62072] = i[62072];
  assign o[62071] = i[62071];
  assign o[62070] = i[62070];
  assign o[62069] = i[62069];
  assign o[62068] = i[62068];
  assign o[62067] = i[62067];
  assign o[62066] = i[62066];
  assign o[62065] = i[62065];
  assign o[62064] = i[62064];
  assign o[62063] = i[62063];
  assign o[62062] = i[62062];
  assign o[62061] = i[62061];
  assign o[62060] = i[62060];
  assign o[62059] = i[62059];
  assign o[62058] = i[62058];
  assign o[62057] = i[62057];
  assign o[62056] = i[62056];
  assign o[62055] = i[62055];
  assign o[62054] = i[62054];
  assign o[62053] = i[62053];
  assign o[62052] = i[62052];
  assign o[62051] = i[62051];
  assign o[62050] = i[62050];
  assign o[62049] = i[62049];
  assign o[62048] = i[62048];
  assign o[62047] = i[62047];
  assign o[62046] = i[62046];
  assign o[62045] = i[62045];
  assign o[62044] = i[62044];
  assign o[62043] = i[62043];
  assign o[62042] = i[62042];
  assign o[62041] = i[62041];
  assign o[62040] = i[62040];
  assign o[62039] = i[62039];
  assign o[62038] = i[62038];
  assign o[62037] = i[62037];
  assign o[62036] = i[62036];
  assign o[62035] = i[62035];
  assign o[62034] = i[62034];
  assign o[62033] = i[62033];
  assign o[62032] = i[62032];
  assign o[62031] = i[62031];
  assign o[62030] = i[62030];
  assign o[62029] = i[62029];
  assign o[62028] = i[62028];
  assign o[62027] = i[62027];
  assign o[62026] = i[62026];
  assign o[62025] = i[62025];
  assign o[62024] = i[62024];
  assign o[62023] = i[62023];
  assign o[62022] = i[62022];
  assign o[62021] = i[62021];
  assign o[62020] = i[62020];
  assign o[62019] = i[62019];
  assign o[62018] = i[62018];
  assign o[62017] = i[62017];
  assign o[62016] = i[62016];
  assign o[62015] = i[62015];
  assign o[62014] = i[62014];
  assign o[62013] = i[62013];
  assign o[62012] = i[62012];
  assign o[62011] = i[62011];
  assign o[62010] = i[62010];
  assign o[62009] = i[62009];
  assign o[62008] = i[62008];
  assign o[62007] = i[62007];
  assign o[62006] = i[62006];
  assign o[62005] = i[62005];
  assign o[62004] = i[62004];
  assign o[62003] = i[62003];
  assign o[62002] = i[62002];
  assign o[62001] = i[62001];
  assign o[62000] = i[62000];
  assign o[61999] = i[61999];
  assign o[61998] = i[61998];
  assign o[61997] = i[61997];
  assign o[61996] = i[61996];
  assign o[61995] = i[61995];
  assign o[61994] = i[61994];
  assign o[61993] = i[61993];
  assign o[61992] = i[61992];
  assign o[61991] = i[61991];
  assign o[61990] = i[61990];
  assign o[61989] = i[61989];
  assign o[61988] = i[61988];
  assign o[61987] = i[61987];
  assign o[61986] = i[61986];
  assign o[61985] = i[61985];
  assign o[61984] = i[61984];
  assign o[61983] = i[61983];
  assign o[61982] = i[61982];
  assign o[61981] = i[61981];
  assign o[61980] = i[61980];
  assign o[61979] = i[61979];
  assign o[61978] = i[61978];
  assign o[61977] = i[61977];
  assign o[61976] = i[61976];
  assign o[61975] = i[61975];
  assign o[61974] = i[61974];
  assign o[61973] = i[61973];
  assign o[61972] = i[61972];
  assign o[61971] = i[61971];
  assign o[61970] = i[61970];
  assign o[61969] = i[61969];
  assign o[61968] = i[61968];
  assign o[61967] = i[61967];
  assign o[61966] = i[61966];
  assign o[61965] = i[61965];
  assign o[61964] = i[61964];
  assign o[61963] = i[61963];
  assign o[61962] = i[61962];
  assign o[61961] = i[61961];
  assign o[61960] = i[61960];
  assign o[61959] = i[61959];
  assign o[61958] = i[61958];
  assign o[61957] = i[61957];
  assign o[61956] = i[61956];
  assign o[61955] = i[61955];
  assign o[61954] = i[61954];
  assign o[61953] = i[61953];
  assign o[61952] = i[61952];
  assign o[61951] = i[61951];
  assign o[61950] = i[61950];
  assign o[61949] = i[61949];
  assign o[61948] = i[61948];
  assign o[61947] = i[61947];
  assign o[61946] = i[61946];
  assign o[61945] = i[61945];
  assign o[61944] = i[61944];
  assign o[61943] = i[61943];
  assign o[61942] = i[61942];
  assign o[61941] = i[61941];
  assign o[61940] = i[61940];
  assign o[61939] = i[61939];
  assign o[61938] = i[61938];
  assign o[61937] = i[61937];
  assign o[61936] = i[61936];
  assign o[61935] = i[61935];
  assign o[61934] = i[61934];
  assign o[61933] = i[61933];
  assign o[61932] = i[61932];
  assign o[61931] = i[61931];
  assign o[61930] = i[61930];
  assign o[61929] = i[61929];
  assign o[61928] = i[61928];
  assign o[61927] = i[61927];
  assign o[61926] = i[61926];
  assign o[61925] = i[61925];
  assign o[61924] = i[61924];
  assign o[61923] = i[61923];
  assign o[61922] = i[61922];
  assign o[61921] = i[61921];
  assign o[61920] = i[61920];
  assign o[61919] = i[61919];
  assign o[61918] = i[61918];
  assign o[61917] = i[61917];
  assign o[61916] = i[61916];
  assign o[61915] = i[61915];
  assign o[61914] = i[61914];
  assign o[61913] = i[61913];
  assign o[61912] = i[61912];
  assign o[61911] = i[61911];
  assign o[61910] = i[61910];
  assign o[61909] = i[61909];
  assign o[61908] = i[61908];
  assign o[61907] = i[61907];
  assign o[61906] = i[61906];
  assign o[61905] = i[61905];
  assign o[61904] = i[61904];
  assign o[61903] = i[61903];
  assign o[61902] = i[61902];
  assign o[61901] = i[61901];
  assign o[61900] = i[61900];
  assign o[61899] = i[61899];
  assign o[61898] = i[61898];
  assign o[61897] = i[61897];
  assign o[61896] = i[61896];
  assign o[61895] = i[61895];
  assign o[61894] = i[61894];
  assign o[61893] = i[61893];
  assign o[61892] = i[61892];
  assign o[61891] = i[61891];
  assign o[61890] = i[61890];
  assign o[61889] = i[61889];
  assign o[61888] = i[61888];
  assign o[61887] = i[61887];
  assign o[61886] = i[61886];
  assign o[61885] = i[61885];
  assign o[61884] = i[61884];
  assign o[61883] = i[61883];
  assign o[61882] = i[61882];
  assign o[61881] = i[61881];
  assign o[61880] = i[61880];
  assign o[61879] = i[61879];
  assign o[61878] = i[61878];
  assign o[61877] = i[61877];
  assign o[61876] = i[61876];
  assign o[61875] = i[61875];
  assign o[61874] = i[61874];
  assign o[61873] = i[61873];
  assign o[61872] = i[61872];
  assign o[61871] = i[61871];
  assign o[61870] = i[61870];
  assign o[61869] = i[61869];
  assign o[61868] = i[61868];
  assign o[61867] = i[61867];
  assign o[61866] = i[61866];
  assign o[61865] = i[61865];
  assign o[61864] = i[61864];
  assign o[61863] = i[61863];
  assign o[61862] = i[61862];
  assign o[61861] = i[61861];
  assign o[61860] = i[61860];
  assign o[61859] = i[61859];
  assign o[61858] = i[61858];
  assign o[61857] = i[61857];
  assign o[61856] = i[61856];
  assign o[61855] = i[61855];
  assign o[61854] = i[61854];
  assign o[61853] = i[61853];
  assign o[61852] = i[61852];
  assign o[61851] = i[61851];
  assign o[61850] = i[61850];
  assign o[61849] = i[61849];
  assign o[61848] = i[61848];
  assign o[61847] = i[61847];
  assign o[61846] = i[61846];
  assign o[61845] = i[61845];
  assign o[61844] = i[61844];
  assign o[61843] = i[61843];
  assign o[61842] = i[61842];
  assign o[61841] = i[61841];
  assign o[61840] = i[61840];
  assign o[61839] = i[61839];
  assign o[61838] = i[61838];
  assign o[61837] = i[61837];
  assign o[61836] = i[61836];
  assign o[61835] = i[61835];
  assign o[61834] = i[61834];
  assign o[61833] = i[61833];
  assign o[61832] = i[61832];
  assign o[61831] = i[61831];
  assign o[61830] = i[61830];
  assign o[61829] = i[61829];
  assign o[61828] = i[61828];
  assign o[61827] = i[61827];
  assign o[61826] = i[61826];
  assign o[61825] = i[61825];
  assign o[61824] = i[61824];
  assign o[61823] = i[61823];
  assign o[61822] = i[61822];
  assign o[61821] = i[61821];
  assign o[61820] = i[61820];
  assign o[61819] = i[61819];
  assign o[61818] = i[61818];
  assign o[61817] = i[61817];
  assign o[61816] = i[61816];
  assign o[61815] = i[61815];
  assign o[61814] = i[61814];
  assign o[61813] = i[61813];
  assign o[61812] = i[61812];
  assign o[61811] = i[61811];
  assign o[61810] = i[61810];
  assign o[61809] = i[61809];
  assign o[61808] = i[61808];
  assign o[61807] = i[61807];
  assign o[61806] = i[61806];
  assign o[61805] = i[61805];
  assign o[61804] = i[61804];
  assign o[61803] = i[61803];
  assign o[61802] = i[61802];
  assign o[61801] = i[61801];
  assign o[61800] = i[61800];
  assign o[61799] = i[61799];
  assign o[61798] = i[61798];
  assign o[61797] = i[61797];
  assign o[61796] = i[61796];
  assign o[61795] = i[61795];
  assign o[61794] = i[61794];
  assign o[61793] = i[61793];
  assign o[61792] = i[61792];
  assign o[61791] = i[61791];
  assign o[61790] = i[61790];
  assign o[61789] = i[61789];
  assign o[61788] = i[61788];
  assign o[61787] = i[61787];
  assign o[61786] = i[61786];
  assign o[61785] = i[61785];
  assign o[61784] = i[61784];
  assign o[61783] = i[61783];
  assign o[61782] = i[61782];
  assign o[61781] = i[61781];
  assign o[61780] = i[61780];
  assign o[61779] = i[61779];
  assign o[61778] = i[61778];
  assign o[61777] = i[61777];
  assign o[61776] = i[61776];
  assign o[61775] = i[61775];
  assign o[61774] = i[61774];
  assign o[61773] = i[61773];
  assign o[61772] = i[61772];
  assign o[61771] = i[61771];
  assign o[61770] = i[61770];
  assign o[61769] = i[61769];
  assign o[61768] = i[61768];
  assign o[61767] = i[61767];
  assign o[61766] = i[61766];
  assign o[61765] = i[61765];
  assign o[61764] = i[61764];
  assign o[61763] = i[61763];
  assign o[61762] = i[61762];
  assign o[61761] = i[61761];
  assign o[61760] = i[61760];
  assign o[61759] = i[61759];
  assign o[61758] = i[61758];
  assign o[61757] = i[61757];
  assign o[61756] = i[61756];
  assign o[61755] = i[61755];
  assign o[61754] = i[61754];
  assign o[61753] = i[61753];
  assign o[61752] = i[61752];
  assign o[61751] = i[61751];
  assign o[61750] = i[61750];
  assign o[61749] = i[61749];
  assign o[61748] = i[61748];
  assign o[61747] = i[61747];
  assign o[61746] = i[61746];
  assign o[61745] = i[61745];
  assign o[61744] = i[61744];
  assign o[61743] = i[61743];
  assign o[61742] = i[61742];
  assign o[61741] = i[61741];
  assign o[61740] = i[61740];
  assign o[61739] = i[61739];
  assign o[61738] = i[61738];
  assign o[61737] = i[61737];
  assign o[61736] = i[61736];
  assign o[61735] = i[61735];
  assign o[61734] = i[61734];
  assign o[61733] = i[61733];
  assign o[61732] = i[61732];
  assign o[61731] = i[61731];
  assign o[61730] = i[61730];
  assign o[61729] = i[61729];
  assign o[61728] = i[61728];
  assign o[61727] = i[61727];
  assign o[61726] = i[61726];
  assign o[61725] = i[61725];
  assign o[61724] = i[61724];
  assign o[61723] = i[61723];
  assign o[61722] = i[61722];
  assign o[61721] = i[61721];
  assign o[61720] = i[61720];
  assign o[61719] = i[61719];
  assign o[61718] = i[61718];
  assign o[61717] = i[61717];
  assign o[61716] = i[61716];
  assign o[61715] = i[61715];
  assign o[61714] = i[61714];
  assign o[61713] = i[61713];
  assign o[61712] = i[61712];
  assign o[61711] = i[61711];
  assign o[61710] = i[61710];
  assign o[61709] = i[61709];
  assign o[61708] = i[61708];
  assign o[61707] = i[61707];
  assign o[61706] = i[61706];
  assign o[61705] = i[61705];
  assign o[61704] = i[61704];
  assign o[61703] = i[61703];
  assign o[61702] = i[61702];
  assign o[61701] = i[61701];
  assign o[61700] = i[61700];
  assign o[61699] = i[61699];
  assign o[61698] = i[61698];
  assign o[61697] = i[61697];
  assign o[61696] = i[61696];
  assign o[61695] = i[61695];
  assign o[61694] = i[61694];
  assign o[61693] = i[61693];
  assign o[61692] = i[61692];
  assign o[61691] = i[61691];
  assign o[61690] = i[61690];
  assign o[61689] = i[61689];
  assign o[61688] = i[61688];
  assign o[61687] = i[61687];
  assign o[61686] = i[61686];
  assign o[61685] = i[61685];
  assign o[61684] = i[61684];
  assign o[61683] = i[61683];
  assign o[61682] = i[61682];
  assign o[61681] = i[61681];
  assign o[61680] = i[61680];
  assign o[61679] = i[61679];
  assign o[61678] = i[61678];
  assign o[61677] = i[61677];
  assign o[61676] = i[61676];
  assign o[61675] = i[61675];
  assign o[61674] = i[61674];
  assign o[61673] = i[61673];
  assign o[61672] = i[61672];
  assign o[61671] = i[61671];
  assign o[61670] = i[61670];
  assign o[61669] = i[61669];
  assign o[61668] = i[61668];
  assign o[61667] = i[61667];
  assign o[61666] = i[61666];
  assign o[61665] = i[61665];
  assign o[61664] = i[61664];
  assign o[61663] = i[61663];
  assign o[61662] = i[61662];
  assign o[61661] = i[61661];
  assign o[61660] = i[61660];
  assign o[61659] = i[61659];
  assign o[61658] = i[61658];
  assign o[61657] = i[61657];
  assign o[61656] = i[61656];
  assign o[61655] = i[61655];
  assign o[61654] = i[61654];
  assign o[61653] = i[61653];
  assign o[61652] = i[61652];
  assign o[61651] = i[61651];
  assign o[61650] = i[61650];
  assign o[61649] = i[61649];
  assign o[61648] = i[61648];
  assign o[61647] = i[61647];
  assign o[61646] = i[61646];
  assign o[61645] = i[61645];
  assign o[61644] = i[61644];
  assign o[61643] = i[61643];
  assign o[61642] = i[61642];
  assign o[61641] = i[61641];
  assign o[61640] = i[61640];
  assign o[61639] = i[61639];
  assign o[61638] = i[61638];
  assign o[61637] = i[61637];
  assign o[61636] = i[61636];
  assign o[61635] = i[61635];
  assign o[61634] = i[61634];
  assign o[61633] = i[61633];
  assign o[61632] = i[61632];
  assign o[61631] = i[61631];
  assign o[61630] = i[61630];
  assign o[61629] = i[61629];
  assign o[61628] = i[61628];
  assign o[61627] = i[61627];
  assign o[61626] = i[61626];
  assign o[61625] = i[61625];
  assign o[61624] = i[61624];
  assign o[61623] = i[61623];
  assign o[61622] = i[61622];
  assign o[61621] = i[61621];
  assign o[61620] = i[61620];
  assign o[61619] = i[61619];
  assign o[61618] = i[61618];
  assign o[61617] = i[61617];
  assign o[61616] = i[61616];
  assign o[61615] = i[61615];
  assign o[61614] = i[61614];
  assign o[61613] = i[61613];
  assign o[61612] = i[61612];
  assign o[61611] = i[61611];
  assign o[61610] = i[61610];
  assign o[61609] = i[61609];
  assign o[61608] = i[61608];
  assign o[61607] = i[61607];
  assign o[61606] = i[61606];
  assign o[61605] = i[61605];
  assign o[61604] = i[61604];
  assign o[61603] = i[61603];
  assign o[61602] = i[61602];
  assign o[61601] = i[61601];
  assign o[61600] = i[61600];
  assign o[61599] = i[61599];
  assign o[61598] = i[61598];
  assign o[61597] = i[61597];
  assign o[61596] = i[61596];
  assign o[61595] = i[61595];
  assign o[61594] = i[61594];
  assign o[61593] = i[61593];
  assign o[61592] = i[61592];
  assign o[61591] = i[61591];
  assign o[61590] = i[61590];
  assign o[61589] = i[61589];
  assign o[61588] = i[61588];
  assign o[61587] = i[61587];
  assign o[61586] = i[61586];
  assign o[61585] = i[61585];
  assign o[61584] = i[61584];
  assign o[61583] = i[61583];
  assign o[61582] = i[61582];
  assign o[61581] = i[61581];
  assign o[61580] = i[61580];
  assign o[61579] = i[61579];
  assign o[61578] = i[61578];
  assign o[61577] = i[61577];
  assign o[61576] = i[61576];
  assign o[61575] = i[61575];
  assign o[61574] = i[61574];
  assign o[61573] = i[61573];
  assign o[61572] = i[61572];
  assign o[61571] = i[61571];
  assign o[61570] = i[61570];
  assign o[61569] = i[61569];
  assign o[61568] = i[61568];
  assign o[61567] = i[61567];
  assign o[61566] = i[61566];
  assign o[61565] = i[61565];
  assign o[61564] = i[61564];
  assign o[61563] = i[61563];
  assign o[61562] = i[61562];
  assign o[61561] = i[61561];
  assign o[61560] = i[61560];
  assign o[61559] = i[61559];
  assign o[61558] = i[61558];
  assign o[61557] = i[61557];
  assign o[61556] = i[61556];
  assign o[61555] = i[61555];
  assign o[61554] = i[61554];
  assign o[61553] = i[61553];
  assign o[61552] = i[61552];
  assign o[61551] = i[61551];
  assign o[61550] = i[61550];
  assign o[61549] = i[61549];
  assign o[61548] = i[61548];
  assign o[61547] = i[61547];
  assign o[61546] = i[61546];
  assign o[61545] = i[61545];
  assign o[61544] = i[61544];
  assign o[61543] = i[61543];
  assign o[61542] = i[61542];
  assign o[61541] = i[61541];
  assign o[61540] = i[61540];
  assign o[61539] = i[61539];
  assign o[61538] = i[61538];
  assign o[61537] = i[61537];
  assign o[61536] = i[61536];
  assign o[61535] = i[61535];
  assign o[61534] = i[61534];
  assign o[61533] = i[61533];
  assign o[61532] = i[61532];
  assign o[61531] = i[61531];
  assign o[61530] = i[61530];
  assign o[61529] = i[61529];
  assign o[61528] = i[61528];
  assign o[61527] = i[61527];
  assign o[61526] = i[61526];
  assign o[61525] = i[61525];
  assign o[61524] = i[61524];
  assign o[61523] = i[61523];
  assign o[61522] = i[61522];
  assign o[61521] = i[61521];
  assign o[61520] = i[61520];
  assign o[61519] = i[61519];
  assign o[61518] = i[61518];
  assign o[61517] = i[61517];
  assign o[61516] = i[61516];
  assign o[61515] = i[61515];
  assign o[61514] = i[61514];
  assign o[61513] = i[61513];
  assign o[61512] = i[61512];
  assign o[61511] = i[61511];
  assign o[61510] = i[61510];
  assign o[61509] = i[61509];
  assign o[61508] = i[61508];
  assign o[61507] = i[61507];
  assign o[61506] = i[61506];
  assign o[61505] = i[61505];
  assign o[61504] = i[61504];
  assign o[61503] = i[61503];
  assign o[61502] = i[61502];
  assign o[61501] = i[61501];
  assign o[61500] = i[61500];
  assign o[61499] = i[61499];
  assign o[61498] = i[61498];
  assign o[61497] = i[61497];
  assign o[61496] = i[61496];
  assign o[61495] = i[61495];
  assign o[61494] = i[61494];
  assign o[61493] = i[61493];
  assign o[61492] = i[61492];
  assign o[61491] = i[61491];
  assign o[61490] = i[61490];
  assign o[61489] = i[61489];
  assign o[61488] = i[61488];
  assign o[61487] = i[61487];
  assign o[61486] = i[61486];
  assign o[61485] = i[61485];
  assign o[61484] = i[61484];
  assign o[61483] = i[61483];
  assign o[61482] = i[61482];
  assign o[61481] = i[61481];
  assign o[61480] = i[61480];
  assign o[61479] = i[61479];
  assign o[61478] = i[61478];
  assign o[61477] = i[61477];
  assign o[61476] = i[61476];
  assign o[61475] = i[61475];
  assign o[61474] = i[61474];
  assign o[61473] = i[61473];
  assign o[61472] = i[61472];
  assign o[61471] = i[61471];
  assign o[61470] = i[61470];
  assign o[61469] = i[61469];
  assign o[61468] = i[61468];
  assign o[61467] = i[61467];
  assign o[61466] = i[61466];
  assign o[61465] = i[61465];
  assign o[61464] = i[61464];
  assign o[61463] = i[61463];
  assign o[61462] = i[61462];
  assign o[61461] = i[61461];
  assign o[61460] = i[61460];
  assign o[61459] = i[61459];
  assign o[61458] = i[61458];
  assign o[61457] = i[61457];
  assign o[61456] = i[61456];
  assign o[61455] = i[61455];
  assign o[61454] = i[61454];
  assign o[61453] = i[61453];
  assign o[61452] = i[61452];
  assign o[61451] = i[61451];
  assign o[61450] = i[61450];
  assign o[61449] = i[61449];
  assign o[61448] = i[61448];
  assign o[61447] = i[61447];
  assign o[61446] = i[61446];
  assign o[61445] = i[61445];
  assign o[61444] = i[61444];
  assign o[61443] = i[61443];
  assign o[61442] = i[61442];
  assign o[61441] = i[61441];
  assign o[61440] = i[61440];
  assign o[61439] = i[61439];
  assign o[61438] = i[61438];
  assign o[61437] = i[61437];
  assign o[61436] = i[61436];
  assign o[61435] = i[61435];
  assign o[61434] = i[61434];
  assign o[61433] = i[61433];
  assign o[61432] = i[61432];
  assign o[61431] = i[61431];
  assign o[61430] = i[61430];
  assign o[61429] = i[61429];
  assign o[61428] = i[61428];
  assign o[61427] = i[61427];
  assign o[61426] = i[61426];
  assign o[61425] = i[61425];
  assign o[61424] = i[61424];
  assign o[61423] = i[61423];
  assign o[61422] = i[61422];
  assign o[61421] = i[61421];
  assign o[61420] = i[61420];
  assign o[61419] = i[61419];
  assign o[61418] = i[61418];
  assign o[61417] = i[61417];
  assign o[61416] = i[61416];
  assign o[61415] = i[61415];
  assign o[61414] = i[61414];
  assign o[61413] = i[61413];
  assign o[61412] = i[61412];
  assign o[61411] = i[61411];
  assign o[61410] = i[61410];
  assign o[61409] = i[61409];
  assign o[61408] = i[61408];
  assign o[61407] = i[61407];
  assign o[61406] = i[61406];
  assign o[61405] = i[61405];
  assign o[61404] = i[61404];
  assign o[61403] = i[61403];
  assign o[61402] = i[61402];
  assign o[61401] = i[61401];
  assign o[61400] = i[61400];
  assign o[61399] = i[61399];
  assign o[61398] = i[61398];
  assign o[61397] = i[61397];
  assign o[61396] = i[61396];
  assign o[61395] = i[61395];
  assign o[61394] = i[61394];
  assign o[61393] = i[61393];
  assign o[61392] = i[61392];
  assign o[61391] = i[61391];
  assign o[61390] = i[61390];
  assign o[61389] = i[61389];
  assign o[61388] = i[61388];
  assign o[61387] = i[61387];
  assign o[61386] = i[61386];
  assign o[61385] = i[61385];
  assign o[61384] = i[61384];
  assign o[61383] = i[61383];
  assign o[61382] = i[61382];
  assign o[61381] = i[61381];
  assign o[61380] = i[61380];
  assign o[61379] = i[61379];
  assign o[61378] = i[61378];
  assign o[61377] = i[61377];
  assign o[61376] = i[61376];
  assign o[61375] = i[61375];
  assign o[61374] = i[61374];
  assign o[61373] = i[61373];
  assign o[61372] = i[61372];
  assign o[61371] = i[61371];
  assign o[61370] = i[61370];
  assign o[61369] = i[61369];
  assign o[61368] = i[61368];
  assign o[61367] = i[61367];
  assign o[61366] = i[61366];
  assign o[61365] = i[61365];
  assign o[61364] = i[61364];
  assign o[61363] = i[61363];
  assign o[61362] = i[61362];
  assign o[61361] = i[61361];
  assign o[61360] = i[61360];
  assign o[61359] = i[61359];
  assign o[61358] = i[61358];
  assign o[61357] = i[61357];
  assign o[61356] = i[61356];
  assign o[61355] = i[61355];
  assign o[61354] = i[61354];
  assign o[61353] = i[61353];
  assign o[61352] = i[61352];
  assign o[61351] = i[61351];
  assign o[61350] = i[61350];
  assign o[61349] = i[61349];
  assign o[61348] = i[61348];
  assign o[61347] = i[61347];
  assign o[61346] = i[61346];
  assign o[61345] = i[61345];
  assign o[61344] = i[61344];
  assign o[61343] = i[61343];
  assign o[61342] = i[61342];
  assign o[61341] = i[61341];
  assign o[61340] = i[61340];
  assign o[61339] = i[61339];
  assign o[61338] = i[61338];
  assign o[61337] = i[61337];
  assign o[61336] = i[61336];
  assign o[61335] = i[61335];
  assign o[61334] = i[61334];
  assign o[61333] = i[61333];
  assign o[61332] = i[61332];
  assign o[61331] = i[61331];
  assign o[61330] = i[61330];
  assign o[61329] = i[61329];
  assign o[61328] = i[61328];
  assign o[61327] = i[61327];
  assign o[61326] = i[61326];
  assign o[61325] = i[61325];
  assign o[61324] = i[61324];
  assign o[61323] = i[61323];
  assign o[61322] = i[61322];
  assign o[61321] = i[61321];
  assign o[61320] = i[61320];
  assign o[61319] = i[61319];
  assign o[61318] = i[61318];
  assign o[61317] = i[61317];
  assign o[61316] = i[61316];
  assign o[61315] = i[61315];
  assign o[61314] = i[61314];
  assign o[61313] = i[61313];
  assign o[61312] = i[61312];
  assign o[61311] = i[61311];
  assign o[61310] = i[61310];
  assign o[61309] = i[61309];
  assign o[61308] = i[61308];
  assign o[61307] = i[61307];
  assign o[61306] = i[61306];
  assign o[61305] = i[61305];
  assign o[61304] = i[61304];
  assign o[61303] = i[61303];
  assign o[61302] = i[61302];
  assign o[61301] = i[61301];
  assign o[61300] = i[61300];
  assign o[61299] = i[61299];
  assign o[61298] = i[61298];
  assign o[61297] = i[61297];
  assign o[61296] = i[61296];
  assign o[61295] = i[61295];
  assign o[61294] = i[61294];
  assign o[61293] = i[61293];
  assign o[61292] = i[61292];
  assign o[61291] = i[61291];
  assign o[61290] = i[61290];
  assign o[61289] = i[61289];
  assign o[61288] = i[61288];
  assign o[61287] = i[61287];
  assign o[61286] = i[61286];
  assign o[61285] = i[61285];
  assign o[61284] = i[61284];
  assign o[61283] = i[61283];
  assign o[61282] = i[61282];
  assign o[61281] = i[61281];
  assign o[61280] = i[61280];
  assign o[61279] = i[61279];
  assign o[61278] = i[61278];
  assign o[61277] = i[61277];
  assign o[61276] = i[61276];
  assign o[61275] = i[61275];
  assign o[61274] = i[61274];
  assign o[61273] = i[61273];
  assign o[61272] = i[61272];
  assign o[61271] = i[61271];
  assign o[61270] = i[61270];
  assign o[61269] = i[61269];
  assign o[61268] = i[61268];
  assign o[61267] = i[61267];
  assign o[61266] = i[61266];
  assign o[61265] = i[61265];
  assign o[61264] = i[61264];
  assign o[61263] = i[61263];
  assign o[61262] = i[61262];
  assign o[61261] = i[61261];
  assign o[61260] = i[61260];
  assign o[61259] = i[61259];
  assign o[61258] = i[61258];
  assign o[61257] = i[61257];
  assign o[61256] = i[61256];
  assign o[61255] = i[61255];
  assign o[61254] = i[61254];
  assign o[61253] = i[61253];
  assign o[61252] = i[61252];
  assign o[61251] = i[61251];
  assign o[61250] = i[61250];
  assign o[61249] = i[61249];
  assign o[61248] = i[61248];
  assign o[61247] = i[61247];
  assign o[61246] = i[61246];
  assign o[61245] = i[61245];
  assign o[61244] = i[61244];
  assign o[61243] = i[61243];
  assign o[61242] = i[61242];
  assign o[61241] = i[61241];
  assign o[61240] = i[61240];
  assign o[61239] = i[61239];
  assign o[61238] = i[61238];
  assign o[61237] = i[61237];
  assign o[61236] = i[61236];
  assign o[61235] = i[61235];
  assign o[61234] = i[61234];
  assign o[61233] = i[61233];
  assign o[61232] = i[61232];
  assign o[61231] = i[61231];
  assign o[61230] = i[61230];
  assign o[61229] = i[61229];
  assign o[61228] = i[61228];
  assign o[61227] = i[61227];
  assign o[61226] = i[61226];
  assign o[61225] = i[61225];
  assign o[61224] = i[61224];
  assign o[61223] = i[61223];
  assign o[61222] = i[61222];
  assign o[61221] = i[61221];
  assign o[61220] = i[61220];
  assign o[61219] = i[61219];
  assign o[61218] = i[61218];
  assign o[61217] = i[61217];
  assign o[61216] = i[61216];
  assign o[61215] = i[61215];
  assign o[61214] = i[61214];
  assign o[61213] = i[61213];
  assign o[61212] = i[61212];
  assign o[61211] = i[61211];
  assign o[61210] = i[61210];
  assign o[61209] = i[61209];
  assign o[61208] = i[61208];
  assign o[61207] = i[61207];
  assign o[61206] = i[61206];
  assign o[61205] = i[61205];
  assign o[61204] = i[61204];
  assign o[61203] = i[61203];
  assign o[61202] = i[61202];
  assign o[61201] = i[61201];
  assign o[61200] = i[61200];
  assign o[61199] = i[61199];
  assign o[61198] = i[61198];
  assign o[61197] = i[61197];
  assign o[61196] = i[61196];
  assign o[61195] = i[61195];
  assign o[61194] = i[61194];
  assign o[61193] = i[61193];
  assign o[61192] = i[61192];
  assign o[61191] = i[61191];
  assign o[61190] = i[61190];
  assign o[61189] = i[61189];
  assign o[61188] = i[61188];
  assign o[61187] = i[61187];
  assign o[61186] = i[61186];
  assign o[61185] = i[61185];
  assign o[61184] = i[61184];
  assign o[61183] = i[61183];
  assign o[61182] = i[61182];
  assign o[61181] = i[61181];
  assign o[61180] = i[61180];
  assign o[61179] = i[61179];
  assign o[61178] = i[61178];
  assign o[61177] = i[61177];
  assign o[61176] = i[61176];
  assign o[61175] = i[61175];
  assign o[61174] = i[61174];
  assign o[61173] = i[61173];
  assign o[61172] = i[61172];
  assign o[61171] = i[61171];
  assign o[61170] = i[61170];
  assign o[61169] = i[61169];
  assign o[61168] = i[61168];
  assign o[61167] = i[61167];
  assign o[61166] = i[61166];
  assign o[61165] = i[61165];
  assign o[61164] = i[61164];
  assign o[61163] = i[61163];
  assign o[61162] = i[61162];
  assign o[61161] = i[61161];
  assign o[61160] = i[61160];
  assign o[61159] = i[61159];
  assign o[61158] = i[61158];
  assign o[61157] = i[61157];
  assign o[61156] = i[61156];
  assign o[61155] = i[61155];
  assign o[61154] = i[61154];
  assign o[61153] = i[61153];
  assign o[61152] = i[61152];
  assign o[61151] = i[61151];
  assign o[61150] = i[61150];
  assign o[61149] = i[61149];
  assign o[61148] = i[61148];
  assign o[61147] = i[61147];
  assign o[61146] = i[61146];
  assign o[61145] = i[61145];
  assign o[61144] = i[61144];
  assign o[61143] = i[61143];
  assign o[61142] = i[61142];
  assign o[61141] = i[61141];
  assign o[61140] = i[61140];
  assign o[61139] = i[61139];
  assign o[61138] = i[61138];
  assign o[61137] = i[61137];
  assign o[61136] = i[61136];
  assign o[61135] = i[61135];
  assign o[61134] = i[61134];
  assign o[61133] = i[61133];
  assign o[61132] = i[61132];
  assign o[61131] = i[61131];
  assign o[61130] = i[61130];
  assign o[61129] = i[61129];
  assign o[61128] = i[61128];
  assign o[61127] = i[61127];
  assign o[61126] = i[61126];
  assign o[61125] = i[61125];
  assign o[61124] = i[61124];
  assign o[61123] = i[61123];
  assign o[61122] = i[61122];
  assign o[61121] = i[61121];
  assign o[61120] = i[61120];
  assign o[61119] = i[61119];
  assign o[61118] = i[61118];
  assign o[61117] = i[61117];
  assign o[61116] = i[61116];
  assign o[61115] = i[61115];
  assign o[61114] = i[61114];
  assign o[61113] = i[61113];
  assign o[61112] = i[61112];
  assign o[61111] = i[61111];
  assign o[61110] = i[61110];
  assign o[61109] = i[61109];
  assign o[61108] = i[61108];
  assign o[61107] = i[61107];
  assign o[61106] = i[61106];
  assign o[61105] = i[61105];
  assign o[61104] = i[61104];
  assign o[61103] = i[61103];
  assign o[61102] = i[61102];
  assign o[61101] = i[61101];
  assign o[61100] = i[61100];
  assign o[61099] = i[61099];
  assign o[61098] = i[61098];
  assign o[61097] = i[61097];
  assign o[61096] = i[61096];
  assign o[61095] = i[61095];
  assign o[61094] = i[61094];
  assign o[61093] = i[61093];
  assign o[61092] = i[61092];
  assign o[61091] = i[61091];
  assign o[61090] = i[61090];
  assign o[61089] = i[61089];
  assign o[61088] = i[61088];
  assign o[61087] = i[61087];
  assign o[61086] = i[61086];
  assign o[61085] = i[61085];
  assign o[61084] = i[61084];
  assign o[61083] = i[61083];
  assign o[61082] = i[61082];
  assign o[61081] = i[61081];
  assign o[61080] = i[61080];
  assign o[61079] = i[61079];
  assign o[61078] = i[61078];
  assign o[61077] = i[61077];
  assign o[61076] = i[61076];
  assign o[61075] = i[61075];
  assign o[61074] = i[61074];
  assign o[61073] = i[61073];
  assign o[61072] = i[61072];
  assign o[61071] = i[61071];
  assign o[61070] = i[61070];
  assign o[61069] = i[61069];
  assign o[61068] = i[61068];
  assign o[61067] = i[61067];
  assign o[61066] = i[61066];
  assign o[61065] = i[61065];
  assign o[61064] = i[61064];
  assign o[61063] = i[61063];
  assign o[61062] = i[61062];
  assign o[61061] = i[61061];
  assign o[61060] = i[61060];
  assign o[61059] = i[61059];
  assign o[61058] = i[61058];
  assign o[61057] = i[61057];
  assign o[61056] = i[61056];
  assign o[61055] = i[61055];
  assign o[61054] = i[61054];
  assign o[61053] = i[61053];
  assign o[61052] = i[61052];
  assign o[61051] = i[61051];
  assign o[61050] = i[61050];
  assign o[61049] = i[61049];
  assign o[61048] = i[61048];
  assign o[61047] = i[61047];
  assign o[61046] = i[61046];
  assign o[61045] = i[61045];
  assign o[61044] = i[61044];
  assign o[61043] = i[61043];
  assign o[61042] = i[61042];
  assign o[61041] = i[61041];
  assign o[61040] = i[61040];
  assign o[61039] = i[61039];
  assign o[61038] = i[61038];
  assign o[61037] = i[61037];
  assign o[61036] = i[61036];
  assign o[61035] = i[61035];
  assign o[61034] = i[61034];
  assign o[61033] = i[61033];
  assign o[61032] = i[61032];
  assign o[61031] = i[61031];
  assign o[61030] = i[61030];
  assign o[61029] = i[61029];
  assign o[61028] = i[61028];
  assign o[61027] = i[61027];
  assign o[61026] = i[61026];
  assign o[61025] = i[61025];
  assign o[61024] = i[61024];
  assign o[61023] = i[61023];
  assign o[61022] = i[61022];
  assign o[61021] = i[61021];
  assign o[61020] = i[61020];
  assign o[61019] = i[61019];
  assign o[61018] = i[61018];
  assign o[61017] = i[61017];
  assign o[61016] = i[61016];
  assign o[61015] = i[61015];
  assign o[61014] = i[61014];
  assign o[61013] = i[61013];
  assign o[61012] = i[61012];
  assign o[61011] = i[61011];
  assign o[61010] = i[61010];
  assign o[61009] = i[61009];
  assign o[61008] = i[61008];
  assign o[61007] = i[61007];
  assign o[61006] = i[61006];
  assign o[61005] = i[61005];
  assign o[61004] = i[61004];
  assign o[61003] = i[61003];
  assign o[61002] = i[61002];
  assign o[61001] = i[61001];
  assign o[61000] = i[61000];
  assign o[60999] = i[60999];
  assign o[60998] = i[60998];
  assign o[60997] = i[60997];
  assign o[60996] = i[60996];
  assign o[60995] = i[60995];
  assign o[60994] = i[60994];
  assign o[60993] = i[60993];
  assign o[60992] = i[60992];
  assign o[60991] = i[60991];
  assign o[60990] = i[60990];
  assign o[60989] = i[60989];
  assign o[60988] = i[60988];
  assign o[60987] = i[60987];
  assign o[60986] = i[60986];
  assign o[60985] = i[60985];
  assign o[60984] = i[60984];
  assign o[60983] = i[60983];
  assign o[60982] = i[60982];
  assign o[60981] = i[60981];
  assign o[60980] = i[60980];
  assign o[60979] = i[60979];
  assign o[60978] = i[60978];
  assign o[60977] = i[60977];
  assign o[60976] = i[60976];
  assign o[60975] = i[60975];
  assign o[60974] = i[60974];
  assign o[60973] = i[60973];
  assign o[60972] = i[60972];
  assign o[60971] = i[60971];
  assign o[60970] = i[60970];
  assign o[60969] = i[60969];
  assign o[60968] = i[60968];
  assign o[60967] = i[60967];
  assign o[60966] = i[60966];
  assign o[60965] = i[60965];
  assign o[60964] = i[60964];
  assign o[60963] = i[60963];
  assign o[60962] = i[60962];
  assign o[60961] = i[60961];
  assign o[60960] = i[60960];
  assign o[60959] = i[60959];
  assign o[60958] = i[60958];
  assign o[60957] = i[60957];
  assign o[60956] = i[60956];
  assign o[60955] = i[60955];
  assign o[60954] = i[60954];
  assign o[60953] = i[60953];
  assign o[60952] = i[60952];
  assign o[60951] = i[60951];
  assign o[60950] = i[60950];
  assign o[60949] = i[60949];
  assign o[60948] = i[60948];
  assign o[60947] = i[60947];
  assign o[60946] = i[60946];
  assign o[60945] = i[60945];
  assign o[60944] = i[60944];
  assign o[60943] = i[60943];
  assign o[60942] = i[60942];
  assign o[60941] = i[60941];
  assign o[60940] = i[60940];
  assign o[60939] = i[60939];
  assign o[60938] = i[60938];
  assign o[60937] = i[60937];
  assign o[60936] = i[60936];
  assign o[60935] = i[60935];
  assign o[60934] = i[60934];
  assign o[60933] = i[60933];
  assign o[60932] = i[60932];
  assign o[60931] = i[60931];
  assign o[60930] = i[60930];
  assign o[60929] = i[60929];
  assign o[60928] = i[60928];
  assign o[60927] = i[60927];
  assign o[60926] = i[60926];
  assign o[60925] = i[60925];
  assign o[60924] = i[60924];
  assign o[60923] = i[60923];
  assign o[60922] = i[60922];
  assign o[60921] = i[60921];
  assign o[60920] = i[60920];
  assign o[60919] = i[60919];
  assign o[60918] = i[60918];
  assign o[60917] = i[60917];
  assign o[60916] = i[60916];
  assign o[60915] = i[60915];
  assign o[60914] = i[60914];
  assign o[60913] = i[60913];
  assign o[60912] = i[60912];
  assign o[60911] = i[60911];
  assign o[60910] = i[60910];
  assign o[60909] = i[60909];
  assign o[60908] = i[60908];
  assign o[60907] = i[60907];
  assign o[60906] = i[60906];
  assign o[60905] = i[60905];
  assign o[60904] = i[60904];
  assign o[60903] = i[60903];
  assign o[60902] = i[60902];
  assign o[60901] = i[60901];
  assign o[60900] = i[60900];
  assign o[60899] = i[60899];
  assign o[60898] = i[60898];
  assign o[60897] = i[60897];
  assign o[60896] = i[60896];
  assign o[60895] = i[60895];
  assign o[60894] = i[60894];
  assign o[60893] = i[60893];
  assign o[60892] = i[60892];
  assign o[60891] = i[60891];
  assign o[60890] = i[60890];
  assign o[60889] = i[60889];
  assign o[60888] = i[60888];
  assign o[60887] = i[60887];
  assign o[60886] = i[60886];
  assign o[60885] = i[60885];
  assign o[60884] = i[60884];
  assign o[60883] = i[60883];
  assign o[60882] = i[60882];
  assign o[60881] = i[60881];
  assign o[60880] = i[60880];
  assign o[60879] = i[60879];
  assign o[60878] = i[60878];
  assign o[60877] = i[60877];
  assign o[60876] = i[60876];
  assign o[60875] = i[60875];
  assign o[60874] = i[60874];
  assign o[60873] = i[60873];
  assign o[60872] = i[60872];
  assign o[60871] = i[60871];
  assign o[60870] = i[60870];
  assign o[60869] = i[60869];
  assign o[60868] = i[60868];
  assign o[60867] = i[60867];
  assign o[60866] = i[60866];
  assign o[60865] = i[60865];
  assign o[60864] = i[60864];
  assign o[60863] = i[60863];
  assign o[60862] = i[60862];
  assign o[60861] = i[60861];
  assign o[60860] = i[60860];
  assign o[60859] = i[60859];
  assign o[60858] = i[60858];
  assign o[60857] = i[60857];
  assign o[60856] = i[60856];
  assign o[60855] = i[60855];
  assign o[60854] = i[60854];
  assign o[60853] = i[60853];
  assign o[60852] = i[60852];
  assign o[60851] = i[60851];
  assign o[60850] = i[60850];
  assign o[60849] = i[60849];
  assign o[60848] = i[60848];
  assign o[60847] = i[60847];
  assign o[60846] = i[60846];
  assign o[60845] = i[60845];
  assign o[60844] = i[60844];
  assign o[60843] = i[60843];
  assign o[60842] = i[60842];
  assign o[60841] = i[60841];
  assign o[60840] = i[60840];
  assign o[60839] = i[60839];
  assign o[60838] = i[60838];
  assign o[60837] = i[60837];
  assign o[60836] = i[60836];
  assign o[60835] = i[60835];
  assign o[60834] = i[60834];
  assign o[60833] = i[60833];
  assign o[60832] = i[60832];
  assign o[60831] = i[60831];
  assign o[60830] = i[60830];
  assign o[60829] = i[60829];
  assign o[60828] = i[60828];
  assign o[60827] = i[60827];
  assign o[60826] = i[60826];
  assign o[60825] = i[60825];
  assign o[60824] = i[60824];
  assign o[60823] = i[60823];
  assign o[60822] = i[60822];
  assign o[60821] = i[60821];
  assign o[60820] = i[60820];
  assign o[60819] = i[60819];
  assign o[60818] = i[60818];
  assign o[60817] = i[60817];
  assign o[60816] = i[60816];
  assign o[60815] = i[60815];
  assign o[60814] = i[60814];
  assign o[60813] = i[60813];
  assign o[60812] = i[60812];
  assign o[60811] = i[60811];
  assign o[60810] = i[60810];
  assign o[60809] = i[60809];
  assign o[60808] = i[60808];
  assign o[60807] = i[60807];
  assign o[60806] = i[60806];
  assign o[60805] = i[60805];
  assign o[60804] = i[60804];
  assign o[60803] = i[60803];
  assign o[60802] = i[60802];
  assign o[60801] = i[60801];
  assign o[60800] = i[60800];
  assign o[60799] = i[60799];
  assign o[60798] = i[60798];
  assign o[60797] = i[60797];
  assign o[60796] = i[60796];
  assign o[60795] = i[60795];
  assign o[60794] = i[60794];
  assign o[60793] = i[60793];
  assign o[60792] = i[60792];
  assign o[60791] = i[60791];
  assign o[60790] = i[60790];
  assign o[60789] = i[60789];
  assign o[60788] = i[60788];
  assign o[60787] = i[60787];
  assign o[60786] = i[60786];
  assign o[60785] = i[60785];
  assign o[60784] = i[60784];
  assign o[60783] = i[60783];
  assign o[60782] = i[60782];
  assign o[60781] = i[60781];
  assign o[60780] = i[60780];
  assign o[60779] = i[60779];
  assign o[60778] = i[60778];
  assign o[60777] = i[60777];
  assign o[60776] = i[60776];
  assign o[60775] = i[60775];
  assign o[60774] = i[60774];
  assign o[60773] = i[60773];
  assign o[60772] = i[60772];
  assign o[60771] = i[60771];
  assign o[60770] = i[60770];
  assign o[60769] = i[60769];
  assign o[60768] = i[60768];
  assign o[60767] = i[60767];
  assign o[60766] = i[60766];
  assign o[60765] = i[60765];
  assign o[60764] = i[60764];
  assign o[60763] = i[60763];
  assign o[60762] = i[60762];
  assign o[60761] = i[60761];
  assign o[60760] = i[60760];
  assign o[60759] = i[60759];
  assign o[60758] = i[60758];
  assign o[60757] = i[60757];
  assign o[60756] = i[60756];
  assign o[60755] = i[60755];
  assign o[60754] = i[60754];
  assign o[60753] = i[60753];
  assign o[60752] = i[60752];
  assign o[60751] = i[60751];
  assign o[60750] = i[60750];
  assign o[60749] = i[60749];
  assign o[60748] = i[60748];
  assign o[60747] = i[60747];
  assign o[60746] = i[60746];
  assign o[60745] = i[60745];
  assign o[60744] = i[60744];
  assign o[60743] = i[60743];
  assign o[60742] = i[60742];
  assign o[60741] = i[60741];
  assign o[60740] = i[60740];
  assign o[60739] = i[60739];
  assign o[60738] = i[60738];
  assign o[60737] = i[60737];
  assign o[60736] = i[60736];
  assign o[60735] = i[60735];
  assign o[60734] = i[60734];
  assign o[60733] = i[60733];
  assign o[60732] = i[60732];
  assign o[60731] = i[60731];
  assign o[60730] = i[60730];
  assign o[60729] = i[60729];
  assign o[60728] = i[60728];
  assign o[60727] = i[60727];
  assign o[60726] = i[60726];
  assign o[60725] = i[60725];
  assign o[60724] = i[60724];
  assign o[60723] = i[60723];
  assign o[60722] = i[60722];
  assign o[60721] = i[60721];
  assign o[60720] = i[60720];
  assign o[60719] = i[60719];
  assign o[60718] = i[60718];
  assign o[60717] = i[60717];
  assign o[60716] = i[60716];
  assign o[60715] = i[60715];
  assign o[60714] = i[60714];
  assign o[60713] = i[60713];
  assign o[60712] = i[60712];
  assign o[60711] = i[60711];
  assign o[60710] = i[60710];
  assign o[60709] = i[60709];
  assign o[60708] = i[60708];
  assign o[60707] = i[60707];
  assign o[60706] = i[60706];
  assign o[60705] = i[60705];
  assign o[60704] = i[60704];
  assign o[60703] = i[60703];
  assign o[60702] = i[60702];
  assign o[60701] = i[60701];
  assign o[60700] = i[60700];
  assign o[60699] = i[60699];
  assign o[60698] = i[60698];
  assign o[60697] = i[60697];
  assign o[60696] = i[60696];
  assign o[60695] = i[60695];
  assign o[60694] = i[60694];
  assign o[60693] = i[60693];
  assign o[60692] = i[60692];
  assign o[60691] = i[60691];
  assign o[60690] = i[60690];
  assign o[60689] = i[60689];
  assign o[60688] = i[60688];
  assign o[60687] = i[60687];
  assign o[60686] = i[60686];
  assign o[60685] = i[60685];
  assign o[60684] = i[60684];
  assign o[60683] = i[60683];
  assign o[60682] = i[60682];
  assign o[60681] = i[60681];
  assign o[60680] = i[60680];
  assign o[60679] = i[60679];
  assign o[60678] = i[60678];
  assign o[60677] = i[60677];
  assign o[60676] = i[60676];
  assign o[60675] = i[60675];
  assign o[60674] = i[60674];
  assign o[60673] = i[60673];
  assign o[60672] = i[60672];
  assign o[60671] = i[60671];
  assign o[60670] = i[60670];
  assign o[60669] = i[60669];
  assign o[60668] = i[60668];
  assign o[60667] = i[60667];
  assign o[60666] = i[60666];
  assign o[60665] = i[60665];
  assign o[60664] = i[60664];
  assign o[60663] = i[60663];
  assign o[60662] = i[60662];
  assign o[60661] = i[60661];
  assign o[60660] = i[60660];
  assign o[60659] = i[60659];
  assign o[60658] = i[60658];
  assign o[60657] = i[60657];
  assign o[60656] = i[60656];
  assign o[60655] = i[60655];
  assign o[60654] = i[60654];
  assign o[60653] = i[60653];
  assign o[60652] = i[60652];
  assign o[60651] = i[60651];
  assign o[60650] = i[60650];
  assign o[60649] = i[60649];
  assign o[60648] = i[60648];
  assign o[60647] = i[60647];
  assign o[60646] = i[60646];
  assign o[60645] = i[60645];
  assign o[60644] = i[60644];
  assign o[60643] = i[60643];
  assign o[60642] = i[60642];
  assign o[60641] = i[60641];
  assign o[60640] = i[60640];
  assign o[60639] = i[60639];
  assign o[60638] = i[60638];
  assign o[60637] = i[60637];
  assign o[60636] = i[60636];
  assign o[60635] = i[60635];
  assign o[60634] = i[60634];
  assign o[60633] = i[60633];
  assign o[60632] = i[60632];
  assign o[60631] = i[60631];
  assign o[60630] = i[60630];
  assign o[60629] = i[60629];
  assign o[60628] = i[60628];
  assign o[60627] = i[60627];
  assign o[60626] = i[60626];
  assign o[60625] = i[60625];
  assign o[60624] = i[60624];
  assign o[60623] = i[60623];
  assign o[60622] = i[60622];
  assign o[60621] = i[60621];
  assign o[60620] = i[60620];
  assign o[60619] = i[60619];
  assign o[60618] = i[60618];
  assign o[60617] = i[60617];
  assign o[60616] = i[60616];
  assign o[60615] = i[60615];
  assign o[60614] = i[60614];
  assign o[60613] = i[60613];
  assign o[60612] = i[60612];
  assign o[60611] = i[60611];
  assign o[60610] = i[60610];
  assign o[60609] = i[60609];
  assign o[60608] = i[60608];
  assign o[60607] = i[60607];
  assign o[60606] = i[60606];
  assign o[60605] = i[60605];
  assign o[60604] = i[60604];
  assign o[60603] = i[60603];
  assign o[60602] = i[60602];
  assign o[60601] = i[60601];
  assign o[60600] = i[60600];
  assign o[60599] = i[60599];
  assign o[60598] = i[60598];
  assign o[60597] = i[60597];
  assign o[60596] = i[60596];
  assign o[60595] = i[60595];
  assign o[60594] = i[60594];
  assign o[60593] = i[60593];
  assign o[60592] = i[60592];
  assign o[60591] = i[60591];
  assign o[60590] = i[60590];
  assign o[60589] = i[60589];
  assign o[60588] = i[60588];
  assign o[60587] = i[60587];
  assign o[60586] = i[60586];
  assign o[60585] = i[60585];
  assign o[60584] = i[60584];
  assign o[60583] = i[60583];
  assign o[60582] = i[60582];
  assign o[60581] = i[60581];
  assign o[60580] = i[60580];
  assign o[60579] = i[60579];
  assign o[60578] = i[60578];
  assign o[60577] = i[60577];
  assign o[60576] = i[60576];
  assign o[60575] = i[60575];
  assign o[60574] = i[60574];
  assign o[60573] = i[60573];
  assign o[60572] = i[60572];
  assign o[60571] = i[60571];
  assign o[60570] = i[60570];
  assign o[60569] = i[60569];
  assign o[60568] = i[60568];
  assign o[60567] = i[60567];
  assign o[60566] = i[60566];
  assign o[60565] = i[60565];
  assign o[60564] = i[60564];
  assign o[60563] = i[60563];
  assign o[60562] = i[60562];
  assign o[60561] = i[60561];
  assign o[60560] = i[60560];
  assign o[60559] = i[60559];
  assign o[60558] = i[60558];
  assign o[60557] = i[60557];
  assign o[60556] = i[60556];
  assign o[60555] = i[60555];
  assign o[60554] = i[60554];
  assign o[60553] = i[60553];
  assign o[60552] = i[60552];
  assign o[60551] = i[60551];
  assign o[60550] = i[60550];
  assign o[60549] = i[60549];
  assign o[60548] = i[60548];
  assign o[60547] = i[60547];
  assign o[60546] = i[60546];
  assign o[60545] = i[60545];
  assign o[60544] = i[60544];
  assign o[60543] = i[60543];
  assign o[60542] = i[60542];
  assign o[60541] = i[60541];
  assign o[60540] = i[60540];
  assign o[60539] = i[60539];
  assign o[60538] = i[60538];
  assign o[60537] = i[60537];
  assign o[60536] = i[60536];
  assign o[60535] = i[60535];
  assign o[60534] = i[60534];
  assign o[60533] = i[60533];
  assign o[60532] = i[60532];
  assign o[60531] = i[60531];
  assign o[60530] = i[60530];
  assign o[60529] = i[60529];
  assign o[60528] = i[60528];
  assign o[60527] = i[60527];
  assign o[60526] = i[60526];
  assign o[60525] = i[60525];
  assign o[60524] = i[60524];
  assign o[60523] = i[60523];
  assign o[60522] = i[60522];
  assign o[60521] = i[60521];
  assign o[60520] = i[60520];
  assign o[60519] = i[60519];
  assign o[60518] = i[60518];
  assign o[60517] = i[60517];
  assign o[60516] = i[60516];
  assign o[60515] = i[60515];
  assign o[60514] = i[60514];
  assign o[60513] = i[60513];
  assign o[60512] = i[60512];
  assign o[60511] = i[60511];
  assign o[60510] = i[60510];
  assign o[60509] = i[60509];
  assign o[60508] = i[60508];
  assign o[60507] = i[60507];
  assign o[60506] = i[60506];
  assign o[60505] = i[60505];
  assign o[60504] = i[60504];
  assign o[60503] = i[60503];
  assign o[60502] = i[60502];
  assign o[60501] = i[60501];
  assign o[60500] = i[60500];
  assign o[60499] = i[60499];
  assign o[60498] = i[60498];
  assign o[60497] = i[60497];
  assign o[60496] = i[60496];
  assign o[60495] = i[60495];
  assign o[60494] = i[60494];
  assign o[60493] = i[60493];
  assign o[60492] = i[60492];
  assign o[60491] = i[60491];
  assign o[60490] = i[60490];
  assign o[60489] = i[60489];
  assign o[60488] = i[60488];
  assign o[60487] = i[60487];
  assign o[60486] = i[60486];
  assign o[60485] = i[60485];
  assign o[60484] = i[60484];
  assign o[60483] = i[60483];
  assign o[60482] = i[60482];
  assign o[60481] = i[60481];
  assign o[60480] = i[60480];
  assign o[60479] = i[60479];
  assign o[60478] = i[60478];
  assign o[60477] = i[60477];
  assign o[60476] = i[60476];
  assign o[60475] = i[60475];
  assign o[60474] = i[60474];
  assign o[60473] = i[60473];
  assign o[60472] = i[60472];
  assign o[60471] = i[60471];
  assign o[60470] = i[60470];
  assign o[60469] = i[60469];
  assign o[60468] = i[60468];
  assign o[60467] = i[60467];
  assign o[60466] = i[60466];
  assign o[60465] = i[60465];
  assign o[60464] = i[60464];
  assign o[60463] = i[60463];
  assign o[60462] = i[60462];
  assign o[60461] = i[60461];
  assign o[60460] = i[60460];
  assign o[60459] = i[60459];
  assign o[60458] = i[60458];
  assign o[60457] = i[60457];
  assign o[60456] = i[60456];
  assign o[60455] = i[60455];
  assign o[60454] = i[60454];
  assign o[60453] = i[60453];
  assign o[60452] = i[60452];
  assign o[60451] = i[60451];
  assign o[60450] = i[60450];
  assign o[60449] = i[60449];
  assign o[60448] = i[60448];
  assign o[60447] = i[60447];
  assign o[60446] = i[60446];
  assign o[60445] = i[60445];
  assign o[60444] = i[60444];
  assign o[60443] = i[60443];
  assign o[60442] = i[60442];
  assign o[60441] = i[60441];
  assign o[60440] = i[60440];
  assign o[60439] = i[60439];
  assign o[60438] = i[60438];
  assign o[60437] = i[60437];
  assign o[60436] = i[60436];
  assign o[60435] = i[60435];
  assign o[60434] = i[60434];
  assign o[60433] = i[60433];
  assign o[60432] = i[60432];
  assign o[60431] = i[60431];
  assign o[60430] = i[60430];
  assign o[60429] = i[60429];
  assign o[60428] = i[60428];
  assign o[60427] = i[60427];
  assign o[60426] = i[60426];
  assign o[60425] = i[60425];
  assign o[60424] = i[60424];
  assign o[60423] = i[60423];
  assign o[60422] = i[60422];
  assign o[60421] = i[60421];
  assign o[60420] = i[60420];
  assign o[60419] = i[60419];
  assign o[60418] = i[60418];
  assign o[60417] = i[60417];
  assign o[60416] = i[60416];
  assign o[60415] = i[60415];
  assign o[60414] = i[60414];
  assign o[60413] = i[60413];
  assign o[60412] = i[60412];
  assign o[60411] = i[60411];
  assign o[60410] = i[60410];
  assign o[60409] = i[60409];
  assign o[60408] = i[60408];
  assign o[60407] = i[60407];
  assign o[60406] = i[60406];
  assign o[60405] = i[60405];
  assign o[60404] = i[60404];
  assign o[60403] = i[60403];
  assign o[60402] = i[60402];
  assign o[60401] = i[60401];
  assign o[60400] = i[60400];
  assign o[60399] = i[60399];
  assign o[60398] = i[60398];
  assign o[60397] = i[60397];
  assign o[60396] = i[60396];
  assign o[60395] = i[60395];
  assign o[60394] = i[60394];
  assign o[60393] = i[60393];
  assign o[60392] = i[60392];
  assign o[60391] = i[60391];
  assign o[60390] = i[60390];
  assign o[60389] = i[60389];
  assign o[60388] = i[60388];
  assign o[60387] = i[60387];
  assign o[60386] = i[60386];
  assign o[60385] = i[60385];
  assign o[60384] = i[60384];
  assign o[60383] = i[60383];
  assign o[60382] = i[60382];
  assign o[60381] = i[60381];
  assign o[60380] = i[60380];
  assign o[60379] = i[60379];
  assign o[60378] = i[60378];
  assign o[60377] = i[60377];
  assign o[60376] = i[60376];
  assign o[60375] = i[60375];
  assign o[60374] = i[60374];
  assign o[60373] = i[60373];
  assign o[60372] = i[60372];
  assign o[60371] = i[60371];
  assign o[60370] = i[60370];
  assign o[60369] = i[60369];
  assign o[60368] = i[60368];
  assign o[60367] = i[60367];
  assign o[60366] = i[60366];
  assign o[60365] = i[60365];
  assign o[60364] = i[60364];
  assign o[60363] = i[60363];
  assign o[60362] = i[60362];
  assign o[60361] = i[60361];
  assign o[60360] = i[60360];
  assign o[60359] = i[60359];
  assign o[60358] = i[60358];
  assign o[60357] = i[60357];
  assign o[60356] = i[60356];
  assign o[60355] = i[60355];
  assign o[60354] = i[60354];
  assign o[60353] = i[60353];
  assign o[60352] = i[60352];
  assign o[60351] = i[60351];
  assign o[60350] = i[60350];
  assign o[60349] = i[60349];
  assign o[60348] = i[60348];
  assign o[60347] = i[60347];
  assign o[60346] = i[60346];
  assign o[60345] = i[60345];
  assign o[60344] = i[60344];
  assign o[60343] = i[60343];
  assign o[60342] = i[60342];
  assign o[60341] = i[60341];
  assign o[60340] = i[60340];
  assign o[60339] = i[60339];
  assign o[60338] = i[60338];
  assign o[60337] = i[60337];
  assign o[60336] = i[60336];
  assign o[60335] = i[60335];
  assign o[60334] = i[60334];
  assign o[60333] = i[60333];
  assign o[60332] = i[60332];
  assign o[60331] = i[60331];
  assign o[60330] = i[60330];
  assign o[60329] = i[60329];
  assign o[60328] = i[60328];
  assign o[60327] = i[60327];
  assign o[60326] = i[60326];
  assign o[60325] = i[60325];
  assign o[60324] = i[60324];
  assign o[60323] = i[60323];
  assign o[60322] = i[60322];
  assign o[60321] = i[60321];
  assign o[60320] = i[60320];
  assign o[60319] = i[60319];
  assign o[60318] = i[60318];
  assign o[60317] = i[60317];
  assign o[60316] = i[60316];
  assign o[60315] = i[60315];
  assign o[60314] = i[60314];
  assign o[60313] = i[60313];
  assign o[60312] = i[60312];
  assign o[60311] = i[60311];
  assign o[60310] = i[60310];
  assign o[60309] = i[60309];
  assign o[60308] = i[60308];
  assign o[60307] = i[60307];
  assign o[60306] = i[60306];
  assign o[60305] = i[60305];
  assign o[60304] = i[60304];
  assign o[60303] = i[60303];
  assign o[60302] = i[60302];
  assign o[60301] = i[60301];
  assign o[60300] = i[60300];
  assign o[60299] = i[60299];
  assign o[60298] = i[60298];
  assign o[60297] = i[60297];
  assign o[60296] = i[60296];
  assign o[60295] = i[60295];
  assign o[60294] = i[60294];
  assign o[60293] = i[60293];
  assign o[60292] = i[60292];
  assign o[60291] = i[60291];
  assign o[60290] = i[60290];
  assign o[60289] = i[60289];
  assign o[60288] = i[60288];
  assign o[60287] = i[60287];
  assign o[60286] = i[60286];
  assign o[60285] = i[60285];
  assign o[60284] = i[60284];
  assign o[60283] = i[60283];
  assign o[60282] = i[60282];
  assign o[60281] = i[60281];
  assign o[60280] = i[60280];
  assign o[60279] = i[60279];
  assign o[60278] = i[60278];
  assign o[60277] = i[60277];
  assign o[60276] = i[60276];
  assign o[60275] = i[60275];
  assign o[60274] = i[60274];
  assign o[60273] = i[60273];
  assign o[60272] = i[60272];
  assign o[60271] = i[60271];
  assign o[60270] = i[60270];
  assign o[60269] = i[60269];
  assign o[60268] = i[60268];
  assign o[60267] = i[60267];
  assign o[60266] = i[60266];
  assign o[60265] = i[60265];
  assign o[60264] = i[60264];
  assign o[60263] = i[60263];
  assign o[60262] = i[60262];
  assign o[60261] = i[60261];
  assign o[60260] = i[60260];
  assign o[60259] = i[60259];
  assign o[60258] = i[60258];
  assign o[60257] = i[60257];
  assign o[60256] = i[60256];
  assign o[60255] = i[60255];
  assign o[60254] = i[60254];
  assign o[60253] = i[60253];
  assign o[60252] = i[60252];
  assign o[60251] = i[60251];
  assign o[60250] = i[60250];
  assign o[60249] = i[60249];
  assign o[60248] = i[60248];
  assign o[60247] = i[60247];
  assign o[60246] = i[60246];
  assign o[60245] = i[60245];
  assign o[60244] = i[60244];
  assign o[60243] = i[60243];
  assign o[60242] = i[60242];
  assign o[60241] = i[60241];
  assign o[60240] = i[60240];
  assign o[60239] = i[60239];
  assign o[60238] = i[60238];
  assign o[60237] = i[60237];
  assign o[60236] = i[60236];
  assign o[60235] = i[60235];
  assign o[60234] = i[60234];
  assign o[60233] = i[60233];
  assign o[60232] = i[60232];
  assign o[60231] = i[60231];
  assign o[60230] = i[60230];
  assign o[60229] = i[60229];
  assign o[60228] = i[60228];
  assign o[60227] = i[60227];
  assign o[60226] = i[60226];
  assign o[60225] = i[60225];
  assign o[60224] = i[60224];
  assign o[60223] = i[60223];
  assign o[60222] = i[60222];
  assign o[60221] = i[60221];
  assign o[60220] = i[60220];
  assign o[60219] = i[60219];
  assign o[60218] = i[60218];
  assign o[60217] = i[60217];
  assign o[60216] = i[60216];
  assign o[60215] = i[60215];
  assign o[60214] = i[60214];
  assign o[60213] = i[60213];
  assign o[60212] = i[60212];
  assign o[60211] = i[60211];
  assign o[60210] = i[60210];
  assign o[60209] = i[60209];
  assign o[60208] = i[60208];
  assign o[60207] = i[60207];
  assign o[60206] = i[60206];
  assign o[60205] = i[60205];
  assign o[60204] = i[60204];
  assign o[60203] = i[60203];
  assign o[60202] = i[60202];
  assign o[60201] = i[60201];
  assign o[60200] = i[60200];
  assign o[60199] = i[60199];
  assign o[60198] = i[60198];
  assign o[60197] = i[60197];
  assign o[60196] = i[60196];
  assign o[60195] = i[60195];
  assign o[60194] = i[60194];
  assign o[60193] = i[60193];
  assign o[60192] = i[60192];
  assign o[60191] = i[60191];
  assign o[60190] = i[60190];
  assign o[60189] = i[60189];
  assign o[60188] = i[60188];
  assign o[60187] = i[60187];
  assign o[60186] = i[60186];
  assign o[60185] = i[60185];
  assign o[60184] = i[60184];
  assign o[60183] = i[60183];
  assign o[60182] = i[60182];
  assign o[60181] = i[60181];
  assign o[60180] = i[60180];
  assign o[60179] = i[60179];
  assign o[60178] = i[60178];
  assign o[60177] = i[60177];
  assign o[60176] = i[60176];
  assign o[60175] = i[60175];
  assign o[60174] = i[60174];
  assign o[60173] = i[60173];
  assign o[60172] = i[60172];
  assign o[60171] = i[60171];
  assign o[60170] = i[60170];
  assign o[60169] = i[60169];
  assign o[60168] = i[60168];
  assign o[60167] = i[60167];
  assign o[60166] = i[60166];
  assign o[60165] = i[60165];
  assign o[60164] = i[60164];
  assign o[60163] = i[60163];
  assign o[60162] = i[60162];
  assign o[60161] = i[60161];
  assign o[60160] = i[60160];
  assign o[60159] = i[60159];
  assign o[60158] = i[60158];
  assign o[60157] = i[60157];
  assign o[60156] = i[60156];
  assign o[60155] = i[60155];
  assign o[60154] = i[60154];
  assign o[60153] = i[60153];
  assign o[60152] = i[60152];
  assign o[60151] = i[60151];
  assign o[60150] = i[60150];
  assign o[60149] = i[60149];
  assign o[60148] = i[60148];
  assign o[60147] = i[60147];
  assign o[60146] = i[60146];
  assign o[60145] = i[60145];
  assign o[60144] = i[60144];
  assign o[60143] = i[60143];
  assign o[60142] = i[60142];
  assign o[60141] = i[60141];
  assign o[60140] = i[60140];
  assign o[60139] = i[60139];
  assign o[60138] = i[60138];
  assign o[60137] = i[60137];
  assign o[60136] = i[60136];
  assign o[60135] = i[60135];
  assign o[60134] = i[60134];
  assign o[60133] = i[60133];
  assign o[60132] = i[60132];
  assign o[60131] = i[60131];
  assign o[60130] = i[60130];
  assign o[60129] = i[60129];
  assign o[60128] = i[60128];
  assign o[60127] = i[60127];
  assign o[60126] = i[60126];
  assign o[60125] = i[60125];
  assign o[60124] = i[60124];
  assign o[60123] = i[60123];
  assign o[60122] = i[60122];
  assign o[60121] = i[60121];
  assign o[60120] = i[60120];
  assign o[60119] = i[60119];
  assign o[60118] = i[60118];
  assign o[60117] = i[60117];
  assign o[60116] = i[60116];
  assign o[60115] = i[60115];
  assign o[60114] = i[60114];
  assign o[60113] = i[60113];
  assign o[60112] = i[60112];
  assign o[60111] = i[60111];
  assign o[60110] = i[60110];
  assign o[60109] = i[60109];
  assign o[60108] = i[60108];
  assign o[60107] = i[60107];
  assign o[60106] = i[60106];
  assign o[60105] = i[60105];
  assign o[60104] = i[60104];
  assign o[60103] = i[60103];
  assign o[60102] = i[60102];
  assign o[60101] = i[60101];
  assign o[60100] = i[60100];
  assign o[60099] = i[60099];
  assign o[60098] = i[60098];
  assign o[60097] = i[60097];
  assign o[60096] = i[60096];
  assign o[60095] = i[60095];
  assign o[60094] = i[60094];
  assign o[60093] = i[60093];
  assign o[60092] = i[60092];
  assign o[60091] = i[60091];
  assign o[60090] = i[60090];
  assign o[60089] = i[60089];
  assign o[60088] = i[60088];
  assign o[60087] = i[60087];
  assign o[60086] = i[60086];
  assign o[60085] = i[60085];
  assign o[60084] = i[60084];
  assign o[60083] = i[60083];
  assign o[60082] = i[60082];
  assign o[60081] = i[60081];
  assign o[60080] = i[60080];
  assign o[60079] = i[60079];
  assign o[60078] = i[60078];
  assign o[60077] = i[60077];
  assign o[60076] = i[60076];
  assign o[60075] = i[60075];
  assign o[60074] = i[60074];
  assign o[60073] = i[60073];
  assign o[60072] = i[60072];
  assign o[60071] = i[60071];
  assign o[60070] = i[60070];
  assign o[60069] = i[60069];
  assign o[60068] = i[60068];
  assign o[60067] = i[60067];
  assign o[60066] = i[60066];
  assign o[60065] = i[60065];
  assign o[60064] = i[60064];
  assign o[60063] = i[60063];
  assign o[60062] = i[60062];
  assign o[60061] = i[60061];
  assign o[60060] = i[60060];
  assign o[60059] = i[60059];
  assign o[60058] = i[60058];
  assign o[60057] = i[60057];
  assign o[60056] = i[60056];
  assign o[60055] = i[60055];
  assign o[60054] = i[60054];
  assign o[60053] = i[60053];
  assign o[60052] = i[60052];
  assign o[60051] = i[60051];
  assign o[60050] = i[60050];
  assign o[60049] = i[60049];
  assign o[60048] = i[60048];
  assign o[60047] = i[60047];
  assign o[60046] = i[60046];
  assign o[60045] = i[60045];
  assign o[60044] = i[60044];
  assign o[60043] = i[60043];
  assign o[60042] = i[60042];
  assign o[60041] = i[60041];
  assign o[60040] = i[60040];
  assign o[60039] = i[60039];
  assign o[60038] = i[60038];
  assign o[60037] = i[60037];
  assign o[60036] = i[60036];
  assign o[60035] = i[60035];
  assign o[60034] = i[60034];
  assign o[60033] = i[60033];
  assign o[60032] = i[60032];
  assign o[60031] = i[60031];
  assign o[60030] = i[60030];
  assign o[60029] = i[60029];
  assign o[60028] = i[60028];
  assign o[60027] = i[60027];
  assign o[60026] = i[60026];
  assign o[60025] = i[60025];
  assign o[60024] = i[60024];
  assign o[60023] = i[60023];
  assign o[60022] = i[60022];
  assign o[60021] = i[60021];
  assign o[60020] = i[60020];
  assign o[60019] = i[60019];
  assign o[60018] = i[60018];
  assign o[60017] = i[60017];
  assign o[60016] = i[60016];
  assign o[60015] = i[60015];
  assign o[60014] = i[60014];
  assign o[60013] = i[60013];
  assign o[60012] = i[60012];
  assign o[60011] = i[60011];
  assign o[60010] = i[60010];
  assign o[60009] = i[60009];
  assign o[60008] = i[60008];
  assign o[60007] = i[60007];
  assign o[60006] = i[60006];
  assign o[60005] = i[60005];
  assign o[60004] = i[60004];
  assign o[60003] = i[60003];
  assign o[60002] = i[60002];
  assign o[60001] = i[60001];
  assign o[60000] = i[60000];
  assign o[59999] = i[59999];
  assign o[59998] = i[59998];
  assign o[59997] = i[59997];
  assign o[59996] = i[59996];
  assign o[59995] = i[59995];
  assign o[59994] = i[59994];
  assign o[59993] = i[59993];
  assign o[59992] = i[59992];
  assign o[59991] = i[59991];
  assign o[59990] = i[59990];
  assign o[59989] = i[59989];
  assign o[59988] = i[59988];
  assign o[59987] = i[59987];
  assign o[59986] = i[59986];
  assign o[59985] = i[59985];
  assign o[59984] = i[59984];
  assign o[59983] = i[59983];
  assign o[59982] = i[59982];
  assign o[59981] = i[59981];
  assign o[59980] = i[59980];
  assign o[59979] = i[59979];
  assign o[59978] = i[59978];
  assign o[59977] = i[59977];
  assign o[59976] = i[59976];
  assign o[59975] = i[59975];
  assign o[59974] = i[59974];
  assign o[59973] = i[59973];
  assign o[59972] = i[59972];
  assign o[59971] = i[59971];
  assign o[59970] = i[59970];
  assign o[59969] = i[59969];
  assign o[59968] = i[59968];
  assign o[59967] = i[59967];
  assign o[59966] = i[59966];
  assign o[59965] = i[59965];
  assign o[59964] = i[59964];
  assign o[59963] = i[59963];
  assign o[59962] = i[59962];
  assign o[59961] = i[59961];
  assign o[59960] = i[59960];
  assign o[59959] = i[59959];
  assign o[59958] = i[59958];
  assign o[59957] = i[59957];
  assign o[59956] = i[59956];
  assign o[59955] = i[59955];
  assign o[59954] = i[59954];
  assign o[59953] = i[59953];
  assign o[59952] = i[59952];
  assign o[59951] = i[59951];
  assign o[59950] = i[59950];
  assign o[59949] = i[59949];
  assign o[59948] = i[59948];
  assign o[59947] = i[59947];
  assign o[59946] = i[59946];
  assign o[59945] = i[59945];
  assign o[59944] = i[59944];
  assign o[59943] = i[59943];
  assign o[59942] = i[59942];
  assign o[59941] = i[59941];
  assign o[59940] = i[59940];
  assign o[59939] = i[59939];
  assign o[59938] = i[59938];
  assign o[59937] = i[59937];
  assign o[59936] = i[59936];
  assign o[59935] = i[59935];
  assign o[59934] = i[59934];
  assign o[59933] = i[59933];
  assign o[59932] = i[59932];
  assign o[59931] = i[59931];
  assign o[59930] = i[59930];
  assign o[59929] = i[59929];
  assign o[59928] = i[59928];
  assign o[59927] = i[59927];
  assign o[59926] = i[59926];
  assign o[59925] = i[59925];
  assign o[59924] = i[59924];
  assign o[59923] = i[59923];
  assign o[59922] = i[59922];
  assign o[59921] = i[59921];
  assign o[59920] = i[59920];
  assign o[59919] = i[59919];
  assign o[59918] = i[59918];
  assign o[59917] = i[59917];
  assign o[59916] = i[59916];
  assign o[59915] = i[59915];
  assign o[59914] = i[59914];
  assign o[59913] = i[59913];
  assign o[59912] = i[59912];
  assign o[59911] = i[59911];
  assign o[59910] = i[59910];
  assign o[59909] = i[59909];
  assign o[59908] = i[59908];
  assign o[59907] = i[59907];
  assign o[59906] = i[59906];
  assign o[59905] = i[59905];
  assign o[59904] = i[59904];
  assign o[59903] = i[59903];
  assign o[59902] = i[59902];
  assign o[59901] = i[59901];
  assign o[59900] = i[59900];
  assign o[59899] = i[59899];
  assign o[59898] = i[59898];
  assign o[59897] = i[59897];
  assign o[59896] = i[59896];
  assign o[59895] = i[59895];
  assign o[59894] = i[59894];
  assign o[59893] = i[59893];
  assign o[59892] = i[59892];
  assign o[59891] = i[59891];
  assign o[59890] = i[59890];
  assign o[59889] = i[59889];
  assign o[59888] = i[59888];
  assign o[59887] = i[59887];
  assign o[59886] = i[59886];
  assign o[59885] = i[59885];
  assign o[59884] = i[59884];
  assign o[59883] = i[59883];
  assign o[59882] = i[59882];
  assign o[59881] = i[59881];
  assign o[59880] = i[59880];
  assign o[59879] = i[59879];
  assign o[59878] = i[59878];
  assign o[59877] = i[59877];
  assign o[59876] = i[59876];
  assign o[59875] = i[59875];
  assign o[59874] = i[59874];
  assign o[59873] = i[59873];
  assign o[59872] = i[59872];
  assign o[59871] = i[59871];
  assign o[59870] = i[59870];
  assign o[59869] = i[59869];
  assign o[59868] = i[59868];
  assign o[59867] = i[59867];
  assign o[59866] = i[59866];
  assign o[59865] = i[59865];
  assign o[59864] = i[59864];
  assign o[59863] = i[59863];
  assign o[59862] = i[59862];
  assign o[59861] = i[59861];
  assign o[59860] = i[59860];
  assign o[59859] = i[59859];
  assign o[59858] = i[59858];
  assign o[59857] = i[59857];
  assign o[59856] = i[59856];
  assign o[59855] = i[59855];
  assign o[59854] = i[59854];
  assign o[59853] = i[59853];
  assign o[59852] = i[59852];
  assign o[59851] = i[59851];
  assign o[59850] = i[59850];
  assign o[59849] = i[59849];
  assign o[59848] = i[59848];
  assign o[59847] = i[59847];
  assign o[59846] = i[59846];
  assign o[59845] = i[59845];
  assign o[59844] = i[59844];
  assign o[59843] = i[59843];
  assign o[59842] = i[59842];
  assign o[59841] = i[59841];
  assign o[59840] = i[59840];
  assign o[59839] = i[59839];
  assign o[59838] = i[59838];
  assign o[59837] = i[59837];
  assign o[59836] = i[59836];
  assign o[59835] = i[59835];
  assign o[59834] = i[59834];
  assign o[59833] = i[59833];
  assign o[59832] = i[59832];
  assign o[59831] = i[59831];
  assign o[59830] = i[59830];
  assign o[59829] = i[59829];
  assign o[59828] = i[59828];
  assign o[59827] = i[59827];
  assign o[59826] = i[59826];
  assign o[59825] = i[59825];
  assign o[59824] = i[59824];
  assign o[59823] = i[59823];
  assign o[59822] = i[59822];
  assign o[59821] = i[59821];
  assign o[59820] = i[59820];
  assign o[59819] = i[59819];
  assign o[59818] = i[59818];
  assign o[59817] = i[59817];
  assign o[59816] = i[59816];
  assign o[59815] = i[59815];
  assign o[59814] = i[59814];
  assign o[59813] = i[59813];
  assign o[59812] = i[59812];
  assign o[59811] = i[59811];
  assign o[59810] = i[59810];
  assign o[59809] = i[59809];
  assign o[59808] = i[59808];
  assign o[59807] = i[59807];
  assign o[59806] = i[59806];
  assign o[59805] = i[59805];
  assign o[59804] = i[59804];
  assign o[59803] = i[59803];
  assign o[59802] = i[59802];
  assign o[59801] = i[59801];
  assign o[59800] = i[59800];
  assign o[59799] = i[59799];
  assign o[59798] = i[59798];
  assign o[59797] = i[59797];
  assign o[59796] = i[59796];
  assign o[59795] = i[59795];
  assign o[59794] = i[59794];
  assign o[59793] = i[59793];
  assign o[59792] = i[59792];
  assign o[59791] = i[59791];
  assign o[59790] = i[59790];
  assign o[59789] = i[59789];
  assign o[59788] = i[59788];
  assign o[59787] = i[59787];
  assign o[59786] = i[59786];
  assign o[59785] = i[59785];
  assign o[59784] = i[59784];
  assign o[59783] = i[59783];
  assign o[59782] = i[59782];
  assign o[59781] = i[59781];
  assign o[59780] = i[59780];
  assign o[59779] = i[59779];
  assign o[59778] = i[59778];
  assign o[59777] = i[59777];
  assign o[59776] = i[59776];
  assign o[59775] = i[59775];
  assign o[59774] = i[59774];
  assign o[59773] = i[59773];
  assign o[59772] = i[59772];
  assign o[59771] = i[59771];
  assign o[59770] = i[59770];
  assign o[59769] = i[59769];
  assign o[59768] = i[59768];
  assign o[59767] = i[59767];
  assign o[59766] = i[59766];
  assign o[59765] = i[59765];
  assign o[59764] = i[59764];
  assign o[59763] = i[59763];
  assign o[59762] = i[59762];
  assign o[59761] = i[59761];
  assign o[59760] = i[59760];
  assign o[59759] = i[59759];
  assign o[59758] = i[59758];
  assign o[59757] = i[59757];
  assign o[59756] = i[59756];
  assign o[59755] = i[59755];
  assign o[59754] = i[59754];
  assign o[59753] = i[59753];
  assign o[59752] = i[59752];
  assign o[59751] = i[59751];
  assign o[59750] = i[59750];
  assign o[59749] = i[59749];
  assign o[59748] = i[59748];
  assign o[59747] = i[59747];
  assign o[59746] = i[59746];
  assign o[59745] = i[59745];
  assign o[59744] = i[59744];
  assign o[59743] = i[59743];
  assign o[59742] = i[59742];
  assign o[59741] = i[59741];
  assign o[59740] = i[59740];
  assign o[59739] = i[59739];
  assign o[59738] = i[59738];
  assign o[59737] = i[59737];
  assign o[59736] = i[59736];
  assign o[59735] = i[59735];
  assign o[59734] = i[59734];
  assign o[59733] = i[59733];
  assign o[59732] = i[59732];
  assign o[59731] = i[59731];
  assign o[59730] = i[59730];
  assign o[59729] = i[59729];
  assign o[59728] = i[59728];
  assign o[59727] = i[59727];
  assign o[59726] = i[59726];
  assign o[59725] = i[59725];
  assign o[59724] = i[59724];
  assign o[59723] = i[59723];
  assign o[59722] = i[59722];
  assign o[59721] = i[59721];
  assign o[59720] = i[59720];
  assign o[59719] = i[59719];
  assign o[59718] = i[59718];
  assign o[59717] = i[59717];
  assign o[59716] = i[59716];
  assign o[59715] = i[59715];
  assign o[59714] = i[59714];
  assign o[59713] = i[59713];
  assign o[59712] = i[59712];
  assign o[59711] = i[59711];
  assign o[59710] = i[59710];
  assign o[59709] = i[59709];
  assign o[59708] = i[59708];
  assign o[59707] = i[59707];
  assign o[59706] = i[59706];
  assign o[59705] = i[59705];
  assign o[59704] = i[59704];
  assign o[59703] = i[59703];
  assign o[59702] = i[59702];
  assign o[59701] = i[59701];
  assign o[59700] = i[59700];
  assign o[59699] = i[59699];
  assign o[59698] = i[59698];
  assign o[59697] = i[59697];
  assign o[59696] = i[59696];
  assign o[59695] = i[59695];
  assign o[59694] = i[59694];
  assign o[59693] = i[59693];
  assign o[59692] = i[59692];
  assign o[59691] = i[59691];
  assign o[59690] = i[59690];
  assign o[59689] = i[59689];
  assign o[59688] = i[59688];
  assign o[59687] = i[59687];
  assign o[59686] = i[59686];
  assign o[59685] = i[59685];
  assign o[59684] = i[59684];
  assign o[59683] = i[59683];
  assign o[59682] = i[59682];
  assign o[59681] = i[59681];
  assign o[59680] = i[59680];
  assign o[59679] = i[59679];
  assign o[59678] = i[59678];
  assign o[59677] = i[59677];
  assign o[59676] = i[59676];
  assign o[59675] = i[59675];
  assign o[59674] = i[59674];
  assign o[59673] = i[59673];
  assign o[59672] = i[59672];
  assign o[59671] = i[59671];
  assign o[59670] = i[59670];
  assign o[59669] = i[59669];
  assign o[59668] = i[59668];
  assign o[59667] = i[59667];
  assign o[59666] = i[59666];
  assign o[59665] = i[59665];
  assign o[59664] = i[59664];
  assign o[59663] = i[59663];
  assign o[59662] = i[59662];
  assign o[59661] = i[59661];
  assign o[59660] = i[59660];
  assign o[59659] = i[59659];
  assign o[59658] = i[59658];
  assign o[59657] = i[59657];
  assign o[59656] = i[59656];
  assign o[59655] = i[59655];
  assign o[59654] = i[59654];
  assign o[59653] = i[59653];
  assign o[59652] = i[59652];
  assign o[59651] = i[59651];
  assign o[59650] = i[59650];
  assign o[59649] = i[59649];
  assign o[59648] = i[59648];
  assign o[59647] = i[59647];
  assign o[59646] = i[59646];
  assign o[59645] = i[59645];
  assign o[59644] = i[59644];
  assign o[59643] = i[59643];
  assign o[59642] = i[59642];
  assign o[59641] = i[59641];
  assign o[59640] = i[59640];
  assign o[59639] = i[59639];
  assign o[59638] = i[59638];
  assign o[59637] = i[59637];
  assign o[59636] = i[59636];
  assign o[59635] = i[59635];
  assign o[59634] = i[59634];
  assign o[59633] = i[59633];
  assign o[59632] = i[59632];
  assign o[59631] = i[59631];
  assign o[59630] = i[59630];
  assign o[59629] = i[59629];
  assign o[59628] = i[59628];
  assign o[59627] = i[59627];
  assign o[59626] = i[59626];
  assign o[59625] = i[59625];
  assign o[59624] = i[59624];
  assign o[59623] = i[59623];
  assign o[59622] = i[59622];
  assign o[59621] = i[59621];
  assign o[59620] = i[59620];
  assign o[59619] = i[59619];
  assign o[59618] = i[59618];
  assign o[59617] = i[59617];
  assign o[59616] = i[59616];
  assign o[59615] = i[59615];
  assign o[59614] = i[59614];
  assign o[59613] = i[59613];
  assign o[59612] = i[59612];
  assign o[59611] = i[59611];
  assign o[59610] = i[59610];
  assign o[59609] = i[59609];
  assign o[59608] = i[59608];
  assign o[59607] = i[59607];
  assign o[59606] = i[59606];
  assign o[59605] = i[59605];
  assign o[59604] = i[59604];
  assign o[59603] = i[59603];
  assign o[59602] = i[59602];
  assign o[59601] = i[59601];
  assign o[59600] = i[59600];
  assign o[59599] = i[59599];
  assign o[59598] = i[59598];
  assign o[59597] = i[59597];
  assign o[59596] = i[59596];
  assign o[59595] = i[59595];
  assign o[59594] = i[59594];
  assign o[59593] = i[59593];
  assign o[59592] = i[59592];
  assign o[59591] = i[59591];
  assign o[59590] = i[59590];
  assign o[59589] = i[59589];
  assign o[59588] = i[59588];
  assign o[59587] = i[59587];
  assign o[59586] = i[59586];
  assign o[59585] = i[59585];
  assign o[59584] = i[59584];
  assign o[59583] = i[59583];
  assign o[59582] = i[59582];
  assign o[59581] = i[59581];
  assign o[59580] = i[59580];
  assign o[59579] = i[59579];
  assign o[59578] = i[59578];
  assign o[59577] = i[59577];
  assign o[59576] = i[59576];
  assign o[59575] = i[59575];
  assign o[59574] = i[59574];
  assign o[59573] = i[59573];
  assign o[59572] = i[59572];
  assign o[59571] = i[59571];
  assign o[59570] = i[59570];
  assign o[59569] = i[59569];
  assign o[59568] = i[59568];
  assign o[59567] = i[59567];
  assign o[59566] = i[59566];
  assign o[59565] = i[59565];
  assign o[59564] = i[59564];
  assign o[59563] = i[59563];
  assign o[59562] = i[59562];
  assign o[59561] = i[59561];
  assign o[59560] = i[59560];
  assign o[59559] = i[59559];
  assign o[59558] = i[59558];
  assign o[59557] = i[59557];
  assign o[59556] = i[59556];
  assign o[59555] = i[59555];
  assign o[59554] = i[59554];
  assign o[59553] = i[59553];
  assign o[59552] = i[59552];
  assign o[59551] = i[59551];
  assign o[59550] = i[59550];
  assign o[59549] = i[59549];
  assign o[59548] = i[59548];
  assign o[59547] = i[59547];
  assign o[59546] = i[59546];
  assign o[59545] = i[59545];
  assign o[59544] = i[59544];
  assign o[59543] = i[59543];
  assign o[59542] = i[59542];
  assign o[59541] = i[59541];
  assign o[59540] = i[59540];
  assign o[59539] = i[59539];
  assign o[59538] = i[59538];
  assign o[59537] = i[59537];
  assign o[59536] = i[59536];
  assign o[59535] = i[59535];
  assign o[59534] = i[59534];
  assign o[59533] = i[59533];
  assign o[59532] = i[59532];
  assign o[59531] = i[59531];
  assign o[59530] = i[59530];
  assign o[59529] = i[59529];
  assign o[59528] = i[59528];
  assign o[59527] = i[59527];
  assign o[59526] = i[59526];
  assign o[59525] = i[59525];
  assign o[59524] = i[59524];
  assign o[59523] = i[59523];
  assign o[59522] = i[59522];
  assign o[59521] = i[59521];
  assign o[59520] = i[59520];
  assign o[59519] = i[59519];
  assign o[59518] = i[59518];
  assign o[59517] = i[59517];
  assign o[59516] = i[59516];
  assign o[59515] = i[59515];
  assign o[59514] = i[59514];
  assign o[59513] = i[59513];
  assign o[59512] = i[59512];
  assign o[59511] = i[59511];
  assign o[59510] = i[59510];
  assign o[59509] = i[59509];
  assign o[59508] = i[59508];
  assign o[59507] = i[59507];
  assign o[59506] = i[59506];
  assign o[59505] = i[59505];
  assign o[59504] = i[59504];
  assign o[59503] = i[59503];
  assign o[59502] = i[59502];
  assign o[59501] = i[59501];
  assign o[59500] = i[59500];
  assign o[59499] = i[59499];
  assign o[59498] = i[59498];
  assign o[59497] = i[59497];
  assign o[59496] = i[59496];
  assign o[59495] = i[59495];
  assign o[59494] = i[59494];
  assign o[59493] = i[59493];
  assign o[59492] = i[59492];
  assign o[59491] = i[59491];
  assign o[59490] = i[59490];
  assign o[59489] = i[59489];
  assign o[59488] = i[59488];
  assign o[59487] = i[59487];
  assign o[59486] = i[59486];
  assign o[59485] = i[59485];
  assign o[59484] = i[59484];
  assign o[59483] = i[59483];
  assign o[59482] = i[59482];
  assign o[59481] = i[59481];
  assign o[59480] = i[59480];
  assign o[59479] = i[59479];
  assign o[59478] = i[59478];
  assign o[59477] = i[59477];
  assign o[59476] = i[59476];
  assign o[59475] = i[59475];
  assign o[59474] = i[59474];
  assign o[59473] = i[59473];
  assign o[59472] = i[59472];
  assign o[59471] = i[59471];
  assign o[59470] = i[59470];
  assign o[59469] = i[59469];
  assign o[59468] = i[59468];
  assign o[59467] = i[59467];
  assign o[59466] = i[59466];
  assign o[59465] = i[59465];
  assign o[59464] = i[59464];
  assign o[59463] = i[59463];
  assign o[59462] = i[59462];
  assign o[59461] = i[59461];
  assign o[59460] = i[59460];
  assign o[59459] = i[59459];
  assign o[59458] = i[59458];
  assign o[59457] = i[59457];
  assign o[59456] = i[59456];
  assign o[59455] = i[59455];
  assign o[59454] = i[59454];
  assign o[59453] = i[59453];
  assign o[59452] = i[59452];
  assign o[59451] = i[59451];
  assign o[59450] = i[59450];
  assign o[59449] = i[59449];
  assign o[59448] = i[59448];
  assign o[59447] = i[59447];
  assign o[59446] = i[59446];
  assign o[59445] = i[59445];
  assign o[59444] = i[59444];
  assign o[59443] = i[59443];
  assign o[59442] = i[59442];
  assign o[59441] = i[59441];
  assign o[59440] = i[59440];
  assign o[59439] = i[59439];
  assign o[59438] = i[59438];
  assign o[59437] = i[59437];
  assign o[59436] = i[59436];
  assign o[59435] = i[59435];
  assign o[59434] = i[59434];
  assign o[59433] = i[59433];
  assign o[59432] = i[59432];
  assign o[59431] = i[59431];
  assign o[59430] = i[59430];
  assign o[59429] = i[59429];
  assign o[59428] = i[59428];
  assign o[59427] = i[59427];
  assign o[59426] = i[59426];
  assign o[59425] = i[59425];
  assign o[59424] = i[59424];
  assign o[59423] = i[59423];
  assign o[59422] = i[59422];
  assign o[59421] = i[59421];
  assign o[59420] = i[59420];
  assign o[59419] = i[59419];
  assign o[59418] = i[59418];
  assign o[59417] = i[59417];
  assign o[59416] = i[59416];
  assign o[59415] = i[59415];
  assign o[59414] = i[59414];
  assign o[59413] = i[59413];
  assign o[59412] = i[59412];
  assign o[59411] = i[59411];
  assign o[59410] = i[59410];
  assign o[59409] = i[59409];
  assign o[59408] = i[59408];
  assign o[59407] = i[59407];
  assign o[59406] = i[59406];
  assign o[59405] = i[59405];
  assign o[59404] = i[59404];
  assign o[59403] = i[59403];
  assign o[59402] = i[59402];
  assign o[59401] = i[59401];
  assign o[59400] = i[59400];
  assign o[59399] = i[59399];
  assign o[59398] = i[59398];
  assign o[59397] = i[59397];
  assign o[59396] = i[59396];
  assign o[59395] = i[59395];
  assign o[59394] = i[59394];
  assign o[59393] = i[59393];
  assign o[59392] = i[59392];
  assign o[59391] = i[59391];
  assign o[59390] = i[59390];
  assign o[59389] = i[59389];
  assign o[59388] = i[59388];
  assign o[59387] = i[59387];
  assign o[59386] = i[59386];
  assign o[59385] = i[59385];
  assign o[59384] = i[59384];
  assign o[59383] = i[59383];
  assign o[59382] = i[59382];
  assign o[59381] = i[59381];
  assign o[59380] = i[59380];
  assign o[59379] = i[59379];
  assign o[59378] = i[59378];
  assign o[59377] = i[59377];
  assign o[59376] = i[59376];
  assign o[59375] = i[59375];
  assign o[59374] = i[59374];
  assign o[59373] = i[59373];
  assign o[59372] = i[59372];
  assign o[59371] = i[59371];
  assign o[59370] = i[59370];
  assign o[59369] = i[59369];
  assign o[59368] = i[59368];
  assign o[59367] = i[59367];
  assign o[59366] = i[59366];
  assign o[59365] = i[59365];
  assign o[59364] = i[59364];
  assign o[59363] = i[59363];
  assign o[59362] = i[59362];
  assign o[59361] = i[59361];
  assign o[59360] = i[59360];
  assign o[59359] = i[59359];
  assign o[59358] = i[59358];
  assign o[59357] = i[59357];
  assign o[59356] = i[59356];
  assign o[59355] = i[59355];
  assign o[59354] = i[59354];
  assign o[59353] = i[59353];
  assign o[59352] = i[59352];
  assign o[59351] = i[59351];
  assign o[59350] = i[59350];
  assign o[59349] = i[59349];
  assign o[59348] = i[59348];
  assign o[59347] = i[59347];
  assign o[59346] = i[59346];
  assign o[59345] = i[59345];
  assign o[59344] = i[59344];
  assign o[59343] = i[59343];
  assign o[59342] = i[59342];
  assign o[59341] = i[59341];
  assign o[59340] = i[59340];
  assign o[59339] = i[59339];
  assign o[59338] = i[59338];
  assign o[59337] = i[59337];
  assign o[59336] = i[59336];
  assign o[59335] = i[59335];
  assign o[59334] = i[59334];
  assign o[59333] = i[59333];
  assign o[59332] = i[59332];
  assign o[59331] = i[59331];
  assign o[59330] = i[59330];
  assign o[59329] = i[59329];
  assign o[59328] = i[59328];
  assign o[59327] = i[59327];
  assign o[59326] = i[59326];
  assign o[59325] = i[59325];
  assign o[59324] = i[59324];
  assign o[59323] = i[59323];
  assign o[59322] = i[59322];
  assign o[59321] = i[59321];
  assign o[59320] = i[59320];
  assign o[59319] = i[59319];
  assign o[59318] = i[59318];
  assign o[59317] = i[59317];
  assign o[59316] = i[59316];
  assign o[59315] = i[59315];
  assign o[59314] = i[59314];
  assign o[59313] = i[59313];
  assign o[59312] = i[59312];
  assign o[59311] = i[59311];
  assign o[59310] = i[59310];
  assign o[59309] = i[59309];
  assign o[59308] = i[59308];
  assign o[59307] = i[59307];
  assign o[59306] = i[59306];
  assign o[59305] = i[59305];
  assign o[59304] = i[59304];
  assign o[59303] = i[59303];
  assign o[59302] = i[59302];
  assign o[59301] = i[59301];
  assign o[59300] = i[59300];
  assign o[59299] = i[59299];
  assign o[59298] = i[59298];
  assign o[59297] = i[59297];
  assign o[59296] = i[59296];
  assign o[59295] = i[59295];
  assign o[59294] = i[59294];
  assign o[59293] = i[59293];
  assign o[59292] = i[59292];
  assign o[59291] = i[59291];
  assign o[59290] = i[59290];
  assign o[59289] = i[59289];
  assign o[59288] = i[59288];
  assign o[59287] = i[59287];
  assign o[59286] = i[59286];
  assign o[59285] = i[59285];
  assign o[59284] = i[59284];
  assign o[59283] = i[59283];
  assign o[59282] = i[59282];
  assign o[59281] = i[59281];
  assign o[59280] = i[59280];
  assign o[59279] = i[59279];
  assign o[59278] = i[59278];
  assign o[59277] = i[59277];
  assign o[59276] = i[59276];
  assign o[59275] = i[59275];
  assign o[59274] = i[59274];
  assign o[59273] = i[59273];
  assign o[59272] = i[59272];
  assign o[59271] = i[59271];
  assign o[59270] = i[59270];
  assign o[59269] = i[59269];
  assign o[59268] = i[59268];
  assign o[59267] = i[59267];
  assign o[59266] = i[59266];
  assign o[59265] = i[59265];
  assign o[59264] = i[59264];
  assign o[59263] = i[59263];
  assign o[59262] = i[59262];
  assign o[59261] = i[59261];
  assign o[59260] = i[59260];
  assign o[59259] = i[59259];
  assign o[59258] = i[59258];
  assign o[59257] = i[59257];
  assign o[59256] = i[59256];
  assign o[59255] = i[59255];
  assign o[59254] = i[59254];
  assign o[59253] = i[59253];
  assign o[59252] = i[59252];
  assign o[59251] = i[59251];
  assign o[59250] = i[59250];
  assign o[59249] = i[59249];
  assign o[59248] = i[59248];
  assign o[59247] = i[59247];
  assign o[59246] = i[59246];
  assign o[59245] = i[59245];
  assign o[59244] = i[59244];
  assign o[59243] = i[59243];
  assign o[59242] = i[59242];
  assign o[59241] = i[59241];
  assign o[59240] = i[59240];
  assign o[59239] = i[59239];
  assign o[59238] = i[59238];
  assign o[59237] = i[59237];
  assign o[59236] = i[59236];
  assign o[59235] = i[59235];
  assign o[59234] = i[59234];
  assign o[59233] = i[59233];
  assign o[59232] = i[59232];
  assign o[59231] = i[59231];
  assign o[59230] = i[59230];
  assign o[59229] = i[59229];
  assign o[59228] = i[59228];
  assign o[59227] = i[59227];
  assign o[59226] = i[59226];
  assign o[59225] = i[59225];
  assign o[59224] = i[59224];
  assign o[59223] = i[59223];
  assign o[59222] = i[59222];
  assign o[59221] = i[59221];
  assign o[59220] = i[59220];
  assign o[59219] = i[59219];
  assign o[59218] = i[59218];
  assign o[59217] = i[59217];
  assign o[59216] = i[59216];
  assign o[59215] = i[59215];
  assign o[59214] = i[59214];
  assign o[59213] = i[59213];
  assign o[59212] = i[59212];
  assign o[59211] = i[59211];
  assign o[59210] = i[59210];
  assign o[59209] = i[59209];
  assign o[59208] = i[59208];
  assign o[59207] = i[59207];
  assign o[59206] = i[59206];
  assign o[59205] = i[59205];
  assign o[59204] = i[59204];
  assign o[59203] = i[59203];
  assign o[59202] = i[59202];
  assign o[59201] = i[59201];
  assign o[59200] = i[59200];
  assign o[59199] = i[59199];
  assign o[59198] = i[59198];
  assign o[59197] = i[59197];
  assign o[59196] = i[59196];
  assign o[59195] = i[59195];
  assign o[59194] = i[59194];
  assign o[59193] = i[59193];
  assign o[59192] = i[59192];
  assign o[59191] = i[59191];
  assign o[59190] = i[59190];
  assign o[59189] = i[59189];
  assign o[59188] = i[59188];
  assign o[59187] = i[59187];
  assign o[59186] = i[59186];
  assign o[59185] = i[59185];
  assign o[59184] = i[59184];
  assign o[59183] = i[59183];
  assign o[59182] = i[59182];
  assign o[59181] = i[59181];
  assign o[59180] = i[59180];
  assign o[59179] = i[59179];
  assign o[59178] = i[59178];
  assign o[59177] = i[59177];
  assign o[59176] = i[59176];
  assign o[59175] = i[59175];
  assign o[59174] = i[59174];
  assign o[59173] = i[59173];
  assign o[59172] = i[59172];
  assign o[59171] = i[59171];
  assign o[59170] = i[59170];
  assign o[59169] = i[59169];
  assign o[59168] = i[59168];
  assign o[59167] = i[59167];
  assign o[59166] = i[59166];
  assign o[59165] = i[59165];
  assign o[59164] = i[59164];
  assign o[59163] = i[59163];
  assign o[59162] = i[59162];
  assign o[59161] = i[59161];
  assign o[59160] = i[59160];
  assign o[59159] = i[59159];
  assign o[59158] = i[59158];
  assign o[59157] = i[59157];
  assign o[59156] = i[59156];
  assign o[59155] = i[59155];
  assign o[59154] = i[59154];
  assign o[59153] = i[59153];
  assign o[59152] = i[59152];
  assign o[59151] = i[59151];
  assign o[59150] = i[59150];
  assign o[59149] = i[59149];
  assign o[59148] = i[59148];
  assign o[59147] = i[59147];
  assign o[59146] = i[59146];
  assign o[59145] = i[59145];
  assign o[59144] = i[59144];
  assign o[59143] = i[59143];
  assign o[59142] = i[59142];
  assign o[59141] = i[59141];
  assign o[59140] = i[59140];
  assign o[59139] = i[59139];
  assign o[59138] = i[59138];
  assign o[59137] = i[59137];
  assign o[59136] = i[59136];
  assign o[59135] = i[59135];
  assign o[59134] = i[59134];
  assign o[59133] = i[59133];
  assign o[59132] = i[59132];
  assign o[59131] = i[59131];
  assign o[59130] = i[59130];
  assign o[59129] = i[59129];
  assign o[59128] = i[59128];
  assign o[59127] = i[59127];
  assign o[59126] = i[59126];
  assign o[59125] = i[59125];
  assign o[59124] = i[59124];
  assign o[59123] = i[59123];
  assign o[59122] = i[59122];
  assign o[59121] = i[59121];
  assign o[59120] = i[59120];
  assign o[59119] = i[59119];
  assign o[59118] = i[59118];
  assign o[59117] = i[59117];
  assign o[59116] = i[59116];
  assign o[59115] = i[59115];
  assign o[59114] = i[59114];
  assign o[59113] = i[59113];
  assign o[59112] = i[59112];
  assign o[59111] = i[59111];
  assign o[59110] = i[59110];
  assign o[59109] = i[59109];
  assign o[59108] = i[59108];
  assign o[59107] = i[59107];
  assign o[59106] = i[59106];
  assign o[59105] = i[59105];
  assign o[59104] = i[59104];
  assign o[59103] = i[59103];
  assign o[59102] = i[59102];
  assign o[59101] = i[59101];
  assign o[59100] = i[59100];
  assign o[59099] = i[59099];
  assign o[59098] = i[59098];
  assign o[59097] = i[59097];
  assign o[59096] = i[59096];
  assign o[59095] = i[59095];
  assign o[59094] = i[59094];
  assign o[59093] = i[59093];
  assign o[59092] = i[59092];
  assign o[59091] = i[59091];
  assign o[59090] = i[59090];
  assign o[59089] = i[59089];
  assign o[59088] = i[59088];
  assign o[59087] = i[59087];
  assign o[59086] = i[59086];
  assign o[59085] = i[59085];
  assign o[59084] = i[59084];
  assign o[59083] = i[59083];
  assign o[59082] = i[59082];
  assign o[59081] = i[59081];
  assign o[59080] = i[59080];
  assign o[59079] = i[59079];
  assign o[59078] = i[59078];
  assign o[59077] = i[59077];
  assign o[59076] = i[59076];
  assign o[59075] = i[59075];
  assign o[59074] = i[59074];
  assign o[59073] = i[59073];
  assign o[59072] = i[59072];
  assign o[59071] = i[59071];
  assign o[59070] = i[59070];
  assign o[59069] = i[59069];
  assign o[59068] = i[59068];
  assign o[59067] = i[59067];
  assign o[59066] = i[59066];
  assign o[59065] = i[59065];
  assign o[59064] = i[59064];
  assign o[59063] = i[59063];
  assign o[59062] = i[59062];
  assign o[59061] = i[59061];
  assign o[59060] = i[59060];
  assign o[59059] = i[59059];
  assign o[59058] = i[59058];
  assign o[59057] = i[59057];
  assign o[59056] = i[59056];
  assign o[59055] = i[59055];
  assign o[59054] = i[59054];
  assign o[59053] = i[59053];
  assign o[59052] = i[59052];
  assign o[59051] = i[59051];
  assign o[59050] = i[59050];
  assign o[59049] = i[59049];
  assign o[59048] = i[59048];
  assign o[59047] = i[59047];
  assign o[59046] = i[59046];
  assign o[59045] = i[59045];
  assign o[59044] = i[59044];
  assign o[59043] = i[59043];
  assign o[59042] = i[59042];
  assign o[59041] = i[59041];
  assign o[59040] = i[59040];
  assign o[59039] = i[59039];
  assign o[59038] = i[59038];
  assign o[59037] = i[59037];
  assign o[59036] = i[59036];
  assign o[59035] = i[59035];
  assign o[59034] = i[59034];
  assign o[59033] = i[59033];
  assign o[59032] = i[59032];
  assign o[59031] = i[59031];
  assign o[59030] = i[59030];
  assign o[59029] = i[59029];
  assign o[59028] = i[59028];
  assign o[59027] = i[59027];
  assign o[59026] = i[59026];
  assign o[59025] = i[59025];
  assign o[59024] = i[59024];
  assign o[59023] = i[59023];
  assign o[59022] = i[59022];
  assign o[59021] = i[59021];
  assign o[59020] = i[59020];
  assign o[59019] = i[59019];
  assign o[59018] = i[59018];
  assign o[59017] = i[59017];
  assign o[59016] = i[59016];
  assign o[59015] = i[59015];
  assign o[59014] = i[59014];
  assign o[59013] = i[59013];
  assign o[59012] = i[59012];
  assign o[59011] = i[59011];
  assign o[59010] = i[59010];
  assign o[59009] = i[59009];
  assign o[59008] = i[59008];
  assign o[59007] = i[59007];
  assign o[59006] = i[59006];
  assign o[59005] = i[59005];
  assign o[59004] = i[59004];
  assign o[59003] = i[59003];
  assign o[59002] = i[59002];
  assign o[59001] = i[59001];
  assign o[59000] = i[59000];
  assign o[58999] = i[58999];
  assign o[58998] = i[58998];
  assign o[58997] = i[58997];
  assign o[58996] = i[58996];
  assign o[58995] = i[58995];
  assign o[58994] = i[58994];
  assign o[58993] = i[58993];
  assign o[58992] = i[58992];
  assign o[58991] = i[58991];
  assign o[58990] = i[58990];
  assign o[58989] = i[58989];
  assign o[58988] = i[58988];
  assign o[58987] = i[58987];
  assign o[58986] = i[58986];
  assign o[58985] = i[58985];
  assign o[58984] = i[58984];
  assign o[58983] = i[58983];
  assign o[58982] = i[58982];
  assign o[58981] = i[58981];
  assign o[58980] = i[58980];
  assign o[58979] = i[58979];
  assign o[58978] = i[58978];
  assign o[58977] = i[58977];
  assign o[58976] = i[58976];
  assign o[58975] = i[58975];
  assign o[58974] = i[58974];
  assign o[58973] = i[58973];
  assign o[58972] = i[58972];
  assign o[58971] = i[58971];
  assign o[58970] = i[58970];
  assign o[58969] = i[58969];
  assign o[58968] = i[58968];
  assign o[58967] = i[58967];
  assign o[58966] = i[58966];
  assign o[58965] = i[58965];
  assign o[58964] = i[58964];
  assign o[58963] = i[58963];
  assign o[58962] = i[58962];
  assign o[58961] = i[58961];
  assign o[58960] = i[58960];
  assign o[58959] = i[58959];
  assign o[58958] = i[58958];
  assign o[58957] = i[58957];
  assign o[58956] = i[58956];
  assign o[58955] = i[58955];
  assign o[58954] = i[58954];
  assign o[58953] = i[58953];
  assign o[58952] = i[58952];
  assign o[58951] = i[58951];
  assign o[58950] = i[58950];
  assign o[58949] = i[58949];
  assign o[58948] = i[58948];
  assign o[58947] = i[58947];
  assign o[58946] = i[58946];
  assign o[58945] = i[58945];
  assign o[58944] = i[58944];
  assign o[58943] = i[58943];
  assign o[58942] = i[58942];
  assign o[58941] = i[58941];
  assign o[58940] = i[58940];
  assign o[58939] = i[58939];
  assign o[58938] = i[58938];
  assign o[58937] = i[58937];
  assign o[58936] = i[58936];
  assign o[58935] = i[58935];
  assign o[58934] = i[58934];
  assign o[58933] = i[58933];
  assign o[58932] = i[58932];
  assign o[58931] = i[58931];
  assign o[58930] = i[58930];
  assign o[58929] = i[58929];
  assign o[58928] = i[58928];
  assign o[58927] = i[58927];
  assign o[58926] = i[58926];
  assign o[58925] = i[58925];
  assign o[58924] = i[58924];
  assign o[58923] = i[58923];
  assign o[58922] = i[58922];
  assign o[58921] = i[58921];
  assign o[58920] = i[58920];
  assign o[58919] = i[58919];
  assign o[58918] = i[58918];
  assign o[58917] = i[58917];
  assign o[58916] = i[58916];
  assign o[58915] = i[58915];
  assign o[58914] = i[58914];
  assign o[58913] = i[58913];
  assign o[58912] = i[58912];
  assign o[58911] = i[58911];
  assign o[58910] = i[58910];
  assign o[58909] = i[58909];
  assign o[58908] = i[58908];
  assign o[58907] = i[58907];
  assign o[58906] = i[58906];
  assign o[58905] = i[58905];
  assign o[58904] = i[58904];
  assign o[58903] = i[58903];
  assign o[58902] = i[58902];
  assign o[58901] = i[58901];
  assign o[58900] = i[58900];
  assign o[58899] = i[58899];
  assign o[58898] = i[58898];
  assign o[58897] = i[58897];
  assign o[58896] = i[58896];
  assign o[58895] = i[58895];
  assign o[58894] = i[58894];
  assign o[58893] = i[58893];
  assign o[58892] = i[58892];
  assign o[58891] = i[58891];
  assign o[58890] = i[58890];
  assign o[58889] = i[58889];
  assign o[58888] = i[58888];
  assign o[58887] = i[58887];
  assign o[58886] = i[58886];
  assign o[58885] = i[58885];
  assign o[58884] = i[58884];
  assign o[58883] = i[58883];
  assign o[58882] = i[58882];
  assign o[58881] = i[58881];
  assign o[58880] = i[58880];
  assign o[58879] = i[58879];
  assign o[58878] = i[58878];
  assign o[58877] = i[58877];
  assign o[58876] = i[58876];
  assign o[58875] = i[58875];
  assign o[58874] = i[58874];
  assign o[58873] = i[58873];
  assign o[58872] = i[58872];
  assign o[58871] = i[58871];
  assign o[58870] = i[58870];
  assign o[58869] = i[58869];
  assign o[58868] = i[58868];
  assign o[58867] = i[58867];
  assign o[58866] = i[58866];
  assign o[58865] = i[58865];
  assign o[58864] = i[58864];
  assign o[58863] = i[58863];
  assign o[58862] = i[58862];
  assign o[58861] = i[58861];
  assign o[58860] = i[58860];
  assign o[58859] = i[58859];
  assign o[58858] = i[58858];
  assign o[58857] = i[58857];
  assign o[58856] = i[58856];
  assign o[58855] = i[58855];
  assign o[58854] = i[58854];
  assign o[58853] = i[58853];
  assign o[58852] = i[58852];
  assign o[58851] = i[58851];
  assign o[58850] = i[58850];
  assign o[58849] = i[58849];
  assign o[58848] = i[58848];
  assign o[58847] = i[58847];
  assign o[58846] = i[58846];
  assign o[58845] = i[58845];
  assign o[58844] = i[58844];
  assign o[58843] = i[58843];
  assign o[58842] = i[58842];
  assign o[58841] = i[58841];
  assign o[58840] = i[58840];
  assign o[58839] = i[58839];
  assign o[58838] = i[58838];
  assign o[58837] = i[58837];
  assign o[58836] = i[58836];
  assign o[58835] = i[58835];
  assign o[58834] = i[58834];
  assign o[58833] = i[58833];
  assign o[58832] = i[58832];
  assign o[58831] = i[58831];
  assign o[58830] = i[58830];
  assign o[58829] = i[58829];
  assign o[58828] = i[58828];
  assign o[58827] = i[58827];
  assign o[58826] = i[58826];
  assign o[58825] = i[58825];
  assign o[58824] = i[58824];
  assign o[58823] = i[58823];
  assign o[58822] = i[58822];
  assign o[58821] = i[58821];
  assign o[58820] = i[58820];
  assign o[58819] = i[58819];
  assign o[58818] = i[58818];
  assign o[58817] = i[58817];
  assign o[58816] = i[58816];
  assign o[58815] = i[58815];
  assign o[58814] = i[58814];
  assign o[58813] = i[58813];
  assign o[58812] = i[58812];
  assign o[58811] = i[58811];
  assign o[58810] = i[58810];
  assign o[58809] = i[58809];
  assign o[58808] = i[58808];
  assign o[58807] = i[58807];
  assign o[58806] = i[58806];
  assign o[58805] = i[58805];
  assign o[58804] = i[58804];
  assign o[58803] = i[58803];
  assign o[58802] = i[58802];
  assign o[58801] = i[58801];
  assign o[58800] = i[58800];
  assign o[58799] = i[58799];
  assign o[58798] = i[58798];
  assign o[58797] = i[58797];
  assign o[58796] = i[58796];
  assign o[58795] = i[58795];
  assign o[58794] = i[58794];
  assign o[58793] = i[58793];
  assign o[58792] = i[58792];
  assign o[58791] = i[58791];
  assign o[58790] = i[58790];
  assign o[58789] = i[58789];
  assign o[58788] = i[58788];
  assign o[58787] = i[58787];
  assign o[58786] = i[58786];
  assign o[58785] = i[58785];
  assign o[58784] = i[58784];
  assign o[58783] = i[58783];
  assign o[58782] = i[58782];
  assign o[58781] = i[58781];
  assign o[58780] = i[58780];
  assign o[58779] = i[58779];
  assign o[58778] = i[58778];
  assign o[58777] = i[58777];
  assign o[58776] = i[58776];
  assign o[58775] = i[58775];
  assign o[58774] = i[58774];
  assign o[58773] = i[58773];
  assign o[58772] = i[58772];
  assign o[58771] = i[58771];
  assign o[58770] = i[58770];
  assign o[58769] = i[58769];
  assign o[58768] = i[58768];
  assign o[58767] = i[58767];
  assign o[58766] = i[58766];
  assign o[58765] = i[58765];
  assign o[58764] = i[58764];
  assign o[58763] = i[58763];
  assign o[58762] = i[58762];
  assign o[58761] = i[58761];
  assign o[58760] = i[58760];
  assign o[58759] = i[58759];
  assign o[58758] = i[58758];
  assign o[58757] = i[58757];
  assign o[58756] = i[58756];
  assign o[58755] = i[58755];
  assign o[58754] = i[58754];
  assign o[58753] = i[58753];
  assign o[58752] = i[58752];
  assign o[58751] = i[58751];
  assign o[58750] = i[58750];
  assign o[58749] = i[58749];
  assign o[58748] = i[58748];
  assign o[58747] = i[58747];
  assign o[58746] = i[58746];
  assign o[58745] = i[58745];
  assign o[58744] = i[58744];
  assign o[58743] = i[58743];
  assign o[58742] = i[58742];
  assign o[58741] = i[58741];
  assign o[58740] = i[58740];
  assign o[58739] = i[58739];
  assign o[58738] = i[58738];
  assign o[58737] = i[58737];
  assign o[58736] = i[58736];
  assign o[58735] = i[58735];
  assign o[58734] = i[58734];
  assign o[58733] = i[58733];
  assign o[58732] = i[58732];
  assign o[58731] = i[58731];
  assign o[58730] = i[58730];
  assign o[58729] = i[58729];
  assign o[58728] = i[58728];
  assign o[58727] = i[58727];
  assign o[58726] = i[58726];
  assign o[58725] = i[58725];
  assign o[58724] = i[58724];
  assign o[58723] = i[58723];
  assign o[58722] = i[58722];
  assign o[58721] = i[58721];
  assign o[58720] = i[58720];
  assign o[58719] = i[58719];
  assign o[58718] = i[58718];
  assign o[58717] = i[58717];
  assign o[58716] = i[58716];
  assign o[58715] = i[58715];
  assign o[58714] = i[58714];
  assign o[58713] = i[58713];
  assign o[58712] = i[58712];
  assign o[58711] = i[58711];
  assign o[58710] = i[58710];
  assign o[58709] = i[58709];
  assign o[58708] = i[58708];
  assign o[58707] = i[58707];
  assign o[58706] = i[58706];
  assign o[58705] = i[58705];
  assign o[58704] = i[58704];
  assign o[58703] = i[58703];
  assign o[58702] = i[58702];
  assign o[58701] = i[58701];
  assign o[58700] = i[58700];
  assign o[58699] = i[58699];
  assign o[58698] = i[58698];
  assign o[58697] = i[58697];
  assign o[58696] = i[58696];
  assign o[58695] = i[58695];
  assign o[58694] = i[58694];
  assign o[58693] = i[58693];
  assign o[58692] = i[58692];
  assign o[58691] = i[58691];
  assign o[58690] = i[58690];
  assign o[58689] = i[58689];
  assign o[58688] = i[58688];
  assign o[58687] = i[58687];
  assign o[58686] = i[58686];
  assign o[58685] = i[58685];
  assign o[58684] = i[58684];
  assign o[58683] = i[58683];
  assign o[58682] = i[58682];
  assign o[58681] = i[58681];
  assign o[58680] = i[58680];
  assign o[58679] = i[58679];
  assign o[58678] = i[58678];
  assign o[58677] = i[58677];
  assign o[58676] = i[58676];
  assign o[58675] = i[58675];
  assign o[58674] = i[58674];
  assign o[58673] = i[58673];
  assign o[58672] = i[58672];
  assign o[58671] = i[58671];
  assign o[58670] = i[58670];
  assign o[58669] = i[58669];
  assign o[58668] = i[58668];
  assign o[58667] = i[58667];
  assign o[58666] = i[58666];
  assign o[58665] = i[58665];
  assign o[58664] = i[58664];
  assign o[58663] = i[58663];
  assign o[58662] = i[58662];
  assign o[58661] = i[58661];
  assign o[58660] = i[58660];
  assign o[58659] = i[58659];
  assign o[58658] = i[58658];
  assign o[58657] = i[58657];
  assign o[58656] = i[58656];
  assign o[58655] = i[58655];
  assign o[58654] = i[58654];
  assign o[58653] = i[58653];
  assign o[58652] = i[58652];
  assign o[58651] = i[58651];
  assign o[58650] = i[58650];
  assign o[58649] = i[58649];
  assign o[58648] = i[58648];
  assign o[58647] = i[58647];
  assign o[58646] = i[58646];
  assign o[58645] = i[58645];
  assign o[58644] = i[58644];
  assign o[58643] = i[58643];
  assign o[58642] = i[58642];
  assign o[58641] = i[58641];
  assign o[58640] = i[58640];
  assign o[58639] = i[58639];
  assign o[58638] = i[58638];
  assign o[58637] = i[58637];
  assign o[58636] = i[58636];
  assign o[58635] = i[58635];
  assign o[58634] = i[58634];
  assign o[58633] = i[58633];
  assign o[58632] = i[58632];
  assign o[58631] = i[58631];
  assign o[58630] = i[58630];
  assign o[58629] = i[58629];
  assign o[58628] = i[58628];
  assign o[58627] = i[58627];
  assign o[58626] = i[58626];
  assign o[58625] = i[58625];
  assign o[58624] = i[58624];
  assign o[58623] = i[58623];
  assign o[58622] = i[58622];
  assign o[58621] = i[58621];
  assign o[58620] = i[58620];
  assign o[58619] = i[58619];
  assign o[58618] = i[58618];
  assign o[58617] = i[58617];
  assign o[58616] = i[58616];
  assign o[58615] = i[58615];
  assign o[58614] = i[58614];
  assign o[58613] = i[58613];
  assign o[58612] = i[58612];
  assign o[58611] = i[58611];
  assign o[58610] = i[58610];
  assign o[58609] = i[58609];
  assign o[58608] = i[58608];
  assign o[58607] = i[58607];
  assign o[58606] = i[58606];
  assign o[58605] = i[58605];
  assign o[58604] = i[58604];
  assign o[58603] = i[58603];
  assign o[58602] = i[58602];
  assign o[58601] = i[58601];
  assign o[58600] = i[58600];
  assign o[58599] = i[58599];
  assign o[58598] = i[58598];
  assign o[58597] = i[58597];
  assign o[58596] = i[58596];
  assign o[58595] = i[58595];
  assign o[58594] = i[58594];
  assign o[58593] = i[58593];
  assign o[58592] = i[58592];
  assign o[58591] = i[58591];
  assign o[58590] = i[58590];
  assign o[58589] = i[58589];
  assign o[58588] = i[58588];
  assign o[58587] = i[58587];
  assign o[58586] = i[58586];
  assign o[58585] = i[58585];
  assign o[58584] = i[58584];
  assign o[58583] = i[58583];
  assign o[58582] = i[58582];
  assign o[58581] = i[58581];
  assign o[58580] = i[58580];
  assign o[58579] = i[58579];
  assign o[58578] = i[58578];
  assign o[58577] = i[58577];
  assign o[58576] = i[58576];
  assign o[58575] = i[58575];
  assign o[58574] = i[58574];
  assign o[58573] = i[58573];
  assign o[58572] = i[58572];
  assign o[58571] = i[58571];
  assign o[58570] = i[58570];
  assign o[58569] = i[58569];
  assign o[58568] = i[58568];
  assign o[58567] = i[58567];
  assign o[58566] = i[58566];
  assign o[58565] = i[58565];
  assign o[58564] = i[58564];
  assign o[58563] = i[58563];
  assign o[58562] = i[58562];
  assign o[58561] = i[58561];
  assign o[58560] = i[58560];
  assign o[58559] = i[58559];
  assign o[58558] = i[58558];
  assign o[58557] = i[58557];
  assign o[58556] = i[58556];
  assign o[58555] = i[58555];
  assign o[58554] = i[58554];
  assign o[58553] = i[58553];
  assign o[58552] = i[58552];
  assign o[58551] = i[58551];
  assign o[58550] = i[58550];
  assign o[58549] = i[58549];
  assign o[58548] = i[58548];
  assign o[58547] = i[58547];
  assign o[58546] = i[58546];
  assign o[58545] = i[58545];
  assign o[58544] = i[58544];
  assign o[58543] = i[58543];
  assign o[58542] = i[58542];
  assign o[58541] = i[58541];
  assign o[58540] = i[58540];
  assign o[58539] = i[58539];
  assign o[58538] = i[58538];
  assign o[58537] = i[58537];
  assign o[58536] = i[58536];
  assign o[58535] = i[58535];
  assign o[58534] = i[58534];
  assign o[58533] = i[58533];
  assign o[58532] = i[58532];
  assign o[58531] = i[58531];
  assign o[58530] = i[58530];
  assign o[58529] = i[58529];
  assign o[58528] = i[58528];
  assign o[58527] = i[58527];
  assign o[58526] = i[58526];
  assign o[58525] = i[58525];
  assign o[58524] = i[58524];
  assign o[58523] = i[58523];
  assign o[58522] = i[58522];
  assign o[58521] = i[58521];
  assign o[58520] = i[58520];
  assign o[58519] = i[58519];
  assign o[58518] = i[58518];
  assign o[58517] = i[58517];
  assign o[58516] = i[58516];
  assign o[58515] = i[58515];
  assign o[58514] = i[58514];
  assign o[58513] = i[58513];
  assign o[58512] = i[58512];
  assign o[58511] = i[58511];
  assign o[58510] = i[58510];
  assign o[58509] = i[58509];
  assign o[58508] = i[58508];
  assign o[58507] = i[58507];
  assign o[58506] = i[58506];
  assign o[58505] = i[58505];
  assign o[58504] = i[58504];
  assign o[58503] = i[58503];
  assign o[58502] = i[58502];
  assign o[58501] = i[58501];
  assign o[58500] = i[58500];
  assign o[58499] = i[58499];
  assign o[58498] = i[58498];
  assign o[58497] = i[58497];
  assign o[58496] = i[58496];
  assign o[58495] = i[58495];
  assign o[58494] = i[58494];
  assign o[58493] = i[58493];
  assign o[58492] = i[58492];
  assign o[58491] = i[58491];
  assign o[58490] = i[58490];
  assign o[58489] = i[58489];
  assign o[58488] = i[58488];
  assign o[58487] = i[58487];
  assign o[58486] = i[58486];
  assign o[58485] = i[58485];
  assign o[58484] = i[58484];
  assign o[58483] = i[58483];
  assign o[58482] = i[58482];
  assign o[58481] = i[58481];
  assign o[58480] = i[58480];
  assign o[58479] = i[58479];
  assign o[58478] = i[58478];
  assign o[58477] = i[58477];
  assign o[58476] = i[58476];
  assign o[58475] = i[58475];
  assign o[58474] = i[58474];
  assign o[58473] = i[58473];
  assign o[58472] = i[58472];
  assign o[58471] = i[58471];
  assign o[58470] = i[58470];
  assign o[58469] = i[58469];
  assign o[58468] = i[58468];
  assign o[58467] = i[58467];
  assign o[58466] = i[58466];
  assign o[58465] = i[58465];
  assign o[58464] = i[58464];
  assign o[58463] = i[58463];
  assign o[58462] = i[58462];
  assign o[58461] = i[58461];
  assign o[58460] = i[58460];
  assign o[58459] = i[58459];
  assign o[58458] = i[58458];
  assign o[58457] = i[58457];
  assign o[58456] = i[58456];
  assign o[58455] = i[58455];
  assign o[58454] = i[58454];
  assign o[58453] = i[58453];
  assign o[58452] = i[58452];
  assign o[58451] = i[58451];
  assign o[58450] = i[58450];
  assign o[58449] = i[58449];
  assign o[58448] = i[58448];
  assign o[58447] = i[58447];
  assign o[58446] = i[58446];
  assign o[58445] = i[58445];
  assign o[58444] = i[58444];
  assign o[58443] = i[58443];
  assign o[58442] = i[58442];
  assign o[58441] = i[58441];
  assign o[58440] = i[58440];
  assign o[58439] = i[58439];
  assign o[58438] = i[58438];
  assign o[58437] = i[58437];
  assign o[58436] = i[58436];
  assign o[58435] = i[58435];
  assign o[58434] = i[58434];
  assign o[58433] = i[58433];
  assign o[58432] = i[58432];
  assign o[58431] = i[58431];
  assign o[58430] = i[58430];
  assign o[58429] = i[58429];
  assign o[58428] = i[58428];
  assign o[58427] = i[58427];
  assign o[58426] = i[58426];
  assign o[58425] = i[58425];
  assign o[58424] = i[58424];
  assign o[58423] = i[58423];
  assign o[58422] = i[58422];
  assign o[58421] = i[58421];
  assign o[58420] = i[58420];
  assign o[58419] = i[58419];
  assign o[58418] = i[58418];
  assign o[58417] = i[58417];
  assign o[58416] = i[58416];
  assign o[58415] = i[58415];
  assign o[58414] = i[58414];
  assign o[58413] = i[58413];
  assign o[58412] = i[58412];
  assign o[58411] = i[58411];
  assign o[58410] = i[58410];
  assign o[58409] = i[58409];
  assign o[58408] = i[58408];
  assign o[58407] = i[58407];
  assign o[58406] = i[58406];
  assign o[58405] = i[58405];
  assign o[58404] = i[58404];
  assign o[58403] = i[58403];
  assign o[58402] = i[58402];
  assign o[58401] = i[58401];
  assign o[58400] = i[58400];
  assign o[58399] = i[58399];
  assign o[58398] = i[58398];
  assign o[58397] = i[58397];
  assign o[58396] = i[58396];
  assign o[58395] = i[58395];
  assign o[58394] = i[58394];
  assign o[58393] = i[58393];
  assign o[58392] = i[58392];
  assign o[58391] = i[58391];
  assign o[58390] = i[58390];
  assign o[58389] = i[58389];
  assign o[58388] = i[58388];
  assign o[58387] = i[58387];
  assign o[58386] = i[58386];
  assign o[58385] = i[58385];
  assign o[58384] = i[58384];
  assign o[58383] = i[58383];
  assign o[58382] = i[58382];
  assign o[58381] = i[58381];
  assign o[58380] = i[58380];
  assign o[58379] = i[58379];
  assign o[58378] = i[58378];
  assign o[58377] = i[58377];
  assign o[58376] = i[58376];
  assign o[58375] = i[58375];
  assign o[58374] = i[58374];
  assign o[58373] = i[58373];
  assign o[58372] = i[58372];
  assign o[58371] = i[58371];
  assign o[58370] = i[58370];
  assign o[58369] = i[58369];
  assign o[58368] = i[58368];
  assign o[58367] = i[58367];
  assign o[58366] = i[58366];
  assign o[58365] = i[58365];
  assign o[58364] = i[58364];
  assign o[58363] = i[58363];
  assign o[58362] = i[58362];
  assign o[58361] = i[58361];
  assign o[58360] = i[58360];
  assign o[58359] = i[58359];
  assign o[58358] = i[58358];
  assign o[58357] = i[58357];
  assign o[58356] = i[58356];
  assign o[58355] = i[58355];
  assign o[58354] = i[58354];
  assign o[58353] = i[58353];
  assign o[58352] = i[58352];
  assign o[58351] = i[58351];
  assign o[58350] = i[58350];
  assign o[58349] = i[58349];
  assign o[58348] = i[58348];
  assign o[58347] = i[58347];
  assign o[58346] = i[58346];
  assign o[58345] = i[58345];
  assign o[58344] = i[58344];
  assign o[58343] = i[58343];
  assign o[58342] = i[58342];
  assign o[58341] = i[58341];
  assign o[58340] = i[58340];
  assign o[58339] = i[58339];
  assign o[58338] = i[58338];
  assign o[58337] = i[58337];
  assign o[58336] = i[58336];
  assign o[58335] = i[58335];
  assign o[58334] = i[58334];
  assign o[58333] = i[58333];
  assign o[58332] = i[58332];
  assign o[58331] = i[58331];
  assign o[58330] = i[58330];
  assign o[58329] = i[58329];
  assign o[58328] = i[58328];
  assign o[58327] = i[58327];
  assign o[58326] = i[58326];
  assign o[58325] = i[58325];
  assign o[58324] = i[58324];
  assign o[58323] = i[58323];
  assign o[58322] = i[58322];
  assign o[58321] = i[58321];
  assign o[58320] = i[58320];
  assign o[58319] = i[58319];
  assign o[58318] = i[58318];
  assign o[58317] = i[58317];
  assign o[58316] = i[58316];
  assign o[58315] = i[58315];
  assign o[58314] = i[58314];
  assign o[58313] = i[58313];
  assign o[58312] = i[58312];
  assign o[58311] = i[58311];
  assign o[58310] = i[58310];
  assign o[58309] = i[58309];
  assign o[58308] = i[58308];
  assign o[58307] = i[58307];
  assign o[58306] = i[58306];
  assign o[58305] = i[58305];
  assign o[58304] = i[58304];
  assign o[58303] = i[58303];
  assign o[58302] = i[58302];
  assign o[58301] = i[58301];
  assign o[58300] = i[58300];
  assign o[58299] = i[58299];
  assign o[58298] = i[58298];
  assign o[58297] = i[58297];
  assign o[58296] = i[58296];
  assign o[58295] = i[58295];
  assign o[58294] = i[58294];
  assign o[58293] = i[58293];
  assign o[58292] = i[58292];
  assign o[58291] = i[58291];
  assign o[58290] = i[58290];
  assign o[58289] = i[58289];
  assign o[58288] = i[58288];
  assign o[58287] = i[58287];
  assign o[58286] = i[58286];
  assign o[58285] = i[58285];
  assign o[58284] = i[58284];
  assign o[58283] = i[58283];
  assign o[58282] = i[58282];
  assign o[58281] = i[58281];
  assign o[58280] = i[58280];
  assign o[58279] = i[58279];
  assign o[58278] = i[58278];
  assign o[58277] = i[58277];
  assign o[58276] = i[58276];
  assign o[58275] = i[58275];
  assign o[58274] = i[58274];
  assign o[58273] = i[58273];
  assign o[58272] = i[58272];
  assign o[58271] = i[58271];
  assign o[58270] = i[58270];
  assign o[58269] = i[58269];
  assign o[58268] = i[58268];
  assign o[58267] = i[58267];
  assign o[58266] = i[58266];
  assign o[58265] = i[58265];
  assign o[58264] = i[58264];
  assign o[58263] = i[58263];
  assign o[58262] = i[58262];
  assign o[58261] = i[58261];
  assign o[58260] = i[58260];
  assign o[58259] = i[58259];
  assign o[58258] = i[58258];
  assign o[58257] = i[58257];
  assign o[58256] = i[58256];
  assign o[58255] = i[58255];
  assign o[58254] = i[58254];
  assign o[58253] = i[58253];
  assign o[58252] = i[58252];
  assign o[58251] = i[58251];
  assign o[58250] = i[58250];
  assign o[58249] = i[58249];
  assign o[58248] = i[58248];
  assign o[58247] = i[58247];
  assign o[58246] = i[58246];
  assign o[58245] = i[58245];
  assign o[58244] = i[58244];
  assign o[58243] = i[58243];
  assign o[58242] = i[58242];
  assign o[58241] = i[58241];
  assign o[58240] = i[58240];
  assign o[58239] = i[58239];
  assign o[58238] = i[58238];
  assign o[58237] = i[58237];
  assign o[58236] = i[58236];
  assign o[58235] = i[58235];
  assign o[58234] = i[58234];
  assign o[58233] = i[58233];
  assign o[58232] = i[58232];
  assign o[58231] = i[58231];
  assign o[58230] = i[58230];
  assign o[58229] = i[58229];
  assign o[58228] = i[58228];
  assign o[58227] = i[58227];
  assign o[58226] = i[58226];
  assign o[58225] = i[58225];
  assign o[58224] = i[58224];
  assign o[58223] = i[58223];
  assign o[58222] = i[58222];
  assign o[58221] = i[58221];
  assign o[58220] = i[58220];
  assign o[58219] = i[58219];
  assign o[58218] = i[58218];
  assign o[58217] = i[58217];
  assign o[58216] = i[58216];
  assign o[58215] = i[58215];
  assign o[58214] = i[58214];
  assign o[58213] = i[58213];
  assign o[58212] = i[58212];
  assign o[58211] = i[58211];
  assign o[58210] = i[58210];
  assign o[58209] = i[58209];
  assign o[58208] = i[58208];
  assign o[58207] = i[58207];
  assign o[58206] = i[58206];
  assign o[58205] = i[58205];
  assign o[58204] = i[58204];
  assign o[58203] = i[58203];
  assign o[58202] = i[58202];
  assign o[58201] = i[58201];
  assign o[58200] = i[58200];
  assign o[58199] = i[58199];
  assign o[58198] = i[58198];
  assign o[58197] = i[58197];
  assign o[58196] = i[58196];
  assign o[58195] = i[58195];
  assign o[58194] = i[58194];
  assign o[58193] = i[58193];
  assign o[58192] = i[58192];
  assign o[58191] = i[58191];
  assign o[58190] = i[58190];
  assign o[58189] = i[58189];
  assign o[58188] = i[58188];
  assign o[58187] = i[58187];
  assign o[58186] = i[58186];
  assign o[58185] = i[58185];
  assign o[58184] = i[58184];
  assign o[58183] = i[58183];
  assign o[58182] = i[58182];
  assign o[58181] = i[58181];
  assign o[58180] = i[58180];
  assign o[58179] = i[58179];
  assign o[58178] = i[58178];
  assign o[58177] = i[58177];
  assign o[58176] = i[58176];
  assign o[58175] = i[58175];
  assign o[58174] = i[58174];
  assign o[58173] = i[58173];
  assign o[58172] = i[58172];
  assign o[58171] = i[58171];
  assign o[58170] = i[58170];
  assign o[58169] = i[58169];
  assign o[58168] = i[58168];
  assign o[58167] = i[58167];
  assign o[58166] = i[58166];
  assign o[58165] = i[58165];
  assign o[58164] = i[58164];
  assign o[58163] = i[58163];
  assign o[58162] = i[58162];
  assign o[58161] = i[58161];
  assign o[58160] = i[58160];
  assign o[58159] = i[58159];
  assign o[58158] = i[58158];
  assign o[58157] = i[58157];
  assign o[58156] = i[58156];
  assign o[58155] = i[58155];
  assign o[58154] = i[58154];
  assign o[58153] = i[58153];
  assign o[58152] = i[58152];
  assign o[58151] = i[58151];
  assign o[58150] = i[58150];
  assign o[58149] = i[58149];
  assign o[58148] = i[58148];
  assign o[58147] = i[58147];
  assign o[58146] = i[58146];
  assign o[58145] = i[58145];
  assign o[58144] = i[58144];
  assign o[58143] = i[58143];
  assign o[58142] = i[58142];
  assign o[58141] = i[58141];
  assign o[58140] = i[58140];
  assign o[58139] = i[58139];
  assign o[58138] = i[58138];
  assign o[58137] = i[58137];
  assign o[58136] = i[58136];
  assign o[58135] = i[58135];
  assign o[58134] = i[58134];
  assign o[58133] = i[58133];
  assign o[58132] = i[58132];
  assign o[58131] = i[58131];
  assign o[58130] = i[58130];
  assign o[58129] = i[58129];
  assign o[58128] = i[58128];
  assign o[58127] = i[58127];
  assign o[58126] = i[58126];
  assign o[58125] = i[58125];
  assign o[58124] = i[58124];
  assign o[58123] = i[58123];
  assign o[58122] = i[58122];
  assign o[58121] = i[58121];
  assign o[58120] = i[58120];
  assign o[58119] = i[58119];
  assign o[58118] = i[58118];
  assign o[58117] = i[58117];
  assign o[58116] = i[58116];
  assign o[58115] = i[58115];
  assign o[58114] = i[58114];
  assign o[58113] = i[58113];
  assign o[58112] = i[58112];
  assign o[58111] = i[58111];
  assign o[58110] = i[58110];
  assign o[58109] = i[58109];
  assign o[58108] = i[58108];
  assign o[58107] = i[58107];
  assign o[58106] = i[58106];
  assign o[58105] = i[58105];
  assign o[58104] = i[58104];
  assign o[58103] = i[58103];
  assign o[58102] = i[58102];
  assign o[58101] = i[58101];
  assign o[58100] = i[58100];
  assign o[58099] = i[58099];
  assign o[58098] = i[58098];
  assign o[58097] = i[58097];
  assign o[58096] = i[58096];
  assign o[58095] = i[58095];
  assign o[58094] = i[58094];
  assign o[58093] = i[58093];
  assign o[58092] = i[58092];
  assign o[58091] = i[58091];
  assign o[58090] = i[58090];
  assign o[58089] = i[58089];
  assign o[58088] = i[58088];
  assign o[58087] = i[58087];
  assign o[58086] = i[58086];
  assign o[58085] = i[58085];
  assign o[58084] = i[58084];
  assign o[58083] = i[58083];
  assign o[58082] = i[58082];
  assign o[58081] = i[58081];
  assign o[58080] = i[58080];
  assign o[58079] = i[58079];
  assign o[58078] = i[58078];
  assign o[58077] = i[58077];
  assign o[58076] = i[58076];
  assign o[58075] = i[58075];
  assign o[58074] = i[58074];
  assign o[58073] = i[58073];
  assign o[58072] = i[58072];
  assign o[58071] = i[58071];
  assign o[58070] = i[58070];
  assign o[58069] = i[58069];
  assign o[58068] = i[58068];
  assign o[58067] = i[58067];
  assign o[58066] = i[58066];
  assign o[58065] = i[58065];
  assign o[58064] = i[58064];
  assign o[58063] = i[58063];
  assign o[58062] = i[58062];
  assign o[58061] = i[58061];
  assign o[58060] = i[58060];
  assign o[58059] = i[58059];
  assign o[58058] = i[58058];
  assign o[58057] = i[58057];
  assign o[58056] = i[58056];
  assign o[58055] = i[58055];
  assign o[58054] = i[58054];
  assign o[58053] = i[58053];
  assign o[58052] = i[58052];
  assign o[58051] = i[58051];
  assign o[58050] = i[58050];
  assign o[58049] = i[58049];
  assign o[58048] = i[58048];
  assign o[58047] = i[58047];
  assign o[58046] = i[58046];
  assign o[58045] = i[58045];
  assign o[58044] = i[58044];
  assign o[58043] = i[58043];
  assign o[58042] = i[58042];
  assign o[58041] = i[58041];
  assign o[58040] = i[58040];
  assign o[58039] = i[58039];
  assign o[58038] = i[58038];
  assign o[58037] = i[58037];
  assign o[58036] = i[58036];
  assign o[58035] = i[58035];
  assign o[58034] = i[58034];
  assign o[58033] = i[58033];
  assign o[58032] = i[58032];
  assign o[58031] = i[58031];
  assign o[58030] = i[58030];
  assign o[58029] = i[58029];
  assign o[58028] = i[58028];
  assign o[58027] = i[58027];
  assign o[58026] = i[58026];
  assign o[58025] = i[58025];
  assign o[58024] = i[58024];
  assign o[58023] = i[58023];
  assign o[58022] = i[58022];
  assign o[58021] = i[58021];
  assign o[58020] = i[58020];
  assign o[58019] = i[58019];
  assign o[58018] = i[58018];
  assign o[58017] = i[58017];
  assign o[58016] = i[58016];
  assign o[58015] = i[58015];
  assign o[58014] = i[58014];
  assign o[58013] = i[58013];
  assign o[58012] = i[58012];
  assign o[58011] = i[58011];
  assign o[58010] = i[58010];
  assign o[58009] = i[58009];
  assign o[58008] = i[58008];
  assign o[58007] = i[58007];
  assign o[58006] = i[58006];
  assign o[58005] = i[58005];
  assign o[58004] = i[58004];
  assign o[58003] = i[58003];
  assign o[58002] = i[58002];
  assign o[58001] = i[58001];
  assign o[58000] = i[58000];
  assign o[57999] = i[57999];
  assign o[57998] = i[57998];
  assign o[57997] = i[57997];
  assign o[57996] = i[57996];
  assign o[57995] = i[57995];
  assign o[57994] = i[57994];
  assign o[57993] = i[57993];
  assign o[57992] = i[57992];
  assign o[57991] = i[57991];
  assign o[57990] = i[57990];
  assign o[57989] = i[57989];
  assign o[57988] = i[57988];
  assign o[57987] = i[57987];
  assign o[57986] = i[57986];
  assign o[57985] = i[57985];
  assign o[57984] = i[57984];
  assign o[57983] = i[57983];
  assign o[57982] = i[57982];
  assign o[57981] = i[57981];
  assign o[57980] = i[57980];
  assign o[57979] = i[57979];
  assign o[57978] = i[57978];
  assign o[57977] = i[57977];
  assign o[57976] = i[57976];
  assign o[57975] = i[57975];
  assign o[57974] = i[57974];
  assign o[57973] = i[57973];
  assign o[57972] = i[57972];
  assign o[57971] = i[57971];
  assign o[57970] = i[57970];
  assign o[57969] = i[57969];
  assign o[57968] = i[57968];
  assign o[57967] = i[57967];
  assign o[57966] = i[57966];
  assign o[57965] = i[57965];
  assign o[57964] = i[57964];
  assign o[57963] = i[57963];
  assign o[57962] = i[57962];
  assign o[57961] = i[57961];
  assign o[57960] = i[57960];
  assign o[57959] = i[57959];
  assign o[57958] = i[57958];
  assign o[57957] = i[57957];
  assign o[57956] = i[57956];
  assign o[57955] = i[57955];
  assign o[57954] = i[57954];
  assign o[57953] = i[57953];
  assign o[57952] = i[57952];
  assign o[57951] = i[57951];
  assign o[57950] = i[57950];
  assign o[57949] = i[57949];
  assign o[57948] = i[57948];
  assign o[57947] = i[57947];
  assign o[57946] = i[57946];
  assign o[57945] = i[57945];
  assign o[57944] = i[57944];
  assign o[57943] = i[57943];
  assign o[57942] = i[57942];
  assign o[57941] = i[57941];
  assign o[57940] = i[57940];
  assign o[57939] = i[57939];
  assign o[57938] = i[57938];
  assign o[57937] = i[57937];
  assign o[57936] = i[57936];
  assign o[57935] = i[57935];
  assign o[57934] = i[57934];
  assign o[57933] = i[57933];
  assign o[57932] = i[57932];
  assign o[57931] = i[57931];
  assign o[57930] = i[57930];
  assign o[57929] = i[57929];
  assign o[57928] = i[57928];
  assign o[57927] = i[57927];
  assign o[57926] = i[57926];
  assign o[57925] = i[57925];
  assign o[57924] = i[57924];
  assign o[57923] = i[57923];
  assign o[57922] = i[57922];
  assign o[57921] = i[57921];
  assign o[57920] = i[57920];
  assign o[57919] = i[57919];
  assign o[57918] = i[57918];
  assign o[57917] = i[57917];
  assign o[57916] = i[57916];
  assign o[57915] = i[57915];
  assign o[57914] = i[57914];
  assign o[57913] = i[57913];
  assign o[57912] = i[57912];
  assign o[57911] = i[57911];
  assign o[57910] = i[57910];
  assign o[57909] = i[57909];
  assign o[57908] = i[57908];
  assign o[57907] = i[57907];
  assign o[57906] = i[57906];
  assign o[57905] = i[57905];
  assign o[57904] = i[57904];
  assign o[57903] = i[57903];
  assign o[57902] = i[57902];
  assign o[57901] = i[57901];
  assign o[57900] = i[57900];
  assign o[57899] = i[57899];
  assign o[57898] = i[57898];
  assign o[57897] = i[57897];
  assign o[57896] = i[57896];
  assign o[57895] = i[57895];
  assign o[57894] = i[57894];
  assign o[57893] = i[57893];
  assign o[57892] = i[57892];
  assign o[57891] = i[57891];
  assign o[57890] = i[57890];
  assign o[57889] = i[57889];
  assign o[57888] = i[57888];
  assign o[57887] = i[57887];
  assign o[57886] = i[57886];
  assign o[57885] = i[57885];
  assign o[57884] = i[57884];
  assign o[57883] = i[57883];
  assign o[57882] = i[57882];
  assign o[57881] = i[57881];
  assign o[57880] = i[57880];
  assign o[57879] = i[57879];
  assign o[57878] = i[57878];
  assign o[57877] = i[57877];
  assign o[57876] = i[57876];
  assign o[57875] = i[57875];
  assign o[57874] = i[57874];
  assign o[57873] = i[57873];
  assign o[57872] = i[57872];
  assign o[57871] = i[57871];
  assign o[57870] = i[57870];
  assign o[57869] = i[57869];
  assign o[57868] = i[57868];
  assign o[57867] = i[57867];
  assign o[57866] = i[57866];
  assign o[57865] = i[57865];
  assign o[57864] = i[57864];
  assign o[57863] = i[57863];
  assign o[57862] = i[57862];
  assign o[57861] = i[57861];
  assign o[57860] = i[57860];
  assign o[57859] = i[57859];
  assign o[57858] = i[57858];
  assign o[57857] = i[57857];
  assign o[57856] = i[57856];
  assign o[57855] = i[57855];
  assign o[57854] = i[57854];
  assign o[57853] = i[57853];
  assign o[57852] = i[57852];
  assign o[57851] = i[57851];
  assign o[57850] = i[57850];
  assign o[57849] = i[57849];
  assign o[57848] = i[57848];
  assign o[57847] = i[57847];
  assign o[57846] = i[57846];
  assign o[57845] = i[57845];
  assign o[57844] = i[57844];
  assign o[57843] = i[57843];
  assign o[57842] = i[57842];
  assign o[57841] = i[57841];
  assign o[57840] = i[57840];
  assign o[57839] = i[57839];
  assign o[57838] = i[57838];
  assign o[57837] = i[57837];
  assign o[57836] = i[57836];
  assign o[57835] = i[57835];
  assign o[57834] = i[57834];
  assign o[57833] = i[57833];
  assign o[57832] = i[57832];
  assign o[57831] = i[57831];
  assign o[57830] = i[57830];
  assign o[57829] = i[57829];
  assign o[57828] = i[57828];
  assign o[57827] = i[57827];
  assign o[57826] = i[57826];
  assign o[57825] = i[57825];
  assign o[57824] = i[57824];
  assign o[57823] = i[57823];
  assign o[57822] = i[57822];
  assign o[57821] = i[57821];
  assign o[57820] = i[57820];
  assign o[57819] = i[57819];
  assign o[57818] = i[57818];
  assign o[57817] = i[57817];
  assign o[57816] = i[57816];
  assign o[57815] = i[57815];
  assign o[57814] = i[57814];
  assign o[57813] = i[57813];
  assign o[57812] = i[57812];
  assign o[57811] = i[57811];
  assign o[57810] = i[57810];
  assign o[57809] = i[57809];
  assign o[57808] = i[57808];
  assign o[57807] = i[57807];
  assign o[57806] = i[57806];
  assign o[57805] = i[57805];
  assign o[57804] = i[57804];
  assign o[57803] = i[57803];
  assign o[57802] = i[57802];
  assign o[57801] = i[57801];
  assign o[57800] = i[57800];
  assign o[57799] = i[57799];
  assign o[57798] = i[57798];
  assign o[57797] = i[57797];
  assign o[57796] = i[57796];
  assign o[57795] = i[57795];
  assign o[57794] = i[57794];
  assign o[57793] = i[57793];
  assign o[57792] = i[57792];
  assign o[57791] = i[57791];
  assign o[57790] = i[57790];
  assign o[57789] = i[57789];
  assign o[57788] = i[57788];
  assign o[57787] = i[57787];
  assign o[57786] = i[57786];
  assign o[57785] = i[57785];
  assign o[57784] = i[57784];
  assign o[57783] = i[57783];
  assign o[57782] = i[57782];
  assign o[57781] = i[57781];
  assign o[57780] = i[57780];
  assign o[57779] = i[57779];
  assign o[57778] = i[57778];
  assign o[57777] = i[57777];
  assign o[57776] = i[57776];
  assign o[57775] = i[57775];
  assign o[57774] = i[57774];
  assign o[57773] = i[57773];
  assign o[57772] = i[57772];
  assign o[57771] = i[57771];
  assign o[57770] = i[57770];
  assign o[57769] = i[57769];
  assign o[57768] = i[57768];
  assign o[57767] = i[57767];
  assign o[57766] = i[57766];
  assign o[57765] = i[57765];
  assign o[57764] = i[57764];
  assign o[57763] = i[57763];
  assign o[57762] = i[57762];
  assign o[57761] = i[57761];
  assign o[57760] = i[57760];
  assign o[57759] = i[57759];
  assign o[57758] = i[57758];
  assign o[57757] = i[57757];
  assign o[57756] = i[57756];
  assign o[57755] = i[57755];
  assign o[57754] = i[57754];
  assign o[57753] = i[57753];
  assign o[57752] = i[57752];
  assign o[57751] = i[57751];
  assign o[57750] = i[57750];
  assign o[57749] = i[57749];
  assign o[57748] = i[57748];
  assign o[57747] = i[57747];
  assign o[57746] = i[57746];
  assign o[57745] = i[57745];
  assign o[57744] = i[57744];
  assign o[57743] = i[57743];
  assign o[57742] = i[57742];
  assign o[57741] = i[57741];
  assign o[57740] = i[57740];
  assign o[57739] = i[57739];
  assign o[57738] = i[57738];
  assign o[57737] = i[57737];
  assign o[57736] = i[57736];
  assign o[57735] = i[57735];
  assign o[57734] = i[57734];
  assign o[57733] = i[57733];
  assign o[57732] = i[57732];
  assign o[57731] = i[57731];
  assign o[57730] = i[57730];
  assign o[57729] = i[57729];
  assign o[57728] = i[57728];
  assign o[57727] = i[57727];
  assign o[57726] = i[57726];
  assign o[57725] = i[57725];
  assign o[57724] = i[57724];
  assign o[57723] = i[57723];
  assign o[57722] = i[57722];
  assign o[57721] = i[57721];
  assign o[57720] = i[57720];
  assign o[57719] = i[57719];
  assign o[57718] = i[57718];
  assign o[57717] = i[57717];
  assign o[57716] = i[57716];
  assign o[57715] = i[57715];
  assign o[57714] = i[57714];
  assign o[57713] = i[57713];
  assign o[57712] = i[57712];
  assign o[57711] = i[57711];
  assign o[57710] = i[57710];
  assign o[57709] = i[57709];
  assign o[57708] = i[57708];
  assign o[57707] = i[57707];
  assign o[57706] = i[57706];
  assign o[57705] = i[57705];
  assign o[57704] = i[57704];
  assign o[57703] = i[57703];
  assign o[57702] = i[57702];
  assign o[57701] = i[57701];
  assign o[57700] = i[57700];
  assign o[57699] = i[57699];
  assign o[57698] = i[57698];
  assign o[57697] = i[57697];
  assign o[57696] = i[57696];
  assign o[57695] = i[57695];
  assign o[57694] = i[57694];
  assign o[57693] = i[57693];
  assign o[57692] = i[57692];
  assign o[57691] = i[57691];
  assign o[57690] = i[57690];
  assign o[57689] = i[57689];
  assign o[57688] = i[57688];
  assign o[57687] = i[57687];
  assign o[57686] = i[57686];
  assign o[57685] = i[57685];
  assign o[57684] = i[57684];
  assign o[57683] = i[57683];
  assign o[57682] = i[57682];
  assign o[57681] = i[57681];
  assign o[57680] = i[57680];
  assign o[57679] = i[57679];
  assign o[57678] = i[57678];
  assign o[57677] = i[57677];
  assign o[57676] = i[57676];
  assign o[57675] = i[57675];
  assign o[57674] = i[57674];
  assign o[57673] = i[57673];
  assign o[57672] = i[57672];
  assign o[57671] = i[57671];
  assign o[57670] = i[57670];
  assign o[57669] = i[57669];
  assign o[57668] = i[57668];
  assign o[57667] = i[57667];
  assign o[57666] = i[57666];
  assign o[57665] = i[57665];
  assign o[57664] = i[57664];
  assign o[57663] = i[57663];
  assign o[57662] = i[57662];
  assign o[57661] = i[57661];
  assign o[57660] = i[57660];
  assign o[57659] = i[57659];
  assign o[57658] = i[57658];
  assign o[57657] = i[57657];
  assign o[57656] = i[57656];
  assign o[57655] = i[57655];
  assign o[57654] = i[57654];
  assign o[57653] = i[57653];
  assign o[57652] = i[57652];
  assign o[57651] = i[57651];
  assign o[57650] = i[57650];
  assign o[57649] = i[57649];
  assign o[57648] = i[57648];
  assign o[57647] = i[57647];
  assign o[57646] = i[57646];
  assign o[57645] = i[57645];
  assign o[57644] = i[57644];
  assign o[57643] = i[57643];
  assign o[57642] = i[57642];
  assign o[57641] = i[57641];
  assign o[57640] = i[57640];
  assign o[57639] = i[57639];
  assign o[57638] = i[57638];
  assign o[57637] = i[57637];
  assign o[57636] = i[57636];
  assign o[57635] = i[57635];
  assign o[57634] = i[57634];
  assign o[57633] = i[57633];
  assign o[57632] = i[57632];
  assign o[57631] = i[57631];
  assign o[57630] = i[57630];
  assign o[57629] = i[57629];
  assign o[57628] = i[57628];
  assign o[57627] = i[57627];
  assign o[57626] = i[57626];
  assign o[57625] = i[57625];
  assign o[57624] = i[57624];
  assign o[57623] = i[57623];
  assign o[57622] = i[57622];
  assign o[57621] = i[57621];
  assign o[57620] = i[57620];
  assign o[57619] = i[57619];
  assign o[57618] = i[57618];
  assign o[57617] = i[57617];
  assign o[57616] = i[57616];
  assign o[57615] = i[57615];
  assign o[57614] = i[57614];
  assign o[57613] = i[57613];
  assign o[57612] = i[57612];
  assign o[57611] = i[57611];
  assign o[57610] = i[57610];
  assign o[57609] = i[57609];
  assign o[57608] = i[57608];
  assign o[57607] = i[57607];
  assign o[57606] = i[57606];
  assign o[57605] = i[57605];
  assign o[57604] = i[57604];
  assign o[57603] = i[57603];
  assign o[57602] = i[57602];
  assign o[57601] = i[57601];
  assign o[57600] = i[57600];
  assign o[57599] = i[57599];
  assign o[57598] = i[57598];
  assign o[57597] = i[57597];
  assign o[57596] = i[57596];
  assign o[57595] = i[57595];
  assign o[57594] = i[57594];
  assign o[57593] = i[57593];
  assign o[57592] = i[57592];
  assign o[57591] = i[57591];
  assign o[57590] = i[57590];
  assign o[57589] = i[57589];
  assign o[57588] = i[57588];
  assign o[57587] = i[57587];
  assign o[57586] = i[57586];
  assign o[57585] = i[57585];
  assign o[57584] = i[57584];
  assign o[57583] = i[57583];
  assign o[57582] = i[57582];
  assign o[57581] = i[57581];
  assign o[57580] = i[57580];
  assign o[57579] = i[57579];
  assign o[57578] = i[57578];
  assign o[57577] = i[57577];
  assign o[57576] = i[57576];
  assign o[57575] = i[57575];
  assign o[57574] = i[57574];
  assign o[57573] = i[57573];
  assign o[57572] = i[57572];
  assign o[57571] = i[57571];
  assign o[57570] = i[57570];
  assign o[57569] = i[57569];
  assign o[57568] = i[57568];
  assign o[57567] = i[57567];
  assign o[57566] = i[57566];
  assign o[57565] = i[57565];
  assign o[57564] = i[57564];
  assign o[57563] = i[57563];
  assign o[57562] = i[57562];
  assign o[57561] = i[57561];
  assign o[57560] = i[57560];
  assign o[57559] = i[57559];
  assign o[57558] = i[57558];
  assign o[57557] = i[57557];
  assign o[57556] = i[57556];
  assign o[57555] = i[57555];
  assign o[57554] = i[57554];
  assign o[57553] = i[57553];
  assign o[57552] = i[57552];
  assign o[57551] = i[57551];
  assign o[57550] = i[57550];
  assign o[57549] = i[57549];
  assign o[57548] = i[57548];
  assign o[57547] = i[57547];
  assign o[57546] = i[57546];
  assign o[57545] = i[57545];
  assign o[57544] = i[57544];
  assign o[57543] = i[57543];
  assign o[57542] = i[57542];
  assign o[57541] = i[57541];
  assign o[57540] = i[57540];
  assign o[57539] = i[57539];
  assign o[57538] = i[57538];
  assign o[57537] = i[57537];
  assign o[57536] = i[57536];
  assign o[57535] = i[57535];
  assign o[57534] = i[57534];
  assign o[57533] = i[57533];
  assign o[57532] = i[57532];
  assign o[57531] = i[57531];
  assign o[57530] = i[57530];
  assign o[57529] = i[57529];
  assign o[57528] = i[57528];
  assign o[57527] = i[57527];
  assign o[57526] = i[57526];
  assign o[57525] = i[57525];
  assign o[57524] = i[57524];
  assign o[57523] = i[57523];
  assign o[57522] = i[57522];
  assign o[57521] = i[57521];
  assign o[57520] = i[57520];
  assign o[57519] = i[57519];
  assign o[57518] = i[57518];
  assign o[57517] = i[57517];
  assign o[57516] = i[57516];
  assign o[57515] = i[57515];
  assign o[57514] = i[57514];
  assign o[57513] = i[57513];
  assign o[57512] = i[57512];
  assign o[57511] = i[57511];
  assign o[57510] = i[57510];
  assign o[57509] = i[57509];
  assign o[57508] = i[57508];
  assign o[57507] = i[57507];
  assign o[57506] = i[57506];
  assign o[57505] = i[57505];
  assign o[57504] = i[57504];
  assign o[57503] = i[57503];
  assign o[57502] = i[57502];
  assign o[57501] = i[57501];
  assign o[57500] = i[57500];
  assign o[57499] = i[57499];
  assign o[57498] = i[57498];
  assign o[57497] = i[57497];
  assign o[57496] = i[57496];
  assign o[57495] = i[57495];
  assign o[57494] = i[57494];
  assign o[57493] = i[57493];
  assign o[57492] = i[57492];
  assign o[57491] = i[57491];
  assign o[57490] = i[57490];
  assign o[57489] = i[57489];
  assign o[57488] = i[57488];
  assign o[57487] = i[57487];
  assign o[57486] = i[57486];
  assign o[57485] = i[57485];
  assign o[57484] = i[57484];
  assign o[57483] = i[57483];
  assign o[57482] = i[57482];
  assign o[57481] = i[57481];
  assign o[57480] = i[57480];
  assign o[57479] = i[57479];
  assign o[57478] = i[57478];
  assign o[57477] = i[57477];
  assign o[57476] = i[57476];
  assign o[57475] = i[57475];
  assign o[57474] = i[57474];
  assign o[57473] = i[57473];
  assign o[57472] = i[57472];
  assign o[57471] = i[57471];
  assign o[57470] = i[57470];
  assign o[57469] = i[57469];
  assign o[57468] = i[57468];
  assign o[57467] = i[57467];
  assign o[57466] = i[57466];
  assign o[57465] = i[57465];
  assign o[57464] = i[57464];
  assign o[57463] = i[57463];
  assign o[57462] = i[57462];
  assign o[57461] = i[57461];
  assign o[57460] = i[57460];
  assign o[57459] = i[57459];
  assign o[57458] = i[57458];
  assign o[57457] = i[57457];
  assign o[57456] = i[57456];
  assign o[57455] = i[57455];
  assign o[57454] = i[57454];
  assign o[57453] = i[57453];
  assign o[57452] = i[57452];
  assign o[57451] = i[57451];
  assign o[57450] = i[57450];
  assign o[57449] = i[57449];
  assign o[57448] = i[57448];
  assign o[57447] = i[57447];
  assign o[57446] = i[57446];
  assign o[57445] = i[57445];
  assign o[57444] = i[57444];
  assign o[57443] = i[57443];
  assign o[57442] = i[57442];
  assign o[57441] = i[57441];
  assign o[57440] = i[57440];
  assign o[57439] = i[57439];
  assign o[57438] = i[57438];
  assign o[57437] = i[57437];
  assign o[57436] = i[57436];
  assign o[57435] = i[57435];
  assign o[57434] = i[57434];
  assign o[57433] = i[57433];
  assign o[57432] = i[57432];
  assign o[57431] = i[57431];
  assign o[57430] = i[57430];
  assign o[57429] = i[57429];
  assign o[57428] = i[57428];
  assign o[57427] = i[57427];
  assign o[57426] = i[57426];
  assign o[57425] = i[57425];
  assign o[57424] = i[57424];
  assign o[57423] = i[57423];
  assign o[57422] = i[57422];
  assign o[57421] = i[57421];
  assign o[57420] = i[57420];
  assign o[57419] = i[57419];
  assign o[57418] = i[57418];
  assign o[57417] = i[57417];
  assign o[57416] = i[57416];
  assign o[57415] = i[57415];
  assign o[57414] = i[57414];
  assign o[57413] = i[57413];
  assign o[57412] = i[57412];
  assign o[57411] = i[57411];
  assign o[57410] = i[57410];
  assign o[57409] = i[57409];
  assign o[57408] = i[57408];
  assign o[57407] = i[57407];
  assign o[57406] = i[57406];
  assign o[57405] = i[57405];
  assign o[57404] = i[57404];
  assign o[57403] = i[57403];
  assign o[57402] = i[57402];
  assign o[57401] = i[57401];
  assign o[57400] = i[57400];
  assign o[57399] = i[57399];
  assign o[57398] = i[57398];
  assign o[57397] = i[57397];
  assign o[57396] = i[57396];
  assign o[57395] = i[57395];
  assign o[57394] = i[57394];
  assign o[57393] = i[57393];
  assign o[57392] = i[57392];
  assign o[57391] = i[57391];
  assign o[57390] = i[57390];
  assign o[57389] = i[57389];
  assign o[57388] = i[57388];
  assign o[57387] = i[57387];
  assign o[57386] = i[57386];
  assign o[57385] = i[57385];
  assign o[57384] = i[57384];
  assign o[57383] = i[57383];
  assign o[57382] = i[57382];
  assign o[57381] = i[57381];
  assign o[57380] = i[57380];
  assign o[57379] = i[57379];
  assign o[57378] = i[57378];
  assign o[57377] = i[57377];
  assign o[57376] = i[57376];
  assign o[57375] = i[57375];
  assign o[57374] = i[57374];
  assign o[57373] = i[57373];
  assign o[57372] = i[57372];
  assign o[57371] = i[57371];
  assign o[57370] = i[57370];
  assign o[57369] = i[57369];
  assign o[57368] = i[57368];
  assign o[57367] = i[57367];
  assign o[57366] = i[57366];
  assign o[57365] = i[57365];
  assign o[57364] = i[57364];
  assign o[57363] = i[57363];
  assign o[57362] = i[57362];
  assign o[57361] = i[57361];
  assign o[57360] = i[57360];
  assign o[57359] = i[57359];
  assign o[57358] = i[57358];
  assign o[57357] = i[57357];
  assign o[57356] = i[57356];
  assign o[57355] = i[57355];
  assign o[57354] = i[57354];
  assign o[57353] = i[57353];
  assign o[57352] = i[57352];
  assign o[57351] = i[57351];
  assign o[57350] = i[57350];
  assign o[57349] = i[57349];
  assign o[57348] = i[57348];
  assign o[57347] = i[57347];
  assign o[57346] = i[57346];
  assign o[57345] = i[57345];
  assign o[57344] = i[57344];
  assign o[57343] = i[57343];
  assign o[57342] = i[57342];
  assign o[57341] = i[57341];
  assign o[57340] = i[57340];
  assign o[57339] = i[57339];
  assign o[57338] = i[57338];
  assign o[57337] = i[57337];
  assign o[57336] = i[57336];
  assign o[57335] = i[57335];
  assign o[57334] = i[57334];
  assign o[57333] = i[57333];
  assign o[57332] = i[57332];
  assign o[57331] = i[57331];
  assign o[57330] = i[57330];
  assign o[57329] = i[57329];
  assign o[57328] = i[57328];
  assign o[57327] = i[57327];
  assign o[57326] = i[57326];
  assign o[57325] = i[57325];
  assign o[57324] = i[57324];
  assign o[57323] = i[57323];
  assign o[57322] = i[57322];
  assign o[57321] = i[57321];
  assign o[57320] = i[57320];
  assign o[57319] = i[57319];
  assign o[57318] = i[57318];
  assign o[57317] = i[57317];
  assign o[57316] = i[57316];
  assign o[57315] = i[57315];
  assign o[57314] = i[57314];
  assign o[57313] = i[57313];
  assign o[57312] = i[57312];
  assign o[57311] = i[57311];
  assign o[57310] = i[57310];
  assign o[57309] = i[57309];
  assign o[57308] = i[57308];
  assign o[57307] = i[57307];
  assign o[57306] = i[57306];
  assign o[57305] = i[57305];
  assign o[57304] = i[57304];
  assign o[57303] = i[57303];
  assign o[57302] = i[57302];
  assign o[57301] = i[57301];
  assign o[57300] = i[57300];
  assign o[57299] = i[57299];
  assign o[57298] = i[57298];
  assign o[57297] = i[57297];
  assign o[57296] = i[57296];
  assign o[57295] = i[57295];
  assign o[57294] = i[57294];
  assign o[57293] = i[57293];
  assign o[57292] = i[57292];
  assign o[57291] = i[57291];
  assign o[57290] = i[57290];
  assign o[57289] = i[57289];
  assign o[57288] = i[57288];
  assign o[57287] = i[57287];
  assign o[57286] = i[57286];
  assign o[57285] = i[57285];
  assign o[57284] = i[57284];
  assign o[57283] = i[57283];
  assign o[57282] = i[57282];
  assign o[57281] = i[57281];
  assign o[57280] = i[57280];
  assign o[57279] = i[57279];
  assign o[57278] = i[57278];
  assign o[57277] = i[57277];
  assign o[57276] = i[57276];
  assign o[57275] = i[57275];
  assign o[57274] = i[57274];
  assign o[57273] = i[57273];
  assign o[57272] = i[57272];
  assign o[57271] = i[57271];
  assign o[57270] = i[57270];
  assign o[57269] = i[57269];
  assign o[57268] = i[57268];
  assign o[57267] = i[57267];
  assign o[57266] = i[57266];
  assign o[57265] = i[57265];
  assign o[57264] = i[57264];
  assign o[57263] = i[57263];
  assign o[57262] = i[57262];
  assign o[57261] = i[57261];
  assign o[57260] = i[57260];
  assign o[57259] = i[57259];
  assign o[57258] = i[57258];
  assign o[57257] = i[57257];
  assign o[57256] = i[57256];
  assign o[57255] = i[57255];
  assign o[57254] = i[57254];
  assign o[57253] = i[57253];
  assign o[57252] = i[57252];
  assign o[57251] = i[57251];
  assign o[57250] = i[57250];
  assign o[57249] = i[57249];
  assign o[57248] = i[57248];
  assign o[57247] = i[57247];
  assign o[57246] = i[57246];
  assign o[57245] = i[57245];
  assign o[57244] = i[57244];
  assign o[57243] = i[57243];
  assign o[57242] = i[57242];
  assign o[57241] = i[57241];
  assign o[57240] = i[57240];
  assign o[57239] = i[57239];
  assign o[57238] = i[57238];
  assign o[57237] = i[57237];
  assign o[57236] = i[57236];
  assign o[57235] = i[57235];
  assign o[57234] = i[57234];
  assign o[57233] = i[57233];
  assign o[57232] = i[57232];
  assign o[57231] = i[57231];
  assign o[57230] = i[57230];
  assign o[57229] = i[57229];
  assign o[57228] = i[57228];
  assign o[57227] = i[57227];
  assign o[57226] = i[57226];
  assign o[57225] = i[57225];
  assign o[57224] = i[57224];
  assign o[57223] = i[57223];
  assign o[57222] = i[57222];
  assign o[57221] = i[57221];
  assign o[57220] = i[57220];
  assign o[57219] = i[57219];
  assign o[57218] = i[57218];
  assign o[57217] = i[57217];
  assign o[57216] = i[57216];
  assign o[57215] = i[57215];
  assign o[57214] = i[57214];
  assign o[57213] = i[57213];
  assign o[57212] = i[57212];
  assign o[57211] = i[57211];
  assign o[57210] = i[57210];
  assign o[57209] = i[57209];
  assign o[57208] = i[57208];
  assign o[57207] = i[57207];
  assign o[57206] = i[57206];
  assign o[57205] = i[57205];
  assign o[57204] = i[57204];
  assign o[57203] = i[57203];
  assign o[57202] = i[57202];
  assign o[57201] = i[57201];
  assign o[57200] = i[57200];
  assign o[57199] = i[57199];
  assign o[57198] = i[57198];
  assign o[57197] = i[57197];
  assign o[57196] = i[57196];
  assign o[57195] = i[57195];
  assign o[57194] = i[57194];
  assign o[57193] = i[57193];
  assign o[57192] = i[57192];
  assign o[57191] = i[57191];
  assign o[57190] = i[57190];
  assign o[57189] = i[57189];
  assign o[57188] = i[57188];
  assign o[57187] = i[57187];
  assign o[57186] = i[57186];
  assign o[57185] = i[57185];
  assign o[57184] = i[57184];
  assign o[57183] = i[57183];
  assign o[57182] = i[57182];
  assign o[57181] = i[57181];
  assign o[57180] = i[57180];
  assign o[57179] = i[57179];
  assign o[57178] = i[57178];
  assign o[57177] = i[57177];
  assign o[57176] = i[57176];
  assign o[57175] = i[57175];
  assign o[57174] = i[57174];
  assign o[57173] = i[57173];
  assign o[57172] = i[57172];
  assign o[57171] = i[57171];
  assign o[57170] = i[57170];
  assign o[57169] = i[57169];
  assign o[57168] = i[57168];
  assign o[57167] = i[57167];
  assign o[57166] = i[57166];
  assign o[57165] = i[57165];
  assign o[57164] = i[57164];
  assign o[57163] = i[57163];
  assign o[57162] = i[57162];
  assign o[57161] = i[57161];
  assign o[57160] = i[57160];
  assign o[57159] = i[57159];
  assign o[57158] = i[57158];
  assign o[57157] = i[57157];
  assign o[57156] = i[57156];
  assign o[57155] = i[57155];
  assign o[57154] = i[57154];
  assign o[57153] = i[57153];
  assign o[57152] = i[57152];
  assign o[57151] = i[57151];
  assign o[57150] = i[57150];
  assign o[57149] = i[57149];
  assign o[57148] = i[57148];
  assign o[57147] = i[57147];
  assign o[57146] = i[57146];
  assign o[57145] = i[57145];
  assign o[57144] = i[57144];
  assign o[57143] = i[57143];
  assign o[57142] = i[57142];
  assign o[57141] = i[57141];
  assign o[57140] = i[57140];
  assign o[57139] = i[57139];
  assign o[57138] = i[57138];
  assign o[57137] = i[57137];
  assign o[57136] = i[57136];
  assign o[57135] = i[57135];
  assign o[57134] = i[57134];
  assign o[57133] = i[57133];
  assign o[57132] = i[57132];
  assign o[57131] = i[57131];
  assign o[57130] = i[57130];
  assign o[57129] = i[57129];
  assign o[57128] = i[57128];
  assign o[57127] = i[57127];
  assign o[57126] = i[57126];
  assign o[57125] = i[57125];
  assign o[57124] = i[57124];
  assign o[57123] = i[57123];
  assign o[57122] = i[57122];
  assign o[57121] = i[57121];
  assign o[57120] = i[57120];
  assign o[57119] = i[57119];
  assign o[57118] = i[57118];
  assign o[57117] = i[57117];
  assign o[57116] = i[57116];
  assign o[57115] = i[57115];
  assign o[57114] = i[57114];
  assign o[57113] = i[57113];
  assign o[57112] = i[57112];
  assign o[57111] = i[57111];
  assign o[57110] = i[57110];
  assign o[57109] = i[57109];
  assign o[57108] = i[57108];
  assign o[57107] = i[57107];
  assign o[57106] = i[57106];
  assign o[57105] = i[57105];
  assign o[57104] = i[57104];
  assign o[57103] = i[57103];
  assign o[57102] = i[57102];
  assign o[57101] = i[57101];
  assign o[57100] = i[57100];
  assign o[57099] = i[57099];
  assign o[57098] = i[57098];
  assign o[57097] = i[57097];
  assign o[57096] = i[57096];
  assign o[57095] = i[57095];
  assign o[57094] = i[57094];
  assign o[57093] = i[57093];
  assign o[57092] = i[57092];
  assign o[57091] = i[57091];
  assign o[57090] = i[57090];
  assign o[57089] = i[57089];
  assign o[57088] = i[57088];
  assign o[57087] = i[57087];
  assign o[57086] = i[57086];
  assign o[57085] = i[57085];
  assign o[57084] = i[57084];
  assign o[57083] = i[57083];
  assign o[57082] = i[57082];
  assign o[57081] = i[57081];
  assign o[57080] = i[57080];
  assign o[57079] = i[57079];
  assign o[57078] = i[57078];
  assign o[57077] = i[57077];
  assign o[57076] = i[57076];
  assign o[57075] = i[57075];
  assign o[57074] = i[57074];
  assign o[57073] = i[57073];
  assign o[57072] = i[57072];
  assign o[57071] = i[57071];
  assign o[57070] = i[57070];
  assign o[57069] = i[57069];
  assign o[57068] = i[57068];
  assign o[57067] = i[57067];
  assign o[57066] = i[57066];
  assign o[57065] = i[57065];
  assign o[57064] = i[57064];
  assign o[57063] = i[57063];
  assign o[57062] = i[57062];
  assign o[57061] = i[57061];
  assign o[57060] = i[57060];
  assign o[57059] = i[57059];
  assign o[57058] = i[57058];
  assign o[57057] = i[57057];
  assign o[57056] = i[57056];
  assign o[57055] = i[57055];
  assign o[57054] = i[57054];
  assign o[57053] = i[57053];
  assign o[57052] = i[57052];
  assign o[57051] = i[57051];
  assign o[57050] = i[57050];
  assign o[57049] = i[57049];
  assign o[57048] = i[57048];
  assign o[57047] = i[57047];
  assign o[57046] = i[57046];
  assign o[57045] = i[57045];
  assign o[57044] = i[57044];
  assign o[57043] = i[57043];
  assign o[57042] = i[57042];
  assign o[57041] = i[57041];
  assign o[57040] = i[57040];
  assign o[57039] = i[57039];
  assign o[57038] = i[57038];
  assign o[57037] = i[57037];
  assign o[57036] = i[57036];
  assign o[57035] = i[57035];
  assign o[57034] = i[57034];
  assign o[57033] = i[57033];
  assign o[57032] = i[57032];
  assign o[57031] = i[57031];
  assign o[57030] = i[57030];
  assign o[57029] = i[57029];
  assign o[57028] = i[57028];
  assign o[57027] = i[57027];
  assign o[57026] = i[57026];
  assign o[57025] = i[57025];
  assign o[57024] = i[57024];
  assign o[57023] = i[57023];
  assign o[57022] = i[57022];
  assign o[57021] = i[57021];
  assign o[57020] = i[57020];
  assign o[57019] = i[57019];
  assign o[57018] = i[57018];
  assign o[57017] = i[57017];
  assign o[57016] = i[57016];
  assign o[57015] = i[57015];
  assign o[57014] = i[57014];
  assign o[57013] = i[57013];
  assign o[57012] = i[57012];
  assign o[57011] = i[57011];
  assign o[57010] = i[57010];
  assign o[57009] = i[57009];
  assign o[57008] = i[57008];
  assign o[57007] = i[57007];
  assign o[57006] = i[57006];
  assign o[57005] = i[57005];
  assign o[57004] = i[57004];
  assign o[57003] = i[57003];
  assign o[57002] = i[57002];
  assign o[57001] = i[57001];
  assign o[57000] = i[57000];
  assign o[56999] = i[56999];
  assign o[56998] = i[56998];
  assign o[56997] = i[56997];
  assign o[56996] = i[56996];
  assign o[56995] = i[56995];
  assign o[56994] = i[56994];
  assign o[56993] = i[56993];
  assign o[56992] = i[56992];
  assign o[56991] = i[56991];
  assign o[56990] = i[56990];
  assign o[56989] = i[56989];
  assign o[56988] = i[56988];
  assign o[56987] = i[56987];
  assign o[56986] = i[56986];
  assign o[56985] = i[56985];
  assign o[56984] = i[56984];
  assign o[56983] = i[56983];
  assign o[56982] = i[56982];
  assign o[56981] = i[56981];
  assign o[56980] = i[56980];
  assign o[56979] = i[56979];
  assign o[56978] = i[56978];
  assign o[56977] = i[56977];
  assign o[56976] = i[56976];
  assign o[56975] = i[56975];
  assign o[56974] = i[56974];
  assign o[56973] = i[56973];
  assign o[56972] = i[56972];
  assign o[56971] = i[56971];
  assign o[56970] = i[56970];
  assign o[56969] = i[56969];
  assign o[56968] = i[56968];
  assign o[56967] = i[56967];
  assign o[56966] = i[56966];
  assign o[56965] = i[56965];
  assign o[56964] = i[56964];
  assign o[56963] = i[56963];
  assign o[56962] = i[56962];
  assign o[56961] = i[56961];
  assign o[56960] = i[56960];
  assign o[56959] = i[56959];
  assign o[56958] = i[56958];
  assign o[56957] = i[56957];
  assign o[56956] = i[56956];
  assign o[56955] = i[56955];
  assign o[56954] = i[56954];
  assign o[56953] = i[56953];
  assign o[56952] = i[56952];
  assign o[56951] = i[56951];
  assign o[56950] = i[56950];
  assign o[56949] = i[56949];
  assign o[56948] = i[56948];
  assign o[56947] = i[56947];
  assign o[56946] = i[56946];
  assign o[56945] = i[56945];
  assign o[56944] = i[56944];
  assign o[56943] = i[56943];
  assign o[56942] = i[56942];
  assign o[56941] = i[56941];
  assign o[56940] = i[56940];
  assign o[56939] = i[56939];
  assign o[56938] = i[56938];
  assign o[56937] = i[56937];
  assign o[56936] = i[56936];
  assign o[56935] = i[56935];
  assign o[56934] = i[56934];
  assign o[56933] = i[56933];
  assign o[56932] = i[56932];
  assign o[56931] = i[56931];
  assign o[56930] = i[56930];
  assign o[56929] = i[56929];
  assign o[56928] = i[56928];
  assign o[56927] = i[56927];
  assign o[56926] = i[56926];
  assign o[56925] = i[56925];
  assign o[56924] = i[56924];
  assign o[56923] = i[56923];
  assign o[56922] = i[56922];
  assign o[56921] = i[56921];
  assign o[56920] = i[56920];
  assign o[56919] = i[56919];
  assign o[56918] = i[56918];
  assign o[56917] = i[56917];
  assign o[56916] = i[56916];
  assign o[56915] = i[56915];
  assign o[56914] = i[56914];
  assign o[56913] = i[56913];
  assign o[56912] = i[56912];
  assign o[56911] = i[56911];
  assign o[56910] = i[56910];
  assign o[56909] = i[56909];
  assign o[56908] = i[56908];
  assign o[56907] = i[56907];
  assign o[56906] = i[56906];
  assign o[56905] = i[56905];
  assign o[56904] = i[56904];
  assign o[56903] = i[56903];
  assign o[56902] = i[56902];
  assign o[56901] = i[56901];
  assign o[56900] = i[56900];
  assign o[56899] = i[56899];
  assign o[56898] = i[56898];
  assign o[56897] = i[56897];
  assign o[56896] = i[56896];
  assign o[56895] = i[56895];
  assign o[56894] = i[56894];
  assign o[56893] = i[56893];
  assign o[56892] = i[56892];
  assign o[56891] = i[56891];
  assign o[56890] = i[56890];
  assign o[56889] = i[56889];
  assign o[56888] = i[56888];
  assign o[56887] = i[56887];
  assign o[56886] = i[56886];
  assign o[56885] = i[56885];
  assign o[56884] = i[56884];
  assign o[56883] = i[56883];
  assign o[56882] = i[56882];
  assign o[56881] = i[56881];
  assign o[56880] = i[56880];
  assign o[56879] = i[56879];
  assign o[56878] = i[56878];
  assign o[56877] = i[56877];
  assign o[56876] = i[56876];
  assign o[56875] = i[56875];
  assign o[56874] = i[56874];
  assign o[56873] = i[56873];
  assign o[56872] = i[56872];
  assign o[56871] = i[56871];
  assign o[56870] = i[56870];
  assign o[56869] = i[56869];
  assign o[56868] = i[56868];
  assign o[56867] = i[56867];
  assign o[56866] = i[56866];
  assign o[56865] = i[56865];
  assign o[56864] = i[56864];
  assign o[56863] = i[56863];
  assign o[56862] = i[56862];
  assign o[56861] = i[56861];
  assign o[56860] = i[56860];
  assign o[56859] = i[56859];
  assign o[56858] = i[56858];
  assign o[56857] = i[56857];
  assign o[56856] = i[56856];
  assign o[56855] = i[56855];
  assign o[56854] = i[56854];
  assign o[56853] = i[56853];
  assign o[56852] = i[56852];
  assign o[56851] = i[56851];
  assign o[56850] = i[56850];
  assign o[56849] = i[56849];
  assign o[56848] = i[56848];
  assign o[56847] = i[56847];
  assign o[56846] = i[56846];
  assign o[56845] = i[56845];
  assign o[56844] = i[56844];
  assign o[56843] = i[56843];
  assign o[56842] = i[56842];
  assign o[56841] = i[56841];
  assign o[56840] = i[56840];
  assign o[56839] = i[56839];
  assign o[56838] = i[56838];
  assign o[56837] = i[56837];
  assign o[56836] = i[56836];
  assign o[56835] = i[56835];
  assign o[56834] = i[56834];
  assign o[56833] = i[56833];
  assign o[56832] = i[56832];
  assign o[56831] = i[56831];
  assign o[56830] = i[56830];
  assign o[56829] = i[56829];
  assign o[56828] = i[56828];
  assign o[56827] = i[56827];
  assign o[56826] = i[56826];
  assign o[56825] = i[56825];
  assign o[56824] = i[56824];
  assign o[56823] = i[56823];
  assign o[56822] = i[56822];
  assign o[56821] = i[56821];
  assign o[56820] = i[56820];
  assign o[56819] = i[56819];
  assign o[56818] = i[56818];
  assign o[56817] = i[56817];
  assign o[56816] = i[56816];
  assign o[56815] = i[56815];
  assign o[56814] = i[56814];
  assign o[56813] = i[56813];
  assign o[56812] = i[56812];
  assign o[56811] = i[56811];
  assign o[56810] = i[56810];
  assign o[56809] = i[56809];
  assign o[56808] = i[56808];
  assign o[56807] = i[56807];
  assign o[56806] = i[56806];
  assign o[56805] = i[56805];
  assign o[56804] = i[56804];
  assign o[56803] = i[56803];
  assign o[56802] = i[56802];
  assign o[56801] = i[56801];
  assign o[56800] = i[56800];
  assign o[56799] = i[56799];
  assign o[56798] = i[56798];
  assign o[56797] = i[56797];
  assign o[56796] = i[56796];
  assign o[56795] = i[56795];
  assign o[56794] = i[56794];
  assign o[56793] = i[56793];
  assign o[56792] = i[56792];
  assign o[56791] = i[56791];
  assign o[56790] = i[56790];
  assign o[56789] = i[56789];
  assign o[56788] = i[56788];
  assign o[56787] = i[56787];
  assign o[56786] = i[56786];
  assign o[56785] = i[56785];
  assign o[56784] = i[56784];
  assign o[56783] = i[56783];
  assign o[56782] = i[56782];
  assign o[56781] = i[56781];
  assign o[56780] = i[56780];
  assign o[56779] = i[56779];
  assign o[56778] = i[56778];
  assign o[56777] = i[56777];
  assign o[56776] = i[56776];
  assign o[56775] = i[56775];
  assign o[56774] = i[56774];
  assign o[56773] = i[56773];
  assign o[56772] = i[56772];
  assign o[56771] = i[56771];
  assign o[56770] = i[56770];
  assign o[56769] = i[56769];
  assign o[56768] = i[56768];
  assign o[56767] = i[56767];
  assign o[56766] = i[56766];
  assign o[56765] = i[56765];
  assign o[56764] = i[56764];
  assign o[56763] = i[56763];
  assign o[56762] = i[56762];
  assign o[56761] = i[56761];
  assign o[56760] = i[56760];
  assign o[56759] = i[56759];
  assign o[56758] = i[56758];
  assign o[56757] = i[56757];
  assign o[56756] = i[56756];
  assign o[56755] = i[56755];
  assign o[56754] = i[56754];
  assign o[56753] = i[56753];
  assign o[56752] = i[56752];
  assign o[56751] = i[56751];
  assign o[56750] = i[56750];
  assign o[56749] = i[56749];
  assign o[56748] = i[56748];
  assign o[56747] = i[56747];
  assign o[56746] = i[56746];
  assign o[56745] = i[56745];
  assign o[56744] = i[56744];
  assign o[56743] = i[56743];
  assign o[56742] = i[56742];
  assign o[56741] = i[56741];
  assign o[56740] = i[56740];
  assign o[56739] = i[56739];
  assign o[56738] = i[56738];
  assign o[56737] = i[56737];
  assign o[56736] = i[56736];
  assign o[56735] = i[56735];
  assign o[56734] = i[56734];
  assign o[56733] = i[56733];
  assign o[56732] = i[56732];
  assign o[56731] = i[56731];
  assign o[56730] = i[56730];
  assign o[56729] = i[56729];
  assign o[56728] = i[56728];
  assign o[56727] = i[56727];
  assign o[56726] = i[56726];
  assign o[56725] = i[56725];
  assign o[56724] = i[56724];
  assign o[56723] = i[56723];
  assign o[56722] = i[56722];
  assign o[56721] = i[56721];
  assign o[56720] = i[56720];
  assign o[56719] = i[56719];
  assign o[56718] = i[56718];
  assign o[56717] = i[56717];
  assign o[56716] = i[56716];
  assign o[56715] = i[56715];
  assign o[56714] = i[56714];
  assign o[56713] = i[56713];
  assign o[56712] = i[56712];
  assign o[56711] = i[56711];
  assign o[56710] = i[56710];
  assign o[56709] = i[56709];
  assign o[56708] = i[56708];
  assign o[56707] = i[56707];
  assign o[56706] = i[56706];
  assign o[56705] = i[56705];
  assign o[56704] = i[56704];
  assign o[56703] = i[56703];
  assign o[56702] = i[56702];
  assign o[56701] = i[56701];
  assign o[56700] = i[56700];
  assign o[56699] = i[56699];
  assign o[56698] = i[56698];
  assign o[56697] = i[56697];
  assign o[56696] = i[56696];
  assign o[56695] = i[56695];
  assign o[56694] = i[56694];
  assign o[56693] = i[56693];
  assign o[56692] = i[56692];
  assign o[56691] = i[56691];
  assign o[56690] = i[56690];
  assign o[56689] = i[56689];
  assign o[56688] = i[56688];
  assign o[56687] = i[56687];
  assign o[56686] = i[56686];
  assign o[56685] = i[56685];
  assign o[56684] = i[56684];
  assign o[56683] = i[56683];
  assign o[56682] = i[56682];
  assign o[56681] = i[56681];
  assign o[56680] = i[56680];
  assign o[56679] = i[56679];
  assign o[56678] = i[56678];
  assign o[56677] = i[56677];
  assign o[56676] = i[56676];
  assign o[56675] = i[56675];
  assign o[56674] = i[56674];
  assign o[56673] = i[56673];
  assign o[56672] = i[56672];
  assign o[56671] = i[56671];
  assign o[56670] = i[56670];
  assign o[56669] = i[56669];
  assign o[56668] = i[56668];
  assign o[56667] = i[56667];
  assign o[56666] = i[56666];
  assign o[56665] = i[56665];
  assign o[56664] = i[56664];
  assign o[56663] = i[56663];
  assign o[56662] = i[56662];
  assign o[56661] = i[56661];
  assign o[56660] = i[56660];
  assign o[56659] = i[56659];
  assign o[56658] = i[56658];
  assign o[56657] = i[56657];
  assign o[56656] = i[56656];
  assign o[56655] = i[56655];
  assign o[56654] = i[56654];
  assign o[56653] = i[56653];
  assign o[56652] = i[56652];
  assign o[56651] = i[56651];
  assign o[56650] = i[56650];
  assign o[56649] = i[56649];
  assign o[56648] = i[56648];
  assign o[56647] = i[56647];
  assign o[56646] = i[56646];
  assign o[56645] = i[56645];
  assign o[56644] = i[56644];
  assign o[56643] = i[56643];
  assign o[56642] = i[56642];
  assign o[56641] = i[56641];
  assign o[56640] = i[56640];
  assign o[56639] = i[56639];
  assign o[56638] = i[56638];
  assign o[56637] = i[56637];
  assign o[56636] = i[56636];
  assign o[56635] = i[56635];
  assign o[56634] = i[56634];
  assign o[56633] = i[56633];
  assign o[56632] = i[56632];
  assign o[56631] = i[56631];
  assign o[56630] = i[56630];
  assign o[56629] = i[56629];
  assign o[56628] = i[56628];
  assign o[56627] = i[56627];
  assign o[56626] = i[56626];
  assign o[56625] = i[56625];
  assign o[56624] = i[56624];
  assign o[56623] = i[56623];
  assign o[56622] = i[56622];
  assign o[56621] = i[56621];
  assign o[56620] = i[56620];
  assign o[56619] = i[56619];
  assign o[56618] = i[56618];
  assign o[56617] = i[56617];
  assign o[56616] = i[56616];
  assign o[56615] = i[56615];
  assign o[56614] = i[56614];
  assign o[56613] = i[56613];
  assign o[56612] = i[56612];
  assign o[56611] = i[56611];
  assign o[56610] = i[56610];
  assign o[56609] = i[56609];
  assign o[56608] = i[56608];
  assign o[56607] = i[56607];
  assign o[56606] = i[56606];
  assign o[56605] = i[56605];
  assign o[56604] = i[56604];
  assign o[56603] = i[56603];
  assign o[56602] = i[56602];
  assign o[56601] = i[56601];
  assign o[56600] = i[56600];
  assign o[56599] = i[56599];
  assign o[56598] = i[56598];
  assign o[56597] = i[56597];
  assign o[56596] = i[56596];
  assign o[56595] = i[56595];
  assign o[56594] = i[56594];
  assign o[56593] = i[56593];
  assign o[56592] = i[56592];
  assign o[56591] = i[56591];
  assign o[56590] = i[56590];
  assign o[56589] = i[56589];
  assign o[56588] = i[56588];
  assign o[56587] = i[56587];
  assign o[56586] = i[56586];
  assign o[56585] = i[56585];
  assign o[56584] = i[56584];
  assign o[56583] = i[56583];
  assign o[56582] = i[56582];
  assign o[56581] = i[56581];
  assign o[56580] = i[56580];
  assign o[56579] = i[56579];
  assign o[56578] = i[56578];
  assign o[56577] = i[56577];
  assign o[56576] = i[56576];
  assign o[56575] = i[56575];
  assign o[56574] = i[56574];
  assign o[56573] = i[56573];
  assign o[56572] = i[56572];
  assign o[56571] = i[56571];
  assign o[56570] = i[56570];
  assign o[56569] = i[56569];
  assign o[56568] = i[56568];
  assign o[56567] = i[56567];
  assign o[56566] = i[56566];
  assign o[56565] = i[56565];
  assign o[56564] = i[56564];
  assign o[56563] = i[56563];
  assign o[56562] = i[56562];
  assign o[56561] = i[56561];
  assign o[56560] = i[56560];
  assign o[56559] = i[56559];
  assign o[56558] = i[56558];
  assign o[56557] = i[56557];
  assign o[56556] = i[56556];
  assign o[56555] = i[56555];
  assign o[56554] = i[56554];
  assign o[56553] = i[56553];
  assign o[56552] = i[56552];
  assign o[56551] = i[56551];
  assign o[56550] = i[56550];
  assign o[56549] = i[56549];
  assign o[56548] = i[56548];
  assign o[56547] = i[56547];
  assign o[56546] = i[56546];
  assign o[56545] = i[56545];
  assign o[56544] = i[56544];
  assign o[56543] = i[56543];
  assign o[56542] = i[56542];
  assign o[56541] = i[56541];
  assign o[56540] = i[56540];
  assign o[56539] = i[56539];
  assign o[56538] = i[56538];
  assign o[56537] = i[56537];
  assign o[56536] = i[56536];
  assign o[56535] = i[56535];
  assign o[56534] = i[56534];
  assign o[56533] = i[56533];
  assign o[56532] = i[56532];
  assign o[56531] = i[56531];
  assign o[56530] = i[56530];
  assign o[56529] = i[56529];
  assign o[56528] = i[56528];
  assign o[56527] = i[56527];
  assign o[56526] = i[56526];
  assign o[56525] = i[56525];
  assign o[56524] = i[56524];
  assign o[56523] = i[56523];
  assign o[56522] = i[56522];
  assign o[56521] = i[56521];
  assign o[56520] = i[56520];
  assign o[56519] = i[56519];
  assign o[56518] = i[56518];
  assign o[56517] = i[56517];
  assign o[56516] = i[56516];
  assign o[56515] = i[56515];
  assign o[56514] = i[56514];
  assign o[56513] = i[56513];
  assign o[56512] = i[56512];
  assign o[56511] = i[56511];
  assign o[56510] = i[56510];
  assign o[56509] = i[56509];
  assign o[56508] = i[56508];
  assign o[56507] = i[56507];
  assign o[56506] = i[56506];
  assign o[56505] = i[56505];
  assign o[56504] = i[56504];
  assign o[56503] = i[56503];
  assign o[56502] = i[56502];
  assign o[56501] = i[56501];
  assign o[56500] = i[56500];
  assign o[56499] = i[56499];
  assign o[56498] = i[56498];
  assign o[56497] = i[56497];
  assign o[56496] = i[56496];
  assign o[56495] = i[56495];
  assign o[56494] = i[56494];
  assign o[56493] = i[56493];
  assign o[56492] = i[56492];
  assign o[56491] = i[56491];
  assign o[56490] = i[56490];
  assign o[56489] = i[56489];
  assign o[56488] = i[56488];
  assign o[56487] = i[56487];
  assign o[56486] = i[56486];
  assign o[56485] = i[56485];
  assign o[56484] = i[56484];
  assign o[56483] = i[56483];
  assign o[56482] = i[56482];
  assign o[56481] = i[56481];
  assign o[56480] = i[56480];
  assign o[56479] = i[56479];
  assign o[56478] = i[56478];
  assign o[56477] = i[56477];
  assign o[56476] = i[56476];
  assign o[56475] = i[56475];
  assign o[56474] = i[56474];
  assign o[56473] = i[56473];
  assign o[56472] = i[56472];
  assign o[56471] = i[56471];
  assign o[56470] = i[56470];
  assign o[56469] = i[56469];
  assign o[56468] = i[56468];
  assign o[56467] = i[56467];
  assign o[56466] = i[56466];
  assign o[56465] = i[56465];
  assign o[56464] = i[56464];
  assign o[56463] = i[56463];
  assign o[56462] = i[56462];
  assign o[56461] = i[56461];
  assign o[56460] = i[56460];
  assign o[56459] = i[56459];
  assign o[56458] = i[56458];
  assign o[56457] = i[56457];
  assign o[56456] = i[56456];
  assign o[56455] = i[56455];
  assign o[56454] = i[56454];
  assign o[56453] = i[56453];
  assign o[56452] = i[56452];
  assign o[56451] = i[56451];
  assign o[56450] = i[56450];
  assign o[56449] = i[56449];
  assign o[56448] = i[56448];
  assign o[56447] = i[56447];
  assign o[56446] = i[56446];
  assign o[56445] = i[56445];
  assign o[56444] = i[56444];
  assign o[56443] = i[56443];
  assign o[56442] = i[56442];
  assign o[56441] = i[56441];
  assign o[56440] = i[56440];
  assign o[56439] = i[56439];
  assign o[56438] = i[56438];
  assign o[56437] = i[56437];
  assign o[56436] = i[56436];
  assign o[56435] = i[56435];
  assign o[56434] = i[56434];
  assign o[56433] = i[56433];
  assign o[56432] = i[56432];
  assign o[56431] = i[56431];
  assign o[56430] = i[56430];
  assign o[56429] = i[56429];
  assign o[56428] = i[56428];
  assign o[56427] = i[56427];
  assign o[56426] = i[56426];
  assign o[56425] = i[56425];
  assign o[56424] = i[56424];
  assign o[56423] = i[56423];
  assign o[56422] = i[56422];
  assign o[56421] = i[56421];
  assign o[56420] = i[56420];
  assign o[56419] = i[56419];
  assign o[56418] = i[56418];
  assign o[56417] = i[56417];
  assign o[56416] = i[56416];
  assign o[56415] = i[56415];
  assign o[56414] = i[56414];
  assign o[56413] = i[56413];
  assign o[56412] = i[56412];
  assign o[56411] = i[56411];
  assign o[56410] = i[56410];
  assign o[56409] = i[56409];
  assign o[56408] = i[56408];
  assign o[56407] = i[56407];
  assign o[56406] = i[56406];
  assign o[56405] = i[56405];
  assign o[56404] = i[56404];
  assign o[56403] = i[56403];
  assign o[56402] = i[56402];
  assign o[56401] = i[56401];
  assign o[56400] = i[56400];
  assign o[56399] = i[56399];
  assign o[56398] = i[56398];
  assign o[56397] = i[56397];
  assign o[56396] = i[56396];
  assign o[56395] = i[56395];
  assign o[56394] = i[56394];
  assign o[56393] = i[56393];
  assign o[56392] = i[56392];
  assign o[56391] = i[56391];
  assign o[56390] = i[56390];
  assign o[56389] = i[56389];
  assign o[56388] = i[56388];
  assign o[56387] = i[56387];
  assign o[56386] = i[56386];
  assign o[56385] = i[56385];
  assign o[56384] = i[56384];
  assign o[56383] = i[56383];
  assign o[56382] = i[56382];
  assign o[56381] = i[56381];
  assign o[56380] = i[56380];
  assign o[56379] = i[56379];
  assign o[56378] = i[56378];
  assign o[56377] = i[56377];
  assign o[56376] = i[56376];
  assign o[56375] = i[56375];
  assign o[56374] = i[56374];
  assign o[56373] = i[56373];
  assign o[56372] = i[56372];
  assign o[56371] = i[56371];
  assign o[56370] = i[56370];
  assign o[56369] = i[56369];
  assign o[56368] = i[56368];
  assign o[56367] = i[56367];
  assign o[56366] = i[56366];
  assign o[56365] = i[56365];
  assign o[56364] = i[56364];
  assign o[56363] = i[56363];
  assign o[56362] = i[56362];
  assign o[56361] = i[56361];
  assign o[56360] = i[56360];
  assign o[56359] = i[56359];
  assign o[56358] = i[56358];
  assign o[56357] = i[56357];
  assign o[56356] = i[56356];
  assign o[56355] = i[56355];
  assign o[56354] = i[56354];
  assign o[56353] = i[56353];
  assign o[56352] = i[56352];
  assign o[56351] = i[56351];
  assign o[56350] = i[56350];
  assign o[56349] = i[56349];
  assign o[56348] = i[56348];
  assign o[56347] = i[56347];
  assign o[56346] = i[56346];
  assign o[56345] = i[56345];
  assign o[56344] = i[56344];
  assign o[56343] = i[56343];
  assign o[56342] = i[56342];
  assign o[56341] = i[56341];
  assign o[56340] = i[56340];
  assign o[56339] = i[56339];
  assign o[56338] = i[56338];
  assign o[56337] = i[56337];
  assign o[56336] = i[56336];
  assign o[56335] = i[56335];
  assign o[56334] = i[56334];
  assign o[56333] = i[56333];
  assign o[56332] = i[56332];
  assign o[56331] = i[56331];
  assign o[56330] = i[56330];
  assign o[56329] = i[56329];
  assign o[56328] = i[56328];
  assign o[56327] = i[56327];
  assign o[56326] = i[56326];
  assign o[56325] = i[56325];
  assign o[56324] = i[56324];
  assign o[56323] = i[56323];
  assign o[56322] = i[56322];
  assign o[56321] = i[56321];
  assign o[56320] = i[56320];
  assign o[56319] = i[56319];
  assign o[56318] = i[56318];
  assign o[56317] = i[56317];
  assign o[56316] = i[56316];
  assign o[56315] = i[56315];
  assign o[56314] = i[56314];
  assign o[56313] = i[56313];
  assign o[56312] = i[56312];
  assign o[56311] = i[56311];
  assign o[56310] = i[56310];
  assign o[56309] = i[56309];
  assign o[56308] = i[56308];
  assign o[56307] = i[56307];
  assign o[56306] = i[56306];
  assign o[56305] = i[56305];
  assign o[56304] = i[56304];
  assign o[56303] = i[56303];
  assign o[56302] = i[56302];
  assign o[56301] = i[56301];
  assign o[56300] = i[56300];
  assign o[56299] = i[56299];
  assign o[56298] = i[56298];
  assign o[56297] = i[56297];
  assign o[56296] = i[56296];
  assign o[56295] = i[56295];
  assign o[56294] = i[56294];
  assign o[56293] = i[56293];
  assign o[56292] = i[56292];
  assign o[56291] = i[56291];
  assign o[56290] = i[56290];
  assign o[56289] = i[56289];
  assign o[56288] = i[56288];
  assign o[56287] = i[56287];
  assign o[56286] = i[56286];
  assign o[56285] = i[56285];
  assign o[56284] = i[56284];
  assign o[56283] = i[56283];
  assign o[56282] = i[56282];
  assign o[56281] = i[56281];
  assign o[56280] = i[56280];
  assign o[56279] = i[56279];
  assign o[56278] = i[56278];
  assign o[56277] = i[56277];
  assign o[56276] = i[56276];
  assign o[56275] = i[56275];
  assign o[56274] = i[56274];
  assign o[56273] = i[56273];
  assign o[56272] = i[56272];
  assign o[56271] = i[56271];
  assign o[56270] = i[56270];
  assign o[56269] = i[56269];
  assign o[56268] = i[56268];
  assign o[56267] = i[56267];
  assign o[56266] = i[56266];
  assign o[56265] = i[56265];
  assign o[56264] = i[56264];
  assign o[56263] = i[56263];
  assign o[56262] = i[56262];
  assign o[56261] = i[56261];
  assign o[56260] = i[56260];
  assign o[56259] = i[56259];
  assign o[56258] = i[56258];
  assign o[56257] = i[56257];
  assign o[56256] = i[56256];
  assign o[56255] = i[56255];
  assign o[56254] = i[56254];
  assign o[56253] = i[56253];
  assign o[56252] = i[56252];
  assign o[56251] = i[56251];
  assign o[56250] = i[56250];
  assign o[56249] = i[56249];
  assign o[56248] = i[56248];
  assign o[56247] = i[56247];
  assign o[56246] = i[56246];
  assign o[56245] = i[56245];
  assign o[56244] = i[56244];
  assign o[56243] = i[56243];
  assign o[56242] = i[56242];
  assign o[56241] = i[56241];
  assign o[56240] = i[56240];
  assign o[56239] = i[56239];
  assign o[56238] = i[56238];
  assign o[56237] = i[56237];
  assign o[56236] = i[56236];
  assign o[56235] = i[56235];
  assign o[56234] = i[56234];
  assign o[56233] = i[56233];
  assign o[56232] = i[56232];
  assign o[56231] = i[56231];
  assign o[56230] = i[56230];
  assign o[56229] = i[56229];
  assign o[56228] = i[56228];
  assign o[56227] = i[56227];
  assign o[56226] = i[56226];
  assign o[56225] = i[56225];
  assign o[56224] = i[56224];
  assign o[56223] = i[56223];
  assign o[56222] = i[56222];
  assign o[56221] = i[56221];
  assign o[56220] = i[56220];
  assign o[56219] = i[56219];
  assign o[56218] = i[56218];
  assign o[56217] = i[56217];
  assign o[56216] = i[56216];
  assign o[56215] = i[56215];
  assign o[56214] = i[56214];
  assign o[56213] = i[56213];
  assign o[56212] = i[56212];
  assign o[56211] = i[56211];
  assign o[56210] = i[56210];
  assign o[56209] = i[56209];
  assign o[56208] = i[56208];
  assign o[56207] = i[56207];
  assign o[56206] = i[56206];
  assign o[56205] = i[56205];
  assign o[56204] = i[56204];
  assign o[56203] = i[56203];
  assign o[56202] = i[56202];
  assign o[56201] = i[56201];
  assign o[56200] = i[56200];
  assign o[56199] = i[56199];
  assign o[56198] = i[56198];
  assign o[56197] = i[56197];
  assign o[56196] = i[56196];
  assign o[56195] = i[56195];
  assign o[56194] = i[56194];
  assign o[56193] = i[56193];
  assign o[56192] = i[56192];
  assign o[56191] = i[56191];
  assign o[56190] = i[56190];
  assign o[56189] = i[56189];
  assign o[56188] = i[56188];
  assign o[56187] = i[56187];
  assign o[56186] = i[56186];
  assign o[56185] = i[56185];
  assign o[56184] = i[56184];
  assign o[56183] = i[56183];
  assign o[56182] = i[56182];
  assign o[56181] = i[56181];
  assign o[56180] = i[56180];
  assign o[56179] = i[56179];
  assign o[56178] = i[56178];
  assign o[56177] = i[56177];
  assign o[56176] = i[56176];
  assign o[56175] = i[56175];
  assign o[56174] = i[56174];
  assign o[56173] = i[56173];
  assign o[56172] = i[56172];
  assign o[56171] = i[56171];
  assign o[56170] = i[56170];
  assign o[56169] = i[56169];
  assign o[56168] = i[56168];
  assign o[56167] = i[56167];
  assign o[56166] = i[56166];
  assign o[56165] = i[56165];
  assign o[56164] = i[56164];
  assign o[56163] = i[56163];
  assign o[56162] = i[56162];
  assign o[56161] = i[56161];
  assign o[56160] = i[56160];
  assign o[56159] = i[56159];
  assign o[56158] = i[56158];
  assign o[56157] = i[56157];
  assign o[56156] = i[56156];
  assign o[56155] = i[56155];
  assign o[56154] = i[56154];
  assign o[56153] = i[56153];
  assign o[56152] = i[56152];
  assign o[56151] = i[56151];
  assign o[56150] = i[56150];
  assign o[56149] = i[56149];
  assign o[56148] = i[56148];
  assign o[56147] = i[56147];
  assign o[56146] = i[56146];
  assign o[56145] = i[56145];
  assign o[56144] = i[56144];
  assign o[56143] = i[56143];
  assign o[56142] = i[56142];
  assign o[56141] = i[56141];
  assign o[56140] = i[56140];
  assign o[56139] = i[56139];
  assign o[56138] = i[56138];
  assign o[56137] = i[56137];
  assign o[56136] = i[56136];
  assign o[56135] = i[56135];
  assign o[56134] = i[56134];
  assign o[56133] = i[56133];
  assign o[56132] = i[56132];
  assign o[56131] = i[56131];
  assign o[56130] = i[56130];
  assign o[56129] = i[56129];
  assign o[56128] = i[56128];
  assign o[56127] = i[56127];
  assign o[56126] = i[56126];
  assign o[56125] = i[56125];
  assign o[56124] = i[56124];
  assign o[56123] = i[56123];
  assign o[56122] = i[56122];
  assign o[56121] = i[56121];
  assign o[56120] = i[56120];
  assign o[56119] = i[56119];
  assign o[56118] = i[56118];
  assign o[56117] = i[56117];
  assign o[56116] = i[56116];
  assign o[56115] = i[56115];
  assign o[56114] = i[56114];
  assign o[56113] = i[56113];
  assign o[56112] = i[56112];
  assign o[56111] = i[56111];
  assign o[56110] = i[56110];
  assign o[56109] = i[56109];
  assign o[56108] = i[56108];
  assign o[56107] = i[56107];
  assign o[56106] = i[56106];
  assign o[56105] = i[56105];
  assign o[56104] = i[56104];
  assign o[56103] = i[56103];
  assign o[56102] = i[56102];
  assign o[56101] = i[56101];
  assign o[56100] = i[56100];
  assign o[56099] = i[56099];
  assign o[56098] = i[56098];
  assign o[56097] = i[56097];
  assign o[56096] = i[56096];
  assign o[56095] = i[56095];
  assign o[56094] = i[56094];
  assign o[56093] = i[56093];
  assign o[56092] = i[56092];
  assign o[56091] = i[56091];
  assign o[56090] = i[56090];
  assign o[56089] = i[56089];
  assign o[56088] = i[56088];
  assign o[56087] = i[56087];
  assign o[56086] = i[56086];
  assign o[56085] = i[56085];
  assign o[56084] = i[56084];
  assign o[56083] = i[56083];
  assign o[56082] = i[56082];
  assign o[56081] = i[56081];
  assign o[56080] = i[56080];
  assign o[56079] = i[56079];
  assign o[56078] = i[56078];
  assign o[56077] = i[56077];
  assign o[56076] = i[56076];
  assign o[56075] = i[56075];
  assign o[56074] = i[56074];
  assign o[56073] = i[56073];
  assign o[56072] = i[56072];
  assign o[56071] = i[56071];
  assign o[56070] = i[56070];
  assign o[56069] = i[56069];
  assign o[56068] = i[56068];
  assign o[56067] = i[56067];
  assign o[56066] = i[56066];
  assign o[56065] = i[56065];
  assign o[56064] = i[56064];
  assign o[56063] = i[56063];
  assign o[56062] = i[56062];
  assign o[56061] = i[56061];
  assign o[56060] = i[56060];
  assign o[56059] = i[56059];
  assign o[56058] = i[56058];
  assign o[56057] = i[56057];
  assign o[56056] = i[56056];
  assign o[56055] = i[56055];
  assign o[56054] = i[56054];
  assign o[56053] = i[56053];
  assign o[56052] = i[56052];
  assign o[56051] = i[56051];
  assign o[56050] = i[56050];
  assign o[56049] = i[56049];
  assign o[56048] = i[56048];
  assign o[56047] = i[56047];
  assign o[56046] = i[56046];
  assign o[56045] = i[56045];
  assign o[56044] = i[56044];
  assign o[56043] = i[56043];
  assign o[56042] = i[56042];
  assign o[56041] = i[56041];
  assign o[56040] = i[56040];
  assign o[56039] = i[56039];
  assign o[56038] = i[56038];
  assign o[56037] = i[56037];
  assign o[56036] = i[56036];
  assign o[56035] = i[56035];
  assign o[56034] = i[56034];
  assign o[56033] = i[56033];
  assign o[56032] = i[56032];
  assign o[56031] = i[56031];
  assign o[56030] = i[56030];
  assign o[56029] = i[56029];
  assign o[56028] = i[56028];
  assign o[56027] = i[56027];
  assign o[56026] = i[56026];
  assign o[56025] = i[56025];
  assign o[56024] = i[56024];
  assign o[56023] = i[56023];
  assign o[56022] = i[56022];
  assign o[56021] = i[56021];
  assign o[56020] = i[56020];
  assign o[56019] = i[56019];
  assign o[56018] = i[56018];
  assign o[56017] = i[56017];
  assign o[56016] = i[56016];
  assign o[56015] = i[56015];
  assign o[56014] = i[56014];
  assign o[56013] = i[56013];
  assign o[56012] = i[56012];
  assign o[56011] = i[56011];
  assign o[56010] = i[56010];
  assign o[56009] = i[56009];
  assign o[56008] = i[56008];
  assign o[56007] = i[56007];
  assign o[56006] = i[56006];
  assign o[56005] = i[56005];
  assign o[56004] = i[56004];
  assign o[56003] = i[56003];
  assign o[56002] = i[56002];
  assign o[56001] = i[56001];
  assign o[56000] = i[56000];
  assign o[55999] = i[55999];
  assign o[55998] = i[55998];
  assign o[55997] = i[55997];
  assign o[55996] = i[55996];
  assign o[55995] = i[55995];
  assign o[55994] = i[55994];
  assign o[55993] = i[55993];
  assign o[55992] = i[55992];
  assign o[55991] = i[55991];
  assign o[55990] = i[55990];
  assign o[55989] = i[55989];
  assign o[55988] = i[55988];
  assign o[55987] = i[55987];
  assign o[55986] = i[55986];
  assign o[55985] = i[55985];
  assign o[55984] = i[55984];
  assign o[55983] = i[55983];
  assign o[55982] = i[55982];
  assign o[55981] = i[55981];
  assign o[55980] = i[55980];
  assign o[55979] = i[55979];
  assign o[55978] = i[55978];
  assign o[55977] = i[55977];
  assign o[55976] = i[55976];
  assign o[55975] = i[55975];
  assign o[55974] = i[55974];
  assign o[55973] = i[55973];
  assign o[55972] = i[55972];
  assign o[55971] = i[55971];
  assign o[55970] = i[55970];
  assign o[55969] = i[55969];
  assign o[55968] = i[55968];
  assign o[55967] = i[55967];
  assign o[55966] = i[55966];
  assign o[55965] = i[55965];
  assign o[55964] = i[55964];
  assign o[55963] = i[55963];
  assign o[55962] = i[55962];
  assign o[55961] = i[55961];
  assign o[55960] = i[55960];
  assign o[55959] = i[55959];
  assign o[55958] = i[55958];
  assign o[55957] = i[55957];
  assign o[55956] = i[55956];
  assign o[55955] = i[55955];
  assign o[55954] = i[55954];
  assign o[55953] = i[55953];
  assign o[55952] = i[55952];
  assign o[55951] = i[55951];
  assign o[55950] = i[55950];
  assign o[55949] = i[55949];
  assign o[55948] = i[55948];
  assign o[55947] = i[55947];
  assign o[55946] = i[55946];
  assign o[55945] = i[55945];
  assign o[55944] = i[55944];
  assign o[55943] = i[55943];
  assign o[55942] = i[55942];
  assign o[55941] = i[55941];
  assign o[55940] = i[55940];
  assign o[55939] = i[55939];
  assign o[55938] = i[55938];
  assign o[55937] = i[55937];
  assign o[55936] = i[55936];
  assign o[55935] = i[55935];
  assign o[55934] = i[55934];
  assign o[55933] = i[55933];
  assign o[55932] = i[55932];
  assign o[55931] = i[55931];
  assign o[55930] = i[55930];
  assign o[55929] = i[55929];
  assign o[55928] = i[55928];
  assign o[55927] = i[55927];
  assign o[55926] = i[55926];
  assign o[55925] = i[55925];
  assign o[55924] = i[55924];
  assign o[55923] = i[55923];
  assign o[55922] = i[55922];
  assign o[55921] = i[55921];
  assign o[55920] = i[55920];
  assign o[55919] = i[55919];
  assign o[55918] = i[55918];
  assign o[55917] = i[55917];
  assign o[55916] = i[55916];
  assign o[55915] = i[55915];
  assign o[55914] = i[55914];
  assign o[55913] = i[55913];
  assign o[55912] = i[55912];
  assign o[55911] = i[55911];
  assign o[55910] = i[55910];
  assign o[55909] = i[55909];
  assign o[55908] = i[55908];
  assign o[55907] = i[55907];
  assign o[55906] = i[55906];
  assign o[55905] = i[55905];
  assign o[55904] = i[55904];
  assign o[55903] = i[55903];
  assign o[55902] = i[55902];
  assign o[55901] = i[55901];
  assign o[55900] = i[55900];
  assign o[55899] = i[55899];
  assign o[55898] = i[55898];
  assign o[55897] = i[55897];
  assign o[55896] = i[55896];
  assign o[55895] = i[55895];
  assign o[55894] = i[55894];
  assign o[55893] = i[55893];
  assign o[55892] = i[55892];
  assign o[55891] = i[55891];
  assign o[55890] = i[55890];
  assign o[55889] = i[55889];
  assign o[55888] = i[55888];
  assign o[55887] = i[55887];
  assign o[55886] = i[55886];
  assign o[55885] = i[55885];
  assign o[55884] = i[55884];
  assign o[55883] = i[55883];
  assign o[55882] = i[55882];
  assign o[55881] = i[55881];
  assign o[55880] = i[55880];
  assign o[55879] = i[55879];
  assign o[55878] = i[55878];
  assign o[55877] = i[55877];
  assign o[55876] = i[55876];
  assign o[55875] = i[55875];
  assign o[55874] = i[55874];
  assign o[55873] = i[55873];
  assign o[55872] = i[55872];
  assign o[55871] = i[55871];
  assign o[55870] = i[55870];
  assign o[55869] = i[55869];
  assign o[55868] = i[55868];
  assign o[55867] = i[55867];
  assign o[55866] = i[55866];
  assign o[55865] = i[55865];
  assign o[55864] = i[55864];
  assign o[55863] = i[55863];
  assign o[55862] = i[55862];
  assign o[55861] = i[55861];
  assign o[55860] = i[55860];
  assign o[55859] = i[55859];
  assign o[55858] = i[55858];
  assign o[55857] = i[55857];
  assign o[55856] = i[55856];
  assign o[55855] = i[55855];
  assign o[55854] = i[55854];
  assign o[55853] = i[55853];
  assign o[55852] = i[55852];
  assign o[55851] = i[55851];
  assign o[55850] = i[55850];
  assign o[55849] = i[55849];
  assign o[55848] = i[55848];
  assign o[55847] = i[55847];
  assign o[55846] = i[55846];
  assign o[55845] = i[55845];
  assign o[55844] = i[55844];
  assign o[55843] = i[55843];
  assign o[55842] = i[55842];
  assign o[55841] = i[55841];
  assign o[55840] = i[55840];
  assign o[55839] = i[55839];
  assign o[55838] = i[55838];
  assign o[55837] = i[55837];
  assign o[55836] = i[55836];
  assign o[55835] = i[55835];
  assign o[55834] = i[55834];
  assign o[55833] = i[55833];
  assign o[55832] = i[55832];
  assign o[55831] = i[55831];
  assign o[55830] = i[55830];
  assign o[55829] = i[55829];
  assign o[55828] = i[55828];
  assign o[55827] = i[55827];
  assign o[55826] = i[55826];
  assign o[55825] = i[55825];
  assign o[55824] = i[55824];
  assign o[55823] = i[55823];
  assign o[55822] = i[55822];
  assign o[55821] = i[55821];
  assign o[55820] = i[55820];
  assign o[55819] = i[55819];
  assign o[55818] = i[55818];
  assign o[55817] = i[55817];
  assign o[55816] = i[55816];
  assign o[55815] = i[55815];
  assign o[55814] = i[55814];
  assign o[55813] = i[55813];
  assign o[55812] = i[55812];
  assign o[55811] = i[55811];
  assign o[55810] = i[55810];
  assign o[55809] = i[55809];
  assign o[55808] = i[55808];
  assign o[55807] = i[55807];
  assign o[55806] = i[55806];
  assign o[55805] = i[55805];
  assign o[55804] = i[55804];
  assign o[55803] = i[55803];
  assign o[55802] = i[55802];
  assign o[55801] = i[55801];
  assign o[55800] = i[55800];
  assign o[55799] = i[55799];
  assign o[55798] = i[55798];
  assign o[55797] = i[55797];
  assign o[55796] = i[55796];
  assign o[55795] = i[55795];
  assign o[55794] = i[55794];
  assign o[55793] = i[55793];
  assign o[55792] = i[55792];
  assign o[55791] = i[55791];
  assign o[55790] = i[55790];
  assign o[55789] = i[55789];
  assign o[55788] = i[55788];
  assign o[55787] = i[55787];
  assign o[55786] = i[55786];
  assign o[55785] = i[55785];
  assign o[55784] = i[55784];
  assign o[55783] = i[55783];
  assign o[55782] = i[55782];
  assign o[55781] = i[55781];
  assign o[55780] = i[55780];
  assign o[55779] = i[55779];
  assign o[55778] = i[55778];
  assign o[55777] = i[55777];
  assign o[55776] = i[55776];
  assign o[55775] = i[55775];
  assign o[55774] = i[55774];
  assign o[55773] = i[55773];
  assign o[55772] = i[55772];
  assign o[55771] = i[55771];
  assign o[55770] = i[55770];
  assign o[55769] = i[55769];
  assign o[55768] = i[55768];
  assign o[55767] = i[55767];
  assign o[55766] = i[55766];
  assign o[55765] = i[55765];
  assign o[55764] = i[55764];
  assign o[55763] = i[55763];
  assign o[55762] = i[55762];
  assign o[55761] = i[55761];
  assign o[55760] = i[55760];
  assign o[55759] = i[55759];
  assign o[55758] = i[55758];
  assign o[55757] = i[55757];
  assign o[55756] = i[55756];
  assign o[55755] = i[55755];
  assign o[55754] = i[55754];
  assign o[55753] = i[55753];
  assign o[55752] = i[55752];
  assign o[55751] = i[55751];
  assign o[55750] = i[55750];
  assign o[55749] = i[55749];
  assign o[55748] = i[55748];
  assign o[55747] = i[55747];
  assign o[55746] = i[55746];
  assign o[55745] = i[55745];
  assign o[55744] = i[55744];
  assign o[55743] = i[55743];
  assign o[55742] = i[55742];
  assign o[55741] = i[55741];
  assign o[55740] = i[55740];
  assign o[55739] = i[55739];
  assign o[55738] = i[55738];
  assign o[55737] = i[55737];
  assign o[55736] = i[55736];
  assign o[55735] = i[55735];
  assign o[55734] = i[55734];
  assign o[55733] = i[55733];
  assign o[55732] = i[55732];
  assign o[55731] = i[55731];
  assign o[55730] = i[55730];
  assign o[55729] = i[55729];
  assign o[55728] = i[55728];
  assign o[55727] = i[55727];
  assign o[55726] = i[55726];
  assign o[55725] = i[55725];
  assign o[55724] = i[55724];
  assign o[55723] = i[55723];
  assign o[55722] = i[55722];
  assign o[55721] = i[55721];
  assign o[55720] = i[55720];
  assign o[55719] = i[55719];
  assign o[55718] = i[55718];
  assign o[55717] = i[55717];
  assign o[55716] = i[55716];
  assign o[55715] = i[55715];
  assign o[55714] = i[55714];
  assign o[55713] = i[55713];
  assign o[55712] = i[55712];
  assign o[55711] = i[55711];
  assign o[55710] = i[55710];
  assign o[55709] = i[55709];
  assign o[55708] = i[55708];
  assign o[55707] = i[55707];
  assign o[55706] = i[55706];
  assign o[55705] = i[55705];
  assign o[55704] = i[55704];
  assign o[55703] = i[55703];
  assign o[55702] = i[55702];
  assign o[55701] = i[55701];
  assign o[55700] = i[55700];
  assign o[55699] = i[55699];
  assign o[55698] = i[55698];
  assign o[55697] = i[55697];
  assign o[55696] = i[55696];
  assign o[55695] = i[55695];
  assign o[55694] = i[55694];
  assign o[55693] = i[55693];
  assign o[55692] = i[55692];
  assign o[55691] = i[55691];
  assign o[55690] = i[55690];
  assign o[55689] = i[55689];
  assign o[55688] = i[55688];
  assign o[55687] = i[55687];
  assign o[55686] = i[55686];
  assign o[55685] = i[55685];
  assign o[55684] = i[55684];
  assign o[55683] = i[55683];
  assign o[55682] = i[55682];
  assign o[55681] = i[55681];
  assign o[55680] = i[55680];
  assign o[55679] = i[55679];
  assign o[55678] = i[55678];
  assign o[55677] = i[55677];
  assign o[55676] = i[55676];
  assign o[55675] = i[55675];
  assign o[55674] = i[55674];
  assign o[55673] = i[55673];
  assign o[55672] = i[55672];
  assign o[55671] = i[55671];
  assign o[55670] = i[55670];
  assign o[55669] = i[55669];
  assign o[55668] = i[55668];
  assign o[55667] = i[55667];
  assign o[55666] = i[55666];
  assign o[55665] = i[55665];
  assign o[55664] = i[55664];
  assign o[55663] = i[55663];
  assign o[55662] = i[55662];
  assign o[55661] = i[55661];
  assign o[55660] = i[55660];
  assign o[55659] = i[55659];
  assign o[55658] = i[55658];
  assign o[55657] = i[55657];
  assign o[55656] = i[55656];
  assign o[55655] = i[55655];
  assign o[55654] = i[55654];
  assign o[55653] = i[55653];
  assign o[55652] = i[55652];
  assign o[55651] = i[55651];
  assign o[55650] = i[55650];
  assign o[55649] = i[55649];
  assign o[55648] = i[55648];
  assign o[55647] = i[55647];
  assign o[55646] = i[55646];
  assign o[55645] = i[55645];
  assign o[55644] = i[55644];
  assign o[55643] = i[55643];
  assign o[55642] = i[55642];
  assign o[55641] = i[55641];
  assign o[55640] = i[55640];
  assign o[55639] = i[55639];
  assign o[55638] = i[55638];
  assign o[55637] = i[55637];
  assign o[55636] = i[55636];
  assign o[55635] = i[55635];
  assign o[55634] = i[55634];
  assign o[55633] = i[55633];
  assign o[55632] = i[55632];
  assign o[55631] = i[55631];
  assign o[55630] = i[55630];
  assign o[55629] = i[55629];
  assign o[55628] = i[55628];
  assign o[55627] = i[55627];
  assign o[55626] = i[55626];
  assign o[55625] = i[55625];
  assign o[55624] = i[55624];
  assign o[55623] = i[55623];
  assign o[55622] = i[55622];
  assign o[55621] = i[55621];
  assign o[55620] = i[55620];
  assign o[55619] = i[55619];
  assign o[55618] = i[55618];
  assign o[55617] = i[55617];
  assign o[55616] = i[55616];
  assign o[55615] = i[55615];
  assign o[55614] = i[55614];
  assign o[55613] = i[55613];
  assign o[55612] = i[55612];
  assign o[55611] = i[55611];
  assign o[55610] = i[55610];
  assign o[55609] = i[55609];
  assign o[55608] = i[55608];
  assign o[55607] = i[55607];
  assign o[55606] = i[55606];
  assign o[55605] = i[55605];
  assign o[55604] = i[55604];
  assign o[55603] = i[55603];
  assign o[55602] = i[55602];
  assign o[55601] = i[55601];
  assign o[55600] = i[55600];
  assign o[55599] = i[55599];
  assign o[55598] = i[55598];
  assign o[55597] = i[55597];
  assign o[55596] = i[55596];
  assign o[55595] = i[55595];
  assign o[55594] = i[55594];
  assign o[55593] = i[55593];
  assign o[55592] = i[55592];
  assign o[55591] = i[55591];
  assign o[55590] = i[55590];
  assign o[55589] = i[55589];
  assign o[55588] = i[55588];
  assign o[55587] = i[55587];
  assign o[55586] = i[55586];
  assign o[55585] = i[55585];
  assign o[55584] = i[55584];
  assign o[55583] = i[55583];
  assign o[55582] = i[55582];
  assign o[55581] = i[55581];
  assign o[55580] = i[55580];
  assign o[55579] = i[55579];
  assign o[55578] = i[55578];
  assign o[55577] = i[55577];
  assign o[55576] = i[55576];
  assign o[55575] = i[55575];
  assign o[55574] = i[55574];
  assign o[55573] = i[55573];
  assign o[55572] = i[55572];
  assign o[55571] = i[55571];
  assign o[55570] = i[55570];
  assign o[55569] = i[55569];
  assign o[55568] = i[55568];
  assign o[55567] = i[55567];
  assign o[55566] = i[55566];
  assign o[55565] = i[55565];
  assign o[55564] = i[55564];
  assign o[55563] = i[55563];
  assign o[55562] = i[55562];
  assign o[55561] = i[55561];
  assign o[55560] = i[55560];
  assign o[55559] = i[55559];
  assign o[55558] = i[55558];
  assign o[55557] = i[55557];
  assign o[55556] = i[55556];
  assign o[55555] = i[55555];
  assign o[55554] = i[55554];
  assign o[55553] = i[55553];
  assign o[55552] = i[55552];
  assign o[55551] = i[55551];
  assign o[55550] = i[55550];
  assign o[55549] = i[55549];
  assign o[55548] = i[55548];
  assign o[55547] = i[55547];
  assign o[55546] = i[55546];
  assign o[55545] = i[55545];
  assign o[55544] = i[55544];
  assign o[55543] = i[55543];
  assign o[55542] = i[55542];
  assign o[55541] = i[55541];
  assign o[55540] = i[55540];
  assign o[55539] = i[55539];
  assign o[55538] = i[55538];
  assign o[55537] = i[55537];
  assign o[55536] = i[55536];
  assign o[55535] = i[55535];
  assign o[55534] = i[55534];
  assign o[55533] = i[55533];
  assign o[55532] = i[55532];
  assign o[55531] = i[55531];
  assign o[55530] = i[55530];
  assign o[55529] = i[55529];
  assign o[55528] = i[55528];
  assign o[55527] = i[55527];
  assign o[55526] = i[55526];
  assign o[55525] = i[55525];
  assign o[55524] = i[55524];
  assign o[55523] = i[55523];
  assign o[55522] = i[55522];
  assign o[55521] = i[55521];
  assign o[55520] = i[55520];
  assign o[55519] = i[55519];
  assign o[55518] = i[55518];
  assign o[55517] = i[55517];
  assign o[55516] = i[55516];
  assign o[55515] = i[55515];
  assign o[55514] = i[55514];
  assign o[55513] = i[55513];
  assign o[55512] = i[55512];
  assign o[55511] = i[55511];
  assign o[55510] = i[55510];
  assign o[55509] = i[55509];
  assign o[55508] = i[55508];
  assign o[55507] = i[55507];
  assign o[55506] = i[55506];
  assign o[55505] = i[55505];
  assign o[55504] = i[55504];
  assign o[55503] = i[55503];
  assign o[55502] = i[55502];
  assign o[55501] = i[55501];
  assign o[55500] = i[55500];
  assign o[55499] = i[55499];
  assign o[55498] = i[55498];
  assign o[55497] = i[55497];
  assign o[55496] = i[55496];
  assign o[55495] = i[55495];
  assign o[55494] = i[55494];
  assign o[55493] = i[55493];
  assign o[55492] = i[55492];
  assign o[55491] = i[55491];
  assign o[55490] = i[55490];
  assign o[55489] = i[55489];
  assign o[55488] = i[55488];
  assign o[55487] = i[55487];
  assign o[55486] = i[55486];
  assign o[55485] = i[55485];
  assign o[55484] = i[55484];
  assign o[55483] = i[55483];
  assign o[55482] = i[55482];
  assign o[55481] = i[55481];
  assign o[55480] = i[55480];
  assign o[55479] = i[55479];
  assign o[55478] = i[55478];
  assign o[55477] = i[55477];
  assign o[55476] = i[55476];
  assign o[55475] = i[55475];
  assign o[55474] = i[55474];
  assign o[55473] = i[55473];
  assign o[55472] = i[55472];
  assign o[55471] = i[55471];
  assign o[55470] = i[55470];
  assign o[55469] = i[55469];
  assign o[55468] = i[55468];
  assign o[55467] = i[55467];
  assign o[55466] = i[55466];
  assign o[55465] = i[55465];
  assign o[55464] = i[55464];
  assign o[55463] = i[55463];
  assign o[55462] = i[55462];
  assign o[55461] = i[55461];
  assign o[55460] = i[55460];
  assign o[55459] = i[55459];
  assign o[55458] = i[55458];
  assign o[55457] = i[55457];
  assign o[55456] = i[55456];
  assign o[55455] = i[55455];
  assign o[55454] = i[55454];
  assign o[55453] = i[55453];
  assign o[55452] = i[55452];
  assign o[55451] = i[55451];
  assign o[55450] = i[55450];
  assign o[55449] = i[55449];
  assign o[55448] = i[55448];
  assign o[55447] = i[55447];
  assign o[55446] = i[55446];
  assign o[55445] = i[55445];
  assign o[55444] = i[55444];
  assign o[55443] = i[55443];
  assign o[55442] = i[55442];
  assign o[55441] = i[55441];
  assign o[55440] = i[55440];
  assign o[55439] = i[55439];
  assign o[55438] = i[55438];
  assign o[55437] = i[55437];
  assign o[55436] = i[55436];
  assign o[55435] = i[55435];
  assign o[55434] = i[55434];
  assign o[55433] = i[55433];
  assign o[55432] = i[55432];
  assign o[55431] = i[55431];
  assign o[55430] = i[55430];
  assign o[55429] = i[55429];
  assign o[55428] = i[55428];
  assign o[55427] = i[55427];
  assign o[55426] = i[55426];
  assign o[55425] = i[55425];
  assign o[55424] = i[55424];
  assign o[55423] = i[55423];
  assign o[55422] = i[55422];
  assign o[55421] = i[55421];
  assign o[55420] = i[55420];
  assign o[55419] = i[55419];
  assign o[55418] = i[55418];
  assign o[55417] = i[55417];
  assign o[55416] = i[55416];
  assign o[55415] = i[55415];
  assign o[55414] = i[55414];
  assign o[55413] = i[55413];
  assign o[55412] = i[55412];
  assign o[55411] = i[55411];
  assign o[55410] = i[55410];
  assign o[55409] = i[55409];
  assign o[55408] = i[55408];
  assign o[55407] = i[55407];
  assign o[55406] = i[55406];
  assign o[55405] = i[55405];
  assign o[55404] = i[55404];
  assign o[55403] = i[55403];
  assign o[55402] = i[55402];
  assign o[55401] = i[55401];
  assign o[55400] = i[55400];
  assign o[55399] = i[55399];
  assign o[55398] = i[55398];
  assign o[55397] = i[55397];
  assign o[55396] = i[55396];
  assign o[55395] = i[55395];
  assign o[55394] = i[55394];
  assign o[55393] = i[55393];
  assign o[55392] = i[55392];
  assign o[55391] = i[55391];
  assign o[55390] = i[55390];
  assign o[55389] = i[55389];
  assign o[55388] = i[55388];
  assign o[55387] = i[55387];
  assign o[55386] = i[55386];
  assign o[55385] = i[55385];
  assign o[55384] = i[55384];
  assign o[55383] = i[55383];
  assign o[55382] = i[55382];
  assign o[55381] = i[55381];
  assign o[55380] = i[55380];
  assign o[55379] = i[55379];
  assign o[55378] = i[55378];
  assign o[55377] = i[55377];
  assign o[55376] = i[55376];
  assign o[55375] = i[55375];
  assign o[55374] = i[55374];
  assign o[55373] = i[55373];
  assign o[55372] = i[55372];
  assign o[55371] = i[55371];
  assign o[55370] = i[55370];
  assign o[55369] = i[55369];
  assign o[55368] = i[55368];
  assign o[55367] = i[55367];
  assign o[55366] = i[55366];
  assign o[55365] = i[55365];
  assign o[55364] = i[55364];
  assign o[55363] = i[55363];
  assign o[55362] = i[55362];
  assign o[55361] = i[55361];
  assign o[55360] = i[55360];
  assign o[55359] = i[55359];
  assign o[55358] = i[55358];
  assign o[55357] = i[55357];
  assign o[55356] = i[55356];
  assign o[55355] = i[55355];
  assign o[55354] = i[55354];
  assign o[55353] = i[55353];
  assign o[55352] = i[55352];
  assign o[55351] = i[55351];
  assign o[55350] = i[55350];
  assign o[55349] = i[55349];
  assign o[55348] = i[55348];
  assign o[55347] = i[55347];
  assign o[55346] = i[55346];
  assign o[55345] = i[55345];
  assign o[55344] = i[55344];
  assign o[55343] = i[55343];
  assign o[55342] = i[55342];
  assign o[55341] = i[55341];
  assign o[55340] = i[55340];
  assign o[55339] = i[55339];
  assign o[55338] = i[55338];
  assign o[55337] = i[55337];
  assign o[55336] = i[55336];
  assign o[55335] = i[55335];
  assign o[55334] = i[55334];
  assign o[55333] = i[55333];
  assign o[55332] = i[55332];
  assign o[55331] = i[55331];
  assign o[55330] = i[55330];
  assign o[55329] = i[55329];
  assign o[55328] = i[55328];
  assign o[55327] = i[55327];
  assign o[55326] = i[55326];
  assign o[55325] = i[55325];
  assign o[55324] = i[55324];
  assign o[55323] = i[55323];
  assign o[55322] = i[55322];
  assign o[55321] = i[55321];
  assign o[55320] = i[55320];
  assign o[55319] = i[55319];
  assign o[55318] = i[55318];
  assign o[55317] = i[55317];
  assign o[55316] = i[55316];
  assign o[55315] = i[55315];
  assign o[55314] = i[55314];
  assign o[55313] = i[55313];
  assign o[55312] = i[55312];
  assign o[55311] = i[55311];
  assign o[55310] = i[55310];
  assign o[55309] = i[55309];
  assign o[55308] = i[55308];
  assign o[55307] = i[55307];
  assign o[55306] = i[55306];
  assign o[55305] = i[55305];
  assign o[55304] = i[55304];
  assign o[55303] = i[55303];
  assign o[55302] = i[55302];
  assign o[55301] = i[55301];
  assign o[55300] = i[55300];
  assign o[55299] = i[55299];
  assign o[55298] = i[55298];
  assign o[55297] = i[55297];
  assign o[55296] = i[55296];
  assign o[55295] = i[55295];
  assign o[55294] = i[55294];
  assign o[55293] = i[55293];
  assign o[55292] = i[55292];
  assign o[55291] = i[55291];
  assign o[55290] = i[55290];
  assign o[55289] = i[55289];
  assign o[55288] = i[55288];
  assign o[55287] = i[55287];
  assign o[55286] = i[55286];
  assign o[55285] = i[55285];
  assign o[55284] = i[55284];
  assign o[55283] = i[55283];
  assign o[55282] = i[55282];
  assign o[55281] = i[55281];
  assign o[55280] = i[55280];
  assign o[55279] = i[55279];
  assign o[55278] = i[55278];
  assign o[55277] = i[55277];
  assign o[55276] = i[55276];
  assign o[55275] = i[55275];
  assign o[55274] = i[55274];
  assign o[55273] = i[55273];
  assign o[55272] = i[55272];
  assign o[55271] = i[55271];
  assign o[55270] = i[55270];
  assign o[55269] = i[55269];
  assign o[55268] = i[55268];
  assign o[55267] = i[55267];
  assign o[55266] = i[55266];
  assign o[55265] = i[55265];
  assign o[55264] = i[55264];
  assign o[55263] = i[55263];
  assign o[55262] = i[55262];
  assign o[55261] = i[55261];
  assign o[55260] = i[55260];
  assign o[55259] = i[55259];
  assign o[55258] = i[55258];
  assign o[55257] = i[55257];
  assign o[55256] = i[55256];
  assign o[55255] = i[55255];
  assign o[55254] = i[55254];
  assign o[55253] = i[55253];
  assign o[55252] = i[55252];
  assign o[55251] = i[55251];
  assign o[55250] = i[55250];
  assign o[55249] = i[55249];
  assign o[55248] = i[55248];
  assign o[55247] = i[55247];
  assign o[55246] = i[55246];
  assign o[55245] = i[55245];
  assign o[55244] = i[55244];
  assign o[55243] = i[55243];
  assign o[55242] = i[55242];
  assign o[55241] = i[55241];
  assign o[55240] = i[55240];
  assign o[55239] = i[55239];
  assign o[55238] = i[55238];
  assign o[55237] = i[55237];
  assign o[55236] = i[55236];
  assign o[55235] = i[55235];
  assign o[55234] = i[55234];
  assign o[55233] = i[55233];
  assign o[55232] = i[55232];
  assign o[55231] = i[55231];
  assign o[55230] = i[55230];
  assign o[55229] = i[55229];
  assign o[55228] = i[55228];
  assign o[55227] = i[55227];
  assign o[55226] = i[55226];
  assign o[55225] = i[55225];
  assign o[55224] = i[55224];
  assign o[55223] = i[55223];
  assign o[55222] = i[55222];
  assign o[55221] = i[55221];
  assign o[55220] = i[55220];
  assign o[55219] = i[55219];
  assign o[55218] = i[55218];
  assign o[55217] = i[55217];
  assign o[55216] = i[55216];
  assign o[55215] = i[55215];
  assign o[55214] = i[55214];
  assign o[55213] = i[55213];
  assign o[55212] = i[55212];
  assign o[55211] = i[55211];
  assign o[55210] = i[55210];
  assign o[55209] = i[55209];
  assign o[55208] = i[55208];
  assign o[55207] = i[55207];
  assign o[55206] = i[55206];
  assign o[55205] = i[55205];
  assign o[55204] = i[55204];
  assign o[55203] = i[55203];
  assign o[55202] = i[55202];
  assign o[55201] = i[55201];
  assign o[55200] = i[55200];
  assign o[55199] = i[55199];
  assign o[55198] = i[55198];
  assign o[55197] = i[55197];
  assign o[55196] = i[55196];
  assign o[55195] = i[55195];
  assign o[55194] = i[55194];
  assign o[55193] = i[55193];
  assign o[55192] = i[55192];
  assign o[55191] = i[55191];
  assign o[55190] = i[55190];
  assign o[55189] = i[55189];
  assign o[55188] = i[55188];
  assign o[55187] = i[55187];
  assign o[55186] = i[55186];
  assign o[55185] = i[55185];
  assign o[55184] = i[55184];
  assign o[55183] = i[55183];
  assign o[55182] = i[55182];
  assign o[55181] = i[55181];
  assign o[55180] = i[55180];
  assign o[55179] = i[55179];
  assign o[55178] = i[55178];
  assign o[55177] = i[55177];
  assign o[55176] = i[55176];
  assign o[55175] = i[55175];
  assign o[55174] = i[55174];
  assign o[55173] = i[55173];
  assign o[55172] = i[55172];
  assign o[55171] = i[55171];
  assign o[55170] = i[55170];
  assign o[55169] = i[55169];
  assign o[55168] = i[55168];
  assign o[55167] = i[55167];
  assign o[55166] = i[55166];
  assign o[55165] = i[55165];
  assign o[55164] = i[55164];
  assign o[55163] = i[55163];
  assign o[55162] = i[55162];
  assign o[55161] = i[55161];
  assign o[55160] = i[55160];
  assign o[55159] = i[55159];
  assign o[55158] = i[55158];
  assign o[55157] = i[55157];
  assign o[55156] = i[55156];
  assign o[55155] = i[55155];
  assign o[55154] = i[55154];
  assign o[55153] = i[55153];
  assign o[55152] = i[55152];
  assign o[55151] = i[55151];
  assign o[55150] = i[55150];
  assign o[55149] = i[55149];
  assign o[55148] = i[55148];
  assign o[55147] = i[55147];
  assign o[55146] = i[55146];
  assign o[55145] = i[55145];
  assign o[55144] = i[55144];
  assign o[55143] = i[55143];
  assign o[55142] = i[55142];
  assign o[55141] = i[55141];
  assign o[55140] = i[55140];
  assign o[55139] = i[55139];
  assign o[55138] = i[55138];
  assign o[55137] = i[55137];
  assign o[55136] = i[55136];
  assign o[55135] = i[55135];
  assign o[55134] = i[55134];
  assign o[55133] = i[55133];
  assign o[55132] = i[55132];
  assign o[55131] = i[55131];
  assign o[55130] = i[55130];
  assign o[55129] = i[55129];
  assign o[55128] = i[55128];
  assign o[55127] = i[55127];
  assign o[55126] = i[55126];
  assign o[55125] = i[55125];
  assign o[55124] = i[55124];
  assign o[55123] = i[55123];
  assign o[55122] = i[55122];
  assign o[55121] = i[55121];
  assign o[55120] = i[55120];
  assign o[55119] = i[55119];
  assign o[55118] = i[55118];
  assign o[55117] = i[55117];
  assign o[55116] = i[55116];
  assign o[55115] = i[55115];
  assign o[55114] = i[55114];
  assign o[55113] = i[55113];
  assign o[55112] = i[55112];
  assign o[55111] = i[55111];
  assign o[55110] = i[55110];
  assign o[55109] = i[55109];
  assign o[55108] = i[55108];
  assign o[55107] = i[55107];
  assign o[55106] = i[55106];
  assign o[55105] = i[55105];
  assign o[55104] = i[55104];
  assign o[55103] = i[55103];
  assign o[55102] = i[55102];
  assign o[55101] = i[55101];
  assign o[55100] = i[55100];
  assign o[55099] = i[55099];
  assign o[55098] = i[55098];
  assign o[55097] = i[55097];
  assign o[55096] = i[55096];
  assign o[55095] = i[55095];
  assign o[55094] = i[55094];
  assign o[55093] = i[55093];
  assign o[55092] = i[55092];
  assign o[55091] = i[55091];
  assign o[55090] = i[55090];
  assign o[55089] = i[55089];
  assign o[55088] = i[55088];
  assign o[55087] = i[55087];
  assign o[55086] = i[55086];
  assign o[55085] = i[55085];
  assign o[55084] = i[55084];
  assign o[55083] = i[55083];
  assign o[55082] = i[55082];
  assign o[55081] = i[55081];
  assign o[55080] = i[55080];
  assign o[55079] = i[55079];
  assign o[55078] = i[55078];
  assign o[55077] = i[55077];
  assign o[55076] = i[55076];
  assign o[55075] = i[55075];
  assign o[55074] = i[55074];
  assign o[55073] = i[55073];
  assign o[55072] = i[55072];
  assign o[55071] = i[55071];
  assign o[55070] = i[55070];
  assign o[55069] = i[55069];
  assign o[55068] = i[55068];
  assign o[55067] = i[55067];
  assign o[55066] = i[55066];
  assign o[55065] = i[55065];
  assign o[55064] = i[55064];
  assign o[55063] = i[55063];
  assign o[55062] = i[55062];
  assign o[55061] = i[55061];
  assign o[55060] = i[55060];
  assign o[55059] = i[55059];
  assign o[55058] = i[55058];
  assign o[55057] = i[55057];
  assign o[55056] = i[55056];
  assign o[55055] = i[55055];
  assign o[55054] = i[55054];
  assign o[55053] = i[55053];
  assign o[55052] = i[55052];
  assign o[55051] = i[55051];
  assign o[55050] = i[55050];
  assign o[55049] = i[55049];
  assign o[55048] = i[55048];
  assign o[55047] = i[55047];
  assign o[55046] = i[55046];
  assign o[55045] = i[55045];
  assign o[55044] = i[55044];
  assign o[55043] = i[55043];
  assign o[55042] = i[55042];
  assign o[55041] = i[55041];
  assign o[55040] = i[55040];
  assign o[55039] = i[55039];
  assign o[55038] = i[55038];
  assign o[55037] = i[55037];
  assign o[55036] = i[55036];
  assign o[55035] = i[55035];
  assign o[55034] = i[55034];
  assign o[55033] = i[55033];
  assign o[55032] = i[55032];
  assign o[55031] = i[55031];
  assign o[55030] = i[55030];
  assign o[55029] = i[55029];
  assign o[55028] = i[55028];
  assign o[55027] = i[55027];
  assign o[55026] = i[55026];
  assign o[55025] = i[55025];
  assign o[55024] = i[55024];
  assign o[55023] = i[55023];
  assign o[55022] = i[55022];
  assign o[55021] = i[55021];
  assign o[55020] = i[55020];
  assign o[55019] = i[55019];
  assign o[55018] = i[55018];
  assign o[55017] = i[55017];
  assign o[55016] = i[55016];
  assign o[55015] = i[55015];
  assign o[55014] = i[55014];
  assign o[55013] = i[55013];
  assign o[55012] = i[55012];
  assign o[55011] = i[55011];
  assign o[55010] = i[55010];
  assign o[55009] = i[55009];
  assign o[55008] = i[55008];
  assign o[55007] = i[55007];
  assign o[55006] = i[55006];
  assign o[55005] = i[55005];
  assign o[55004] = i[55004];
  assign o[55003] = i[55003];
  assign o[55002] = i[55002];
  assign o[55001] = i[55001];
  assign o[55000] = i[55000];
  assign o[54999] = i[54999];
  assign o[54998] = i[54998];
  assign o[54997] = i[54997];
  assign o[54996] = i[54996];
  assign o[54995] = i[54995];
  assign o[54994] = i[54994];
  assign o[54993] = i[54993];
  assign o[54992] = i[54992];
  assign o[54991] = i[54991];
  assign o[54990] = i[54990];
  assign o[54989] = i[54989];
  assign o[54988] = i[54988];
  assign o[54987] = i[54987];
  assign o[54986] = i[54986];
  assign o[54985] = i[54985];
  assign o[54984] = i[54984];
  assign o[54983] = i[54983];
  assign o[54982] = i[54982];
  assign o[54981] = i[54981];
  assign o[54980] = i[54980];
  assign o[54979] = i[54979];
  assign o[54978] = i[54978];
  assign o[54977] = i[54977];
  assign o[54976] = i[54976];
  assign o[54975] = i[54975];
  assign o[54974] = i[54974];
  assign o[54973] = i[54973];
  assign o[54972] = i[54972];
  assign o[54971] = i[54971];
  assign o[54970] = i[54970];
  assign o[54969] = i[54969];
  assign o[54968] = i[54968];
  assign o[54967] = i[54967];
  assign o[54966] = i[54966];
  assign o[54965] = i[54965];
  assign o[54964] = i[54964];
  assign o[54963] = i[54963];
  assign o[54962] = i[54962];
  assign o[54961] = i[54961];
  assign o[54960] = i[54960];
  assign o[54959] = i[54959];
  assign o[54958] = i[54958];
  assign o[54957] = i[54957];
  assign o[54956] = i[54956];
  assign o[54955] = i[54955];
  assign o[54954] = i[54954];
  assign o[54953] = i[54953];
  assign o[54952] = i[54952];
  assign o[54951] = i[54951];
  assign o[54950] = i[54950];
  assign o[54949] = i[54949];
  assign o[54948] = i[54948];
  assign o[54947] = i[54947];
  assign o[54946] = i[54946];
  assign o[54945] = i[54945];
  assign o[54944] = i[54944];
  assign o[54943] = i[54943];
  assign o[54942] = i[54942];
  assign o[54941] = i[54941];
  assign o[54940] = i[54940];
  assign o[54939] = i[54939];
  assign o[54938] = i[54938];
  assign o[54937] = i[54937];
  assign o[54936] = i[54936];
  assign o[54935] = i[54935];
  assign o[54934] = i[54934];
  assign o[54933] = i[54933];
  assign o[54932] = i[54932];
  assign o[54931] = i[54931];
  assign o[54930] = i[54930];
  assign o[54929] = i[54929];
  assign o[54928] = i[54928];
  assign o[54927] = i[54927];
  assign o[54926] = i[54926];
  assign o[54925] = i[54925];
  assign o[54924] = i[54924];
  assign o[54923] = i[54923];
  assign o[54922] = i[54922];
  assign o[54921] = i[54921];
  assign o[54920] = i[54920];
  assign o[54919] = i[54919];
  assign o[54918] = i[54918];
  assign o[54917] = i[54917];
  assign o[54916] = i[54916];
  assign o[54915] = i[54915];
  assign o[54914] = i[54914];
  assign o[54913] = i[54913];
  assign o[54912] = i[54912];
  assign o[54911] = i[54911];
  assign o[54910] = i[54910];
  assign o[54909] = i[54909];
  assign o[54908] = i[54908];
  assign o[54907] = i[54907];
  assign o[54906] = i[54906];
  assign o[54905] = i[54905];
  assign o[54904] = i[54904];
  assign o[54903] = i[54903];
  assign o[54902] = i[54902];
  assign o[54901] = i[54901];
  assign o[54900] = i[54900];
  assign o[54899] = i[54899];
  assign o[54898] = i[54898];
  assign o[54897] = i[54897];
  assign o[54896] = i[54896];
  assign o[54895] = i[54895];
  assign o[54894] = i[54894];
  assign o[54893] = i[54893];
  assign o[54892] = i[54892];
  assign o[54891] = i[54891];
  assign o[54890] = i[54890];
  assign o[54889] = i[54889];
  assign o[54888] = i[54888];
  assign o[54887] = i[54887];
  assign o[54886] = i[54886];
  assign o[54885] = i[54885];
  assign o[54884] = i[54884];
  assign o[54883] = i[54883];
  assign o[54882] = i[54882];
  assign o[54881] = i[54881];
  assign o[54880] = i[54880];
  assign o[54879] = i[54879];
  assign o[54878] = i[54878];
  assign o[54877] = i[54877];
  assign o[54876] = i[54876];
  assign o[54875] = i[54875];
  assign o[54874] = i[54874];
  assign o[54873] = i[54873];
  assign o[54872] = i[54872];
  assign o[54871] = i[54871];
  assign o[54870] = i[54870];
  assign o[54869] = i[54869];
  assign o[54868] = i[54868];
  assign o[54867] = i[54867];
  assign o[54866] = i[54866];
  assign o[54865] = i[54865];
  assign o[54864] = i[54864];
  assign o[54863] = i[54863];
  assign o[54862] = i[54862];
  assign o[54861] = i[54861];
  assign o[54860] = i[54860];
  assign o[54859] = i[54859];
  assign o[54858] = i[54858];
  assign o[54857] = i[54857];
  assign o[54856] = i[54856];
  assign o[54855] = i[54855];
  assign o[54854] = i[54854];
  assign o[54853] = i[54853];
  assign o[54852] = i[54852];
  assign o[54851] = i[54851];
  assign o[54850] = i[54850];
  assign o[54849] = i[54849];
  assign o[54848] = i[54848];
  assign o[54847] = i[54847];
  assign o[54846] = i[54846];
  assign o[54845] = i[54845];
  assign o[54844] = i[54844];
  assign o[54843] = i[54843];
  assign o[54842] = i[54842];
  assign o[54841] = i[54841];
  assign o[54840] = i[54840];
  assign o[54839] = i[54839];
  assign o[54838] = i[54838];
  assign o[54837] = i[54837];
  assign o[54836] = i[54836];
  assign o[54835] = i[54835];
  assign o[54834] = i[54834];
  assign o[54833] = i[54833];
  assign o[54832] = i[54832];
  assign o[54831] = i[54831];
  assign o[54830] = i[54830];
  assign o[54829] = i[54829];
  assign o[54828] = i[54828];
  assign o[54827] = i[54827];
  assign o[54826] = i[54826];
  assign o[54825] = i[54825];
  assign o[54824] = i[54824];
  assign o[54823] = i[54823];
  assign o[54822] = i[54822];
  assign o[54821] = i[54821];
  assign o[54820] = i[54820];
  assign o[54819] = i[54819];
  assign o[54818] = i[54818];
  assign o[54817] = i[54817];
  assign o[54816] = i[54816];
  assign o[54815] = i[54815];
  assign o[54814] = i[54814];
  assign o[54813] = i[54813];
  assign o[54812] = i[54812];
  assign o[54811] = i[54811];
  assign o[54810] = i[54810];
  assign o[54809] = i[54809];
  assign o[54808] = i[54808];
  assign o[54807] = i[54807];
  assign o[54806] = i[54806];
  assign o[54805] = i[54805];
  assign o[54804] = i[54804];
  assign o[54803] = i[54803];
  assign o[54802] = i[54802];
  assign o[54801] = i[54801];
  assign o[54800] = i[54800];
  assign o[54799] = i[54799];
  assign o[54798] = i[54798];
  assign o[54797] = i[54797];
  assign o[54796] = i[54796];
  assign o[54795] = i[54795];
  assign o[54794] = i[54794];
  assign o[54793] = i[54793];
  assign o[54792] = i[54792];
  assign o[54791] = i[54791];
  assign o[54790] = i[54790];
  assign o[54789] = i[54789];
  assign o[54788] = i[54788];
  assign o[54787] = i[54787];
  assign o[54786] = i[54786];
  assign o[54785] = i[54785];
  assign o[54784] = i[54784];
  assign o[54783] = i[54783];
  assign o[54782] = i[54782];
  assign o[54781] = i[54781];
  assign o[54780] = i[54780];
  assign o[54779] = i[54779];
  assign o[54778] = i[54778];
  assign o[54777] = i[54777];
  assign o[54776] = i[54776];
  assign o[54775] = i[54775];
  assign o[54774] = i[54774];
  assign o[54773] = i[54773];
  assign o[54772] = i[54772];
  assign o[54771] = i[54771];
  assign o[54770] = i[54770];
  assign o[54769] = i[54769];
  assign o[54768] = i[54768];
  assign o[54767] = i[54767];
  assign o[54766] = i[54766];
  assign o[54765] = i[54765];
  assign o[54764] = i[54764];
  assign o[54763] = i[54763];
  assign o[54762] = i[54762];
  assign o[54761] = i[54761];
  assign o[54760] = i[54760];
  assign o[54759] = i[54759];
  assign o[54758] = i[54758];
  assign o[54757] = i[54757];
  assign o[54756] = i[54756];
  assign o[54755] = i[54755];
  assign o[54754] = i[54754];
  assign o[54753] = i[54753];
  assign o[54752] = i[54752];
  assign o[54751] = i[54751];
  assign o[54750] = i[54750];
  assign o[54749] = i[54749];
  assign o[54748] = i[54748];
  assign o[54747] = i[54747];
  assign o[54746] = i[54746];
  assign o[54745] = i[54745];
  assign o[54744] = i[54744];
  assign o[54743] = i[54743];
  assign o[54742] = i[54742];
  assign o[54741] = i[54741];
  assign o[54740] = i[54740];
  assign o[54739] = i[54739];
  assign o[54738] = i[54738];
  assign o[54737] = i[54737];
  assign o[54736] = i[54736];
  assign o[54735] = i[54735];
  assign o[54734] = i[54734];
  assign o[54733] = i[54733];
  assign o[54732] = i[54732];
  assign o[54731] = i[54731];
  assign o[54730] = i[54730];
  assign o[54729] = i[54729];
  assign o[54728] = i[54728];
  assign o[54727] = i[54727];
  assign o[54726] = i[54726];
  assign o[54725] = i[54725];
  assign o[54724] = i[54724];
  assign o[54723] = i[54723];
  assign o[54722] = i[54722];
  assign o[54721] = i[54721];
  assign o[54720] = i[54720];
  assign o[54719] = i[54719];
  assign o[54718] = i[54718];
  assign o[54717] = i[54717];
  assign o[54716] = i[54716];
  assign o[54715] = i[54715];
  assign o[54714] = i[54714];
  assign o[54713] = i[54713];
  assign o[54712] = i[54712];
  assign o[54711] = i[54711];
  assign o[54710] = i[54710];
  assign o[54709] = i[54709];
  assign o[54708] = i[54708];
  assign o[54707] = i[54707];
  assign o[54706] = i[54706];
  assign o[54705] = i[54705];
  assign o[54704] = i[54704];
  assign o[54703] = i[54703];
  assign o[54702] = i[54702];
  assign o[54701] = i[54701];
  assign o[54700] = i[54700];
  assign o[54699] = i[54699];
  assign o[54698] = i[54698];
  assign o[54697] = i[54697];
  assign o[54696] = i[54696];
  assign o[54695] = i[54695];
  assign o[54694] = i[54694];
  assign o[54693] = i[54693];
  assign o[54692] = i[54692];
  assign o[54691] = i[54691];
  assign o[54690] = i[54690];
  assign o[54689] = i[54689];
  assign o[54688] = i[54688];
  assign o[54687] = i[54687];
  assign o[54686] = i[54686];
  assign o[54685] = i[54685];
  assign o[54684] = i[54684];
  assign o[54683] = i[54683];
  assign o[54682] = i[54682];
  assign o[54681] = i[54681];
  assign o[54680] = i[54680];
  assign o[54679] = i[54679];
  assign o[54678] = i[54678];
  assign o[54677] = i[54677];
  assign o[54676] = i[54676];
  assign o[54675] = i[54675];
  assign o[54674] = i[54674];
  assign o[54673] = i[54673];
  assign o[54672] = i[54672];
  assign o[54671] = i[54671];
  assign o[54670] = i[54670];
  assign o[54669] = i[54669];
  assign o[54668] = i[54668];
  assign o[54667] = i[54667];
  assign o[54666] = i[54666];
  assign o[54665] = i[54665];
  assign o[54664] = i[54664];
  assign o[54663] = i[54663];
  assign o[54662] = i[54662];
  assign o[54661] = i[54661];
  assign o[54660] = i[54660];
  assign o[54659] = i[54659];
  assign o[54658] = i[54658];
  assign o[54657] = i[54657];
  assign o[54656] = i[54656];
  assign o[54655] = i[54655];
  assign o[54654] = i[54654];
  assign o[54653] = i[54653];
  assign o[54652] = i[54652];
  assign o[54651] = i[54651];
  assign o[54650] = i[54650];
  assign o[54649] = i[54649];
  assign o[54648] = i[54648];
  assign o[54647] = i[54647];
  assign o[54646] = i[54646];
  assign o[54645] = i[54645];
  assign o[54644] = i[54644];
  assign o[54643] = i[54643];
  assign o[54642] = i[54642];
  assign o[54641] = i[54641];
  assign o[54640] = i[54640];
  assign o[54639] = i[54639];
  assign o[54638] = i[54638];
  assign o[54637] = i[54637];
  assign o[54636] = i[54636];
  assign o[54635] = i[54635];
  assign o[54634] = i[54634];
  assign o[54633] = i[54633];
  assign o[54632] = i[54632];
  assign o[54631] = i[54631];
  assign o[54630] = i[54630];
  assign o[54629] = i[54629];
  assign o[54628] = i[54628];
  assign o[54627] = i[54627];
  assign o[54626] = i[54626];
  assign o[54625] = i[54625];
  assign o[54624] = i[54624];
  assign o[54623] = i[54623];
  assign o[54622] = i[54622];
  assign o[54621] = i[54621];
  assign o[54620] = i[54620];
  assign o[54619] = i[54619];
  assign o[54618] = i[54618];
  assign o[54617] = i[54617];
  assign o[54616] = i[54616];
  assign o[54615] = i[54615];
  assign o[54614] = i[54614];
  assign o[54613] = i[54613];
  assign o[54612] = i[54612];
  assign o[54611] = i[54611];
  assign o[54610] = i[54610];
  assign o[54609] = i[54609];
  assign o[54608] = i[54608];
  assign o[54607] = i[54607];
  assign o[54606] = i[54606];
  assign o[54605] = i[54605];
  assign o[54604] = i[54604];
  assign o[54603] = i[54603];
  assign o[54602] = i[54602];
  assign o[54601] = i[54601];
  assign o[54600] = i[54600];
  assign o[54599] = i[54599];
  assign o[54598] = i[54598];
  assign o[54597] = i[54597];
  assign o[54596] = i[54596];
  assign o[54595] = i[54595];
  assign o[54594] = i[54594];
  assign o[54593] = i[54593];
  assign o[54592] = i[54592];
  assign o[54591] = i[54591];
  assign o[54590] = i[54590];
  assign o[54589] = i[54589];
  assign o[54588] = i[54588];
  assign o[54587] = i[54587];
  assign o[54586] = i[54586];
  assign o[54585] = i[54585];
  assign o[54584] = i[54584];
  assign o[54583] = i[54583];
  assign o[54582] = i[54582];
  assign o[54581] = i[54581];
  assign o[54580] = i[54580];
  assign o[54579] = i[54579];
  assign o[54578] = i[54578];
  assign o[54577] = i[54577];
  assign o[54576] = i[54576];
  assign o[54575] = i[54575];
  assign o[54574] = i[54574];
  assign o[54573] = i[54573];
  assign o[54572] = i[54572];
  assign o[54571] = i[54571];
  assign o[54570] = i[54570];
  assign o[54569] = i[54569];
  assign o[54568] = i[54568];
  assign o[54567] = i[54567];
  assign o[54566] = i[54566];
  assign o[54565] = i[54565];
  assign o[54564] = i[54564];
  assign o[54563] = i[54563];
  assign o[54562] = i[54562];
  assign o[54561] = i[54561];
  assign o[54560] = i[54560];
  assign o[54559] = i[54559];
  assign o[54558] = i[54558];
  assign o[54557] = i[54557];
  assign o[54556] = i[54556];
  assign o[54555] = i[54555];
  assign o[54554] = i[54554];
  assign o[54553] = i[54553];
  assign o[54552] = i[54552];
  assign o[54551] = i[54551];
  assign o[54550] = i[54550];
  assign o[54549] = i[54549];
  assign o[54548] = i[54548];
  assign o[54547] = i[54547];
  assign o[54546] = i[54546];
  assign o[54545] = i[54545];
  assign o[54544] = i[54544];
  assign o[54543] = i[54543];
  assign o[54542] = i[54542];
  assign o[54541] = i[54541];
  assign o[54540] = i[54540];
  assign o[54539] = i[54539];
  assign o[54538] = i[54538];
  assign o[54537] = i[54537];
  assign o[54536] = i[54536];
  assign o[54535] = i[54535];
  assign o[54534] = i[54534];
  assign o[54533] = i[54533];
  assign o[54532] = i[54532];
  assign o[54531] = i[54531];
  assign o[54530] = i[54530];
  assign o[54529] = i[54529];
  assign o[54528] = i[54528];
  assign o[54527] = i[54527];
  assign o[54526] = i[54526];
  assign o[54525] = i[54525];
  assign o[54524] = i[54524];
  assign o[54523] = i[54523];
  assign o[54522] = i[54522];
  assign o[54521] = i[54521];
  assign o[54520] = i[54520];
  assign o[54519] = i[54519];
  assign o[54518] = i[54518];
  assign o[54517] = i[54517];
  assign o[54516] = i[54516];
  assign o[54515] = i[54515];
  assign o[54514] = i[54514];
  assign o[54513] = i[54513];
  assign o[54512] = i[54512];
  assign o[54511] = i[54511];
  assign o[54510] = i[54510];
  assign o[54509] = i[54509];
  assign o[54508] = i[54508];
  assign o[54507] = i[54507];
  assign o[54506] = i[54506];
  assign o[54505] = i[54505];
  assign o[54504] = i[54504];
  assign o[54503] = i[54503];
  assign o[54502] = i[54502];
  assign o[54501] = i[54501];
  assign o[54500] = i[54500];
  assign o[54499] = i[54499];
  assign o[54498] = i[54498];
  assign o[54497] = i[54497];
  assign o[54496] = i[54496];
  assign o[54495] = i[54495];
  assign o[54494] = i[54494];
  assign o[54493] = i[54493];
  assign o[54492] = i[54492];
  assign o[54491] = i[54491];
  assign o[54490] = i[54490];
  assign o[54489] = i[54489];
  assign o[54488] = i[54488];
  assign o[54487] = i[54487];
  assign o[54486] = i[54486];
  assign o[54485] = i[54485];
  assign o[54484] = i[54484];
  assign o[54483] = i[54483];
  assign o[54482] = i[54482];
  assign o[54481] = i[54481];
  assign o[54480] = i[54480];
  assign o[54479] = i[54479];
  assign o[54478] = i[54478];
  assign o[54477] = i[54477];
  assign o[54476] = i[54476];
  assign o[54475] = i[54475];
  assign o[54474] = i[54474];
  assign o[54473] = i[54473];
  assign o[54472] = i[54472];
  assign o[54471] = i[54471];
  assign o[54470] = i[54470];
  assign o[54469] = i[54469];
  assign o[54468] = i[54468];
  assign o[54467] = i[54467];
  assign o[54466] = i[54466];
  assign o[54465] = i[54465];
  assign o[54464] = i[54464];
  assign o[54463] = i[54463];
  assign o[54462] = i[54462];
  assign o[54461] = i[54461];
  assign o[54460] = i[54460];
  assign o[54459] = i[54459];
  assign o[54458] = i[54458];
  assign o[54457] = i[54457];
  assign o[54456] = i[54456];
  assign o[54455] = i[54455];
  assign o[54454] = i[54454];
  assign o[54453] = i[54453];
  assign o[54452] = i[54452];
  assign o[54451] = i[54451];
  assign o[54450] = i[54450];
  assign o[54449] = i[54449];
  assign o[54448] = i[54448];
  assign o[54447] = i[54447];
  assign o[54446] = i[54446];
  assign o[54445] = i[54445];
  assign o[54444] = i[54444];
  assign o[54443] = i[54443];
  assign o[54442] = i[54442];
  assign o[54441] = i[54441];
  assign o[54440] = i[54440];
  assign o[54439] = i[54439];
  assign o[54438] = i[54438];
  assign o[54437] = i[54437];
  assign o[54436] = i[54436];
  assign o[54435] = i[54435];
  assign o[54434] = i[54434];
  assign o[54433] = i[54433];
  assign o[54432] = i[54432];
  assign o[54431] = i[54431];
  assign o[54430] = i[54430];
  assign o[54429] = i[54429];
  assign o[54428] = i[54428];
  assign o[54427] = i[54427];
  assign o[54426] = i[54426];
  assign o[54425] = i[54425];
  assign o[54424] = i[54424];
  assign o[54423] = i[54423];
  assign o[54422] = i[54422];
  assign o[54421] = i[54421];
  assign o[54420] = i[54420];
  assign o[54419] = i[54419];
  assign o[54418] = i[54418];
  assign o[54417] = i[54417];
  assign o[54416] = i[54416];
  assign o[54415] = i[54415];
  assign o[54414] = i[54414];
  assign o[54413] = i[54413];
  assign o[54412] = i[54412];
  assign o[54411] = i[54411];
  assign o[54410] = i[54410];
  assign o[54409] = i[54409];
  assign o[54408] = i[54408];
  assign o[54407] = i[54407];
  assign o[54406] = i[54406];
  assign o[54405] = i[54405];
  assign o[54404] = i[54404];
  assign o[54403] = i[54403];
  assign o[54402] = i[54402];
  assign o[54401] = i[54401];
  assign o[54400] = i[54400];
  assign o[54399] = i[54399];
  assign o[54398] = i[54398];
  assign o[54397] = i[54397];
  assign o[54396] = i[54396];
  assign o[54395] = i[54395];
  assign o[54394] = i[54394];
  assign o[54393] = i[54393];
  assign o[54392] = i[54392];
  assign o[54391] = i[54391];
  assign o[54390] = i[54390];
  assign o[54389] = i[54389];
  assign o[54388] = i[54388];
  assign o[54387] = i[54387];
  assign o[54386] = i[54386];
  assign o[54385] = i[54385];
  assign o[54384] = i[54384];
  assign o[54383] = i[54383];
  assign o[54382] = i[54382];
  assign o[54381] = i[54381];
  assign o[54380] = i[54380];
  assign o[54379] = i[54379];
  assign o[54378] = i[54378];
  assign o[54377] = i[54377];
  assign o[54376] = i[54376];
  assign o[54375] = i[54375];
  assign o[54374] = i[54374];
  assign o[54373] = i[54373];
  assign o[54372] = i[54372];
  assign o[54371] = i[54371];
  assign o[54370] = i[54370];
  assign o[54369] = i[54369];
  assign o[54368] = i[54368];
  assign o[54367] = i[54367];
  assign o[54366] = i[54366];
  assign o[54365] = i[54365];
  assign o[54364] = i[54364];
  assign o[54363] = i[54363];
  assign o[54362] = i[54362];
  assign o[54361] = i[54361];
  assign o[54360] = i[54360];
  assign o[54359] = i[54359];
  assign o[54358] = i[54358];
  assign o[54357] = i[54357];
  assign o[54356] = i[54356];
  assign o[54355] = i[54355];
  assign o[54354] = i[54354];
  assign o[54353] = i[54353];
  assign o[54352] = i[54352];
  assign o[54351] = i[54351];
  assign o[54350] = i[54350];
  assign o[54349] = i[54349];
  assign o[54348] = i[54348];
  assign o[54347] = i[54347];
  assign o[54346] = i[54346];
  assign o[54345] = i[54345];
  assign o[54344] = i[54344];
  assign o[54343] = i[54343];
  assign o[54342] = i[54342];
  assign o[54341] = i[54341];
  assign o[54340] = i[54340];
  assign o[54339] = i[54339];
  assign o[54338] = i[54338];
  assign o[54337] = i[54337];
  assign o[54336] = i[54336];
  assign o[54335] = i[54335];
  assign o[54334] = i[54334];
  assign o[54333] = i[54333];
  assign o[54332] = i[54332];
  assign o[54331] = i[54331];
  assign o[54330] = i[54330];
  assign o[54329] = i[54329];
  assign o[54328] = i[54328];
  assign o[54327] = i[54327];
  assign o[54326] = i[54326];
  assign o[54325] = i[54325];
  assign o[54324] = i[54324];
  assign o[54323] = i[54323];
  assign o[54322] = i[54322];
  assign o[54321] = i[54321];
  assign o[54320] = i[54320];
  assign o[54319] = i[54319];
  assign o[54318] = i[54318];
  assign o[54317] = i[54317];
  assign o[54316] = i[54316];
  assign o[54315] = i[54315];
  assign o[54314] = i[54314];
  assign o[54313] = i[54313];
  assign o[54312] = i[54312];
  assign o[54311] = i[54311];
  assign o[54310] = i[54310];
  assign o[54309] = i[54309];
  assign o[54308] = i[54308];
  assign o[54307] = i[54307];
  assign o[54306] = i[54306];
  assign o[54305] = i[54305];
  assign o[54304] = i[54304];
  assign o[54303] = i[54303];
  assign o[54302] = i[54302];
  assign o[54301] = i[54301];
  assign o[54300] = i[54300];
  assign o[54299] = i[54299];
  assign o[54298] = i[54298];
  assign o[54297] = i[54297];
  assign o[54296] = i[54296];
  assign o[54295] = i[54295];
  assign o[54294] = i[54294];
  assign o[54293] = i[54293];
  assign o[54292] = i[54292];
  assign o[54291] = i[54291];
  assign o[54290] = i[54290];
  assign o[54289] = i[54289];
  assign o[54288] = i[54288];
  assign o[54287] = i[54287];
  assign o[54286] = i[54286];
  assign o[54285] = i[54285];
  assign o[54284] = i[54284];
  assign o[54283] = i[54283];
  assign o[54282] = i[54282];
  assign o[54281] = i[54281];
  assign o[54280] = i[54280];
  assign o[54279] = i[54279];
  assign o[54278] = i[54278];
  assign o[54277] = i[54277];
  assign o[54276] = i[54276];
  assign o[54275] = i[54275];
  assign o[54274] = i[54274];
  assign o[54273] = i[54273];
  assign o[54272] = i[54272];
  assign o[54271] = i[54271];
  assign o[54270] = i[54270];
  assign o[54269] = i[54269];
  assign o[54268] = i[54268];
  assign o[54267] = i[54267];
  assign o[54266] = i[54266];
  assign o[54265] = i[54265];
  assign o[54264] = i[54264];
  assign o[54263] = i[54263];
  assign o[54262] = i[54262];
  assign o[54261] = i[54261];
  assign o[54260] = i[54260];
  assign o[54259] = i[54259];
  assign o[54258] = i[54258];
  assign o[54257] = i[54257];
  assign o[54256] = i[54256];
  assign o[54255] = i[54255];
  assign o[54254] = i[54254];
  assign o[54253] = i[54253];
  assign o[54252] = i[54252];
  assign o[54251] = i[54251];
  assign o[54250] = i[54250];
  assign o[54249] = i[54249];
  assign o[54248] = i[54248];
  assign o[54247] = i[54247];
  assign o[54246] = i[54246];
  assign o[54245] = i[54245];
  assign o[54244] = i[54244];
  assign o[54243] = i[54243];
  assign o[54242] = i[54242];
  assign o[54241] = i[54241];
  assign o[54240] = i[54240];
  assign o[54239] = i[54239];
  assign o[54238] = i[54238];
  assign o[54237] = i[54237];
  assign o[54236] = i[54236];
  assign o[54235] = i[54235];
  assign o[54234] = i[54234];
  assign o[54233] = i[54233];
  assign o[54232] = i[54232];
  assign o[54231] = i[54231];
  assign o[54230] = i[54230];
  assign o[54229] = i[54229];
  assign o[54228] = i[54228];
  assign o[54227] = i[54227];
  assign o[54226] = i[54226];
  assign o[54225] = i[54225];
  assign o[54224] = i[54224];
  assign o[54223] = i[54223];
  assign o[54222] = i[54222];
  assign o[54221] = i[54221];
  assign o[54220] = i[54220];
  assign o[54219] = i[54219];
  assign o[54218] = i[54218];
  assign o[54217] = i[54217];
  assign o[54216] = i[54216];
  assign o[54215] = i[54215];
  assign o[54214] = i[54214];
  assign o[54213] = i[54213];
  assign o[54212] = i[54212];
  assign o[54211] = i[54211];
  assign o[54210] = i[54210];
  assign o[54209] = i[54209];
  assign o[54208] = i[54208];
  assign o[54207] = i[54207];
  assign o[54206] = i[54206];
  assign o[54205] = i[54205];
  assign o[54204] = i[54204];
  assign o[54203] = i[54203];
  assign o[54202] = i[54202];
  assign o[54201] = i[54201];
  assign o[54200] = i[54200];
  assign o[54199] = i[54199];
  assign o[54198] = i[54198];
  assign o[54197] = i[54197];
  assign o[54196] = i[54196];
  assign o[54195] = i[54195];
  assign o[54194] = i[54194];
  assign o[54193] = i[54193];
  assign o[54192] = i[54192];
  assign o[54191] = i[54191];
  assign o[54190] = i[54190];
  assign o[54189] = i[54189];
  assign o[54188] = i[54188];
  assign o[54187] = i[54187];
  assign o[54186] = i[54186];
  assign o[54185] = i[54185];
  assign o[54184] = i[54184];
  assign o[54183] = i[54183];
  assign o[54182] = i[54182];
  assign o[54181] = i[54181];
  assign o[54180] = i[54180];
  assign o[54179] = i[54179];
  assign o[54178] = i[54178];
  assign o[54177] = i[54177];
  assign o[54176] = i[54176];
  assign o[54175] = i[54175];
  assign o[54174] = i[54174];
  assign o[54173] = i[54173];
  assign o[54172] = i[54172];
  assign o[54171] = i[54171];
  assign o[54170] = i[54170];
  assign o[54169] = i[54169];
  assign o[54168] = i[54168];
  assign o[54167] = i[54167];
  assign o[54166] = i[54166];
  assign o[54165] = i[54165];
  assign o[54164] = i[54164];
  assign o[54163] = i[54163];
  assign o[54162] = i[54162];
  assign o[54161] = i[54161];
  assign o[54160] = i[54160];
  assign o[54159] = i[54159];
  assign o[54158] = i[54158];
  assign o[54157] = i[54157];
  assign o[54156] = i[54156];
  assign o[54155] = i[54155];
  assign o[54154] = i[54154];
  assign o[54153] = i[54153];
  assign o[54152] = i[54152];
  assign o[54151] = i[54151];
  assign o[54150] = i[54150];
  assign o[54149] = i[54149];
  assign o[54148] = i[54148];
  assign o[54147] = i[54147];
  assign o[54146] = i[54146];
  assign o[54145] = i[54145];
  assign o[54144] = i[54144];
  assign o[54143] = i[54143];
  assign o[54142] = i[54142];
  assign o[54141] = i[54141];
  assign o[54140] = i[54140];
  assign o[54139] = i[54139];
  assign o[54138] = i[54138];
  assign o[54137] = i[54137];
  assign o[54136] = i[54136];
  assign o[54135] = i[54135];
  assign o[54134] = i[54134];
  assign o[54133] = i[54133];
  assign o[54132] = i[54132];
  assign o[54131] = i[54131];
  assign o[54130] = i[54130];
  assign o[54129] = i[54129];
  assign o[54128] = i[54128];
  assign o[54127] = i[54127];
  assign o[54126] = i[54126];
  assign o[54125] = i[54125];
  assign o[54124] = i[54124];
  assign o[54123] = i[54123];
  assign o[54122] = i[54122];
  assign o[54121] = i[54121];
  assign o[54120] = i[54120];
  assign o[54119] = i[54119];
  assign o[54118] = i[54118];
  assign o[54117] = i[54117];
  assign o[54116] = i[54116];
  assign o[54115] = i[54115];
  assign o[54114] = i[54114];
  assign o[54113] = i[54113];
  assign o[54112] = i[54112];
  assign o[54111] = i[54111];
  assign o[54110] = i[54110];
  assign o[54109] = i[54109];
  assign o[54108] = i[54108];
  assign o[54107] = i[54107];
  assign o[54106] = i[54106];
  assign o[54105] = i[54105];
  assign o[54104] = i[54104];
  assign o[54103] = i[54103];
  assign o[54102] = i[54102];
  assign o[54101] = i[54101];
  assign o[54100] = i[54100];
  assign o[54099] = i[54099];
  assign o[54098] = i[54098];
  assign o[54097] = i[54097];
  assign o[54096] = i[54096];
  assign o[54095] = i[54095];
  assign o[54094] = i[54094];
  assign o[54093] = i[54093];
  assign o[54092] = i[54092];
  assign o[54091] = i[54091];
  assign o[54090] = i[54090];
  assign o[54089] = i[54089];
  assign o[54088] = i[54088];
  assign o[54087] = i[54087];
  assign o[54086] = i[54086];
  assign o[54085] = i[54085];
  assign o[54084] = i[54084];
  assign o[54083] = i[54083];
  assign o[54082] = i[54082];
  assign o[54081] = i[54081];
  assign o[54080] = i[54080];
  assign o[54079] = i[54079];
  assign o[54078] = i[54078];
  assign o[54077] = i[54077];
  assign o[54076] = i[54076];
  assign o[54075] = i[54075];
  assign o[54074] = i[54074];
  assign o[54073] = i[54073];
  assign o[54072] = i[54072];
  assign o[54071] = i[54071];
  assign o[54070] = i[54070];
  assign o[54069] = i[54069];
  assign o[54068] = i[54068];
  assign o[54067] = i[54067];
  assign o[54066] = i[54066];
  assign o[54065] = i[54065];
  assign o[54064] = i[54064];
  assign o[54063] = i[54063];
  assign o[54062] = i[54062];
  assign o[54061] = i[54061];
  assign o[54060] = i[54060];
  assign o[54059] = i[54059];
  assign o[54058] = i[54058];
  assign o[54057] = i[54057];
  assign o[54056] = i[54056];
  assign o[54055] = i[54055];
  assign o[54054] = i[54054];
  assign o[54053] = i[54053];
  assign o[54052] = i[54052];
  assign o[54051] = i[54051];
  assign o[54050] = i[54050];
  assign o[54049] = i[54049];
  assign o[54048] = i[54048];
  assign o[54047] = i[54047];
  assign o[54046] = i[54046];
  assign o[54045] = i[54045];
  assign o[54044] = i[54044];
  assign o[54043] = i[54043];
  assign o[54042] = i[54042];
  assign o[54041] = i[54041];
  assign o[54040] = i[54040];
  assign o[54039] = i[54039];
  assign o[54038] = i[54038];
  assign o[54037] = i[54037];
  assign o[54036] = i[54036];
  assign o[54035] = i[54035];
  assign o[54034] = i[54034];
  assign o[54033] = i[54033];
  assign o[54032] = i[54032];
  assign o[54031] = i[54031];
  assign o[54030] = i[54030];
  assign o[54029] = i[54029];
  assign o[54028] = i[54028];
  assign o[54027] = i[54027];
  assign o[54026] = i[54026];
  assign o[54025] = i[54025];
  assign o[54024] = i[54024];
  assign o[54023] = i[54023];
  assign o[54022] = i[54022];
  assign o[54021] = i[54021];
  assign o[54020] = i[54020];
  assign o[54019] = i[54019];
  assign o[54018] = i[54018];
  assign o[54017] = i[54017];
  assign o[54016] = i[54016];
  assign o[54015] = i[54015];
  assign o[54014] = i[54014];
  assign o[54013] = i[54013];
  assign o[54012] = i[54012];
  assign o[54011] = i[54011];
  assign o[54010] = i[54010];
  assign o[54009] = i[54009];
  assign o[54008] = i[54008];
  assign o[54007] = i[54007];
  assign o[54006] = i[54006];
  assign o[54005] = i[54005];
  assign o[54004] = i[54004];
  assign o[54003] = i[54003];
  assign o[54002] = i[54002];
  assign o[54001] = i[54001];
  assign o[54000] = i[54000];
  assign o[53999] = i[53999];
  assign o[53998] = i[53998];
  assign o[53997] = i[53997];
  assign o[53996] = i[53996];
  assign o[53995] = i[53995];
  assign o[53994] = i[53994];
  assign o[53993] = i[53993];
  assign o[53992] = i[53992];
  assign o[53991] = i[53991];
  assign o[53990] = i[53990];
  assign o[53989] = i[53989];
  assign o[53988] = i[53988];
  assign o[53987] = i[53987];
  assign o[53986] = i[53986];
  assign o[53985] = i[53985];
  assign o[53984] = i[53984];
  assign o[53983] = i[53983];
  assign o[53982] = i[53982];
  assign o[53981] = i[53981];
  assign o[53980] = i[53980];
  assign o[53979] = i[53979];
  assign o[53978] = i[53978];
  assign o[53977] = i[53977];
  assign o[53976] = i[53976];
  assign o[53975] = i[53975];
  assign o[53974] = i[53974];
  assign o[53973] = i[53973];
  assign o[53972] = i[53972];
  assign o[53971] = i[53971];
  assign o[53970] = i[53970];
  assign o[53969] = i[53969];
  assign o[53968] = i[53968];
  assign o[53967] = i[53967];
  assign o[53966] = i[53966];
  assign o[53965] = i[53965];
  assign o[53964] = i[53964];
  assign o[53963] = i[53963];
  assign o[53962] = i[53962];
  assign o[53961] = i[53961];
  assign o[53960] = i[53960];
  assign o[53959] = i[53959];
  assign o[53958] = i[53958];
  assign o[53957] = i[53957];
  assign o[53956] = i[53956];
  assign o[53955] = i[53955];
  assign o[53954] = i[53954];
  assign o[53953] = i[53953];
  assign o[53952] = i[53952];
  assign o[53951] = i[53951];
  assign o[53950] = i[53950];
  assign o[53949] = i[53949];
  assign o[53948] = i[53948];
  assign o[53947] = i[53947];
  assign o[53946] = i[53946];
  assign o[53945] = i[53945];
  assign o[53944] = i[53944];
  assign o[53943] = i[53943];
  assign o[53942] = i[53942];
  assign o[53941] = i[53941];
  assign o[53940] = i[53940];
  assign o[53939] = i[53939];
  assign o[53938] = i[53938];
  assign o[53937] = i[53937];
  assign o[53936] = i[53936];
  assign o[53935] = i[53935];
  assign o[53934] = i[53934];
  assign o[53933] = i[53933];
  assign o[53932] = i[53932];
  assign o[53931] = i[53931];
  assign o[53930] = i[53930];
  assign o[53929] = i[53929];
  assign o[53928] = i[53928];
  assign o[53927] = i[53927];
  assign o[53926] = i[53926];
  assign o[53925] = i[53925];
  assign o[53924] = i[53924];
  assign o[53923] = i[53923];
  assign o[53922] = i[53922];
  assign o[53921] = i[53921];
  assign o[53920] = i[53920];
  assign o[53919] = i[53919];
  assign o[53918] = i[53918];
  assign o[53917] = i[53917];
  assign o[53916] = i[53916];
  assign o[53915] = i[53915];
  assign o[53914] = i[53914];
  assign o[53913] = i[53913];
  assign o[53912] = i[53912];
  assign o[53911] = i[53911];
  assign o[53910] = i[53910];
  assign o[53909] = i[53909];
  assign o[53908] = i[53908];
  assign o[53907] = i[53907];
  assign o[53906] = i[53906];
  assign o[53905] = i[53905];
  assign o[53904] = i[53904];
  assign o[53903] = i[53903];
  assign o[53902] = i[53902];
  assign o[53901] = i[53901];
  assign o[53900] = i[53900];
  assign o[53899] = i[53899];
  assign o[53898] = i[53898];
  assign o[53897] = i[53897];
  assign o[53896] = i[53896];
  assign o[53895] = i[53895];
  assign o[53894] = i[53894];
  assign o[53893] = i[53893];
  assign o[53892] = i[53892];
  assign o[53891] = i[53891];
  assign o[53890] = i[53890];
  assign o[53889] = i[53889];
  assign o[53888] = i[53888];
  assign o[53887] = i[53887];
  assign o[53886] = i[53886];
  assign o[53885] = i[53885];
  assign o[53884] = i[53884];
  assign o[53883] = i[53883];
  assign o[53882] = i[53882];
  assign o[53881] = i[53881];
  assign o[53880] = i[53880];
  assign o[53879] = i[53879];
  assign o[53878] = i[53878];
  assign o[53877] = i[53877];
  assign o[53876] = i[53876];
  assign o[53875] = i[53875];
  assign o[53874] = i[53874];
  assign o[53873] = i[53873];
  assign o[53872] = i[53872];
  assign o[53871] = i[53871];
  assign o[53870] = i[53870];
  assign o[53869] = i[53869];
  assign o[53868] = i[53868];
  assign o[53867] = i[53867];
  assign o[53866] = i[53866];
  assign o[53865] = i[53865];
  assign o[53864] = i[53864];
  assign o[53863] = i[53863];
  assign o[53862] = i[53862];
  assign o[53861] = i[53861];
  assign o[53860] = i[53860];
  assign o[53859] = i[53859];
  assign o[53858] = i[53858];
  assign o[53857] = i[53857];
  assign o[53856] = i[53856];
  assign o[53855] = i[53855];
  assign o[53854] = i[53854];
  assign o[53853] = i[53853];
  assign o[53852] = i[53852];
  assign o[53851] = i[53851];
  assign o[53850] = i[53850];
  assign o[53849] = i[53849];
  assign o[53848] = i[53848];
  assign o[53847] = i[53847];
  assign o[53846] = i[53846];
  assign o[53845] = i[53845];
  assign o[53844] = i[53844];
  assign o[53843] = i[53843];
  assign o[53842] = i[53842];
  assign o[53841] = i[53841];
  assign o[53840] = i[53840];
  assign o[53839] = i[53839];
  assign o[53838] = i[53838];
  assign o[53837] = i[53837];
  assign o[53836] = i[53836];
  assign o[53835] = i[53835];
  assign o[53834] = i[53834];
  assign o[53833] = i[53833];
  assign o[53832] = i[53832];
  assign o[53831] = i[53831];
  assign o[53830] = i[53830];
  assign o[53829] = i[53829];
  assign o[53828] = i[53828];
  assign o[53827] = i[53827];
  assign o[53826] = i[53826];
  assign o[53825] = i[53825];
  assign o[53824] = i[53824];
  assign o[53823] = i[53823];
  assign o[53822] = i[53822];
  assign o[53821] = i[53821];
  assign o[53820] = i[53820];
  assign o[53819] = i[53819];
  assign o[53818] = i[53818];
  assign o[53817] = i[53817];
  assign o[53816] = i[53816];
  assign o[53815] = i[53815];
  assign o[53814] = i[53814];
  assign o[53813] = i[53813];
  assign o[53812] = i[53812];
  assign o[53811] = i[53811];
  assign o[53810] = i[53810];
  assign o[53809] = i[53809];
  assign o[53808] = i[53808];
  assign o[53807] = i[53807];
  assign o[53806] = i[53806];
  assign o[53805] = i[53805];
  assign o[53804] = i[53804];
  assign o[53803] = i[53803];
  assign o[53802] = i[53802];
  assign o[53801] = i[53801];
  assign o[53800] = i[53800];
  assign o[53799] = i[53799];
  assign o[53798] = i[53798];
  assign o[53797] = i[53797];
  assign o[53796] = i[53796];
  assign o[53795] = i[53795];
  assign o[53794] = i[53794];
  assign o[53793] = i[53793];
  assign o[53792] = i[53792];
  assign o[53791] = i[53791];
  assign o[53790] = i[53790];
  assign o[53789] = i[53789];
  assign o[53788] = i[53788];
  assign o[53787] = i[53787];
  assign o[53786] = i[53786];
  assign o[53785] = i[53785];
  assign o[53784] = i[53784];
  assign o[53783] = i[53783];
  assign o[53782] = i[53782];
  assign o[53781] = i[53781];
  assign o[53780] = i[53780];
  assign o[53779] = i[53779];
  assign o[53778] = i[53778];
  assign o[53777] = i[53777];
  assign o[53776] = i[53776];
  assign o[53775] = i[53775];
  assign o[53774] = i[53774];
  assign o[53773] = i[53773];
  assign o[53772] = i[53772];
  assign o[53771] = i[53771];
  assign o[53770] = i[53770];
  assign o[53769] = i[53769];
  assign o[53768] = i[53768];
  assign o[53767] = i[53767];
  assign o[53766] = i[53766];
  assign o[53765] = i[53765];
  assign o[53764] = i[53764];
  assign o[53763] = i[53763];
  assign o[53762] = i[53762];
  assign o[53761] = i[53761];
  assign o[53760] = i[53760];
  assign o[53759] = i[53759];
  assign o[53758] = i[53758];
  assign o[53757] = i[53757];
  assign o[53756] = i[53756];
  assign o[53755] = i[53755];
  assign o[53754] = i[53754];
  assign o[53753] = i[53753];
  assign o[53752] = i[53752];
  assign o[53751] = i[53751];
  assign o[53750] = i[53750];
  assign o[53749] = i[53749];
  assign o[53748] = i[53748];
  assign o[53747] = i[53747];
  assign o[53746] = i[53746];
  assign o[53745] = i[53745];
  assign o[53744] = i[53744];
  assign o[53743] = i[53743];
  assign o[53742] = i[53742];
  assign o[53741] = i[53741];
  assign o[53740] = i[53740];
  assign o[53739] = i[53739];
  assign o[53738] = i[53738];
  assign o[53737] = i[53737];
  assign o[53736] = i[53736];
  assign o[53735] = i[53735];
  assign o[53734] = i[53734];
  assign o[53733] = i[53733];
  assign o[53732] = i[53732];
  assign o[53731] = i[53731];
  assign o[53730] = i[53730];
  assign o[53729] = i[53729];
  assign o[53728] = i[53728];
  assign o[53727] = i[53727];
  assign o[53726] = i[53726];
  assign o[53725] = i[53725];
  assign o[53724] = i[53724];
  assign o[53723] = i[53723];
  assign o[53722] = i[53722];
  assign o[53721] = i[53721];
  assign o[53720] = i[53720];
  assign o[53719] = i[53719];
  assign o[53718] = i[53718];
  assign o[53717] = i[53717];
  assign o[53716] = i[53716];
  assign o[53715] = i[53715];
  assign o[53714] = i[53714];
  assign o[53713] = i[53713];
  assign o[53712] = i[53712];
  assign o[53711] = i[53711];
  assign o[53710] = i[53710];
  assign o[53709] = i[53709];
  assign o[53708] = i[53708];
  assign o[53707] = i[53707];
  assign o[53706] = i[53706];
  assign o[53705] = i[53705];
  assign o[53704] = i[53704];
  assign o[53703] = i[53703];
  assign o[53702] = i[53702];
  assign o[53701] = i[53701];
  assign o[53700] = i[53700];
  assign o[53699] = i[53699];
  assign o[53698] = i[53698];
  assign o[53697] = i[53697];
  assign o[53696] = i[53696];
  assign o[53695] = i[53695];
  assign o[53694] = i[53694];
  assign o[53693] = i[53693];
  assign o[53692] = i[53692];
  assign o[53691] = i[53691];
  assign o[53690] = i[53690];
  assign o[53689] = i[53689];
  assign o[53688] = i[53688];
  assign o[53687] = i[53687];
  assign o[53686] = i[53686];
  assign o[53685] = i[53685];
  assign o[53684] = i[53684];
  assign o[53683] = i[53683];
  assign o[53682] = i[53682];
  assign o[53681] = i[53681];
  assign o[53680] = i[53680];
  assign o[53679] = i[53679];
  assign o[53678] = i[53678];
  assign o[53677] = i[53677];
  assign o[53676] = i[53676];
  assign o[53675] = i[53675];
  assign o[53674] = i[53674];
  assign o[53673] = i[53673];
  assign o[53672] = i[53672];
  assign o[53671] = i[53671];
  assign o[53670] = i[53670];
  assign o[53669] = i[53669];
  assign o[53668] = i[53668];
  assign o[53667] = i[53667];
  assign o[53666] = i[53666];
  assign o[53665] = i[53665];
  assign o[53664] = i[53664];
  assign o[53663] = i[53663];
  assign o[53662] = i[53662];
  assign o[53661] = i[53661];
  assign o[53660] = i[53660];
  assign o[53659] = i[53659];
  assign o[53658] = i[53658];
  assign o[53657] = i[53657];
  assign o[53656] = i[53656];
  assign o[53655] = i[53655];
  assign o[53654] = i[53654];
  assign o[53653] = i[53653];
  assign o[53652] = i[53652];
  assign o[53651] = i[53651];
  assign o[53650] = i[53650];
  assign o[53649] = i[53649];
  assign o[53648] = i[53648];
  assign o[53647] = i[53647];
  assign o[53646] = i[53646];
  assign o[53645] = i[53645];
  assign o[53644] = i[53644];
  assign o[53643] = i[53643];
  assign o[53642] = i[53642];
  assign o[53641] = i[53641];
  assign o[53640] = i[53640];
  assign o[53639] = i[53639];
  assign o[53638] = i[53638];
  assign o[53637] = i[53637];
  assign o[53636] = i[53636];
  assign o[53635] = i[53635];
  assign o[53634] = i[53634];
  assign o[53633] = i[53633];
  assign o[53632] = i[53632];
  assign o[53631] = i[53631];
  assign o[53630] = i[53630];
  assign o[53629] = i[53629];
  assign o[53628] = i[53628];
  assign o[53627] = i[53627];
  assign o[53626] = i[53626];
  assign o[53625] = i[53625];
  assign o[53624] = i[53624];
  assign o[53623] = i[53623];
  assign o[53622] = i[53622];
  assign o[53621] = i[53621];
  assign o[53620] = i[53620];
  assign o[53619] = i[53619];
  assign o[53618] = i[53618];
  assign o[53617] = i[53617];
  assign o[53616] = i[53616];
  assign o[53615] = i[53615];
  assign o[53614] = i[53614];
  assign o[53613] = i[53613];
  assign o[53612] = i[53612];
  assign o[53611] = i[53611];
  assign o[53610] = i[53610];
  assign o[53609] = i[53609];
  assign o[53608] = i[53608];
  assign o[53607] = i[53607];
  assign o[53606] = i[53606];
  assign o[53605] = i[53605];
  assign o[53604] = i[53604];
  assign o[53603] = i[53603];
  assign o[53602] = i[53602];
  assign o[53601] = i[53601];
  assign o[53600] = i[53600];
  assign o[53599] = i[53599];
  assign o[53598] = i[53598];
  assign o[53597] = i[53597];
  assign o[53596] = i[53596];
  assign o[53595] = i[53595];
  assign o[53594] = i[53594];
  assign o[53593] = i[53593];
  assign o[53592] = i[53592];
  assign o[53591] = i[53591];
  assign o[53590] = i[53590];
  assign o[53589] = i[53589];
  assign o[53588] = i[53588];
  assign o[53587] = i[53587];
  assign o[53586] = i[53586];
  assign o[53585] = i[53585];
  assign o[53584] = i[53584];
  assign o[53583] = i[53583];
  assign o[53582] = i[53582];
  assign o[53581] = i[53581];
  assign o[53580] = i[53580];
  assign o[53579] = i[53579];
  assign o[53578] = i[53578];
  assign o[53577] = i[53577];
  assign o[53576] = i[53576];
  assign o[53575] = i[53575];
  assign o[53574] = i[53574];
  assign o[53573] = i[53573];
  assign o[53572] = i[53572];
  assign o[53571] = i[53571];
  assign o[53570] = i[53570];
  assign o[53569] = i[53569];
  assign o[53568] = i[53568];
  assign o[53567] = i[53567];
  assign o[53566] = i[53566];
  assign o[53565] = i[53565];
  assign o[53564] = i[53564];
  assign o[53563] = i[53563];
  assign o[53562] = i[53562];
  assign o[53561] = i[53561];
  assign o[53560] = i[53560];
  assign o[53559] = i[53559];
  assign o[53558] = i[53558];
  assign o[53557] = i[53557];
  assign o[53556] = i[53556];
  assign o[53555] = i[53555];
  assign o[53554] = i[53554];
  assign o[53553] = i[53553];
  assign o[53552] = i[53552];
  assign o[53551] = i[53551];
  assign o[53550] = i[53550];
  assign o[53549] = i[53549];
  assign o[53548] = i[53548];
  assign o[53547] = i[53547];
  assign o[53546] = i[53546];
  assign o[53545] = i[53545];
  assign o[53544] = i[53544];
  assign o[53543] = i[53543];
  assign o[53542] = i[53542];
  assign o[53541] = i[53541];
  assign o[53540] = i[53540];
  assign o[53539] = i[53539];
  assign o[53538] = i[53538];
  assign o[53537] = i[53537];
  assign o[53536] = i[53536];
  assign o[53535] = i[53535];
  assign o[53534] = i[53534];
  assign o[53533] = i[53533];
  assign o[53532] = i[53532];
  assign o[53531] = i[53531];
  assign o[53530] = i[53530];
  assign o[53529] = i[53529];
  assign o[53528] = i[53528];
  assign o[53527] = i[53527];
  assign o[53526] = i[53526];
  assign o[53525] = i[53525];
  assign o[53524] = i[53524];
  assign o[53523] = i[53523];
  assign o[53522] = i[53522];
  assign o[53521] = i[53521];
  assign o[53520] = i[53520];
  assign o[53519] = i[53519];
  assign o[53518] = i[53518];
  assign o[53517] = i[53517];
  assign o[53516] = i[53516];
  assign o[53515] = i[53515];
  assign o[53514] = i[53514];
  assign o[53513] = i[53513];
  assign o[53512] = i[53512];
  assign o[53511] = i[53511];
  assign o[53510] = i[53510];
  assign o[53509] = i[53509];
  assign o[53508] = i[53508];
  assign o[53507] = i[53507];
  assign o[53506] = i[53506];
  assign o[53505] = i[53505];
  assign o[53504] = i[53504];
  assign o[53503] = i[53503];
  assign o[53502] = i[53502];
  assign o[53501] = i[53501];
  assign o[53500] = i[53500];
  assign o[53499] = i[53499];
  assign o[53498] = i[53498];
  assign o[53497] = i[53497];
  assign o[53496] = i[53496];
  assign o[53495] = i[53495];
  assign o[53494] = i[53494];
  assign o[53493] = i[53493];
  assign o[53492] = i[53492];
  assign o[53491] = i[53491];
  assign o[53490] = i[53490];
  assign o[53489] = i[53489];
  assign o[53488] = i[53488];
  assign o[53487] = i[53487];
  assign o[53486] = i[53486];
  assign o[53485] = i[53485];
  assign o[53484] = i[53484];
  assign o[53483] = i[53483];
  assign o[53482] = i[53482];
  assign o[53481] = i[53481];
  assign o[53480] = i[53480];
  assign o[53479] = i[53479];
  assign o[53478] = i[53478];
  assign o[53477] = i[53477];
  assign o[53476] = i[53476];
  assign o[53475] = i[53475];
  assign o[53474] = i[53474];
  assign o[53473] = i[53473];
  assign o[53472] = i[53472];
  assign o[53471] = i[53471];
  assign o[53470] = i[53470];
  assign o[53469] = i[53469];
  assign o[53468] = i[53468];
  assign o[53467] = i[53467];
  assign o[53466] = i[53466];
  assign o[53465] = i[53465];
  assign o[53464] = i[53464];
  assign o[53463] = i[53463];
  assign o[53462] = i[53462];
  assign o[53461] = i[53461];
  assign o[53460] = i[53460];
  assign o[53459] = i[53459];
  assign o[53458] = i[53458];
  assign o[53457] = i[53457];
  assign o[53456] = i[53456];
  assign o[53455] = i[53455];
  assign o[53454] = i[53454];
  assign o[53453] = i[53453];
  assign o[53452] = i[53452];
  assign o[53451] = i[53451];
  assign o[53450] = i[53450];
  assign o[53449] = i[53449];
  assign o[53448] = i[53448];
  assign o[53447] = i[53447];
  assign o[53446] = i[53446];
  assign o[53445] = i[53445];
  assign o[53444] = i[53444];
  assign o[53443] = i[53443];
  assign o[53442] = i[53442];
  assign o[53441] = i[53441];
  assign o[53440] = i[53440];
  assign o[53439] = i[53439];
  assign o[53438] = i[53438];
  assign o[53437] = i[53437];
  assign o[53436] = i[53436];
  assign o[53435] = i[53435];
  assign o[53434] = i[53434];
  assign o[53433] = i[53433];
  assign o[53432] = i[53432];
  assign o[53431] = i[53431];
  assign o[53430] = i[53430];
  assign o[53429] = i[53429];
  assign o[53428] = i[53428];
  assign o[53427] = i[53427];
  assign o[53426] = i[53426];
  assign o[53425] = i[53425];
  assign o[53424] = i[53424];
  assign o[53423] = i[53423];
  assign o[53422] = i[53422];
  assign o[53421] = i[53421];
  assign o[53420] = i[53420];
  assign o[53419] = i[53419];
  assign o[53418] = i[53418];
  assign o[53417] = i[53417];
  assign o[53416] = i[53416];
  assign o[53415] = i[53415];
  assign o[53414] = i[53414];
  assign o[53413] = i[53413];
  assign o[53412] = i[53412];
  assign o[53411] = i[53411];
  assign o[53410] = i[53410];
  assign o[53409] = i[53409];
  assign o[53408] = i[53408];
  assign o[53407] = i[53407];
  assign o[53406] = i[53406];
  assign o[53405] = i[53405];
  assign o[53404] = i[53404];
  assign o[53403] = i[53403];
  assign o[53402] = i[53402];
  assign o[53401] = i[53401];
  assign o[53400] = i[53400];
  assign o[53399] = i[53399];
  assign o[53398] = i[53398];
  assign o[53397] = i[53397];
  assign o[53396] = i[53396];
  assign o[53395] = i[53395];
  assign o[53394] = i[53394];
  assign o[53393] = i[53393];
  assign o[53392] = i[53392];
  assign o[53391] = i[53391];
  assign o[53390] = i[53390];
  assign o[53389] = i[53389];
  assign o[53388] = i[53388];
  assign o[53387] = i[53387];
  assign o[53386] = i[53386];
  assign o[53385] = i[53385];
  assign o[53384] = i[53384];
  assign o[53383] = i[53383];
  assign o[53382] = i[53382];
  assign o[53381] = i[53381];
  assign o[53380] = i[53380];
  assign o[53379] = i[53379];
  assign o[53378] = i[53378];
  assign o[53377] = i[53377];
  assign o[53376] = i[53376];
  assign o[53375] = i[53375];
  assign o[53374] = i[53374];
  assign o[53373] = i[53373];
  assign o[53372] = i[53372];
  assign o[53371] = i[53371];
  assign o[53370] = i[53370];
  assign o[53369] = i[53369];
  assign o[53368] = i[53368];
  assign o[53367] = i[53367];
  assign o[53366] = i[53366];
  assign o[53365] = i[53365];
  assign o[53364] = i[53364];
  assign o[53363] = i[53363];
  assign o[53362] = i[53362];
  assign o[53361] = i[53361];
  assign o[53360] = i[53360];
  assign o[53359] = i[53359];
  assign o[53358] = i[53358];
  assign o[53357] = i[53357];
  assign o[53356] = i[53356];
  assign o[53355] = i[53355];
  assign o[53354] = i[53354];
  assign o[53353] = i[53353];
  assign o[53352] = i[53352];
  assign o[53351] = i[53351];
  assign o[53350] = i[53350];
  assign o[53349] = i[53349];
  assign o[53348] = i[53348];
  assign o[53347] = i[53347];
  assign o[53346] = i[53346];
  assign o[53345] = i[53345];
  assign o[53344] = i[53344];
  assign o[53343] = i[53343];
  assign o[53342] = i[53342];
  assign o[53341] = i[53341];
  assign o[53340] = i[53340];
  assign o[53339] = i[53339];
  assign o[53338] = i[53338];
  assign o[53337] = i[53337];
  assign o[53336] = i[53336];
  assign o[53335] = i[53335];
  assign o[53334] = i[53334];
  assign o[53333] = i[53333];
  assign o[53332] = i[53332];
  assign o[53331] = i[53331];
  assign o[53330] = i[53330];
  assign o[53329] = i[53329];
  assign o[53328] = i[53328];
  assign o[53327] = i[53327];
  assign o[53326] = i[53326];
  assign o[53325] = i[53325];
  assign o[53324] = i[53324];
  assign o[53323] = i[53323];
  assign o[53322] = i[53322];
  assign o[53321] = i[53321];
  assign o[53320] = i[53320];
  assign o[53319] = i[53319];
  assign o[53318] = i[53318];
  assign o[53317] = i[53317];
  assign o[53316] = i[53316];
  assign o[53315] = i[53315];
  assign o[53314] = i[53314];
  assign o[53313] = i[53313];
  assign o[53312] = i[53312];
  assign o[53311] = i[53311];
  assign o[53310] = i[53310];
  assign o[53309] = i[53309];
  assign o[53308] = i[53308];
  assign o[53307] = i[53307];
  assign o[53306] = i[53306];
  assign o[53305] = i[53305];
  assign o[53304] = i[53304];
  assign o[53303] = i[53303];
  assign o[53302] = i[53302];
  assign o[53301] = i[53301];
  assign o[53300] = i[53300];
  assign o[53299] = i[53299];
  assign o[53298] = i[53298];
  assign o[53297] = i[53297];
  assign o[53296] = i[53296];
  assign o[53295] = i[53295];
  assign o[53294] = i[53294];
  assign o[53293] = i[53293];
  assign o[53292] = i[53292];
  assign o[53291] = i[53291];
  assign o[53290] = i[53290];
  assign o[53289] = i[53289];
  assign o[53288] = i[53288];
  assign o[53287] = i[53287];
  assign o[53286] = i[53286];
  assign o[53285] = i[53285];
  assign o[53284] = i[53284];
  assign o[53283] = i[53283];
  assign o[53282] = i[53282];
  assign o[53281] = i[53281];
  assign o[53280] = i[53280];
  assign o[53279] = i[53279];
  assign o[53278] = i[53278];
  assign o[53277] = i[53277];
  assign o[53276] = i[53276];
  assign o[53275] = i[53275];
  assign o[53274] = i[53274];
  assign o[53273] = i[53273];
  assign o[53272] = i[53272];
  assign o[53271] = i[53271];
  assign o[53270] = i[53270];
  assign o[53269] = i[53269];
  assign o[53268] = i[53268];
  assign o[53267] = i[53267];
  assign o[53266] = i[53266];
  assign o[53265] = i[53265];
  assign o[53264] = i[53264];
  assign o[53263] = i[53263];
  assign o[53262] = i[53262];
  assign o[53261] = i[53261];
  assign o[53260] = i[53260];
  assign o[53259] = i[53259];
  assign o[53258] = i[53258];
  assign o[53257] = i[53257];
  assign o[53256] = i[53256];
  assign o[53255] = i[53255];
  assign o[53254] = i[53254];
  assign o[53253] = i[53253];
  assign o[53252] = i[53252];
  assign o[53251] = i[53251];
  assign o[53250] = i[53250];
  assign o[53249] = i[53249];
  assign o[53248] = i[53248];
  assign o[53247] = i[53247];
  assign o[53246] = i[53246];
  assign o[53245] = i[53245];
  assign o[53244] = i[53244];
  assign o[53243] = i[53243];
  assign o[53242] = i[53242];
  assign o[53241] = i[53241];
  assign o[53240] = i[53240];
  assign o[53239] = i[53239];
  assign o[53238] = i[53238];
  assign o[53237] = i[53237];
  assign o[53236] = i[53236];
  assign o[53235] = i[53235];
  assign o[53234] = i[53234];
  assign o[53233] = i[53233];
  assign o[53232] = i[53232];
  assign o[53231] = i[53231];
  assign o[53230] = i[53230];
  assign o[53229] = i[53229];
  assign o[53228] = i[53228];
  assign o[53227] = i[53227];
  assign o[53226] = i[53226];
  assign o[53225] = i[53225];
  assign o[53224] = i[53224];
  assign o[53223] = i[53223];
  assign o[53222] = i[53222];
  assign o[53221] = i[53221];
  assign o[53220] = i[53220];
  assign o[53219] = i[53219];
  assign o[53218] = i[53218];
  assign o[53217] = i[53217];
  assign o[53216] = i[53216];
  assign o[53215] = i[53215];
  assign o[53214] = i[53214];
  assign o[53213] = i[53213];
  assign o[53212] = i[53212];
  assign o[53211] = i[53211];
  assign o[53210] = i[53210];
  assign o[53209] = i[53209];
  assign o[53208] = i[53208];
  assign o[53207] = i[53207];
  assign o[53206] = i[53206];
  assign o[53205] = i[53205];
  assign o[53204] = i[53204];
  assign o[53203] = i[53203];
  assign o[53202] = i[53202];
  assign o[53201] = i[53201];
  assign o[53200] = i[53200];
  assign o[53199] = i[53199];
  assign o[53198] = i[53198];
  assign o[53197] = i[53197];
  assign o[53196] = i[53196];
  assign o[53195] = i[53195];
  assign o[53194] = i[53194];
  assign o[53193] = i[53193];
  assign o[53192] = i[53192];
  assign o[53191] = i[53191];
  assign o[53190] = i[53190];
  assign o[53189] = i[53189];
  assign o[53188] = i[53188];
  assign o[53187] = i[53187];
  assign o[53186] = i[53186];
  assign o[53185] = i[53185];
  assign o[53184] = i[53184];
  assign o[53183] = i[53183];
  assign o[53182] = i[53182];
  assign o[53181] = i[53181];
  assign o[53180] = i[53180];
  assign o[53179] = i[53179];
  assign o[53178] = i[53178];
  assign o[53177] = i[53177];
  assign o[53176] = i[53176];
  assign o[53175] = i[53175];
  assign o[53174] = i[53174];
  assign o[53173] = i[53173];
  assign o[53172] = i[53172];
  assign o[53171] = i[53171];
  assign o[53170] = i[53170];
  assign o[53169] = i[53169];
  assign o[53168] = i[53168];
  assign o[53167] = i[53167];
  assign o[53166] = i[53166];
  assign o[53165] = i[53165];
  assign o[53164] = i[53164];
  assign o[53163] = i[53163];
  assign o[53162] = i[53162];
  assign o[53161] = i[53161];
  assign o[53160] = i[53160];
  assign o[53159] = i[53159];
  assign o[53158] = i[53158];
  assign o[53157] = i[53157];
  assign o[53156] = i[53156];
  assign o[53155] = i[53155];
  assign o[53154] = i[53154];
  assign o[53153] = i[53153];
  assign o[53152] = i[53152];
  assign o[53151] = i[53151];
  assign o[53150] = i[53150];
  assign o[53149] = i[53149];
  assign o[53148] = i[53148];
  assign o[53147] = i[53147];
  assign o[53146] = i[53146];
  assign o[53145] = i[53145];
  assign o[53144] = i[53144];
  assign o[53143] = i[53143];
  assign o[53142] = i[53142];
  assign o[53141] = i[53141];
  assign o[53140] = i[53140];
  assign o[53139] = i[53139];
  assign o[53138] = i[53138];
  assign o[53137] = i[53137];
  assign o[53136] = i[53136];
  assign o[53135] = i[53135];
  assign o[53134] = i[53134];
  assign o[53133] = i[53133];
  assign o[53132] = i[53132];
  assign o[53131] = i[53131];
  assign o[53130] = i[53130];
  assign o[53129] = i[53129];
  assign o[53128] = i[53128];
  assign o[53127] = i[53127];
  assign o[53126] = i[53126];
  assign o[53125] = i[53125];
  assign o[53124] = i[53124];
  assign o[53123] = i[53123];
  assign o[53122] = i[53122];
  assign o[53121] = i[53121];
  assign o[53120] = i[53120];
  assign o[53119] = i[53119];
  assign o[53118] = i[53118];
  assign o[53117] = i[53117];
  assign o[53116] = i[53116];
  assign o[53115] = i[53115];
  assign o[53114] = i[53114];
  assign o[53113] = i[53113];
  assign o[53112] = i[53112];
  assign o[53111] = i[53111];
  assign o[53110] = i[53110];
  assign o[53109] = i[53109];
  assign o[53108] = i[53108];
  assign o[53107] = i[53107];
  assign o[53106] = i[53106];
  assign o[53105] = i[53105];
  assign o[53104] = i[53104];
  assign o[53103] = i[53103];
  assign o[53102] = i[53102];
  assign o[53101] = i[53101];
  assign o[53100] = i[53100];
  assign o[53099] = i[53099];
  assign o[53098] = i[53098];
  assign o[53097] = i[53097];
  assign o[53096] = i[53096];
  assign o[53095] = i[53095];
  assign o[53094] = i[53094];
  assign o[53093] = i[53093];
  assign o[53092] = i[53092];
  assign o[53091] = i[53091];
  assign o[53090] = i[53090];
  assign o[53089] = i[53089];
  assign o[53088] = i[53088];
  assign o[53087] = i[53087];
  assign o[53086] = i[53086];
  assign o[53085] = i[53085];
  assign o[53084] = i[53084];
  assign o[53083] = i[53083];
  assign o[53082] = i[53082];
  assign o[53081] = i[53081];
  assign o[53080] = i[53080];
  assign o[53079] = i[53079];
  assign o[53078] = i[53078];
  assign o[53077] = i[53077];
  assign o[53076] = i[53076];
  assign o[53075] = i[53075];
  assign o[53074] = i[53074];
  assign o[53073] = i[53073];
  assign o[53072] = i[53072];
  assign o[53071] = i[53071];
  assign o[53070] = i[53070];
  assign o[53069] = i[53069];
  assign o[53068] = i[53068];
  assign o[53067] = i[53067];
  assign o[53066] = i[53066];
  assign o[53065] = i[53065];
  assign o[53064] = i[53064];
  assign o[53063] = i[53063];
  assign o[53062] = i[53062];
  assign o[53061] = i[53061];
  assign o[53060] = i[53060];
  assign o[53059] = i[53059];
  assign o[53058] = i[53058];
  assign o[53057] = i[53057];
  assign o[53056] = i[53056];
  assign o[53055] = i[53055];
  assign o[53054] = i[53054];
  assign o[53053] = i[53053];
  assign o[53052] = i[53052];
  assign o[53051] = i[53051];
  assign o[53050] = i[53050];
  assign o[53049] = i[53049];
  assign o[53048] = i[53048];
  assign o[53047] = i[53047];
  assign o[53046] = i[53046];
  assign o[53045] = i[53045];
  assign o[53044] = i[53044];
  assign o[53043] = i[53043];
  assign o[53042] = i[53042];
  assign o[53041] = i[53041];
  assign o[53040] = i[53040];
  assign o[53039] = i[53039];
  assign o[53038] = i[53038];
  assign o[53037] = i[53037];
  assign o[53036] = i[53036];
  assign o[53035] = i[53035];
  assign o[53034] = i[53034];
  assign o[53033] = i[53033];
  assign o[53032] = i[53032];
  assign o[53031] = i[53031];
  assign o[53030] = i[53030];
  assign o[53029] = i[53029];
  assign o[53028] = i[53028];
  assign o[53027] = i[53027];
  assign o[53026] = i[53026];
  assign o[53025] = i[53025];
  assign o[53024] = i[53024];
  assign o[53023] = i[53023];
  assign o[53022] = i[53022];
  assign o[53021] = i[53021];
  assign o[53020] = i[53020];
  assign o[53019] = i[53019];
  assign o[53018] = i[53018];
  assign o[53017] = i[53017];
  assign o[53016] = i[53016];
  assign o[53015] = i[53015];
  assign o[53014] = i[53014];
  assign o[53013] = i[53013];
  assign o[53012] = i[53012];
  assign o[53011] = i[53011];
  assign o[53010] = i[53010];
  assign o[53009] = i[53009];
  assign o[53008] = i[53008];
  assign o[53007] = i[53007];
  assign o[53006] = i[53006];
  assign o[53005] = i[53005];
  assign o[53004] = i[53004];
  assign o[53003] = i[53003];
  assign o[53002] = i[53002];
  assign o[53001] = i[53001];
  assign o[53000] = i[53000];
  assign o[52999] = i[52999];
  assign o[52998] = i[52998];
  assign o[52997] = i[52997];
  assign o[52996] = i[52996];
  assign o[52995] = i[52995];
  assign o[52994] = i[52994];
  assign o[52993] = i[52993];
  assign o[52992] = i[52992];
  assign o[52991] = i[52991];
  assign o[52990] = i[52990];
  assign o[52989] = i[52989];
  assign o[52988] = i[52988];
  assign o[52987] = i[52987];
  assign o[52986] = i[52986];
  assign o[52985] = i[52985];
  assign o[52984] = i[52984];
  assign o[52983] = i[52983];
  assign o[52982] = i[52982];
  assign o[52981] = i[52981];
  assign o[52980] = i[52980];
  assign o[52979] = i[52979];
  assign o[52978] = i[52978];
  assign o[52977] = i[52977];
  assign o[52976] = i[52976];
  assign o[52975] = i[52975];
  assign o[52974] = i[52974];
  assign o[52973] = i[52973];
  assign o[52972] = i[52972];
  assign o[52971] = i[52971];
  assign o[52970] = i[52970];
  assign o[52969] = i[52969];
  assign o[52968] = i[52968];
  assign o[52967] = i[52967];
  assign o[52966] = i[52966];
  assign o[52965] = i[52965];
  assign o[52964] = i[52964];
  assign o[52963] = i[52963];
  assign o[52962] = i[52962];
  assign o[52961] = i[52961];
  assign o[52960] = i[52960];
  assign o[52959] = i[52959];
  assign o[52958] = i[52958];
  assign o[52957] = i[52957];
  assign o[52956] = i[52956];
  assign o[52955] = i[52955];
  assign o[52954] = i[52954];
  assign o[52953] = i[52953];
  assign o[52952] = i[52952];
  assign o[52951] = i[52951];
  assign o[52950] = i[52950];
  assign o[52949] = i[52949];
  assign o[52948] = i[52948];
  assign o[52947] = i[52947];
  assign o[52946] = i[52946];
  assign o[52945] = i[52945];
  assign o[52944] = i[52944];
  assign o[52943] = i[52943];
  assign o[52942] = i[52942];
  assign o[52941] = i[52941];
  assign o[52940] = i[52940];
  assign o[52939] = i[52939];
  assign o[52938] = i[52938];
  assign o[52937] = i[52937];
  assign o[52936] = i[52936];
  assign o[52935] = i[52935];
  assign o[52934] = i[52934];
  assign o[52933] = i[52933];
  assign o[52932] = i[52932];
  assign o[52931] = i[52931];
  assign o[52930] = i[52930];
  assign o[52929] = i[52929];
  assign o[52928] = i[52928];
  assign o[52927] = i[52927];
  assign o[52926] = i[52926];
  assign o[52925] = i[52925];
  assign o[52924] = i[52924];
  assign o[52923] = i[52923];
  assign o[52922] = i[52922];
  assign o[52921] = i[52921];
  assign o[52920] = i[52920];
  assign o[52919] = i[52919];
  assign o[52918] = i[52918];
  assign o[52917] = i[52917];
  assign o[52916] = i[52916];
  assign o[52915] = i[52915];
  assign o[52914] = i[52914];
  assign o[52913] = i[52913];
  assign o[52912] = i[52912];
  assign o[52911] = i[52911];
  assign o[52910] = i[52910];
  assign o[52909] = i[52909];
  assign o[52908] = i[52908];
  assign o[52907] = i[52907];
  assign o[52906] = i[52906];
  assign o[52905] = i[52905];
  assign o[52904] = i[52904];
  assign o[52903] = i[52903];
  assign o[52902] = i[52902];
  assign o[52901] = i[52901];
  assign o[52900] = i[52900];
  assign o[52899] = i[52899];
  assign o[52898] = i[52898];
  assign o[52897] = i[52897];
  assign o[52896] = i[52896];
  assign o[52895] = i[52895];
  assign o[52894] = i[52894];
  assign o[52893] = i[52893];
  assign o[52892] = i[52892];
  assign o[52891] = i[52891];
  assign o[52890] = i[52890];
  assign o[52889] = i[52889];
  assign o[52888] = i[52888];
  assign o[52887] = i[52887];
  assign o[52886] = i[52886];
  assign o[52885] = i[52885];
  assign o[52884] = i[52884];
  assign o[52883] = i[52883];
  assign o[52882] = i[52882];
  assign o[52881] = i[52881];
  assign o[52880] = i[52880];
  assign o[52879] = i[52879];
  assign o[52878] = i[52878];
  assign o[52877] = i[52877];
  assign o[52876] = i[52876];
  assign o[52875] = i[52875];
  assign o[52874] = i[52874];
  assign o[52873] = i[52873];
  assign o[52872] = i[52872];
  assign o[52871] = i[52871];
  assign o[52870] = i[52870];
  assign o[52869] = i[52869];
  assign o[52868] = i[52868];
  assign o[52867] = i[52867];
  assign o[52866] = i[52866];
  assign o[52865] = i[52865];
  assign o[52864] = i[52864];
  assign o[52863] = i[52863];
  assign o[52862] = i[52862];
  assign o[52861] = i[52861];
  assign o[52860] = i[52860];
  assign o[52859] = i[52859];
  assign o[52858] = i[52858];
  assign o[52857] = i[52857];
  assign o[52856] = i[52856];
  assign o[52855] = i[52855];
  assign o[52854] = i[52854];
  assign o[52853] = i[52853];
  assign o[52852] = i[52852];
  assign o[52851] = i[52851];
  assign o[52850] = i[52850];
  assign o[52849] = i[52849];
  assign o[52848] = i[52848];
  assign o[52847] = i[52847];
  assign o[52846] = i[52846];
  assign o[52845] = i[52845];
  assign o[52844] = i[52844];
  assign o[52843] = i[52843];
  assign o[52842] = i[52842];
  assign o[52841] = i[52841];
  assign o[52840] = i[52840];
  assign o[52839] = i[52839];
  assign o[52838] = i[52838];
  assign o[52837] = i[52837];
  assign o[52836] = i[52836];
  assign o[52835] = i[52835];
  assign o[52834] = i[52834];
  assign o[52833] = i[52833];
  assign o[52832] = i[52832];
  assign o[52831] = i[52831];
  assign o[52830] = i[52830];
  assign o[52829] = i[52829];
  assign o[52828] = i[52828];
  assign o[52827] = i[52827];
  assign o[52826] = i[52826];
  assign o[52825] = i[52825];
  assign o[52824] = i[52824];
  assign o[52823] = i[52823];
  assign o[52822] = i[52822];
  assign o[52821] = i[52821];
  assign o[52820] = i[52820];
  assign o[52819] = i[52819];
  assign o[52818] = i[52818];
  assign o[52817] = i[52817];
  assign o[52816] = i[52816];
  assign o[52815] = i[52815];
  assign o[52814] = i[52814];
  assign o[52813] = i[52813];
  assign o[52812] = i[52812];
  assign o[52811] = i[52811];
  assign o[52810] = i[52810];
  assign o[52809] = i[52809];
  assign o[52808] = i[52808];
  assign o[52807] = i[52807];
  assign o[52806] = i[52806];
  assign o[52805] = i[52805];
  assign o[52804] = i[52804];
  assign o[52803] = i[52803];
  assign o[52802] = i[52802];
  assign o[52801] = i[52801];
  assign o[52800] = i[52800];
  assign o[52799] = i[52799];
  assign o[52798] = i[52798];
  assign o[52797] = i[52797];
  assign o[52796] = i[52796];
  assign o[52795] = i[52795];
  assign o[52794] = i[52794];
  assign o[52793] = i[52793];
  assign o[52792] = i[52792];
  assign o[52791] = i[52791];
  assign o[52790] = i[52790];
  assign o[52789] = i[52789];
  assign o[52788] = i[52788];
  assign o[52787] = i[52787];
  assign o[52786] = i[52786];
  assign o[52785] = i[52785];
  assign o[52784] = i[52784];
  assign o[52783] = i[52783];
  assign o[52782] = i[52782];
  assign o[52781] = i[52781];
  assign o[52780] = i[52780];
  assign o[52779] = i[52779];
  assign o[52778] = i[52778];
  assign o[52777] = i[52777];
  assign o[52776] = i[52776];
  assign o[52775] = i[52775];
  assign o[52774] = i[52774];
  assign o[52773] = i[52773];
  assign o[52772] = i[52772];
  assign o[52771] = i[52771];
  assign o[52770] = i[52770];
  assign o[52769] = i[52769];
  assign o[52768] = i[52768];
  assign o[52767] = i[52767];
  assign o[52766] = i[52766];
  assign o[52765] = i[52765];
  assign o[52764] = i[52764];
  assign o[52763] = i[52763];
  assign o[52762] = i[52762];
  assign o[52761] = i[52761];
  assign o[52760] = i[52760];
  assign o[52759] = i[52759];
  assign o[52758] = i[52758];
  assign o[52757] = i[52757];
  assign o[52756] = i[52756];
  assign o[52755] = i[52755];
  assign o[52754] = i[52754];
  assign o[52753] = i[52753];
  assign o[52752] = i[52752];
  assign o[52751] = i[52751];
  assign o[52750] = i[52750];
  assign o[52749] = i[52749];
  assign o[52748] = i[52748];
  assign o[52747] = i[52747];
  assign o[52746] = i[52746];
  assign o[52745] = i[52745];
  assign o[52744] = i[52744];
  assign o[52743] = i[52743];
  assign o[52742] = i[52742];
  assign o[52741] = i[52741];
  assign o[52740] = i[52740];
  assign o[52739] = i[52739];
  assign o[52738] = i[52738];
  assign o[52737] = i[52737];
  assign o[52736] = i[52736];
  assign o[52735] = i[52735];
  assign o[52734] = i[52734];
  assign o[52733] = i[52733];
  assign o[52732] = i[52732];
  assign o[52731] = i[52731];
  assign o[52730] = i[52730];
  assign o[52729] = i[52729];
  assign o[52728] = i[52728];
  assign o[52727] = i[52727];
  assign o[52726] = i[52726];
  assign o[52725] = i[52725];
  assign o[52724] = i[52724];
  assign o[52723] = i[52723];
  assign o[52722] = i[52722];
  assign o[52721] = i[52721];
  assign o[52720] = i[52720];
  assign o[52719] = i[52719];
  assign o[52718] = i[52718];
  assign o[52717] = i[52717];
  assign o[52716] = i[52716];
  assign o[52715] = i[52715];
  assign o[52714] = i[52714];
  assign o[52713] = i[52713];
  assign o[52712] = i[52712];
  assign o[52711] = i[52711];
  assign o[52710] = i[52710];
  assign o[52709] = i[52709];
  assign o[52708] = i[52708];
  assign o[52707] = i[52707];
  assign o[52706] = i[52706];
  assign o[52705] = i[52705];
  assign o[52704] = i[52704];
  assign o[52703] = i[52703];
  assign o[52702] = i[52702];
  assign o[52701] = i[52701];
  assign o[52700] = i[52700];
  assign o[52699] = i[52699];
  assign o[52698] = i[52698];
  assign o[52697] = i[52697];
  assign o[52696] = i[52696];
  assign o[52695] = i[52695];
  assign o[52694] = i[52694];
  assign o[52693] = i[52693];
  assign o[52692] = i[52692];
  assign o[52691] = i[52691];
  assign o[52690] = i[52690];
  assign o[52689] = i[52689];
  assign o[52688] = i[52688];
  assign o[52687] = i[52687];
  assign o[52686] = i[52686];
  assign o[52685] = i[52685];
  assign o[52684] = i[52684];
  assign o[52683] = i[52683];
  assign o[52682] = i[52682];
  assign o[52681] = i[52681];
  assign o[52680] = i[52680];
  assign o[52679] = i[52679];
  assign o[52678] = i[52678];
  assign o[52677] = i[52677];
  assign o[52676] = i[52676];
  assign o[52675] = i[52675];
  assign o[52674] = i[52674];
  assign o[52673] = i[52673];
  assign o[52672] = i[52672];
  assign o[52671] = i[52671];
  assign o[52670] = i[52670];
  assign o[52669] = i[52669];
  assign o[52668] = i[52668];
  assign o[52667] = i[52667];
  assign o[52666] = i[52666];
  assign o[52665] = i[52665];
  assign o[52664] = i[52664];
  assign o[52663] = i[52663];
  assign o[52662] = i[52662];
  assign o[52661] = i[52661];
  assign o[52660] = i[52660];
  assign o[52659] = i[52659];
  assign o[52658] = i[52658];
  assign o[52657] = i[52657];
  assign o[52656] = i[52656];
  assign o[52655] = i[52655];
  assign o[52654] = i[52654];
  assign o[52653] = i[52653];
  assign o[52652] = i[52652];
  assign o[52651] = i[52651];
  assign o[52650] = i[52650];
  assign o[52649] = i[52649];
  assign o[52648] = i[52648];
  assign o[52647] = i[52647];
  assign o[52646] = i[52646];
  assign o[52645] = i[52645];
  assign o[52644] = i[52644];
  assign o[52643] = i[52643];
  assign o[52642] = i[52642];
  assign o[52641] = i[52641];
  assign o[52640] = i[52640];
  assign o[52639] = i[52639];
  assign o[52638] = i[52638];
  assign o[52637] = i[52637];
  assign o[52636] = i[52636];
  assign o[52635] = i[52635];
  assign o[52634] = i[52634];
  assign o[52633] = i[52633];
  assign o[52632] = i[52632];
  assign o[52631] = i[52631];
  assign o[52630] = i[52630];
  assign o[52629] = i[52629];
  assign o[52628] = i[52628];
  assign o[52627] = i[52627];
  assign o[52626] = i[52626];
  assign o[52625] = i[52625];
  assign o[52624] = i[52624];
  assign o[52623] = i[52623];
  assign o[52622] = i[52622];
  assign o[52621] = i[52621];
  assign o[52620] = i[52620];
  assign o[52619] = i[52619];
  assign o[52618] = i[52618];
  assign o[52617] = i[52617];
  assign o[52616] = i[52616];
  assign o[52615] = i[52615];
  assign o[52614] = i[52614];
  assign o[52613] = i[52613];
  assign o[52612] = i[52612];
  assign o[52611] = i[52611];
  assign o[52610] = i[52610];
  assign o[52609] = i[52609];
  assign o[52608] = i[52608];
  assign o[52607] = i[52607];
  assign o[52606] = i[52606];
  assign o[52605] = i[52605];
  assign o[52604] = i[52604];
  assign o[52603] = i[52603];
  assign o[52602] = i[52602];
  assign o[52601] = i[52601];
  assign o[52600] = i[52600];
  assign o[52599] = i[52599];
  assign o[52598] = i[52598];
  assign o[52597] = i[52597];
  assign o[52596] = i[52596];
  assign o[52595] = i[52595];
  assign o[52594] = i[52594];
  assign o[52593] = i[52593];
  assign o[52592] = i[52592];
  assign o[52591] = i[52591];
  assign o[52590] = i[52590];
  assign o[52589] = i[52589];
  assign o[52588] = i[52588];
  assign o[52587] = i[52587];
  assign o[52586] = i[52586];
  assign o[52585] = i[52585];
  assign o[52584] = i[52584];
  assign o[52583] = i[52583];
  assign o[52582] = i[52582];
  assign o[52581] = i[52581];
  assign o[52580] = i[52580];
  assign o[52579] = i[52579];
  assign o[52578] = i[52578];
  assign o[52577] = i[52577];
  assign o[52576] = i[52576];
  assign o[52575] = i[52575];
  assign o[52574] = i[52574];
  assign o[52573] = i[52573];
  assign o[52572] = i[52572];
  assign o[52571] = i[52571];
  assign o[52570] = i[52570];
  assign o[52569] = i[52569];
  assign o[52568] = i[52568];
  assign o[52567] = i[52567];
  assign o[52566] = i[52566];
  assign o[52565] = i[52565];
  assign o[52564] = i[52564];
  assign o[52563] = i[52563];
  assign o[52562] = i[52562];
  assign o[52561] = i[52561];
  assign o[52560] = i[52560];
  assign o[52559] = i[52559];
  assign o[52558] = i[52558];
  assign o[52557] = i[52557];
  assign o[52556] = i[52556];
  assign o[52555] = i[52555];
  assign o[52554] = i[52554];
  assign o[52553] = i[52553];
  assign o[52552] = i[52552];
  assign o[52551] = i[52551];
  assign o[52550] = i[52550];
  assign o[52549] = i[52549];
  assign o[52548] = i[52548];
  assign o[52547] = i[52547];
  assign o[52546] = i[52546];
  assign o[52545] = i[52545];
  assign o[52544] = i[52544];
  assign o[52543] = i[52543];
  assign o[52542] = i[52542];
  assign o[52541] = i[52541];
  assign o[52540] = i[52540];
  assign o[52539] = i[52539];
  assign o[52538] = i[52538];
  assign o[52537] = i[52537];
  assign o[52536] = i[52536];
  assign o[52535] = i[52535];
  assign o[52534] = i[52534];
  assign o[52533] = i[52533];
  assign o[52532] = i[52532];
  assign o[52531] = i[52531];
  assign o[52530] = i[52530];
  assign o[52529] = i[52529];
  assign o[52528] = i[52528];
  assign o[52527] = i[52527];
  assign o[52526] = i[52526];
  assign o[52525] = i[52525];
  assign o[52524] = i[52524];
  assign o[52523] = i[52523];
  assign o[52522] = i[52522];
  assign o[52521] = i[52521];
  assign o[52520] = i[52520];
  assign o[52519] = i[52519];
  assign o[52518] = i[52518];
  assign o[52517] = i[52517];
  assign o[52516] = i[52516];
  assign o[52515] = i[52515];
  assign o[52514] = i[52514];
  assign o[52513] = i[52513];
  assign o[52512] = i[52512];
  assign o[52511] = i[52511];
  assign o[52510] = i[52510];
  assign o[52509] = i[52509];
  assign o[52508] = i[52508];
  assign o[52507] = i[52507];
  assign o[52506] = i[52506];
  assign o[52505] = i[52505];
  assign o[52504] = i[52504];
  assign o[52503] = i[52503];
  assign o[52502] = i[52502];
  assign o[52501] = i[52501];
  assign o[52500] = i[52500];
  assign o[52499] = i[52499];
  assign o[52498] = i[52498];
  assign o[52497] = i[52497];
  assign o[52496] = i[52496];
  assign o[52495] = i[52495];
  assign o[52494] = i[52494];
  assign o[52493] = i[52493];
  assign o[52492] = i[52492];
  assign o[52491] = i[52491];
  assign o[52490] = i[52490];
  assign o[52489] = i[52489];
  assign o[52488] = i[52488];
  assign o[52487] = i[52487];
  assign o[52486] = i[52486];
  assign o[52485] = i[52485];
  assign o[52484] = i[52484];
  assign o[52483] = i[52483];
  assign o[52482] = i[52482];
  assign o[52481] = i[52481];
  assign o[52480] = i[52480];
  assign o[52479] = i[52479];
  assign o[52478] = i[52478];
  assign o[52477] = i[52477];
  assign o[52476] = i[52476];
  assign o[52475] = i[52475];
  assign o[52474] = i[52474];
  assign o[52473] = i[52473];
  assign o[52472] = i[52472];
  assign o[52471] = i[52471];
  assign o[52470] = i[52470];
  assign o[52469] = i[52469];
  assign o[52468] = i[52468];
  assign o[52467] = i[52467];
  assign o[52466] = i[52466];
  assign o[52465] = i[52465];
  assign o[52464] = i[52464];
  assign o[52463] = i[52463];
  assign o[52462] = i[52462];
  assign o[52461] = i[52461];
  assign o[52460] = i[52460];
  assign o[52459] = i[52459];
  assign o[52458] = i[52458];
  assign o[52457] = i[52457];
  assign o[52456] = i[52456];
  assign o[52455] = i[52455];
  assign o[52454] = i[52454];
  assign o[52453] = i[52453];
  assign o[52452] = i[52452];
  assign o[52451] = i[52451];
  assign o[52450] = i[52450];
  assign o[52449] = i[52449];
  assign o[52448] = i[52448];
  assign o[52447] = i[52447];
  assign o[52446] = i[52446];
  assign o[52445] = i[52445];
  assign o[52444] = i[52444];
  assign o[52443] = i[52443];
  assign o[52442] = i[52442];
  assign o[52441] = i[52441];
  assign o[52440] = i[52440];
  assign o[52439] = i[52439];
  assign o[52438] = i[52438];
  assign o[52437] = i[52437];
  assign o[52436] = i[52436];
  assign o[52435] = i[52435];
  assign o[52434] = i[52434];
  assign o[52433] = i[52433];
  assign o[52432] = i[52432];
  assign o[52431] = i[52431];
  assign o[52430] = i[52430];
  assign o[52429] = i[52429];
  assign o[52428] = i[52428];
  assign o[52427] = i[52427];
  assign o[52426] = i[52426];
  assign o[52425] = i[52425];
  assign o[52424] = i[52424];
  assign o[52423] = i[52423];
  assign o[52422] = i[52422];
  assign o[52421] = i[52421];
  assign o[52420] = i[52420];
  assign o[52419] = i[52419];
  assign o[52418] = i[52418];
  assign o[52417] = i[52417];
  assign o[52416] = i[52416];
  assign o[52415] = i[52415];
  assign o[52414] = i[52414];
  assign o[52413] = i[52413];
  assign o[52412] = i[52412];
  assign o[52411] = i[52411];
  assign o[52410] = i[52410];
  assign o[52409] = i[52409];
  assign o[52408] = i[52408];
  assign o[52407] = i[52407];
  assign o[52406] = i[52406];
  assign o[52405] = i[52405];
  assign o[52404] = i[52404];
  assign o[52403] = i[52403];
  assign o[52402] = i[52402];
  assign o[52401] = i[52401];
  assign o[52400] = i[52400];
  assign o[52399] = i[52399];
  assign o[52398] = i[52398];
  assign o[52397] = i[52397];
  assign o[52396] = i[52396];
  assign o[52395] = i[52395];
  assign o[52394] = i[52394];
  assign o[52393] = i[52393];
  assign o[52392] = i[52392];
  assign o[52391] = i[52391];
  assign o[52390] = i[52390];
  assign o[52389] = i[52389];
  assign o[52388] = i[52388];
  assign o[52387] = i[52387];
  assign o[52386] = i[52386];
  assign o[52385] = i[52385];
  assign o[52384] = i[52384];
  assign o[52383] = i[52383];
  assign o[52382] = i[52382];
  assign o[52381] = i[52381];
  assign o[52380] = i[52380];
  assign o[52379] = i[52379];
  assign o[52378] = i[52378];
  assign o[52377] = i[52377];
  assign o[52376] = i[52376];
  assign o[52375] = i[52375];
  assign o[52374] = i[52374];
  assign o[52373] = i[52373];
  assign o[52372] = i[52372];
  assign o[52371] = i[52371];
  assign o[52370] = i[52370];
  assign o[52369] = i[52369];
  assign o[52368] = i[52368];
  assign o[52367] = i[52367];
  assign o[52366] = i[52366];
  assign o[52365] = i[52365];
  assign o[52364] = i[52364];
  assign o[52363] = i[52363];
  assign o[52362] = i[52362];
  assign o[52361] = i[52361];
  assign o[52360] = i[52360];
  assign o[52359] = i[52359];
  assign o[52358] = i[52358];
  assign o[52357] = i[52357];
  assign o[52356] = i[52356];
  assign o[52355] = i[52355];
  assign o[52354] = i[52354];
  assign o[52353] = i[52353];
  assign o[52352] = i[52352];
  assign o[52351] = i[52351];
  assign o[52350] = i[52350];
  assign o[52349] = i[52349];
  assign o[52348] = i[52348];
  assign o[52347] = i[52347];
  assign o[52346] = i[52346];
  assign o[52345] = i[52345];
  assign o[52344] = i[52344];
  assign o[52343] = i[52343];
  assign o[52342] = i[52342];
  assign o[52341] = i[52341];
  assign o[52340] = i[52340];
  assign o[52339] = i[52339];
  assign o[52338] = i[52338];
  assign o[52337] = i[52337];
  assign o[52336] = i[52336];
  assign o[52335] = i[52335];
  assign o[52334] = i[52334];
  assign o[52333] = i[52333];
  assign o[52332] = i[52332];
  assign o[52331] = i[52331];
  assign o[52330] = i[52330];
  assign o[52329] = i[52329];
  assign o[52328] = i[52328];
  assign o[52327] = i[52327];
  assign o[52326] = i[52326];
  assign o[52325] = i[52325];
  assign o[52324] = i[52324];
  assign o[52323] = i[52323];
  assign o[52322] = i[52322];
  assign o[52321] = i[52321];
  assign o[52320] = i[52320];
  assign o[52319] = i[52319];
  assign o[52318] = i[52318];
  assign o[52317] = i[52317];
  assign o[52316] = i[52316];
  assign o[52315] = i[52315];
  assign o[52314] = i[52314];
  assign o[52313] = i[52313];
  assign o[52312] = i[52312];
  assign o[52311] = i[52311];
  assign o[52310] = i[52310];
  assign o[52309] = i[52309];
  assign o[52308] = i[52308];
  assign o[52307] = i[52307];
  assign o[52306] = i[52306];
  assign o[52305] = i[52305];
  assign o[52304] = i[52304];
  assign o[52303] = i[52303];
  assign o[52302] = i[52302];
  assign o[52301] = i[52301];
  assign o[52300] = i[52300];
  assign o[52299] = i[52299];
  assign o[52298] = i[52298];
  assign o[52297] = i[52297];
  assign o[52296] = i[52296];
  assign o[52295] = i[52295];
  assign o[52294] = i[52294];
  assign o[52293] = i[52293];
  assign o[52292] = i[52292];
  assign o[52291] = i[52291];
  assign o[52290] = i[52290];
  assign o[52289] = i[52289];
  assign o[52288] = i[52288];
  assign o[52287] = i[52287];
  assign o[52286] = i[52286];
  assign o[52285] = i[52285];
  assign o[52284] = i[52284];
  assign o[52283] = i[52283];
  assign o[52282] = i[52282];
  assign o[52281] = i[52281];
  assign o[52280] = i[52280];
  assign o[52279] = i[52279];
  assign o[52278] = i[52278];
  assign o[52277] = i[52277];
  assign o[52276] = i[52276];
  assign o[52275] = i[52275];
  assign o[52274] = i[52274];
  assign o[52273] = i[52273];
  assign o[52272] = i[52272];
  assign o[52271] = i[52271];
  assign o[52270] = i[52270];
  assign o[52269] = i[52269];
  assign o[52268] = i[52268];
  assign o[52267] = i[52267];
  assign o[52266] = i[52266];
  assign o[52265] = i[52265];
  assign o[52264] = i[52264];
  assign o[52263] = i[52263];
  assign o[52262] = i[52262];
  assign o[52261] = i[52261];
  assign o[52260] = i[52260];
  assign o[52259] = i[52259];
  assign o[52258] = i[52258];
  assign o[52257] = i[52257];
  assign o[52256] = i[52256];
  assign o[52255] = i[52255];
  assign o[52254] = i[52254];
  assign o[52253] = i[52253];
  assign o[52252] = i[52252];
  assign o[52251] = i[52251];
  assign o[52250] = i[52250];
  assign o[52249] = i[52249];
  assign o[52248] = i[52248];
  assign o[52247] = i[52247];
  assign o[52246] = i[52246];
  assign o[52245] = i[52245];
  assign o[52244] = i[52244];
  assign o[52243] = i[52243];
  assign o[52242] = i[52242];
  assign o[52241] = i[52241];
  assign o[52240] = i[52240];
  assign o[52239] = i[52239];
  assign o[52238] = i[52238];
  assign o[52237] = i[52237];
  assign o[52236] = i[52236];
  assign o[52235] = i[52235];
  assign o[52234] = i[52234];
  assign o[52233] = i[52233];
  assign o[52232] = i[52232];
  assign o[52231] = i[52231];
  assign o[52230] = i[52230];
  assign o[52229] = i[52229];
  assign o[52228] = i[52228];
  assign o[52227] = i[52227];
  assign o[52226] = i[52226];
  assign o[52225] = i[52225];
  assign o[52224] = i[52224];
  assign o[52223] = i[52223];
  assign o[52222] = i[52222];
  assign o[52221] = i[52221];
  assign o[52220] = i[52220];
  assign o[52219] = i[52219];
  assign o[52218] = i[52218];
  assign o[52217] = i[52217];
  assign o[52216] = i[52216];
  assign o[52215] = i[52215];
  assign o[52214] = i[52214];
  assign o[52213] = i[52213];
  assign o[52212] = i[52212];
  assign o[52211] = i[52211];
  assign o[52210] = i[52210];
  assign o[52209] = i[52209];
  assign o[52208] = i[52208];
  assign o[52207] = i[52207];
  assign o[52206] = i[52206];
  assign o[52205] = i[52205];
  assign o[52204] = i[52204];
  assign o[52203] = i[52203];
  assign o[52202] = i[52202];
  assign o[52201] = i[52201];
  assign o[52200] = i[52200];
  assign o[52199] = i[52199];
  assign o[52198] = i[52198];
  assign o[52197] = i[52197];
  assign o[52196] = i[52196];
  assign o[52195] = i[52195];
  assign o[52194] = i[52194];
  assign o[52193] = i[52193];
  assign o[52192] = i[52192];
  assign o[52191] = i[52191];
  assign o[52190] = i[52190];
  assign o[52189] = i[52189];
  assign o[52188] = i[52188];
  assign o[52187] = i[52187];
  assign o[52186] = i[52186];
  assign o[52185] = i[52185];
  assign o[52184] = i[52184];
  assign o[52183] = i[52183];
  assign o[52182] = i[52182];
  assign o[52181] = i[52181];
  assign o[52180] = i[52180];
  assign o[52179] = i[52179];
  assign o[52178] = i[52178];
  assign o[52177] = i[52177];
  assign o[52176] = i[52176];
  assign o[52175] = i[52175];
  assign o[52174] = i[52174];
  assign o[52173] = i[52173];
  assign o[52172] = i[52172];
  assign o[52171] = i[52171];
  assign o[52170] = i[52170];
  assign o[52169] = i[52169];
  assign o[52168] = i[52168];
  assign o[52167] = i[52167];
  assign o[52166] = i[52166];
  assign o[52165] = i[52165];
  assign o[52164] = i[52164];
  assign o[52163] = i[52163];
  assign o[52162] = i[52162];
  assign o[52161] = i[52161];
  assign o[52160] = i[52160];
  assign o[52159] = i[52159];
  assign o[52158] = i[52158];
  assign o[52157] = i[52157];
  assign o[52156] = i[52156];
  assign o[52155] = i[52155];
  assign o[52154] = i[52154];
  assign o[52153] = i[52153];
  assign o[52152] = i[52152];
  assign o[52151] = i[52151];
  assign o[52150] = i[52150];
  assign o[52149] = i[52149];
  assign o[52148] = i[52148];
  assign o[52147] = i[52147];
  assign o[52146] = i[52146];
  assign o[52145] = i[52145];
  assign o[52144] = i[52144];
  assign o[52143] = i[52143];
  assign o[52142] = i[52142];
  assign o[52141] = i[52141];
  assign o[52140] = i[52140];
  assign o[52139] = i[52139];
  assign o[52138] = i[52138];
  assign o[52137] = i[52137];
  assign o[52136] = i[52136];
  assign o[52135] = i[52135];
  assign o[52134] = i[52134];
  assign o[52133] = i[52133];
  assign o[52132] = i[52132];
  assign o[52131] = i[52131];
  assign o[52130] = i[52130];
  assign o[52129] = i[52129];
  assign o[52128] = i[52128];
  assign o[52127] = i[52127];
  assign o[52126] = i[52126];
  assign o[52125] = i[52125];
  assign o[52124] = i[52124];
  assign o[52123] = i[52123];
  assign o[52122] = i[52122];
  assign o[52121] = i[52121];
  assign o[52120] = i[52120];
  assign o[52119] = i[52119];
  assign o[52118] = i[52118];
  assign o[52117] = i[52117];
  assign o[52116] = i[52116];
  assign o[52115] = i[52115];
  assign o[52114] = i[52114];
  assign o[52113] = i[52113];
  assign o[52112] = i[52112];
  assign o[52111] = i[52111];
  assign o[52110] = i[52110];
  assign o[52109] = i[52109];
  assign o[52108] = i[52108];
  assign o[52107] = i[52107];
  assign o[52106] = i[52106];
  assign o[52105] = i[52105];
  assign o[52104] = i[52104];
  assign o[52103] = i[52103];
  assign o[52102] = i[52102];
  assign o[52101] = i[52101];
  assign o[52100] = i[52100];
  assign o[52099] = i[52099];
  assign o[52098] = i[52098];
  assign o[52097] = i[52097];
  assign o[52096] = i[52096];
  assign o[52095] = i[52095];
  assign o[52094] = i[52094];
  assign o[52093] = i[52093];
  assign o[52092] = i[52092];
  assign o[52091] = i[52091];
  assign o[52090] = i[52090];
  assign o[52089] = i[52089];
  assign o[52088] = i[52088];
  assign o[52087] = i[52087];
  assign o[52086] = i[52086];
  assign o[52085] = i[52085];
  assign o[52084] = i[52084];
  assign o[52083] = i[52083];
  assign o[52082] = i[52082];
  assign o[52081] = i[52081];
  assign o[52080] = i[52080];
  assign o[52079] = i[52079];
  assign o[52078] = i[52078];
  assign o[52077] = i[52077];
  assign o[52076] = i[52076];
  assign o[52075] = i[52075];
  assign o[52074] = i[52074];
  assign o[52073] = i[52073];
  assign o[52072] = i[52072];
  assign o[52071] = i[52071];
  assign o[52070] = i[52070];
  assign o[52069] = i[52069];
  assign o[52068] = i[52068];
  assign o[52067] = i[52067];
  assign o[52066] = i[52066];
  assign o[52065] = i[52065];
  assign o[52064] = i[52064];
  assign o[52063] = i[52063];
  assign o[52062] = i[52062];
  assign o[52061] = i[52061];
  assign o[52060] = i[52060];
  assign o[52059] = i[52059];
  assign o[52058] = i[52058];
  assign o[52057] = i[52057];
  assign o[52056] = i[52056];
  assign o[52055] = i[52055];
  assign o[52054] = i[52054];
  assign o[52053] = i[52053];
  assign o[52052] = i[52052];
  assign o[52051] = i[52051];
  assign o[52050] = i[52050];
  assign o[52049] = i[52049];
  assign o[52048] = i[52048];
  assign o[52047] = i[52047];
  assign o[52046] = i[52046];
  assign o[52045] = i[52045];
  assign o[52044] = i[52044];
  assign o[52043] = i[52043];
  assign o[52042] = i[52042];
  assign o[52041] = i[52041];
  assign o[52040] = i[52040];
  assign o[52039] = i[52039];
  assign o[52038] = i[52038];
  assign o[52037] = i[52037];
  assign o[52036] = i[52036];
  assign o[52035] = i[52035];
  assign o[52034] = i[52034];
  assign o[52033] = i[52033];
  assign o[52032] = i[52032];
  assign o[52031] = i[52031];
  assign o[52030] = i[52030];
  assign o[52029] = i[52029];
  assign o[52028] = i[52028];
  assign o[52027] = i[52027];
  assign o[52026] = i[52026];
  assign o[52025] = i[52025];
  assign o[52024] = i[52024];
  assign o[52023] = i[52023];
  assign o[52022] = i[52022];
  assign o[52021] = i[52021];
  assign o[52020] = i[52020];
  assign o[52019] = i[52019];
  assign o[52018] = i[52018];
  assign o[52017] = i[52017];
  assign o[52016] = i[52016];
  assign o[52015] = i[52015];
  assign o[52014] = i[52014];
  assign o[52013] = i[52013];
  assign o[52012] = i[52012];
  assign o[52011] = i[52011];
  assign o[52010] = i[52010];
  assign o[52009] = i[52009];
  assign o[52008] = i[52008];
  assign o[52007] = i[52007];
  assign o[52006] = i[52006];
  assign o[52005] = i[52005];
  assign o[52004] = i[52004];
  assign o[52003] = i[52003];
  assign o[52002] = i[52002];
  assign o[52001] = i[52001];
  assign o[52000] = i[52000];
  assign o[51999] = i[51999];
  assign o[51998] = i[51998];
  assign o[51997] = i[51997];
  assign o[51996] = i[51996];
  assign o[51995] = i[51995];
  assign o[51994] = i[51994];
  assign o[51993] = i[51993];
  assign o[51992] = i[51992];
  assign o[51991] = i[51991];
  assign o[51990] = i[51990];
  assign o[51989] = i[51989];
  assign o[51988] = i[51988];
  assign o[51987] = i[51987];
  assign o[51986] = i[51986];
  assign o[51985] = i[51985];
  assign o[51984] = i[51984];
  assign o[51983] = i[51983];
  assign o[51982] = i[51982];
  assign o[51981] = i[51981];
  assign o[51980] = i[51980];
  assign o[51979] = i[51979];
  assign o[51978] = i[51978];
  assign o[51977] = i[51977];
  assign o[51976] = i[51976];
  assign o[51975] = i[51975];
  assign o[51974] = i[51974];
  assign o[51973] = i[51973];
  assign o[51972] = i[51972];
  assign o[51971] = i[51971];
  assign o[51970] = i[51970];
  assign o[51969] = i[51969];
  assign o[51968] = i[51968];
  assign o[51967] = i[51967];
  assign o[51966] = i[51966];
  assign o[51965] = i[51965];
  assign o[51964] = i[51964];
  assign o[51963] = i[51963];
  assign o[51962] = i[51962];
  assign o[51961] = i[51961];
  assign o[51960] = i[51960];
  assign o[51959] = i[51959];
  assign o[51958] = i[51958];
  assign o[51957] = i[51957];
  assign o[51956] = i[51956];
  assign o[51955] = i[51955];
  assign o[51954] = i[51954];
  assign o[51953] = i[51953];
  assign o[51952] = i[51952];
  assign o[51951] = i[51951];
  assign o[51950] = i[51950];
  assign o[51949] = i[51949];
  assign o[51948] = i[51948];
  assign o[51947] = i[51947];
  assign o[51946] = i[51946];
  assign o[51945] = i[51945];
  assign o[51944] = i[51944];
  assign o[51943] = i[51943];
  assign o[51942] = i[51942];
  assign o[51941] = i[51941];
  assign o[51940] = i[51940];
  assign o[51939] = i[51939];
  assign o[51938] = i[51938];
  assign o[51937] = i[51937];
  assign o[51936] = i[51936];
  assign o[51935] = i[51935];
  assign o[51934] = i[51934];
  assign o[51933] = i[51933];
  assign o[51932] = i[51932];
  assign o[51931] = i[51931];
  assign o[51930] = i[51930];
  assign o[51929] = i[51929];
  assign o[51928] = i[51928];
  assign o[51927] = i[51927];
  assign o[51926] = i[51926];
  assign o[51925] = i[51925];
  assign o[51924] = i[51924];
  assign o[51923] = i[51923];
  assign o[51922] = i[51922];
  assign o[51921] = i[51921];
  assign o[51920] = i[51920];
  assign o[51919] = i[51919];
  assign o[51918] = i[51918];
  assign o[51917] = i[51917];
  assign o[51916] = i[51916];
  assign o[51915] = i[51915];
  assign o[51914] = i[51914];
  assign o[51913] = i[51913];
  assign o[51912] = i[51912];
  assign o[51911] = i[51911];
  assign o[51910] = i[51910];
  assign o[51909] = i[51909];
  assign o[51908] = i[51908];
  assign o[51907] = i[51907];
  assign o[51906] = i[51906];
  assign o[51905] = i[51905];
  assign o[51904] = i[51904];
  assign o[51903] = i[51903];
  assign o[51902] = i[51902];
  assign o[51901] = i[51901];
  assign o[51900] = i[51900];
  assign o[51899] = i[51899];
  assign o[51898] = i[51898];
  assign o[51897] = i[51897];
  assign o[51896] = i[51896];
  assign o[51895] = i[51895];
  assign o[51894] = i[51894];
  assign o[51893] = i[51893];
  assign o[51892] = i[51892];
  assign o[51891] = i[51891];
  assign o[51890] = i[51890];
  assign o[51889] = i[51889];
  assign o[51888] = i[51888];
  assign o[51887] = i[51887];
  assign o[51886] = i[51886];
  assign o[51885] = i[51885];
  assign o[51884] = i[51884];
  assign o[51883] = i[51883];
  assign o[51882] = i[51882];
  assign o[51881] = i[51881];
  assign o[51880] = i[51880];
  assign o[51879] = i[51879];
  assign o[51878] = i[51878];
  assign o[51877] = i[51877];
  assign o[51876] = i[51876];
  assign o[51875] = i[51875];
  assign o[51874] = i[51874];
  assign o[51873] = i[51873];
  assign o[51872] = i[51872];
  assign o[51871] = i[51871];
  assign o[51870] = i[51870];
  assign o[51869] = i[51869];
  assign o[51868] = i[51868];
  assign o[51867] = i[51867];
  assign o[51866] = i[51866];
  assign o[51865] = i[51865];
  assign o[51864] = i[51864];
  assign o[51863] = i[51863];
  assign o[51862] = i[51862];
  assign o[51861] = i[51861];
  assign o[51860] = i[51860];
  assign o[51859] = i[51859];
  assign o[51858] = i[51858];
  assign o[51857] = i[51857];
  assign o[51856] = i[51856];
  assign o[51855] = i[51855];
  assign o[51854] = i[51854];
  assign o[51853] = i[51853];
  assign o[51852] = i[51852];
  assign o[51851] = i[51851];
  assign o[51850] = i[51850];
  assign o[51849] = i[51849];
  assign o[51848] = i[51848];
  assign o[51847] = i[51847];
  assign o[51846] = i[51846];
  assign o[51845] = i[51845];
  assign o[51844] = i[51844];
  assign o[51843] = i[51843];
  assign o[51842] = i[51842];
  assign o[51841] = i[51841];
  assign o[51840] = i[51840];
  assign o[51839] = i[51839];
  assign o[51838] = i[51838];
  assign o[51837] = i[51837];
  assign o[51836] = i[51836];
  assign o[51835] = i[51835];
  assign o[51834] = i[51834];
  assign o[51833] = i[51833];
  assign o[51832] = i[51832];
  assign o[51831] = i[51831];
  assign o[51830] = i[51830];
  assign o[51829] = i[51829];
  assign o[51828] = i[51828];
  assign o[51827] = i[51827];
  assign o[51826] = i[51826];
  assign o[51825] = i[51825];
  assign o[51824] = i[51824];
  assign o[51823] = i[51823];
  assign o[51822] = i[51822];
  assign o[51821] = i[51821];
  assign o[51820] = i[51820];
  assign o[51819] = i[51819];
  assign o[51818] = i[51818];
  assign o[51817] = i[51817];
  assign o[51816] = i[51816];
  assign o[51815] = i[51815];
  assign o[51814] = i[51814];
  assign o[51813] = i[51813];
  assign o[51812] = i[51812];
  assign o[51811] = i[51811];
  assign o[51810] = i[51810];
  assign o[51809] = i[51809];
  assign o[51808] = i[51808];
  assign o[51807] = i[51807];
  assign o[51806] = i[51806];
  assign o[51805] = i[51805];
  assign o[51804] = i[51804];
  assign o[51803] = i[51803];
  assign o[51802] = i[51802];
  assign o[51801] = i[51801];
  assign o[51800] = i[51800];
  assign o[51799] = i[51799];
  assign o[51798] = i[51798];
  assign o[51797] = i[51797];
  assign o[51796] = i[51796];
  assign o[51795] = i[51795];
  assign o[51794] = i[51794];
  assign o[51793] = i[51793];
  assign o[51792] = i[51792];
  assign o[51791] = i[51791];
  assign o[51790] = i[51790];
  assign o[51789] = i[51789];
  assign o[51788] = i[51788];
  assign o[51787] = i[51787];
  assign o[51786] = i[51786];
  assign o[51785] = i[51785];
  assign o[51784] = i[51784];
  assign o[51783] = i[51783];
  assign o[51782] = i[51782];
  assign o[51781] = i[51781];
  assign o[51780] = i[51780];
  assign o[51779] = i[51779];
  assign o[51778] = i[51778];
  assign o[51777] = i[51777];
  assign o[51776] = i[51776];
  assign o[51775] = i[51775];
  assign o[51774] = i[51774];
  assign o[51773] = i[51773];
  assign o[51772] = i[51772];
  assign o[51771] = i[51771];
  assign o[51770] = i[51770];
  assign o[51769] = i[51769];
  assign o[51768] = i[51768];
  assign o[51767] = i[51767];
  assign o[51766] = i[51766];
  assign o[51765] = i[51765];
  assign o[51764] = i[51764];
  assign o[51763] = i[51763];
  assign o[51762] = i[51762];
  assign o[51761] = i[51761];
  assign o[51760] = i[51760];
  assign o[51759] = i[51759];
  assign o[51758] = i[51758];
  assign o[51757] = i[51757];
  assign o[51756] = i[51756];
  assign o[51755] = i[51755];
  assign o[51754] = i[51754];
  assign o[51753] = i[51753];
  assign o[51752] = i[51752];
  assign o[51751] = i[51751];
  assign o[51750] = i[51750];
  assign o[51749] = i[51749];
  assign o[51748] = i[51748];
  assign o[51747] = i[51747];
  assign o[51746] = i[51746];
  assign o[51745] = i[51745];
  assign o[51744] = i[51744];
  assign o[51743] = i[51743];
  assign o[51742] = i[51742];
  assign o[51741] = i[51741];
  assign o[51740] = i[51740];
  assign o[51739] = i[51739];
  assign o[51738] = i[51738];
  assign o[51737] = i[51737];
  assign o[51736] = i[51736];
  assign o[51735] = i[51735];
  assign o[51734] = i[51734];
  assign o[51733] = i[51733];
  assign o[51732] = i[51732];
  assign o[51731] = i[51731];
  assign o[51730] = i[51730];
  assign o[51729] = i[51729];
  assign o[51728] = i[51728];
  assign o[51727] = i[51727];
  assign o[51726] = i[51726];
  assign o[51725] = i[51725];
  assign o[51724] = i[51724];
  assign o[51723] = i[51723];
  assign o[51722] = i[51722];
  assign o[51721] = i[51721];
  assign o[51720] = i[51720];
  assign o[51719] = i[51719];
  assign o[51718] = i[51718];
  assign o[51717] = i[51717];
  assign o[51716] = i[51716];
  assign o[51715] = i[51715];
  assign o[51714] = i[51714];
  assign o[51713] = i[51713];
  assign o[51712] = i[51712];
  assign o[51711] = i[51711];
  assign o[51710] = i[51710];
  assign o[51709] = i[51709];
  assign o[51708] = i[51708];
  assign o[51707] = i[51707];
  assign o[51706] = i[51706];
  assign o[51705] = i[51705];
  assign o[51704] = i[51704];
  assign o[51703] = i[51703];
  assign o[51702] = i[51702];
  assign o[51701] = i[51701];
  assign o[51700] = i[51700];
  assign o[51699] = i[51699];
  assign o[51698] = i[51698];
  assign o[51697] = i[51697];
  assign o[51696] = i[51696];
  assign o[51695] = i[51695];
  assign o[51694] = i[51694];
  assign o[51693] = i[51693];
  assign o[51692] = i[51692];
  assign o[51691] = i[51691];
  assign o[51690] = i[51690];
  assign o[51689] = i[51689];
  assign o[51688] = i[51688];
  assign o[51687] = i[51687];
  assign o[51686] = i[51686];
  assign o[51685] = i[51685];
  assign o[51684] = i[51684];
  assign o[51683] = i[51683];
  assign o[51682] = i[51682];
  assign o[51681] = i[51681];
  assign o[51680] = i[51680];
  assign o[51679] = i[51679];
  assign o[51678] = i[51678];
  assign o[51677] = i[51677];
  assign o[51676] = i[51676];
  assign o[51675] = i[51675];
  assign o[51674] = i[51674];
  assign o[51673] = i[51673];
  assign o[51672] = i[51672];
  assign o[51671] = i[51671];
  assign o[51670] = i[51670];
  assign o[51669] = i[51669];
  assign o[51668] = i[51668];
  assign o[51667] = i[51667];
  assign o[51666] = i[51666];
  assign o[51665] = i[51665];
  assign o[51664] = i[51664];
  assign o[51663] = i[51663];
  assign o[51662] = i[51662];
  assign o[51661] = i[51661];
  assign o[51660] = i[51660];
  assign o[51659] = i[51659];
  assign o[51658] = i[51658];
  assign o[51657] = i[51657];
  assign o[51656] = i[51656];
  assign o[51655] = i[51655];
  assign o[51654] = i[51654];
  assign o[51653] = i[51653];
  assign o[51652] = i[51652];
  assign o[51651] = i[51651];
  assign o[51650] = i[51650];
  assign o[51649] = i[51649];
  assign o[51648] = i[51648];
  assign o[51647] = i[51647];
  assign o[51646] = i[51646];
  assign o[51645] = i[51645];
  assign o[51644] = i[51644];
  assign o[51643] = i[51643];
  assign o[51642] = i[51642];
  assign o[51641] = i[51641];
  assign o[51640] = i[51640];
  assign o[51639] = i[51639];
  assign o[51638] = i[51638];
  assign o[51637] = i[51637];
  assign o[51636] = i[51636];
  assign o[51635] = i[51635];
  assign o[51634] = i[51634];
  assign o[51633] = i[51633];
  assign o[51632] = i[51632];
  assign o[51631] = i[51631];
  assign o[51630] = i[51630];
  assign o[51629] = i[51629];
  assign o[51628] = i[51628];
  assign o[51627] = i[51627];
  assign o[51626] = i[51626];
  assign o[51625] = i[51625];
  assign o[51624] = i[51624];
  assign o[51623] = i[51623];
  assign o[51622] = i[51622];
  assign o[51621] = i[51621];
  assign o[51620] = i[51620];
  assign o[51619] = i[51619];
  assign o[51618] = i[51618];
  assign o[51617] = i[51617];
  assign o[51616] = i[51616];
  assign o[51615] = i[51615];
  assign o[51614] = i[51614];
  assign o[51613] = i[51613];
  assign o[51612] = i[51612];
  assign o[51611] = i[51611];
  assign o[51610] = i[51610];
  assign o[51609] = i[51609];
  assign o[51608] = i[51608];
  assign o[51607] = i[51607];
  assign o[51606] = i[51606];
  assign o[51605] = i[51605];
  assign o[51604] = i[51604];
  assign o[51603] = i[51603];
  assign o[51602] = i[51602];
  assign o[51601] = i[51601];
  assign o[51600] = i[51600];
  assign o[51599] = i[51599];
  assign o[51598] = i[51598];
  assign o[51597] = i[51597];
  assign o[51596] = i[51596];
  assign o[51595] = i[51595];
  assign o[51594] = i[51594];
  assign o[51593] = i[51593];
  assign o[51592] = i[51592];
  assign o[51591] = i[51591];
  assign o[51590] = i[51590];
  assign o[51589] = i[51589];
  assign o[51588] = i[51588];
  assign o[51587] = i[51587];
  assign o[51586] = i[51586];
  assign o[51585] = i[51585];
  assign o[51584] = i[51584];
  assign o[51583] = i[51583];
  assign o[51582] = i[51582];
  assign o[51581] = i[51581];
  assign o[51580] = i[51580];
  assign o[51579] = i[51579];
  assign o[51578] = i[51578];
  assign o[51577] = i[51577];
  assign o[51576] = i[51576];
  assign o[51575] = i[51575];
  assign o[51574] = i[51574];
  assign o[51573] = i[51573];
  assign o[51572] = i[51572];
  assign o[51571] = i[51571];
  assign o[51570] = i[51570];
  assign o[51569] = i[51569];
  assign o[51568] = i[51568];
  assign o[51567] = i[51567];
  assign o[51566] = i[51566];
  assign o[51565] = i[51565];
  assign o[51564] = i[51564];
  assign o[51563] = i[51563];
  assign o[51562] = i[51562];
  assign o[51561] = i[51561];
  assign o[51560] = i[51560];
  assign o[51559] = i[51559];
  assign o[51558] = i[51558];
  assign o[51557] = i[51557];
  assign o[51556] = i[51556];
  assign o[51555] = i[51555];
  assign o[51554] = i[51554];
  assign o[51553] = i[51553];
  assign o[51552] = i[51552];
  assign o[51551] = i[51551];
  assign o[51550] = i[51550];
  assign o[51549] = i[51549];
  assign o[51548] = i[51548];
  assign o[51547] = i[51547];
  assign o[51546] = i[51546];
  assign o[51545] = i[51545];
  assign o[51544] = i[51544];
  assign o[51543] = i[51543];
  assign o[51542] = i[51542];
  assign o[51541] = i[51541];
  assign o[51540] = i[51540];
  assign o[51539] = i[51539];
  assign o[51538] = i[51538];
  assign o[51537] = i[51537];
  assign o[51536] = i[51536];
  assign o[51535] = i[51535];
  assign o[51534] = i[51534];
  assign o[51533] = i[51533];
  assign o[51532] = i[51532];
  assign o[51531] = i[51531];
  assign o[51530] = i[51530];
  assign o[51529] = i[51529];
  assign o[51528] = i[51528];
  assign o[51527] = i[51527];
  assign o[51526] = i[51526];
  assign o[51525] = i[51525];
  assign o[51524] = i[51524];
  assign o[51523] = i[51523];
  assign o[51522] = i[51522];
  assign o[51521] = i[51521];
  assign o[51520] = i[51520];
  assign o[51519] = i[51519];
  assign o[51518] = i[51518];
  assign o[51517] = i[51517];
  assign o[51516] = i[51516];
  assign o[51515] = i[51515];
  assign o[51514] = i[51514];
  assign o[51513] = i[51513];
  assign o[51512] = i[51512];
  assign o[51511] = i[51511];
  assign o[51510] = i[51510];
  assign o[51509] = i[51509];
  assign o[51508] = i[51508];
  assign o[51507] = i[51507];
  assign o[51506] = i[51506];
  assign o[51505] = i[51505];
  assign o[51504] = i[51504];
  assign o[51503] = i[51503];
  assign o[51502] = i[51502];
  assign o[51501] = i[51501];
  assign o[51500] = i[51500];
  assign o[51499] = i[51499];
  assign o[51498] = i[51498];
  assign o[51497] = i[51497];
  assign o[51496] = i[51496];
  assign o[51495] = i[51495];
  assign o[51494] = i[51494];
  assign o[51493] = i[51493];
  assign o[51492] = i[51492];
  assign o[51491] = i[51491];
  assign o[51490] = i[51490];
  assign o[51489] = i[51489];
  assign o[51488] = i[51488];
  assign o[51487] = i[51487];
  assign o[51486] = i[51486];
  assign o[51485] = i[51485];
  assign o[51484] = i[51484];
  assign o[51483] = i[51483];
  assign o[51482] = i[51482];
  assign o[51481] = i[51481];
  assign o[51480] = i[51480];
  assign o[51479] = i[51479];
  assign o[51478] = i[51478];
  assign o[51477] = i[51477];
  assign o[51476] = i[51476];
  assign o[51475] = i[51475];
  assign o[51474] = i[51474];
  assign o[51473] = i[51473];
  assign o[51472] = i[51472];
  assign o[51471] = i[51471];
  assign o[51470] = i[51470];
  assign o[51469] = i[51469];
  assign o[51468] = i[51468];
  assign o[51467] = i[51467];
  assign o[51466] = i[51466];
  assign o[51465] = i[51465];
  assign o[51464] = i[51464];
  assign o[51463] = i[51463];
  assign o[51462] = i[51462];
  assign o[51461] = i[51461];
  assign o[51460] = i[51460];
  assign o[51459] = i[51459];
  assign o[51458] = i[51458];
  assign o[51457] = i[51457];
  assign o[51456] = i[51456];
  assign o[51455] = i[51455];
  assign o[51454] = i[51454];
  assign o[51453] = i[51453];
  assign o[51452] = i[51452];
  assign o[51451] = i[51451];
  assign o[51450] = i[51450];
  assign o[51449] = i[51449];
  assign o[51448] = i[51448];
  assign o[51447] = i[51447];
  assign o[51446] = i[51446];
  assign o[51445] = i[51445];
  assign o[51444] = i[51444];
  assign o[51443] = i[51443];
  assign o[51442] = i[51442];
  assign o[51441] = i[51441];
  assign o[51440] = i[51440];
  assign o[51439] = i[51439];
  assign o[51438] = i[51438];
  assign o[51437] = i[51437];
  assign o[51436] = i[51436];
  assign o[51435] = i[51435];
  assign o[51434] = i[51434];
  assign o[51433] = i[51433];
  assign o[51432] = i[51432];
  assign o[51431] = i[51431];
  assign o[51430] = i[51430];
  assign o[51429] = i[51429];
  assign o[51428] = i[51428];
  assign o[51427] = i[51427];
  assign o[51426] = i[51426];
  assign o[51425] = i[51425];
  assign o[51424] = i[51424];
  assign o[51423] = i[51423];
  assign o[51422] = i[51422];
  assign o[51421] = i[51421];
  assign o[51420] = i[51420];
  assign o[51419] = i[51419];
  assign o[51418] = i[51418];
  assign o[51417] = i[51417];
  assign o[51416] = i[51416];
  assign o[51415] = i[51415];
  assign o[51414] = i[51414];
  assign o[51413] = i[51413];
  assign o[51412] = i[51412];
  assign o[51411] = i[51411];
  assign o[51410] = i[51410];
  assign o[51409] = i[51409];
  assign o[51408] = i[51408];
  assign o[51407] = i[51407];
  assign o[51406] = i[51406];
  assign o[51405] = i[51405];
  assign o[51404] = i[51404];
  assign o[51403] = i[51403];
  assign o[51402] = i[51402];
  assign o[51401] = i[51401];
  assign o[51400] = i[51400];
  assign o[51399] = i[51399];
  assign o[51398] = i[51398];
  assign o[51397] = i[51397];
  assign o[51396] = i[51396];
  assign o[51395] = i[51395];
  assign o[51394] = i[51394];
  assign o[51393] = i[51393];
  assign o[51392] = i[51392];
  assign o[51391] = i[51391];
  assign o[51390] = i[51390];
  assign o[51389] = i[51389];
  assign o[51388] = i[51388];
  assign o[51387] = i[51387];
  assign o[51386] = i[51386];
  assign o[51385] = i[51385];
  assign o[51384] = i[51384];
  assign o[51383] = i[51383];
  assign o[51382] = i[51382];
  assign o[51381] = i[51381];
  assign o[51380] = i[51380];
  assign o[51379] = i[51379];
  assign o[51378] = i[51378];
  assign o[51377] = i[51377];
  assign o[51376] = i[51376];
  assign o[51375] = i[51375];
  assign o[51374] = i[51374];
  assign o[51373] = i[51373];
  assign o[51372] = i[51372];
  assign o[51371] = i[51371];
  assign o[51370] = i[51370];
  assign o[51369] = i[51369];
  assign o[51368] = i[51368];
  assign o[51367] = i[51367];
  assign o[51366] = i[51366];
  assign o[51365] = i[51365];
  assign o[51364] = i[51364];
  assign o[51363] = i[51363];
  assign o[51362] = i[51362];
  assign o[51361] = i[51361];
  assign o[51360] = i[51360];
  assign o[51359] = i[51359];
  assign o[51358] = i[51358];
  assign o[51357] = i[51357];
  assign o[51356] = i[51356];
  assign o[51355] = i[51355];
  assign o[51354] = i[51354];
  assign o[51353] = i[51353];
  assign o[51352] = i[51352];
  assign o[51351] = i[51351];
  assign o[51350] = i[51350];
  assign o[51349] = i[51349];
  assign o[51348] = i[51348];
  assign o[51347] = i[51347];
  assign o[51346] = i[51346];
  assign o[51345] = i[51345];
  assign o[51344] = i[51344];
  assign o[51343] = i[51343];
  assign o[51342] = i[51342];
  assign o[51341] = i[51341];
  assign o[51340] = i[51340];
  assign o[51339] = i[51339];
  assign o[51338] = i[51338];
  assign o[51337] = i[51337];
  assign o[51336] = i[51336];
  assign o[51335] = i[51335];
  assign o[51334] = i[51334];
  assign o[51333] = i[51333];
  assign o[51332] = i[51332];
  assign o[51331] = i[51331];
  assign o[51330] = i[51330];
  assign o[51329] = i[51329];
  assign o[51328] = i[51328];
  assign o[51327] = i[51327];
  assign o[51326] = i[51326];
  assign o[51325] = i[51325];
  assign o[51324] = i[51324];
  assign o[51323] = i[51323];
  assign o[51322] = i[51322];
  assign o[51321] = i[51321];
  assign o[51320] = i[51320];
  assign o[51319] = i[51319];
  assign o[51318] = i[51318];
  assign o[51317] = i[51317];
  assign o[51316] = i[51316];
  assign o[51315] = i[51315];
  assign o[51314] = i[51314];
  assign o[51313] = i[51313];
  assign o[51312] = i[51312];
  assign o[51311] = i[51311];
  assign o[51310] = i[51310];
  assign o[51309] = i[51309];
  assign o[51308] = i[51308];
  assign o[51307] = i[51307];
  assign o[51306] = i[51306];
  assign o[51305] = i[51305];
  assign o[51304] = i[51304];
  assign o[51303] = i[51303];
  assign o[51302] = i[51302];
  assign o[51301] = i[51301];
  assign o[51300] = i[51300];
  assign o[51299] = i[51299];
  assign o[51298] = i[51298];
  assign o[51297] = i[51297];
  assign o[51296] = i[51296];
  assign o[51295] = i[51295];
  assign o[51294] = i[51294];
  assign o[51293] = i[51293];
  assign o[51292] = i[51292];
  assign o[51291] = i[51291];
  assign o[51290] = i[51290];
  assign o[51289] = i[51289];
  assign o[51288] = i[51288];
  assign o[51287] = i[51287];
  assign o[51286] = i[51286];
  assign o[51285] = i[51285];
  assign o[51284] = i[51284];
  assign o[51283] = i[51283];
  assign o[51282] = i[51282];
  assign o[51281] = i[51281];
  assign o[51280] = i[51280];
  assign o[51279] = i[51279];
  assign o[51278] = i[51278];
  assign o[51277] = i[51277];
  assign o[51276] = i[51276];
  assign o[51275] = i[51275];
  assign o[51274] = i[51274];
  assign o[51273] = i[51273];
  assign o[51272] = i[51272];
  assign o[51271] = i[51271];
  assign o[51270] = i[51270];
  assign o[51269] = i[51269];
  assign o[51268] = i[51268];
  assign o[51267] = i[51267];
  assign o[51266] = i[51266];
  assign o[51265] = i[51265];
  assign o[51264] = i[51264];
  assign o[51263] = i[51263];
  assign o[51262] = i[51262];
  assign o[51261] = i[51261];
  assign o[51260] = i[51260];
  assign o[51259] = i[51259];
  assign o[51258] = i[51258];
  assign o[51257] = i[51257];
  assign o[51256] = i[51256];
  assign o[51255] = i[51255];
  assign o[51254] = i[51254];
  assign o[51253] = i[51253];
  assign o[51252] = i[51252];
  assign o[51251] = i[51251];
  assign o[51250] = i[51250];
  assign o[51249] = i[51249];
  assign o[51248] = i[51248];
  assign o[51247] = i[51247];
  assign o[51246] = i[51246];
  assign o[51245] = i[51245];
  assign o[51244] = i[51244];
  assign o[51243] = i[51243];
  assign o[51242] = i[51242];
  assign o[51241] = i[51241];
  assign o[51240] = i[51240];
  assign o[51239] = i[51239];
  assign o[51238] = i[51238];
  assign o[51237] = i[51237];
  assign o[51236] = i[51236];
  assign o[51235] = i[51235];
  assign o[51234] = i[51234];
  assign o[51233] = i[51233];
  assign o[51232] = i[51232];
  assign o[51231] = i[51231];
  assign o[51230] = i[51230];
  assign o[51229] = i[51229];
  assign o[51228] = i[51228];
  assign o[51227] = i[51227];
  assign o[51226] = i[51226];
  assign o[51225] = i[51225];
  assign o[51224] = i[51224];
  assign o[51223] = i[51223];
  assign o[51222] = i[51222];
  assign o[51221] = i[51221];
  assign o[51220] = i[51220];
  assign o[51219] = i[51219];
  assign o[51218] = i[51218];
  assign o[51217] = i[51217];
  assign o[51216] = i[51216];
  assign o[51215] = i[51215];
  assign o[51214] = i[51214];
  assign o[51213] = i[51213];
  assign o[51212] = i[51212];
  assign o[51211] = i[51211];
  assign o[51210] = i[51210];
  assign o[51209] = i[51209];
  assign o[51208] = i[51208];
  assign o[51207] = i[51207];
  assign o[51206] = i[51206];
  assign o[51205] = i[51205];
  assign o[51204] = i[51204];
  assign o[51203] = i[51203];
  assign o[51202] = i[51202];
  assign o[51201] = i[51201];
  assign o[51200] = i[51200];
  assign o[51199] = i[51199];
  assign o[51198] = i[51198];
  assign o[51197] = i[51197];
  assign o[51196] = i[51196];
  assign o[51195] = i[51195];
  assign o[51194] = i[51194];
  assign o[51193] = i[51193];
  assign o[51192] = i[51192];
  assign o[51191] = i[51191];
  assign o[51190] = i[51190];
  assign o[51189] = i[51189];
  assign o[51188] = i[51188];
  assign o[51187] = i[51187];
  assign o[51186] = i[51186];
  assign o[51185] = i[51185];
  assign o[51184] = i[51184];
  assign o[51183] = i[51183];
  assign o[51182] = i[51182];
  assign o[51181] = i[51181];
  assign o[51180] = i[51180];
  assign o[51179] = i[51179];
  assign o[51178] = i[51178];
  assign o[51177] = i[51177];
  assign o[51176] = i[51176];
  assign o[51175] = i[51175];
  assign o[51174] = i[51174];
  assign o[51173] = i[51173];
  assign o[51172] = i[51172];
  assign o[51171] = i[51171];
  assign o[51170] = i[51170];
  assign o[51169] = i[51169];
  assign o[51168] = i[51168];
  assign o[51167] = i[51167];
  assign o[51166] = i[51166];
  assign o[51165] = i[51165];
  assign o[51164] = i[51164];
  assign o[51163] = i[51163];
  assign o[51162] = i[51162];
  assign o[51161] = i[51161];
  assign o[51160] = i[51160];
  assign o[51159] = i[51159];
  assign o[51158] = i[51158];
  assign o[51157] = i[51157];
  assign o[51156] = i[51156];
  assign o[51155] = i[51155];
  assign o[51154] = i[51154];
  assign o[51153] = i[51153];
  assign o[51152] = i[51152];
  assign o[51151] = i[51151];
  assign o[51150] = i[51150];
  assign o[51149] = i[51149];
  assign o[51148] = i[51148];
  assign o[51147] = i[51147];
  assign o[51146] = i[51146];
  assign o[51145] = i[51145];
  assign o[51144] = i[51144];
  assign o[51143] = i[51143];
  assign o[51142] = i[51142];
  assign o[51141] = i[51141];
  assign o[51140] = i[51140];
  assign o[51139] = i[51139];
  assign o[51138] = i[51138];
  assign o[51137] = i[51137];
  assign o[51136] = i[51136];
  assign o[51135] = i[51135];
  assign o[51134] = i[51134];
  assign o[51133] = i[51133];
  assign o[51132] = i[51132];
  assign o[51131] = i[51131];
  assign o[51130] = i[51130];
  assign o[51129] = i[51129];
  assign o[51128] = i[51128];
  assign o[51127] = i[51127];
  assign o[51126] = i[51126];
  assign o[51125] = i[51125];
  assign o[51124] = i[51124];
  assign o[51123] = i[51123];
  assign o[51122] = i[51122];
  assign o[51121] = i[51121];
  assign o[51120] = i[51120];
  assign o[51119] = i[51119];
  assign o[51118] = i[51118];
  assign o[51117] = i[51117];
  assign o[51116] = i[51116];
  assign o[51115] = i[51115];
  assign o[51114] = i[51114];
  assign o[51113] = i[51113];
  assign o[51112] = i[51112];
  assign o[51111] = i[51111];
  assign o[51110] = i[51110];
  assign o[51109] = i[51109];
  assign o[51108] = i[51108];
  assign o[51107] = i[51107];
  assign o[51106] = i[51106];
  assign o[51105] = i[51105];
  assign o[51104] = i[51104];
  assign o[51103] = i[51103];
  assign o[51102] = i[51102];
  assign o[51101] = i[51101];
  assign o[51100] = i[51100];
  assign o[51099] = i[51099];
  assign o[51098] = i[51098];
  assign o[51097] = i[51097];
  assign o[51096] = i[51096];
  assign o[51095] = i[51095];
  assign o[51094] = i[51094];
  assign o[51093] = i[51093];
  assign o[51092] = i[51092];
  assign o[51091] = i[51091];
  assign o[51090] = i[51090];
  assign o[51089] = i[51089];
  assign o[51088] = i[51088];
  assign o[51087] = i[51087];
  assign o[51086] = i[51086];
  assign o[51085] = i[51085];
  assign o[51084] = i[51084];
  assign o[51083] = i[51083];
  assign o[51082] = i[51082];
  assign o[51081] = i[51081];
  assign o[51080] = i[51080];
  assign o[51079] = i[51079];
  assign o[51078] = i[51078];
  assign o[51077] = i[51077];
  assign o[51076] = i[51076];
  assign o[51075] = i[51075];
  assign o[51074] = i[51074];
  assign o[51073] = i[51073];
  assign o[51072] = i[51072];
  assign o[51071] = i[51071];
  assign o[51070] = i[51070];
  assign o[51069] = i[51069];
  assign o[51068] = i[51068];
  assign o[51067] = i[51067];
  assign o[51066] = i[51066];
  assign o[51065] = i[51065];
  assign o[51064] = i[51064];
  assign o[51063] = i[51063];
  assign o[51062] = i[51062];
  assign o[51061] = i[51061];
  assign o[51060] = i[51060];
  assign o[51059] = i[51059];
  assign o[51058] = i[51058];
  assign o[51057] = i[51057];
  assign o[51056] = i[51056];
  assign o[51055] = i[51055];
  assign o[51054] = i[51054];
  assign o[51053] = i[51053];
  assign o[51052] = i[51052];
  assign o[51051] = i[51051];
  assign o[51050] = i[51050];
  assign o[51049] = i[51049];
  assign o[51048] = i[51048];
  assign o[51047] = i[51047];
  assign o[51046] = i[51046];
  assign o[51045] = i[51045];
  assign o[51044] = i[51044];
  assign o[51043] = i[51043];
  assign o[51042] = i[51042];
  assign o[51041] = i[51041];
  assign o[51040] = i[51040];
  assign o[51039] = i[51039];
  assign o[51038] = i[51038];
  assign o[51037] = i[51037];
  assign o[51036] = i[51036];
  assign o[51035] = i[51035];
  assign o[51034] = i[51034];
  assign o[51033] = i[51033];
  assign o[51032] = i[51032];
  assign o[51031] = i[51031];
  assign o[51030] = i[51030];
  assign o[51029] = i[51029];
  assign o[51028] = i[51028];
  assign o[51027] = i[51027];
  assign o[51026] = i[51026];
  assign o[51025] = i[51025];
  assign o[51024] = i[51024];
  assign o[51023] = i[51023];
  assign o[51022] = i[51022];
  assign o[51021] = i[51021];
  assign o[51020] = i[51020];
  assign o[51019] = i[51019];
  assign o[51018] = i[51018];
  assign o[51017] = i[51017];
  assign o[51016] = i[51016];
  assign o[51015] = i[51015];
  assign o[51014] = i[51014];
  assign o[51013] = i[51013];
  assign o[51012] = i[51012];
  assign o[51011] = i[51011];
  assign o[51010] = i[51010];
  assign o[51009] = i[51009];
  assign o[51008] = i[51008];
  assign o[51007] = i[51007];
  assign o[51006] = i[51006];
  assign o[51005] = i[51005];
  assign o[51004] = i[51004];
  assign o[51003] = i[51003];
  assign o[51002] = i[51002];
  assign o[51001] = i[51001];
  assign o[51000] = i[51000];
  assign o[50999] = i[50999];
  assign o[50998] = i[50998];
  assign o[50997] = i[50997];
  assign o[50996] = i[50996];
  assign o[50995] = i[50995];
  assign o[50994] = i[50994];
  assign o[50993] = i[50993];
  assign o[50992] = i[50992];
  assign o[50991] = i[50991];
  assign o[50990] = i[50990];
  assign o[50989] = i[50989];
  assign o[50988] = i[50988];
  assign o[50987] = i[50987];
  assign o[50986] = i[50986];
  assign o[50985] = i[50985];
  assign o[50984] = i[50984];
  assign o[50983] = i[50983];
  assign o[50982] = i[50982];
  assign o[50981] = i[50981];
  assign o[50980] = i[50980];
  assign o[50979] = i[50979];
  assign o[50978] = i[50978];
  assign o[50977] = i[50977];
  assign o[50976] = i[50976];
  assign o[50975] = i[50975];
  assign o[50974] = i[50974];
  assign o[50973] = i[50973];
  assign o[50972] = i[50972];
  assign o[50971] = i[50971];
  assign o[50970] = i[50970];
  assign o[50969] = i[50969];
  assign o[50968] = i[50968];
  assign o[50967] = i[50967];
  assign o[50966] = i[50966];
  assign o[50965] = i[50965];
  assign o[50964] = i[50964];
  assign o[50963] = i[50963];
  assign o[50962] = i[50962];
  assign o[50961] = i[50961];
  assign o[50960] = i[50960];
  assign o[50959] = i[50959];
  assign o[50958] = i[50958];
  assign o[50957] = i[50957];
  assign o[50956] = i[50956];
  assign o[50955] = i[50955];
  assign o[50954] = i[50954];
  assign o[50953] = i[50953];
  assign o[50952] = i[50952];
  assign o[50951] = i[50951];
  assign o[50950] = i[50950];
  assign o[50949] = i[50949];
  assign o[50948] = i[50948];
  assign o[50947] = i[50947];
  assign o[50946] = i[50946];
  assign o[50945] = i[50945];
  assign o[50944] = i[50944];
  assign o[50943] = i[50943];
  assign o[50942] = i[50942];
  assign o[50941] = i[50941];
  assign o[50940] = i[50940];
  assign o[50939] = i[50939];
  assign o[50938] = i[50938];
  assign o[50937] = i[50937];
  assign o[50936] = i[50936];
  assign o[50935] = i[50935];
  assign o[50934] = i[50934];
  assign o[50933] = i[50933];
  assign o[50932] = i[50932];
  assign o[50931] = i[50931];
  assign o[50930] = i[50930];
  assign o[50929] = i[50929];
  assign o[50928] = i[50928];
  assign o[50927] = i[50927];
  assign o[50926] = i[50926];
  assign o[50925] = i[50925];
  assign o[50924] = i[50924];
  assign o[50923] = i[50923];
  assign o[50922] = i[50922];
  assign o[50921] = i[50921];
  assign o[50920] = i[50920];
  assign o[50919] = i[50919];
  assign o[50918] = i[50918];
  assign o[50917] = i[50917];
  assign o[50916] = i[50916];
  assign o[50915] = i[50915];
  assign o[50914] = i[50914];
  assign o[50913] = i[50913];
  assign o[50912] = i[50912];
  assign o[50911] = i[50911];
  assign o[50910] = i[50910];
  assign o[50909] = i[50909];
  assign o[50908] = i[50908];
  assign o[50907] = i[50907];
  assign o[50906] = i[50906];
  assign o[50905] = i[50905];
  assign o[50904] = i[50904];
  assign o[50903] = i[50903];
  assign o[50902] = i[50902];
  assign o[50901] = i[50901];
  assign o[50900] = i[50900];
  assign o[50899] = i[50899];
  assign o[50898] = i[50898];
  assign o[50897] = i[50897];
  assign o[50896] = i[50896];
  assign o[50895] = i[50895];
  assign o[50894] = i[50894];
  assign o[50893] = i[50893];
  assign o[50892] = i[50892];
  assign o[50891] = i[50891];
  assign o[50890] = i[50890];
  assign o[50889] = i[50889];
  assign o[50888] = i[50888];
  assign o[50887] = i[50887];
  assign o[50886] = i[50886];
  assign o[50885] = i[50885];
  assign o[50884] = i[50884];
  assign o[50883] = i[50883];
  assign o[50882] = i[50882];
  assign o[50881] = i[50881];
  assign o[50880] = i[50880];
  assign o[50879] = i[50879];
  assign o[50878] = i[50878];
  assign o[50877] = i[50877];
  assign o[50876] = i[50876];
  assign o[50875] = i[50875];
  assign o[50874] = i[50874];
  assign o[50873] = i[50873];
  assign o[50872] = i[50872];
  assign o[50871] = i[50871];
  assign o[50870] = i[50870];
  assign o[50869] = i[50869];
  assign o[50868] = i[50868];
  assign o[50867] = i[50867];
  assign o[50866] = i[50866];
  assign o[50865] = i[50865];
  assign o[50864] = i[50864];
  assign o[50863] = i[50863];
  assign o[50862] = i[50862];
  assign o[50861] = i[50861];
  assign o[50860] = i[50860];
  assign o[50859] = i[50859];
  assign o[50858] = i[50858];
  assign o[50857] = i[50857];
  assign o[50856] = i[50856];
  assign o[50855] = i[50855];
  assign o[50854] = i[50854];
  assign o[50853] = i[50853];
  assign o[50852] = i[50852];
  assign o[50851] = i[50851];
  assign o[50850] = i[50850];
  assign o[50849] = i[50849];
  assign o[50848] = i[50848];
  assign o[50847] = i[50847];
  assign o[50846] = i[50846];
  assign o[50845] = i[50845];
  assign o[50844] = i[50844];
  assign o[50843] = i[50843];
  assign o[50842] = i[50842];
  assign o[50841] = i[50841];
  assign o[50840] = i[50840];
  assign o[50839] = i[50839];
  assign o[50838] = i[50838];
  assign o[50837] = i[50837];
  assign o[50836] = i[50836];
  assign o[50835] = i[50835];
  assign o[50834] = i[50834];
  assign o[50833] = i[50833];
  assign o[50832] = i[50832];
  assign o[50831] = i[50831];
  assign o[50830] = i[50830];
  assign o[50829] = i[50829];
  assign o[50828] = i[50828];
  assign o[50827] = i[50827];
  assign o[50826] = i[50826];
  assign o[50825] = i[50825];
  assign o[50824] = i[50824];
  assign o[50823] = i[50823];
  assign o[50822] = i[50822];
  assign o[50821] = i[50821];
  assign o[50820] = i[50820];
  assign o[50819] = i[50819];
  assign o[50818] = i[50818];
  assign o[50817] = i[50817];
  assign o[50816] = i[50816];
  assign o[50815] = i[50815];
  assign o[50814] = i[50814];
  assign o[50813] = i[50813];
  assign o[50812] = i[50812];
  assign o[50811] = i[50811];
  assign o[50810] = i[50810];
  assign o[50809] = i[50809];
  assign o[50808] = i[50808];
  assign o[50807] = i[50807];
  assign o[50806] = i[50806];
  assign o[50805] = i[50805];
  assign o[50804] = i[50804];
  assign o[50803] = i[50803];
  assign o[50802] = i[50802];
  assign o[50801] = i[50801];
  assign o[50800] = i[50800];
  assign o[50799] = i[50799];
  assign o[50798] = i[50798];
  assign o[50797] = i[50797];
  assign o[50796] = i[50796];
  assign o[50795] = i[50795];
  assign o[50794] = i[50794];
  assign o[50793] = i[50793];
  assign o[50792] = i[50792];
  assign o[50791] = i[50791];
  assign o[50790] = i[50790];
  assign o[50789] = i[50789];
  assign o[50788] = i[50788];
  assign o[50787] = i[50787];
  assign o[50786] = i[50786];
  assign o[50785] = i[50785];
  assign o[50784] = i[50784];
  assign o[50783] = i[50783];
  assign o[50782] = i[50782];
  assign o[50781] = i[50781];
  assign o[50780] = i[50780];
  assign o[50779] = i[50779];
  assign o[50778] = i[50778];
  assign o[50777] = i[50777];
  assign o[50776] = i[50776];
  assign o[50775] = i[50775];
  assign o[50774] = i[50774];
  assign o[50773] = i[50773];
  assign o[50772] = i[50772];
  assign o[50771] = i[50771];
  assign o[50770] = i[50770];
  assign o[50769] = i[50769];
  assign o[50768] = i[50768];
  assign o[50767] = i[50767];
  assign o[50766] = i[50766];
  assign o[50765] = i[50765];
  assign o[50764] = i[50764];
  assign o[50763] = i[50763];
  assign o[50762] = i[50762];
  assign o[50761] = i[50761];
  assign o[50760] = i[50760];
  assign o[50759] = i[50759];
  assign o[50758] = i[50758];
  assign o[50757] = i[50757];
  assign o[50756] = i[50756];
  assign o[50755] = i[50755];
  assign o[50754] = i[50754];
  assign o[50753] = i[50753];
  assign o[50752] = i[50752];
  assign o[50751] = i[50751];
  assign o[50750] = i[50750];
  assign o[50749] = i[50749];
  assign o[50748] = i[50748];
  assign o[50747] = i[50747];
  assign o[50746] = i[50746];
  assign o[50745] = i[50745];
  assign o[50744] = i[50744];
  assign o[50743] = i[50743];
  assign o[50742] = i[50742];
  assign o[50741] = i[50741];
  assign o[50740] = i[50740];
  assign o[50739] = i[50739];
  assign o[50738] = i[50738];
  assign o[50737] = i[50737];
  assign o[50736] = i[50736];
  assign o[50735] = i[50735];
  assign o[50734] = i[50734];
  assign o[50733] = i[50733];
  assign o[50732] = i[50732];
  assign o[50731] = i[50731];
  assign o[50730] = i[50730];
  assign o[50729] = i[50729];
  assign o[50728] = i[50728];
  assign o[50727] = i[50727];
  assign o[50726] = i[50726];
  assign o[50725] = i[50725];
  assign o[50724] = i[50724];
  assign o[50723] = i[50723];
  assign o[50722] = i[50722];
  assign o[50721] = i[50721];
  assign o[50720] = i[50720];
  assign o[50719] = i[50719];
  assign o[50718] = i[50718];
  assign o[50717] = i[50717];
  assign o[50716] = i[50716];
  assign o[50715] = i[50715];
  assign o[50714] = i[50714];
  assign o[50713] = i[50713];
  assign o[50712] = i[50712];
  assign o[50711] = i[50711];
  assign o[50710] = i[50710];
  assign o[50709] = i[50709];
  assign o[50708] = i[50708];
  assign o[50707] = i[50707];
  assign o[50706] = i[50706];
  assign o[50705] = i[50705];
  assign o[50704] = i[50704];
  assign o[50703] = i[50703];
  assign o[50702] = i[50702];
  assign o[50701] = i[50701];
  assign o[50700] = i[50700];
  assign o[50699] = i[50699];
  assign o[50698] = i[50698];
  assign o[50697] = i[50697];
  assign o[50696] = i[50696];
  assign o[50695] = i[50695];
  assign o[50694] = i[50694];
  assign o[50693] = i[50693];
  assign o[50692] = i[50692];
  assign o[50691] = i[50691];
  assign o[50690] = i[50690];
  assign o[50689] = i[50689];
  assign o[50688] = i[50688];
  assign o[50687] = i[50687];
  assign o[50686] = i[50686];
  assign o[50685] = i[50685];
  assign o[50684] = i[50684];
  assign o[50683] = i[50683];
  assign o[50682] = i[50682];
  assign o[50681] = i[50681];
  assign o[50680] = i[50680];
  assign o[50679] = i[50679];
  assign o[50678] = i[50678];
  assign o[50677] = i[50677];
  assign o[50676] = i[50676];
  assign o[50675] = i[50675];
  assign o[50674] = i[50674];
  assign o[50673] = i[50673];
  assign o[50672] = i[50672];
  assign o[50671] = i[50671];
  assign o[50670] = i[50670];
  assign o[50669] = i[50669];
  assign o[50668] = i[50668];
  assign o[50667] = i[50667];
  assign o[50666] = i[50666];
  assign o[50665] = i[50665];
  assign o[50664] = i[50664];
  assign o[50663] = i[50663];
  assign o[50662] = i[50662];
  assign o[50661] = i[50661];
  assign o[50660] = i[50660];
  assign o[50659] = i[50659];
  assign o[50658] = i[50658];
  assign o[50657] = i[50657];
  assign o[50656] = i[50656];
  assign o[50655] = i[50655];
  assign o[50654] = i[50654];
  assign o[50653] = i[50653];
  assign o[50652] = i[50652];
  assign o[50651] = i[50651];
  assign o[50650] = i[50650];
  assign o[50649] = i[50649];
  assign o[50648] = i[50648];
  assign o[50647] = i[50647];
  assign o[50646] = i[50646];
  assign o[50645] = i[50645];
  assign o[50644] = i[50644];
  assign o[50643] = i[50643];
  assign o[50642] = i[50642];
  assign o[50641] = i[50641];
  assign o[50640] = i[50640];
  assign o[50639] = i[50639];
  assign o[50638] = i[50638];
  assign o[50637] = i[50637];
  assign o[50636] = i[50636];
  assign o[50635] = i[50635];
  assign o[50634] = i[50634];
  assign o[50633] = i[50633];
  assign o[50632] = i[50632];
  assign o[50631] = i[50631];
  assign o[50630] = i[50630];
  assign o[50629] = i[50629];
  assign o[50628] = i[50628];
  assign o[50627] = i[50627];
  assign o[50626] = i[50626];
  assign o[50625] = i[50625];
  assign o[50624] = i[50624];
  assign o[50623] = i[50623];
  assign o[50622] = i[50622];
  assign o[50621] = i[50621];
  assign o[50620] = i[50620];
  assign o[50619] = i[50619];
  assign o[50618] = i[50618];
  assign o[50617] = i[50617];
  assign o[50616] = i[50616];
  assign o[50615] = i[50615];
  assign o[50614] = i[50614];
  assign o[50613] = i[50613];
  assign o[50612] = i[50612];
  assign o[50611] = i[50611];
  assign o[50610] = i[50610];
  assign o[50609] = i[50609];
  assign o[50608] = i[50608];
  assign o[50607] = i[50607];
  assign o[50606] = i[50606];
  assign o[50605] = i[50605];
  assign o[50604] = i[50604];
  assign o[50603] = i[50603];
  assign o[50602] = i[50602];
  assign o[50601] = i[50601];
  assign o[50600] = i[50600];
  assign o[50599] = i[50599];
  assign o[50598] = i[50598];
  assign o[50597] = i[50597];
  assign o[50596] = i[50596];
  assign o[50595] = i[50595];
  assign o[50594] = i[50594];
  assign o[50593] = i[50593];
  assign o[50592] = i[50592];
  assign o[50591] = i[50591];
  assign o[50590] = i[50590];
  assign o[50589] = i[50589];
  assign o[50588] = i[50588];
  assign o[50587] = i[50587];
  assign o[50586] = i[50586];
  assign o[50585] = i[50585];
  assign o[50584] = i[50584];
  assign o[50583] = i[50583];
  assign o[50582] = i[50582];
  assign o[50581] = i[50581];
  assign o[50580] = i[50580];
  assign o[50579] = i[50579];
  assign o[50578] = i[50578];
  assign o[50577] = i[50577];
  assign o[50576] = i[50576];
  assign o[50575] = i[50575];
  assign o[50574] = i[50574];
  assign o[50573] = i[50573];
  assign o[50572] = i[50572];
  assign o[50571] = i[50571];
  assign o[50570] = i[50570];
  assign o[50569] = i[50569];
  assign o[50568] = i[50568];
  assign o[50567] = i[50567];
  assign o[50566] = i[50566];
  assign o[50565] = i[50565];
  assign o[50564] = i[50564];
  assign o[50563] = i[50563];
  assign o[50562] = i[50562];
  assign o[50561] = i[50561];
  assign o[50560] = i[50560];
  assign o[50559] = i[50559];
  assign o[50558] = i[50558];
  assign o[50557] = i[50557];
  assign o[50556] = i[50556];
  assign o[50555] = i[50555];
  assign o[50554] = i[50554];
  assign o[50553] = i[50553];
  assign o[50552] = i[50552];
  assign o[50551] = i[50551];
  assign o[50550] = i[50550];
  assign o[50549] = i[50549];
  assign o[50548] = i[50548];
  assign o[50547] = i[50547];
  assign o[50546] = i[50546];
  assign o[50545] = i[50545];
  assign o[50544] = i[50544];
  assign o[50543] = i[50543];
  assign o[50542] = i[50542];
  assign o[50541] = i[50541];
  assign o[50540] = i[50540];
  assign o[50539] = i[50539];
  assign o[50538] = i[50538];
  assign o[50537] = i[50537];
  assign o[50536] = i[50536];
  assign o[50535] = i[50535];
  assign o[50534] = i[50534];
  assign o[50533] = i[50533];
  assign o[50532] = i[50532];
  assign o[50531] = i[50531];
  assign o[50530] = i[50530];
  assign o[50529] = i[50529];
  assign o[50528] = i[50528];
  assign o[50527] = i[50527];
  assign o[50526] = i[50526];
  assign o[50525] = i[50525];
  assign o[50524] = i[50524];
  assign o[50523] = i[50523];
  assign o[50522] = i[50522];
  assign o[50521] = i[50521];
  assign o[50520] = i[50520];
  assign o[50519] = i[50519];
  assign o[50518] = i[50518];
  assign o[50517] = i[50517];
  assign o[50516] = i[50516];
  assign o[50515] = i[50515];
  assign o[50514] = i[50514];
  assign o[50513] = i[50513];
  assign o[50512] = i[50512];
  assign o[50511] = i[50511];
  assign o[50510] = i[50510];
  assign o[50509] = i[50509];
  assign o[50508] = i[50508];
  assign o[50507] = i[50507];
  assign o[50506] = i[50506];
  assign o[50505] = i[50505];
  assign o[50504] = i[50504];
  assign o[50503] = i[50503];
  assign o[50502] = i[50502];
  assign o[50501] = i[50501];
  assign o[50500] = i[50500];
  assign o[50499] = i[50499];
  assign o[50498] = i[50498];
  assign o[50497] = i[50497];
  assign o[50496] = i[50496];
  assign o[50495] = i[50495];
  assign o[50494] = i[50494];
  assign o[50493] = i[50493];
  assign o[50492] = i[50492];
  assign o[50491] = i[50491];
  assign o[50490] = i[50490];
  assign o[50489] = i[50489];
  assign o[50488] = i[50488];
  assign o[50487] = i[50487];
  assign o[50486] = i[50486];
  assign o[50485] = i[50485];
  assign o[50484] = i[50484];
  assign o[50483] = i[50483];
  assign o[50482] = i[50482];
  assign o[50481] = i[50481];
  assign o[50480] = i[50480];
  assign o[50479] = i[50479];
  assign o[50478] = i[50478];
  assign o[50477] = i[50477];
  assign o[50476] = i[50476];
  assign o[50475] = i[50475];
  assign o[50474] = i[50474];
  assign o[50473] = i[50473];
  assign o[50472] = i[50472];
  assign o[50471] = i[50471];
  assign o[50470] = i[50470];
  assign o[50469] = i[50469];
  assign o[50468] = i[50468];
  assign o[50467] = i[50467];
  assign o[50466] = i[50466];
  assign o[50465] = i[50465];
  assign o[50464] = i[50464];
  assign o[50463] = i[50463];
  assign o[50462] = i[50462];
  assign o[50461] = i[50461];
  assign o[50460] = i[50460];
  assign o[50459] = i[50459];
  assign o[50458] = i[50458];
  assign o[50457] = i[50457];
  assign o[50456] = i[50456];
  assign o[50455] = i[50455];
  assign o[50454] = i[50454];
  assign o[50453] = i[50453];
  assign o[50452] = i[50452];
  assign o[50451] = i[50451];
  assign o[50450] = i[50450];
  assign o[50449] = i[50449];
  assign o[50448] = i[50448];
  assign o[50447] = i[50447];
  assign o[50446] = i[50446];
  assign o[50445] = i[50445];
  assign o[50444] = i[50444];
  assign o[50443] = i[50443];
  assign o[50442] = i[50442];
  assign o[50441] = i[50441];
  assign o[50440] = i[50440];
  assign o[50439] = i[50439];
  assign o[50438] = i[50438];
  assign o[50437] = i[50437];
  assign o[50436] = i[50436];
  assign o[50435] = i[50435];
  assign o[50434] = i[50434];
  assign o[50433] = i[50433];
  assign o[50432] = i[50432];
  assign o[50431] = i[50431];
  assign o[50430] = i[50430];
  assign o[50429] = i[50429];
  assign o[50428] = i[50428];
  assign o[50427] = i[50427];
  assign o[50426] = i[50426];
  assign o[50425] = i[50425];
  assign o[50424] = i[50424];
  assign o[50423] = i[50423];
  assign o[50422] = i[50422];
  assign o[50421] = i[50421];
  assign o[50420] = i[50420];
  assign o[50419] = i[50419];
  assign o[50418] = i[50418];
  assign o[50417] = i[50417];
  assign o[50416] = i[50416];
  assign o[50415] = i[50415];
  assign o[50414] = i[50414];
  assign o[50413] = i[50413];
  assign o[50412] = i[50412];
  assign o[50411] = i[50411];
  assign o[50410] = i[50410];
  assign o[50409] = i[50409];
  assign o[50408] = i[50408];
  assign o[50407] = i[50407];
  assign o[50406] = i[50406];
  assign o[50405] = i[50405];
  assign o[50404] = i[50404];
  assign o[50403] = i[50403];
  assign o[50402] = i[50402];
  assign o[50401] = i[50401];
  assign o[50400] = i[50400];
  assign o[50399] = i[50399];
  assign o[50398] = i[50398];
  assign o[50397] = i[50397];
  assign o[50396] = i[50396];
  assign o[50395] = i[50395];
  assign o[50394] = i[50394];
  assign o[50393] = i[50393];
  assign o[50392] = i[50392];
  assign o[50391] = i[50391];
  assign o[50390] = i[50390];
  assign o[50389] = i[50389];
  assign o[50388] = i[50388];
  assign o[50387] = i[50387];
  assign o[50386] = i[50386];
  assign o[50385] = i[50385];
  assign o[50384] = i[50384];
  assign o[50383] = i[50383];
  assign o[50382] = i[50382];
  assign o[50381] = i[50381];
  assign o[50380] = i[50380];
  assign o[50379] = i[50379];
  assign o[50378] = i[50378];
  assign o[50377] = i[50377];
  assign o[50376] = i[50376];
  assign o[50375] = i[50375];
  assign o[50374] = i[50374];
  assign o[50373] = i[50373];
  assign o[50372] = i[50372];
  assign o[50371] = i[50371];
  assign o[50370] = i[50370];
  assign o[50369] = i[50369];
  assign o[50368] = i[50368];
  assign o[50367] = i[50367];
  assign o[50366] = i[50366];
  assign o[50365] = i[50365];
  assign o[50364] = i[50364];
  assign o[50363] = i[50363];
  assign o[50362] = i[50362];
  assign o[50361] = i[50361];
  assign o[50360] = i[50360];
  assign o[50359] = i[50359];
  assign o[50358] = i[50358];
  assign o[50357] = i[50357];
  assign o[50356] = i[50356];
  assign o[50355] = i[50355];
  assign o[50354] = i[50354];
  assign o[50353] = i[50353];
  assign o[50352] = i[50352];
  assign o[50351] = i[50351];
  assign o[50350] = i[50350];
  assign o[50349] = i[50349];
  assign o[50348] = i[50348];
  assign o[50347] = i[50347];
  assign o[50346] = i[50346];
  assign o[50345] = i[50345];
  assign o[50344] = i[50344];
  assign o[50343] = i[50343];
  assign o[50342] = i[50342];
  assign o[50341] = i[50341];
  assign o[50340] = i[50340];
  assign o[50339] = i[50339];
  assign o[50338] = i[50338];
  assign o[50337] = i[50337];
  assign o[50336] = i[50336];
  assign o[50335] = i[50335];
  assign o[50334] = i[50334];
  assign o[50333] = i[50333];
  assign o[50332] = i[50332];
  assign o[50331] = i[50331];
  assign o[50330] = i[50330];
  assign o[50329] = i[50329];
  assign o[50328] = i[50328];
  assign o[50327] = i[50327];
  assign o[50326] = i[50326];
  assign o[50325] = i[50325];
  assign o[50324] = i[50324];
  assign o[50323] = i[50323];
  assign o[50322] = i[50322];
  assign o[50321] = i[50321];
  assign o[50320] = i[50320];
  assign o[50319] = i[50319];
  assign o[50318] = i[50318];
  assign o[50317] = i[50317];
  assign o[50316] = i[50316];
  assign o[50315] = i[50315];
  assign o[50314] = i[50314];
  assign o[50313] = i[50313];
  assign o[50312] = i[50312];
  assign o[50311] = i[50311];
  assign o[50310] = i[50310];
  assign o[50309] = i[50309];
  assign o[50308] = i[50308];
  assign o[50307] = i[50307];
  assign o[50306] = i[50306];
  assign o[50305] = i[50305];
  assign o[50304] = i[50304];
  assign o[50303] = i[50303];
  assign o[50302] = i[50302];
  assign o[50301] = i[50301];
  assign o[50300] = i[50300];
  assign o[50299] = i[50299];
  assign o[50298] = i[50298];
  assign o[50297] = i[50297];
  assign o[50296] = i[50296];
  assign o[50295] = i[50295];
  assign o[50294] = i[50294];
  assign o[50293] = i[50293];
  assign o[50292] = i[50292];
  assign o[50291] = i[50291];
  assign o[50290] = i[50290];
  assign o[50289] = i[50289];
  assign o[50288] = i[50288];
  assign o[50287] = i[50287];
  assign o[50286] = i[50286];
  assign o[50285] = i[50285];
  assign o[50284] = i[50284];
  assign o[50283] = i[50283];
  assign o[50282] = i[50282];
  assign o[50281] = i[50281];
  assign o[50280] = i[50280];
  assign o[50279] = i[50279];
  assign o[50278] = i[50278];
  assign o[50277] = i[50277];
  assign o[50276] = i[50276];
  assign o[50275] = i[50275];
  assign o[50274] = i[50274];
  assign o[50273] = i[50273];
  assign o[50272] = i[50272];
  assign o[50271] = i[50271];
  assign o[50270] = i[50270];
  assign o[50269] = i[50269];
  assign o[50268] = i[50268];
  assign o[50267] = i[50267];
  assign o[50266] = i[50266];
  assign o[50265] = i[50265];
  assign o[50264] = i[50264];
  assign o[50263] = i[50263];
  assign o[50262] = i[50262];
  assign o[50261] = i[50261];
  assign o[50260] = i[50260];
  assign o[50259] = i[50259];
  assign o[50258] = i[50258];
  assign o[50257] = i[50257];
  assign o[50256] = i[50256];
  assign o[50255] = i[50255];
  assign o[50254] = i[50254];
  assign o[50253] = i[50253];
  assign o[50252] = i[50252];
  assign o[50251] = i[50251];
  assign o[50250] = i[50250];
  assign o[50249] = i[50249];
  assign o[50248] = i[50248];
  assign o[50247] = i[50247];
  assign o[50246] = i[50246];
  assign o[50245] = i[50245];
  assign o[50244] = i[50244];
  assign o[50243] = i[50243];
  assign o[50242] = i[50242];
  assign o[50241] = i[50241];
  assign o[50240] = i[50240];
  assign o[50239] = i[50239];
  assign o[50238] = i[50238];
  assign o[50237] = i[50237];
  assign o[50236] = i[50236];
  assign o[50235] = i[50235];
  assign o[50234] = i[50234];
  assign o[50233] = i[50233];
  assign o[50232] = i[50232];
  assign o[50231] = i[50231];
  assign o[50230] = i[50230];
  assign o[50229] = i[50229];
  assign o[50228] = i[50228];
  assign o[50227] = i[50227];
  assign o[50226] = i[50226];
  assign o[50225] = i[50225];
  assign o[50224] = i[50224];
  assign o[50223] = i[50223];
  assign o[50222] = i[50222];
  assign o[50221] = i[50221];
  assign o[50220] = i[50220];
  assign o[50219] = i[50219];
  assign o[50218] = i[50218];
  assign o[50217] = i[50217];
  assign o[50216] = i[50216];
  assign o[50215] = i[50215];
  assign o[50214] = i[50214];
  assign o[50213] = i[50213];
  assign o[50212] = i[50212];
  assign o[50211] = i[50211];
  assign o[50210] = i[50210];
  assign o[50209] = i[50209];
  assign o[50208] = i[50208];
  assign o[50207] = i[50207];
  assign o[50206] = i[50206];
  assign o[50205] = i[50205];
  assign o[50204] = i[50204];
  assign o[50203] = i[50203];
  assign o[50202] = i[50202];
  assign o[50201] = i[50201];
  assign o[50200] = i[50200];
  assign o[50199] = i[50199];
  assign o[50198] = i[50198];
  assign o[50197] = i[50197];
  assign o[50196] = i[50196];
  assign o[50195] = i[50195];
  assign o[50194] = i[50194];
  assign o[50193] = i[50193];
  assign o[50192] = i[50192];
  assign o[50191] = i[50191];
  assign o[50190] = i[50190];
  assign o[50189] = i[50189];
  assign o[50188] = i[50188];
  assign o[50187] = i[50187];
  assign o[50186] = i[50186];
  assign o[50185] = i[50185];
  assign o[50184] = i[50184];
  assign o[50183] = i[50183];
  assign o[50182] = i[50182];
  assign o[50181] = i[50181];
  assign o[50180] = i[50180];
  assign o[50179] = i[50179];
  assign o[50178] = i[50178];
  assign o[50177] = i[50177];
  assign o[50176] = i[50176];
  assign o[50175] = i[50175];
  assign o[50174] = i[50174];
  assign o[50173] = i[50173];
  assign o[50172] = i[50172];
  assign o[50171] = i[50171];
  assign o[50170] = i[50170];
  assign o[50169] = i[50169];
  assign o[50168] = i[50168];
  assign o[50167] = i[50167];
  assign o[50166] = i[50166];
  assign o[50165] = i[50165];
  assign o[50164] = i[50164];
  assign o[50163] = i[50163];
  assign o[50162] = i[50162];
  assign o[50161] = i[50161];
  assign o[50160] = i[50160];
  assign o[50159] = i[50159];
  assign o[50158] = i[50158];
  assign o[50157] = i[50157];
  assign o[50156] = i[50156];
  assign o[50155] = i[50155];
  assign o[50154] = i[50154];
  assign o[50153] = i[50153];
  assign o[50152] = i[50152];
  assign o[50151] = i[50151];
  assign o[50150] = i[50150];
  assign o[50149] = i[50149];
  assign o[50148] = i[50148];
  assign o[50147] = i[50147];
  assign o[50146] = i[50146];
  assign o[50145] = i[50145];
  assign o[50144] = i[50144];
  assign o[50143] = i[50143];
  assign o[50142] = i[50142];
  assign o[50141] = i[50141];
  assign o[50140] = i[50140];
  assign o[50139] = i[50139];
  assign o[50138] = i[50138];
  assign o[50137] = i[50137];
  assign o[50136] = i[50136];
  assign o[50135] = i[50135];
  assign o[50134] = i[50134];
  assign o[50133] = i[50133];
  assign o[50132] = i[50132];
  assign o[50131] = i[50131];
  assign o[50130] = i[50130];
  assign o[50129] = i[50129];
  assign o[50128] = i[50128];
  assign o[50127] = i[50127];
  assign o[50126] = i[50126];
  assign o[50125] = i[50125];
  assign o[50124] = i[50124];
  assign o[50123] = i[50123];
  assign o[50122] = i[50122];
  assign o[50121] = i[50121];
  assign o[50120] = i[50120];
  assign o[50119] = i[50119];
  assign o[50118] = i[50118];
  assign o[50117] = i[50117];
  assign o[50116] = i[50116];
  assign o[50115] = i[50115];
  assign o[50114] = i[50114];
  assign o[50113] = i[50113];
  assign o[50112] = i[50112];
  assign o[50111] = i[50111];
  assign o[50110] = i[50110];
  assign o[50109] = i[50109];
  assign o[50108] = i[50108];
  assign o[50107] = i[50107];
  assign o[50106] = i[50106];
  assign o[50105] = i[50105];
  assign o[50104] = i[50104];
  assign o[50103] = i[50103];
  assign o[50102] = i[50102];
  assign o[50101] = i[50101];
  assign o[50100] = i[50100];
  assign o[50099] = i[50099];
  assign o[50098] = i[50098];
  assign o[50097] = i[50097];
  assign o[50096] = i[50096];
  assign o[50095] = i[50095];
  assign o[50094] = i[50094];
  assign o[50093] = i[50093];
  assign o[50092] = i[50092];
  assign o[50091] = i[50091];
  assign o[50090] = i[50090];
  assign o[50089] = i[50089];
  assign o[50088] = i[50088];
  assign o[50087] = i[50087];
  assign o[50086] = i[50086];
  assign o[50085] = i[50085];
  assign o[50084] = i[50084];
  assign o[50083] = i[50083];
  assign o[50082] = i[50082];
  assign o[50081] = i[50081];
  assign o[50080] = i[50080];
  assign o[50079] = i[50079];
  assign o[50078] = i[50078];
  assign o[50077] = i[50077];
  assign o[50076] = i[50076];
  assign o[50075] = i[50075];
  assign o[50074] = i[50074];
  assign o[50073] = i[50073];
  assign o[50072] = i[50072];
  assign o[50071] = i[50071];
  assign o[50070] = i[50070];
  assign o[50069] = i[50069];
  assign o[50068] = i[50068];
  assign o[50067] = i[50067];
  assign o[50066] = i[50066];
  assign o[50065] = i[50065];
  assign o[50064] = i[50064];
  assign o[50063] = i[50063];
  assign o[50062] = i[50062];
  assign o[50061] = i[50061];
  assign o[50060] = i[50060];
  assign o[50059] = i[50059];
  assign o[50058] = i[50058];
  assign o[50057] = i[50057];
  assign o[50056] = i[50056];
  assign o[50055] = i[50055];
  assign o[50054] = i[50054];
  assign o[50053] = i[50053];
  assign o[50052] = i[50052];
  assign o[50051] = i[50051];
  assign o[50050] = i[50050];
  assign o[50049] = i[50049];
  assign o[50048] = i[50048];
  assign o[50047] = i[50047];
  assign o[50046] = i[50046];
  assign o[50045] = i[50045];
  assign o[50044] = i[50044];
  assign o[50043] = i[50043];
  assign o[50042] = i[50042];
  assign o[50041] = i[50041];
  assign o[50040] = i[50040];
  assign o[50039] = i[50039];
  assign o[50038] = i[50038];
  assign o[50037] = i[50037];
  assign o[50036] = i[50036];
  assign o[50035] = i[50035];
  assign o[50034] = i[50034];
  assign o[50033] = i[50033];
  assign o[50032] = i[50032];
  assign o[50031] = i[50031];
  assign o[50030] = i[50030];
  assign o[50029] = i[50029];
  assign o[50028] = i[50028];
  assign o[50027] = i[50027];
  assign o[50026] = i[50026];
  assign o[50025] = i[50025];
  assign o[50024] = i[50024];
  assign o[50023] = i[50023];
  assign o[50022] = i[50022];
  assign o[50021] = i[50021];
  assign o[50020] = i[50020];
  assign o[50019] = i[50019];
  assign o[50018] = i[50018];
  assign o[50017] = i[50017];
  assign o[50016] = i[50016];
  assign o[50015] = i[50015];
  assign o[50014] = i[50014];
  assign o[50013] = i[50013];
  assign o[50012] = i[50012];
  assign o[50011] = i[50011];
  assign o[50010] = i[50010];
  assign o[50009] = i[50009];
  assign o[50008] = i[50008];
  assign o[50007] = i[50007];
  assign o[50006] = i[50006];
  assign o[50005] = i[50005];
  assign o[50004] = i[50004];
  assign o[50003] = i[50003];
  assign o[50002] = i[50002];
  assign o[50001] = i[50001];
  assign o[50000] = i[50000];
  assign o[49999] = i[49999];
  assign o[49998] = i[49998];
  assign o[49997] = i[49997];
  assign o[49996] = i[49996];
  assign o[49995] = i[49995];
  assign o[49994] = i[49994];
  assign o[49993] = i[49993];
  assign o[49992] = i[49992];
  assign o[49991] = i[49991];
  assign o[49990] = i[49990];
  assign o[49989] = i[49989];
  assign o[49988] = i[49988];
  assign o[49987] = i[49987];
  assign o[49986] = i[49986];
  assign o[49985] = i[49985];
  assign o[49984] = i[49984];
  assign o[49983] = i[49983];
  assign o[49982] = i[49982];
  assign o[49981] = i[49981];
  assign o[49980] = i[49980];
  assign o[49979] = i[49979];
  assign o[49978] = i[49978];
  assign o[49977] = i[49977];
  assign o[49976] = i[49976];
  assign o[49975] = i[49975];
  assign o[49974] = i[49974];
  assign o[49973] = i[49973];
  assign o[49972] = i[49972];
  assign o[49971] = i[49971];
  assign o[49970] = i[49970];
  assign o[49969] = i[49969];
  assign o[49968] = i[49968];
  assign o[49967] = i[49967];
  assign o[49966] = i[49966];
  assign o[49965] = i[49965];
  assign o[49964] = i[49964];
  assign o[49963] = i[49963];
  assign o[49962] = i[49962];
  assign o[49961] = i[49961];
  assign o[49960] = i[49960];
  assign o[49959] = i[49959];
  assign o[49958] = i[49958];
  assign o[49957] = i[49957];
  assign o[49956] = i[49956];
  assign o[49955] = i[49955];
  assign o[49954] = i[49954];
  assign o[49953] = i[49953];
  assign o[49952] = i[49952];
  assign o[49951] = i[49951];
  assign o[49950] = i[49950];
  assign o[49949] = i[49949];
  assign o[49948] = i[49948];
  assign o[49947] = i[49947];
  assign o[49946] = i[49946];
  assign o[49945] = i[49945];
  assign o[49944] = i[49944];
  assign o[49943] = i[49943];
  assign o[49942] = i[49942];
  assign o[49941] = i[49941];
  assign o[49940] = i[49940];
  assign o[49939] = i[49939];
  assign o[49938] = i[49938];
  assign o[49937] = i[49937];
  assign o[49936] = i[49936];
  assign o[49935] = i[49935];
  assign o[49934] = i[49934];
  assign o[49933] = i[49933];
  assign o[49932] = i[49932];
  assign o[49931] = i[49931];
  assign o[49930] = i[49930];
  assign o[49929] = i[49929];
  assign o[49928] = i[49928];
  assign o[49927] = i[49927];
  assign o[49926] = i[49926];
  assign o[49925] = i[49925];
  assign o[49924] = i[49924];
  assign o[49923] = i[49923];
  assign o[49922] = i[49922];
  assign o[49921] = i[49921];
  assign o[49920] = i[49920];
  assign o[49919] = i[49919];
  assign o[49918] = i[49918];
  assign o[49917] = i[49917];
  assign o[49916] = i[49916];
  assign o[49915] = i[49915];
  assign o[49914] = i[49914];
  assign o[49913] = i[49913];
  assign o[49912] = i[49912];
  assign o[49911] = i[49911];
  assign o[49910] = i[49910];
  assign o[49909] = i[49909];
  assign o[49908] = i[49908];
  assign o[49907] = i[49907];
  assign o[49906] = i[49906];
  assign o[49905] = i[49905];
  assign o[49904] = i[49904];
  assign o[49903] = i[49903];
  assign o[49902] = i[49902];
  assign o[49901] = i[49901];
  assign o[49900] = i[49900];
  assign o[49899] = i[49899];
  assign o[49898] = i[49898];
  assign o[49897] = i[49897];
  assign o[49896] = i[49896];
  assign o[49895] = i[49895];
  assign o[49894] = i[49894];
  assign o[49893] = i[49893];
  assign o[49892] = i[49892];
  assign o[49891] = i[49891];
  assign o[49890] = i[49890];
  assign o[49889] = i[49889];
  assign o[49888] = i[49888];
  assign o[49887] = i[49887];
  assign o[49886] = i[49886];
  assign o[49885] = i[49885];
  assign o[49884] = i[49884];
  assign o[49883] = i[49883];
  assign o[49882] = i[49882];
  assign o[49881] = i[49881];
  assign o[49880] = i[49880];
  assign o[49879] = i[49879];
  assign o[49878] = i[49878];
  assign o[49877] = i[49877];
  assign o[49876] = i[49876];
  assign o[49875] = i[49875];
  assign o[49874] = i[49874];
  assign o[49873] = i[49873];
  assign o[49872] = i[49872];
  assign o[49871] = i[49871];
  assign o[49870] = i[49870];
  assign o[49869] = i[49869];
  assign o[49868] = i[49868];
  assign o[49867] = i[49867];
  assign o[49866] = i[49866];
  assign o[49865] = i[49865];
  assign o[49864] = i[49864];
  assign o[49863] = i[49863];
  assign o[49862] = i[49862];
  assign o[49861] = i[49861];
  assign o[49860] = i[49860];
  assign o[49859] = i[49859];
  assign o[49858] = i[49858];
  assign o[49857] = i[49857];
  assign o[49856] = i[49856];
  assign o[49855] = i[49855];
  assign o[49854] = i[49854];
  assign o[49853] = i[49853];
  assign o[49852] = i[49852];
  assign o[49851] = i[49851];
  assign o[49850] = i[49850];
  assign o[49849] = i[49849];
  assign o[49848] = i[49848];
  assign o[49847] = i[49847];
  assign o[49846] = i[49846];
  assign o[49845] = i[49845];
  assign o[49844] = i[49844];
  assign o[49843] = i[49843];
  assign o[49842] = i[49842];
  assign o[49841] = i[49841];
  assign o[49840] = i[49840];
  assign o[49839] = i[49839];
  assign o[49838] = i[49838];
  assign o[49837] = i[49837];
  assign o[49836] = i[49836];
  assign o[49835] = i[49835];
  assign o[49834] = i[49834];
  assign o[49833] = i[49833];
  assign o[49832] = i[49832];
  assign o[49831] = i[49831];
  assign o[49830] = i[49830];
  assign o[49829] = i[49829];
  assign o[49828] = i[49828];
  assign o[49827] = i[49827];
  assign o[49826] = i[49826];
  assign o[49825] = i[49825];
  assign o[49824] = i[49824];
  assign o[49823] = i[49823];
  assign o[49822] = i[49822];
  assign o[49821] = i[49821];
  assign o[49820] = i[49820];
  assign o[49819] = i[49819];
  assign o[49818] = i[49818];
  assign o[49817] = i[49817];
  assign o[49816] = i[49816];
  assign o[49815] = i[49815];
  assign o[49814] = i[49814];
  assign o[49813] = i[49813];
  assign o[49812] = i[49812];
  assign o[49811] = i[49811];
  assign o[49810] = i[49810];
  assign o[49809] = i[49809];
  assign o[49808] = i[49808];
  assign o[49807] = i[49807];
  assign o[49806] = i[49806];
  assign o[49805] = i[49805];
  assign o[49804] = i[49804];
  assign o[49803] = i[49803];
  assign o[49802] = i[49802];
  assign o[49801] = i[49801];
  assign o[49800] = i[49800];
  assign o[49799] = i[49799];
  assign o[49798] = i[49798];
  assign o[49797] = i[49797];
  assign o[49796] = i[49796];
  assign o[49795] = i[49795];
  assign o[49794] = i[49794];
  assign o[49793] = i[49793];
  assign o[49792] = i[49792];
  assign o[49791] = i[49791];
  assign o[49790] = i[49790];
  assign o[49789] = i[49789];
  assign o[49788] = i[49788];
  assign o[49787] = i[49787];
  assign o[49786] = i[49786];
  assign o[49785] = i[49785];
  assign o[49784] = i[49784];
  assign o[49783] = i[49783];
  assign o[49782] = i[49782];
  assign o[49781] = i[49781];
  assign o[49780] = i[49780];
  assign o[49779] = i[49779];
  assign o[49778] = i[49778];
  assign o[49777] = i[49777];
  assign o[49776] = i[49776];
  assign o[49775] = i[49775];
  assign o[49774] = i[49774];
  assign o[49773] = i[49773];
  assign o[49772] = i[49772];
  assign o[49771] = i[49771];
  assign o[49770] = i[49770];
  assign o[49769] = i[49769];
  assign o[49768] = i[49768];
  assign o[49767] = i[49767];
  assign o[49766] = i[49766];
  assign o[49765] = i[49765];
  assign o[49764] = i[49764];
  assign o[49763] = i[49763];
  assign o[49762] = i[49762];
  assign o[49761] = i[49761];
  assign o[49760] = i[49760];
  assign o[49759] = i[49759];
  assign o[49758] = i[49758];
  assign o[49757] = i[49757];
  assign o[49756] = i[49756];
  assign o[49755] = i[49755];
  assign o[49754] = i[49754];
  assign o[49753] = i[49753];
  assign o[49752] = i[49752];
  assign o[49751] = i[49751];
  assign o[49750] = i[49750];
  assign o[49749] = i[49749];
  assign o[49748] = i[49748];
  assign o[49747] = i[49747];
  assign o[49746] = i[49746];
  assign o[49745] = i[49745];
  assign o[49744] = i[49744];
  assign o[49743] = i[49743];
  assign o[49742] = i[49742];
  assign o[49741] = i[49741];
  assign o[49740] = i[49740];
  assign o[49739] = i[49739];
  assign o[49738] = i[49738];
  assign o[49737] = i[49737];
  assign o[49736] = i[49736];
  assign o[49735] = i[49735];
  assign o[49734] = i[49734];
  assign o[49733] = i[49733];
  assign o[49732] = i[49732];
  assign o[49731] = i[49731];
  assign o[49730] = i[49730];
  assign o[49729] = i[49729];
  assign o[49728] = i[49728];
  assign o[49727] = i[49727];
  assign o[49726] = i[49726];
  assign o[49725] = i[49725];
  assign o[49724] = i[49724];
  assign o[49723] = i[49723];
  assign o[49722] = i[49722];
  assign o[49721] = i[49721];
  assign o[49720] = i[49720];
  assign o[49719] = i[49719];
  assign o[49718] = i[49718];
  assign o[49717] = i[49717];
  assign o[49716] = i[49716];
  assign o[49715] = i[49715];
  assign o[49714] = i[49714];
  assign o[49713] = i[49713];
  assign o[49712] = i[49712];
  assign o[49711] = i[49711];
  assign o[49710] = i[49710];
  assign o[49709] = i[49709];
  assign o[49708] = i[49708];
  assign o[49707] = i[49707];
  assign o[49706] = i[49706];
  assign o[49705] = i[49705];
  assign o[49704] = i[49704];
  assign o[49703] = i[49703];
  assign o[49702] = i[49702];
  assign o[49701] = i[49701];
  assign o[49700] = i[49700];
  assign o[49699] = i[49699];
  assign o[49698] = i[49698];
  assign o[49697] = i[49697];
  assign o[49696] = i[49696];
  assign o[49695] = i[49695];
  assign o[49694] = i[49694];
  assign o[49693] = i[49693];
  assign o[49692] = i[49692];
  assign o[49691] = i[49691];
  assign o[49690] = i[49690];
  assign o[49689] = i[49689];
  assign o[49688] = i[49688];
  assign o[49687] = i[49687];
  assign o[49686] = i[49686];
  assign o[49685] = i[49685];
  assign o[49684] = i[49684];
  assign o[49683] = i[49683];
  assign o[49682] = i[49682];
  assign o[49681] = i[49681];
  assign o[49680] = i[49680];
  assign o[49679] = i[49679];
  assign o[49678] = i[49678];
  assign o[49677] = i[49677];
  assign o[49676] = i[49676];
  assign o[49675] = i[49675];
  assign o[49674] = i[49674];
  assign o[49673] = i[49673];
  assign o[49672] = i[49672];
  assign o[49671] = i[49671];
  assign o[49670] = i[49670];
  assign o[49669] = i[49669];
  assign o[49668] = i[49668];
  assign o[49667] = i[49667];
  assign o[49666] = i[49666];
  assign o[49665] = i[49665];
  assign o[49664] = i[49664];
  assign o[49663] = i[49663];
  assign o[49662] = i[49662];
  assign o[49661] = i[49661];
  assign o[49660] = i[49660];
  assign o[49659] = i[49659];
  assign o[49658] = i[49658];
  assign o[49657] = i[49657];
  assign o[49656] = i[49656];
  assign o[49655] = i[49655];
  assign o[49654] = i[49654];
  assign o[49653] = i[49653];
  assign o[49652] = i[49652];
  assign o[49651] = i[49651];
  assign o[49650] = i[49650];
  assign o[49649] = i[49649];
  assign o[49648] = i[49648];
  assign o[49647] = i[49647];
  assign o[49646] = i[49646];
  assign o[49645] = i[49645];
  assign o[49644] = i[49644];
  assign o[49643] = i[49643];
  assign o[49642] = i[49642];
  assign o[49641] = i[49641];
  assign o[49640] = i[49640];
  assign o[49639] = i[49639];
  assign o[49638] = i[49638];
  assign o[49637] = i[49637];
  assign o[49636] = i[49636];
  assign o[49635] = i[49635];
  assign o[49634] = i[49634];
  assign o[49633] = i[49633];
  assign o[49632] = i[49632];
  assign o[49631] = i[49631];
  assign o[49630] = i[49630];
  assign o[49629] = i[49629];
  assign o[49628] = i[49628];
  assign o[49627] = i[49627];
  assign o[49626] = i[49626];
  assign o[49625] = i[49625];
  assign o[49624] = i[49624];
  assign o[49623] = i[49623];
  assign o[49622] = i[49622];
  assign o[49621] = i[49621];
  assign o[49620] = i[49620];
  assign o[49619] = i[49619];
  assign o[49618] = i[49618];
  assign o[49617] = i[49617];
  assign o[49616] = i[49616];
  assign o[49615] = i[49615];
  assign o[49614] = i[49614];
  assign o[49613] = i[49613];
  assign o[49612] = i[49612];
  assign o[49611] = i[49611];
  assign o[49610] = i[49610];
  assign o[49609] = i[49609];
  assign o[49608] = i[49608];
  assign o[49607] = i[49607];
  assign o[49606] = i[49606];
  assign o[49605] = i[49605];
  assign o[49604] = i[49604];
  assign o[49603] = i[49603];
  assign o[49602] = i[49602];
  assign o[49601] = i[49601];
  assign o[49600] = i[49600];
  assign o[49599] = i[49599];
  assign o[49598] = i[49598];
  assign o[49597] = i[49597];
  assign o[49596] = i[49596];
  assign o[49595] = i[49595];
  assign o[49594] = i[49594];
  assign o[49593] = i[49593];
  assign o[49592] = i[49592];
  assign o[49591] = i[49591];
  assign o[49590] = i[49590];
  assign o[49589] = i[49589];
  assign o[49588] = i[49588];
  assign o[49587] = i[49587];
  assign o[49586] = i[49586];
  assign o[49585] = i[49585];
  assign o[49584] = i[49584];
  assign o[49583] = i[49583];
  assign o[49582] = i[49582];
  assign o[49581] = i[49581];
  assign o[49580] = i[49580];
  assign o[49579] = i[49579];
  assign o[49578] = i[49578];
  assign o[49577] = i[49577];
  assign o[49576] = i[49576];
  assign o[49575] = i[49575];
  assign o[49574] = i[49574];
  assign o[49573] = i[49573];
  assign o[49572] = i[49572];
  assign o[49571] = i[49571];
  assign o[49570] = i[49570];
  assign o[49569] = i[49569];
  assign o[49568] = i[49568];
  assign o[49567] = i[49567];
  assign o[49566] = i[49566];
  assign o[49565] = i[49565];
  assign o[49564] = i[49564];
  assign o[49563] = i[49563];
  assign o[49562] = i[49562];
  assign o[49561] = i[49561];
  assign o[49560] = i[49560];
  assign o[49559] = i[49559];
  assign o[49558] = i[49558];
  assign o[49557] = i[49557];
  assign o[49556] = i[49556];
  assign o[49555] = i[49555];
  assign o[49554] = i[49554];
  assign o[49553] = i[49553];
  assign o[49552] = i[49552];
  assign o[49551] = i[49551];
  assign o[49550] = i[49550];
  assign o[49549] = i[49549];
  assign o[49548] = i[49548];
  assign o[49547] = i[49547];
  assign o[49546] = i[49546];
  assign o[49545] = i[49545];
  assign o[49544] = i[49544];
  assign o[49543] = i[49543];
  assign o[49542] = i[49542];
  assign o[49541] = i[49541];
  assign o[49540] = i[49540];
  assign o[49539] = i[49539];
  assign o[49538] = i[49538];
  assign o[49537] = i[49537];
  assign o[49536] = i[49536];
  assign o[49535] = i[49535];
  assign o[49534] = i[49534];
  assign o[49533] = i[49533];
  assign o[49532] = i[49532];
  assign o[49531] = i[49531];
  assign o[49530] = i[49530];
  assign o[49529] = i[49529];
  assign o[49528] = i[49528];
  assign o[49527] = i[49527];
  assign o[49526] = i[49526];
  assign o[49525] = i[49525];
  assign o[49524] = i[49524];
  assign o[49523] = i[49523];
  assign o[49522] = i[49522];
  assign o[49521] = i[49521];
  assign o[49520] = i[49520];
  assign o[49519] = i[49519];
  assign o[49518] = i[49518];
  assign o[49517] = i[49517];
  assign o[49516] = i[49516];
  assign o[49515] = i[49515];
  assign o[49514] = i[49514];
  assign o[49513] = i[49513];
  assign o[49512] = i[49512];
  assign o[49511] = i[49511];
  assign o[49510] = i[49510];
  assign o[49509] = i[49509];
  assign o[49508] = i[49508];
  assign o[49507] = i[49507];
  assign o[49506] = i[49506];
  assign o[49505] = i[49505];
  assign o[49504] = i[49504];
  assign o[49503] = i[49503];
  assign o[49502] = i[49502];
  assign o[49501] = i[49501];
  assign o[49500] = i[49500];
  assign o[49499] = i[49499];
  assign o[49498] = i[49498];
  assign o[49497] = i[49497];
  assign o[49496] = i[49496];
  assign o[49495] = i[49495];
  assign o[49494] = i[49494];
  assign o[49493] = i[49493];
  assign o[49492] = i[49492];
  assign o[49491] = i[49491];
  assign o[49490] = i[49490];
  assign o[49489] = i[49489];
  assign o[49488] = i[49488];
  assign o[49487] = i[49487];
  assign o[49486] = i[49486];
  assign o[49485] = i[49485];
  assign o[49484] = i[49484];
  assign o[49483] = i[49483];
  assign o[49482] = i[49482];
  assign o[49481] = i[49481];
  assign o[49480] = i[49480];
  assign o[49479] = i[49479];
  assign o[49478] = i[49478];
  assign o[49477] = i[49477];
  assign o[49476] = i[49476];
  assign o[49475] = i[49475];
  assign o[49474] = i[49474];
  assign o[49473] = i[49473];
  assign o[49472] = i[49472];
  assign o[49471] = i[49471];
  assign o[49470] = i[49470];
  assign o[49469] = i[49469];
  assign o[49468] = i[49468];
  assign o[49467] = i[49467];
  assign o[49466] = i[49466];
  assign o[49465] = i[49465];
  assign o[49464] = i[49464];
  assign o[49463] = i[49463];
  assign o[49462] = i[49462];
  assign o[49461] = i[49461];
  assign o[49460] = i[49460];
  assign o[49459] = i[49459];
  assign o[49458] = i[49458];
  assign o[49457] = i[49457];
  assign o[49456] = i[49456];
  assign o[49455] = i[49455];
  assign o[49454] = i[49454];
  assign o[49453] = i[49453];
  assign o[49452] = i[49452];
  assign o[49451] = i[49451];
  assign o[49450] = i[49450];
  assign o[49449] = i[49449];
  assign o[49448] = i[49448];
  assign o[49447] = i[49447];
  assign o[49446] = i[49446];
  assign o[49445] = i[49445];
  assign o[49444] = i[49444];
  assign o[49443] = i[49443];
  assign o[49442] = i[49442];
  assign o[49441] = i[49441];
  assign o[49440] = i[49440];
  assign o[49439] = i[49439];
  assign o[49438] = i[49438];
  assign o[49437] = i[49437];
  assign o[49436] = i[49436];
  assign o[49435] = i[49435];
  assign o[49434] = i[49434];
  assign o[49433] = i[49433];
  assign o[49432] = i[49432];
  assign o[49431] = i[49431];
  assign o[49430] = i[49430];
  assign o[49429] = i[49429];
  assign o[49428] = i[49428];
  assign o[49427] = i[49427];
  assign o[49426] = i[49426];
  assign o[49425] = i[49425];
  assign o[49424] = i[49424];
  assign o[49423] = i[49423];
  assign o[49422] = i[49422];
  assign o[49421] = i[49421];
  assign o[49420] = i[49420];
  assign o[49419] = i[49419];
  assign o[49418] = i[49418];
  assign o[49417] = i[49417];
  assign o[49416] = i[49416];
  assign o[49415] = i[49415];
  assign o[49414] = i[49414];
  assign o[49413] = i[49413];
  assign o[49412] = i[49412];
  assign o[49411] = i[49411];
  assign o[49410] = i[49410];
  assign o[49409] = i[49409];
  assign o[49408] = i[49408];
  assign o[49407] = i[49407];
  assign o[49406] = i[49406];
  assign o[49405] = i[49405];
  assign o[49404] = i[49404];
  assign o[49403] = i[49403];
  assign o[49402] = i[49402];
  assign o[49401] = i[49401];
  assign o[49400] = i[49400];
  assign o[49399] = i[49399];
  assign o[49398] = i[49398];
  assign o[49397] = i[49397];
  assign o[49396] = i[49396];
  assign o[49395] = i[49395];
  assign o[49394] = i[49394];
  assign o[49393] = i[49393];
  assign o[49392] = i[49392];
  assign o[49391] = i[49391];
  assign o[49390] = i[49390];
  assign o[49389] = i[49389];
  assign o[49388] = i[49388];
  assign o[49387] = i[49387];
  assign o[49386] = i[49386];
  assign o[49385] = i[49385];
  assign o[49384] = i[49384];
  assign o[49383] = i[49383];
  assign o[49382] = i[49382];
  assign o[49381] = i[49381];
  assign o[49380] = i[49380];
  assign o[49379] = i[49379];
  assign o[49378] = i[49378];
  assign o[49377] = i[49377];
  assign o[49376] = i[49376];
  assign o[49375] = i[49375];
  assign o[49374] = i[49374];
  assign o[49373] = i[49373];
  assign o[49372] = i[49372];
  assign o[49371] = i[49371];
  assign o[49370] = i[49370];
  assign o[49369] = i[49369];
  assign o[49368] = i[49368];
  assign o[49367] = i[49367];
  assign o[49366] = i[49366];
  assign o[49365] = i[49365];
  assign o[49364] = i[49364];
  assign o[49363] = i[49363];
  assign o[49362] = i[49362];
  assign o[49361] = i[49361];
  assign o[49360] = i[49360];
  assign o[49359] = i[49359];
  assign o[49358] = i[49358];
  assign o[49357] = i[49357];
  assign o[49356] = i[49356];
  assign o[49355] = i[49355];
  assign o[49354] = i[49354];
  assign o[49353] = i[49353];
  assign o[49352] = i[49352];
  assign o[49351] = i[49351];
  assign o[49350] = i[49350];
  assign o[49349] = i[49349];
  assign o[49348] = i[49348];
  assign o[49347] = i[49347];
  assign o[49346] = i[49346];
  assign o[49345] = i[49345];
  assign o[49344] = i[49344];
  assign o[49343] = i[49343];
  assign o[49342] = i[49342];
  assign o[49341] = i[49341];
  assign o[49340] = i[49340];
  assign o[49339] = i[49339];
  assign o[49338] = i[49338];
  assign o[49337] = i[49337];
  assign o[49336] = i[49336];
  assign o[49335] = i[49335];
  assign o[49334] = i[49334];
  assign o[49333] = i[49333];
  assign o[49332] = i[49332];
  assign o[49331] = i[49331];
  assign o[49330] = i[49330];
  assign o[49329] = i[49329];
  assign o[49328] = i[49328];
  assign o[49327] = i[49327];
  assign o[49326] = i[49326];
  assign o[49325] = i[49325];
  assign o[49324] = i[49324];
  assign o[49323] = i[49323];
  assign o[49322] = i[49322];
  assign o[49321] = i[49321];
  assign o[49320] = i[49320];
  assign o[49319] = i[49319];
  assign o[49318] = i[49318];
  assign o[49317] = i[49317];
  assign o[49316] = i[49316];
  assign o[49315] = i[49315];
  assign o[49314] = i[49314];
  assign o[49313] = i[49313];
  assign o[49312] = i[49312];
  assign o[49311] = i[49311];
  assign o[49310] = i[49310];
  assign o[49309] = i[49309];
  assign o[49308] = i[49308];
  assign o[49307] = i[49307];
  assign o[49306] = i[49306];
  assign o[49305] = i[49305];
  assign o[49304] = i[49304];
  assign o[49303] = i[49303];
  assign o[49302] = i[49302];
  assign o[49301] = i[49301];
  assign o[49300] = i[49300];
  assign o[49299] = i[49299];
  assign o[49298] = i[49298];
  assign o[49297] = i[49297];
  assign o[49296] = i[49296];
  assign o[49295] = i[49295];
  assign o[49294] = i[49294];
  assign o[49293] = i[49293];
  assign o[49292] = i[49292];
  assign o[49291] = i[49291];
  assign o[49290] = i[49290];
  assign o[49289] = i[49289];
  assign o[49288] = i[49288];
  assign o[49287] = i[49287];
  assign o[49286] = i[49286];
  assign o[49285] = i[49285];
  assign o[49284] = i[49284];
  assign o[49283] = i[49283];
  assign o[49282] = i[49282];
  assign o[49281] = i[49281];
  assign o[49280] = i[49280];
  assign o[49279] = i[49279];
  assign o[49278] = i[49278];
  assign o[49277] = i[49277];
  assign o[49276] = i[49276];
  assign o[49275] = i[49275];
  assign o[49274] = i[49274];
  assign o[49273] = i[49273];
  assign o[49272] = i[49272];
  assign o[49271] = i[49271];
  assign o[49270] = i[49270];
  assign o[49269] = i[49269];
  assign o[49268] = i[49268];
  assign o[49267] = i[49267];
  assign o[49266] = i[49266];
  assign o[49265] = i[49265];
  assign o[49264] = i[49264];
  assign o[49263] = i[49263];
  assign o[49262] = i[49262];
  assign o[49261] = i[49261];
  assign o[49260] = i[49260];
  assign o[49259] = i[49259];
  assign o[49258] = i[49258];
  assign o[49257] = i[49257];
  assign o[49256] = i[49256];
  assign o[49255] = i[49255];
  assign o[49254] = i[49254];
  assign o[49253] = i[49253];
  assign o[49252] = i[49252];
  assign o[49251] = i[49251];
  assign o[49250] = i[49250];
  assign o[49249] = i[49249];
  assign o[49248] = i[49248];
  assign o[49247] = i[49247];
  assign o[49246] = i[49246];
  assign o[49245] = i[49245];
  assign o[49244] = i[49244];
  assign o[49243] = i[49243];
  assign o[49242] = i[49242];
  assign o[49241] = i[49241];
  assign o[49240] = i[49240];
  assign o[49239] = i[49239];
  assign o[49238] = i[49238];
  assign o[49237] = i[49237];
  assign o[49236] = i[49236];
  assign o[49235] = i[49235];
  assign o[49234] = i[49234];
  assign o[49233] = i[49233];
  assign o[49232] = i[49232];
  assign o[49231] = i[49231];
  assign o[49230] = i[49230];
  assign o[49229] = i[49229];
  assign o[49228] = i[49228];
  assign o[49227] = i[49227];
  assign o[49226] = i[49226];
  assign o[49225] = i[49225];
  assign o[49224] = i[49224];
  assign o[49223] = i[49223];
  assign o[49222] = i[49222];
  assign o[49221] = i[49221];
  assign o[49220] = i[49220];
  assign o[49219] = i[49219];
  assign o[49218] = i[49218];
  assign o[49217] = i[49217];
  assign o[49216] = i[49216];
  assign o[49215] = i[49215];
  assign o[49214] = i[49214];
  assign o[49213] = i[49213];
  assign o[49212] = i[49212];
  assign o[49211] = i[49211];
  assign o[49210] = i[49210];
  assign o[49209] = i[49209];
  assign o[49208] = i[49208];
  assign o[49207] = i[49207];
  assign o[49206] = i[49206];
  assign o[49205] = i[49205];
  assign o[49204] = i[49204];
  assign o[49203] = i[49203];
  assign o[49202] = i[49202];
  assign o[49201] = i[49201];
  assign o[49200] = i[49200];
  assign o[49199] = i[49199];
  assign o[49198] = i[49198];
  assign o[49197] = i[49197];
  assign o[49196] = i[49196];
  assign o[49195] = i[49195];
  assign o[49194] = i[49194];
  assign o[49193] = i[49193];
  assign o[49192] = i[49192];
  assign o[49191] = i[49191];
  assign o[49190] = i[49190];
  assign o[49189] = i[49189];
  assign o[49188] = i[49188];
  assign o[49187] = i[49187];
  assign o[49186] = i[49186];
  assign o[49185] = i[49185];
  assign o[49184] = i[49184];
  assign o[49183] = i[49183];
  assign o[49182] = i[49182];
  assign o[49181] = i[49181];
  assign o[49180] = i[49180];
  assign o[49179] = i[49179];
  assign o[49178] = i[49178];
  assign o[49177] = i[49177];
  assign o[49176] = i[49176];
  assign o[49175] = i[49175];
  assign o[49174] = i[49174];
  assign o[49173] = i[49173];
  assign o[49172] = i[49172];
  assign o[49171] = i[49171];
  assign o[49170] = i[49170];
  assign o[49169] = i[49169];
  assign o[49168] = i[49168];
  assign o[49167] = i[49167];
  assign o[49166] = i[49166];
  assign o[49165] = i[49165];
  assign o[49164] = i[49164];
  assign o[49163] = i[49163];
  assign o[49162] = i[49162];
  assign o[49161] = i[49161];
  assign o[49160] = i[49160];
  assign o[49159] = i[49159];
  assign o[49158] = i[49158];
  assign o[49157] = i[49157];
  assign o[49156] = i[49156];
  assign o[49155] = i[49155];
  assign o[49154] = i[49154];
  assign o[49153] = i[49153];
  assign o[49152] = i[49152];
  assign o[49151] = i[49151];
  assign o[49150] = i[49150];
  assign o[49149] = i[49149];
  assign o[49148] = i[49148];
  assign o[49147] = i[49147];
  assign o[49146] = i[49146];
  assign o[49145] = i[49145];
  assign o[49144] = i[49144];
  assign o[49143] = i[49143];
  assign o[49142] = i[49142];
  assign o[49141] = i[49141];
  assign o[49140] = i[49140];
  assign o[49139] = i[49139];
  assign o[49138] = i[49138];
  assign o[49137] = i[49137];
  assign o[49136] = i[49136];
  assign o[49135] = i[49135];
  assign o[49134] = i[49134];
  assign o[49133] = i[49133];
  assign o[49132] = i[49132];
  assign o[49131] = i[49131];
  assign o[49130] = i[49130];
  assign o[49129] = i[49129];
  assign o[49128] = i[49128];
  assign o[49127] = i[49127];
  assign o[49126] = i[49126];
  assign o[49125] = i[49125];
  assign o[49124] = i[49124];
  assign o[49123] = i[49123];
  assign o[49122] = i[49122];
  assign o[49121] = i[49121];
  assign o[49120] = i[49120];
  assign o[49119] = i[49119];
  assign o[49118] = i[49118];
  assign o[49117] = i[49117];
  assign o[49116] = i[49116];
  assign o[49115] = i[49115];
  assign o[49114] = i[49114];
  assign o[49113] = i[49113];
  assign o[49112] = i[49112];
  assign o[49111] = i[49111];
  assign o[49110] = i[49110];
  assign o[49109] = i[49109];
  assign o[49108] = i[49108];
  assign o[49107] = i[49107];
  assign o[49106] = i[49106];
  assign o[49105] = i[49105];
  assign o[49104] = i[49104];
  assign o[49103] = i[49103];
  assign o[49102] = i[49102];
  assign o[49101] = i[49101];
  assign o[49100] = i[49100];
  assign o[49099] = i[49099];
  assign o[49098] = i[49098];
  assign o[49097] = i[49097];
  assign o[49096] = i[49096];
  assign o[49095] = i[49095];
  assign o[49094] = i[49094];
  assign o[49093] = i[49093];
  assign o[49092] = i[49092];
  assign o[49091] = i[49091];
  assign o[49090] = i[49090];
  assign o[49089] = i[49089];
  assign o[49088] = i[49088];
  assign o[49087] = i[49087];
  assign o[49086] = i[49086];
  assign o[49085] = i[49085];
  assign o[49084] = i[49084];
  assign o[49083] = i[49083];
  assign o[49082] = i[49082];
  assign o[49081] = i[49081];
  assign o[49080] = i[49080];
  assign o[49079] = i[49079];
  assign o[49078] = i[49078];
  assign o[49077] = i[49077];
  assign o[49076] = i[49076];
  assign o[49075] = i[49075];
  assign o[49074] = i[49074];
  assign o[49073] = i[49073];
  assign o[49072] = i[49072];
  assign o[49071] = i[49071];
  assign o[49070] = i[49070];
  assign o[49069] = i[49069];
  assign o[49068] = i[49068];
  assign o[49067] = i[49067];
  assign o[49066] = i[49066];
  assign o[49065] = i[49065];
  assign o[49064] = i[49064];
  assign o[49063] = i[49063];
  assign o[49062] = i[49062];
  assign o[49061] = i[49061];
  assign o[49060] = i[49060];
  assign o[49059] = i[49059];
  assign o[49058] = i[49058];
  assign o[49057] = i[49057];
  assign o[49056] = i[49056];
  assign o[49055] = i[49055];
  assign o[49054] = i[49054];
  assign o[49053] = i[49053];
  assign o[49052] = i[49052];
  assign o[49051] = i[49051];
  assign o[49050] = i[49050];
  assign o[49049] = i[49049];
  assign o[49048] = i[49048];
  assign o[49047] = i[49047];
  assign o[49046] = i[49046];
  assign o[49045] = i[49045];
  assign o[49044] = i[49044];
  assign o[49043] = i[49043];
  assign o[49042] = i[49042];
  assign o[49041] = i[49041];
  assign o[49040] = i[49040];
  assign o[49039] = i[49039];
  assign o[49038] = i[49038];
  assign o[49037] = i[49037];
  assign o[49036] = i[49036];
  assign o[49035] = i[49035];
  assign o[49034] = i[49034];
  assign o[49033] = i[49033];
  assign o[49032] = i[49032];
  assign o[49031] = i[49031];
  assign o[49030] = i[49030];
  assign o[49029] = i[49029];
  assign o[49028] = i[49028];
  assign o[49027] = i[49027];
  assign o[49026] = i[49026];
  assign o[49025] = i[49025];
  assign o[49024] = i[49024];
  assign o[49023] = i[49023];
  assign o[49022] = i[49022];
  assign o[49021] = i[49021];
  assign o[49020] = i[49020];
  assign o[49019] = i[49019];
  assign o[49018] = i[49018];
  assign o[49017] = i[49017];
  assign o[49016] = i[49016];
  assign o[49015] = i[49015];
  assign o[49014] = i[49014];
  assign o[49013] = i[49013];
  assign o[49012] = i[49012];
  assign o[49011] = i[49011];
  assign o[49010] = i[49010];
  assign o[49009] = i[49009];
  assign o[49008] = i[49008];
  assign o[49007] = i[49007];
  assign o[49006] = i[49006];
  assign o[49005] = i[49005];
  assign o[49004] = i[49004];
  assign o[49003] = i[49003];
  assign o[49002] = i[49002];
  assign o[49001] = i[49001];
  assign o[49000] = i[49000];
  assign o[48999] = i[48999];
  assign o[48998] = i[48998];
  assign o[48997] = i[48997];
  assign o[48996] = i[48996];
  assign o[48995] = i[48995];
  assign o[48994] = i[48994];
  assign o[48993] = i[48993];
  assign o[48992] = i[48992];
  assign o[48991] = i[48991];
  assign o[48990] = i[48990];
  assign o[48989] = i[48989];
  assign o[48988] = i[48988];
  assign o[48987] = i[48987];
  assign o[48986] = i[48986];
  assign o[48985] = i[48985];
  assign o[48984] = i[48984];
  assign o[48983] = i[48983];
  assign o[48982] = i[48982];
  assign o[48981] = i[48981];
  assign o[48980] = i[48980];
  assign o[48979] = i[48979];
  assign o[48978] = i[48978];
  assign o[48977] = i[48977];
  assign o[48976] = i[48976];
  assign o[48975] = i[48975];
  assign o[48974] = i[48974];
  assign o[48973] = i[48973];
  assign o[48972] = i[48972];
  assign o[48971] = i[48971];
  assign o[48970] = i[48970];
  assign o[48969] = i[48969];
  assign o[48968] = i[48968];
  assign o[48967] = i[48967];
  assign o[48966] = i[48966];
  assign o[48965] = i[48965];
  assign o[48964] = i[48964];
  assign o[48963] = i[48963];
  assign o[48962] = i[48962];
  assign o[48961] = i[48961];
  assign o[48960] = i[48960];
  assign o[48959] = i[48959];
  assign o[48958] = i[48958];
  assign o[48957] = i[48957];
  assign o[48956] = i[48956];
  assign o[48955] = i[48955];
  assign o[48954] = i[48954];
  assign o[48953] = i[48953];
  assign o[48952] = i[48952];
  assign o[48951] = i[48951];
  assign o[48950] = i[48950];
  assign o[48949] = i[48949];
  assign o[48948] = i[48948];
  assign o[48947] = i[48947];
  assign o[48946] = i[48946];
  assign o[48945] = i[48945];
  assign o[48944] = i[48944];
  assign o[48943] = i[48943];
  assign o[48942] = i[48942];
  assign o[48941] = i[48941];
  assign o[48940] = i[48940];
  assign o[48939] = i[48939];
  assign o[48938] = i[48938];
  assign o[48937] = i[48937];
  assign o[48936] = i[48936];
  assign o[48935] = i[48935];
  assign o[48934] = i[48934];
  assign o[48933] = i[48933];
  assign o[48932] = i[48932];
  assign o[48931] = i[48931];
  assign o[48930] = i[48930];
  assign o[48929] = i[48929];
  assign o[48928] = i[48928];
  assign o[48927] = i[48927];
  assign o[48926] = i[48926];
  assign o[48925] = i[48925];
  assign o[48924] = i[48924];
  assign o[48923] = i[48923];
  assign o[48922] = i[48922];
  assign o[48921] = i[48921];
  assign o[48920] = i[48920];
  assign o[48919] = i[48919];
  assign o[48918] = i[48918];
  assign o[48917] = i[48917];
  assign o[48916] = i[48916];
  assign o[48915] = i[48915];
  assign o[48914] = i[48914];
  assign o[48913] = i[48913];
  assign o[48912] = i[48912];
  assign o[48911] = i[48911];
  assign o[48910] = i[48910];
  assign o[48909] = i[48909];
  assign o[48908] = i[48908];
  assign o[48907] = i[48907];
  assign o[48906] = i[48906];
  assign o[48905] = i[48905];
  assign o[48904] = i[48904];
  assign o[48903] = i[48903];
  assign o[48902] = i[48902];
  assign o[48901] = i[48901];
  assign o[48900] = i[48900];
  assign o[48899] = i[48899];
  assign o[48898] = i[48898];
  assign o[48897] = i[48897];
  assign o[48896] = i[48896];
  assign o[48895] = i[48895];
  assign o[48894] = i[48894];
  assign o[48893] = i[48893];
  assign o[48892] = i[48892];
  assign o[48891] = i[48891];
  assign o[48890] = i[48890];
  assign o[48889] = i[48889];
  assign o[48888] = i[48888];
  assign o[48887] = i[48887];
  assign o[48886] = i[48886];
  assign o[48885] = i[48885];
  assign o[48884] = i[48884];
  assign o[48883] = i[48883];
  assign o[48882] = i[48882];
  assign o[48881] = i[48881];
  assign o[48880] = i[48880];
  assign o[48879] = i[48879];
  assign o[48878] = i[48878];
  assign o[48877] = i[48877];
  assign o[48876] = i[48876];
  assign o[48875] = i[48875];
  assign o[48874] = i[48874];
  assign o[48873] = i[48873];
  assign o[48872] = i[48872];
  assign o[48871] = i[48871];
  assign o[48870] = i[48870];
  assign o[48869] = i[48869];
  assign o[48868] = i[48868];
  assign o[48867] = i[48867];
  assign o[48866] = i[48866];
  assign o[48865] = i[48865];
  assign o[48864] = i[48864];
  assign o[48863] = i[48863];
  assign o[48862] = i[48862];
  assign o[48861] = i[48861];
  assign o[48860] = i[48860];
  assign o[48859] = i[48859];
  assign o[48858] = i[48858];
  assign o[48857] = i[48857];
  assign o[48856] = i[48856];
  assign o[48855] = i[48855];
  assign o[48854] = i[48854];
  assign o[48853] = i[48853];
  assign o[48852] = i[48852];
  assign o[48851] = i[48851];
  assign o[48850] = i[48850];
  assign o[48849] = i[48849];
  assign o[48848] = i[48848];
  assign o[48847] = i[48847];
  assign o[48846] = i[48846];
  assign o[48845] = i[48845];
  assign o[48844] = i[48844];
  assign o[48843] = i[48843];
  assign o[48842] = i[48842];
  assign o[48841] = i[48841];
  assign o[48840] = i[48840];
  assign o[48839] = i[48839];
  assign o[48838] = i[48838];
  assign o[48837] = i[48837];
  assign o[48836] = i[48836];
  assign o[48835] = i[48835];
  assign o[48834] = i[48834];
  assign o[48833] = i[48833];
  assign o[48832] = i[48832];
  assign o[48831] = i[48831];
  assign o[48830] = i[48830];
  assign o[48829] = i[48829];
  assign o[48828] = i[48828];
  assign o[48827] = i[48827];
  assign o[48826] = i[48826];
  assign o[48825] = i[48825];
  assign o[48824] = i[48824];
  assign o[48823] = i[48823];
  assign o[48822] = i[48822];
  assign o[48821] = i[48821];
  assign o[48820] = i[48820];
  assign o[48819] = i[48819];
  assign o[48818] = i[48818];
  assign o[48817] = i[48817];
  assign o[48816] = i[48816];
  assign o[48815] = i[48815];
  assign o[48814] = i[48814];
  assign o[48813] = i[48813];
  assign o[48812] = i[48812];
  assign o[48811] = i[48811];
  assign o[48810] = i[48810];
  assign o[48809] = i[48809];
  assign o[48808] = i[48808];
  assign o[48807] = i[48807];
  assign o[48806] = i[48806];
  assign o[48805] = i[48805];
  assign o[48804] = i[48804];
  assign o[48803] = i[48803];
  assign o[48802] = i[48802];
  assign o[48801] = i[48801];
  assign o[48800] = i[48800];
  assign o[48799] = i[48799];
  assign o[48798] = i[48798];
  assign o[48797] = i[48797];
  assign o[48796] = i[48796];
  assign o[48795] = i[48795];
  assign o[48794] = i[48794];
  assign o[48793] = i[48793];
  assign o[48792] = i[48792];
  assign o[48791] = i[48791];
  assign o[48790] = i[48790];
  assign o[48789] = i[48789];
  assign o[48788] = i[48788];
  assign o[48787] = i[48787];
  assign o[48786] = i[48786];
  assign o[48785] = i[48785];
  assign o[48784] = i[48784];
  assign o[48783] = i[48783];
  assign o[48782] = i[48782];
  assign o[48781] = i[48781];
  assign o[48780] = i[48780];
  assign o[48779] = i[48779];
  assign o[48778] = i[48778];
  assign o[48777] = i[48777];
  assign o[48776] = i[48776];
  assign o[48775] = i[48775];
  assign o[48774] = i[48774];
  assign o[48773] = i[48773];
  assign o[48772] = i[48772];
  assign o[48771] = i[48771];
  assign o[48770] = i[48770];
  assign o[48769] = i[48769];
  assign o[48768] = i[48768];
  assign o[48767] = i[48767];
  assign o[48766] = i[48766];
  assign o[48765] = i[48765];
  assign o[48764] = i[48764];
  assign o[48763] = i[48763];
  assign o[48762] = i[48762];
  assign o[48761] = i[48761];
  assign o[48760] = i[48760];
  assign o[48759] = i[48759];
  assign o[48758] = i[48758];
  assign o[48757] = i[48757];
  assign o[48756] = i[48756];
  assign o[48755] = i[48755];
  assign o[48754] = i[48754];
  assign o[48753] = i[48753];
  assign o[48752] = i[48752];
  assign o[48751] = i[48751];
  assign o[48750] = i[48750];
  assign o[48749] = i[48749];
  assign o[48748] = i[48748];
  assign o[48747] = i[48747];
  assign o[48746] = i[48746];
  assign o[48745] = i[48745];
  assign o[48744] = i[48744];
  assign o[48743] = i[48743];
  assign o[48742] = i[48742];
  assign o[48741] = i[48741];
  assign o[48740] = i[48740];
  assign o[48739] = i[48739];
  assign o[48738] = i[48738];
  assign o[48737] = i[48737];
  assign o[48736] = i[48736];
  assign o[48735] = i[48735];
  assign o[48734] = i[48734];
  assign o[48733] = i[48733];
  assign o[48732] = i[48732];
  assign o[48731] = i[48731];
  assign o[48730] = i[48730];
  assign o[48729] = i[48729];
  assign o[48728] = i[48728];
  assign o[48727] = i[48727];
  assign o[48726] = i[48726];
  assign o[48725] = i[48725];
  assign o[48724] = i[48724];
  assign o[48723] = i[48723];
  assign o[48722] = i[48722];
  assign o[48721] = i[48721];
  assign o[48720] = i[48720];
  assign o[48719] = i[48719];
  assign o[48718] = i[48718];
  assign o[48717] = i[48717];
  assign o[48716] = i[48716];
  assign o[48715] = i[48715];
  assign o[48714] = i[48714];
  assign o[48713] = i[48713];
  assign o[48712] = i[48712];
  assign o[48711] = i[48711];
  assign o[48710] = i[48710];
  assign o[48709] = i[48709];
  assign o[48708] = i[48708];
  assign o[48707] = i[48707];
  assign o[48706] = i[48706];
  assign o[48705] = i[48705];
  assign o[48704] = i[48704];
  assign o[48703] = i[48703];
  assign o[48702] = i[48702];
  assign o[48701] = i[48701];
  assign o[48700] = i[48700];
  assign o[48699] = i[48699];
  assign o[48698] = i[48698];
  assign o[48697] = i[48697];
  assign o[48696] = i[48696];
  assign o[48695] = i[48695];
  assign o[48694] = i[48694];
  assign o[48693] = i[48693];
  assign o[48692] = i[48692];
  assign o[48691] = i[48691];
  assign o[48690] = i[48690];
  assign o[48689] = i[48689];
  assign o[48688] = i[48688];
  assign o[48687] = i[48687];
  assign o[48686] = i[48686];
  assign o[48685] = i[48685];
  assign o[48684] = i[48684];
  assign o[48683] = i[48683];
  assign o[48682] = i[48682];
  assign o[48681] = i[48681];
  assign o[48680] = i[48680];
  assign o[48679] = i[48679];
  assign o[48678] = i[48678];
  assign o[48677] = i[48677];
  assign o[48676] = i[48676];
  assign o[48675] = i[48675];
  assign o[48674] = i[48674];
  assign o[48673] = i[48673];
  assign o[48672] = i[48672];
  assign o[48671] = i[48671];
  assign o[48670] = i[48670];
  assign o[48669] = i[48669];
  assign o[48668] = i[48668];
  assign o[48667] = i[48667];
  assign o[48666] = i[48666];
  assign o[48665] = i[48665];
  assign o[48664] = i[48664];
  assign o[48663] = i[48663];
  assign o[48662] = i[48662];
  assign o[48661] = i[48661];
  assign o[48660] = i[48660];
  assign o[48659] = i[48659];
  assign o[48658] = i[48658];
  assign o[48657] = i[48657];
  assign o[48656] = i[48656];
  assign o[48655] = i[48655];
  assign o[48654] = i[48654];
  assign o[48653] = i[48653];
  assign o[48652] = i[48652];
  assign o[48651] = i[48651];
  assign o[48650] = i[48650];
  assign o[48649] = i[48649];
  assign o[48648] = i[48648];
  assign o[48647] = i[48647];
  assign o[48646] = i[48646];
  assign o[48645] = i[48645];
  assign o[48644] = i[48644];
  assign o[48643] = i[48643];
  assign o[48642] = i[48642];
  assign o[48641] = i[48641];
  assign o[48640] = i[48640];
  assign o[48639] = i[48639];
  assign o[48638] = i[48638];
  assign o[48637] = i[48637];
  assign o[48636] = i[48636];
  assign o[48635] = i[48635];
  assign o[48634] = i[48634];
  assign o[48633] = i[48633];
  assign o[48632] = i[48632];
  assign o[48631] = i[48631];
  assign o[48630] = i[48630];
  assign o[48629] = i[48629];
  assign o[48628] = i[48628];
  assign o[48627] = i[48627];
  assign o[48626] = i[48626];
  assign o[48625] = i[48625];
  assign o[48624] = i[48624];
  assign o[48623] = i[48623];
  assign o[48622] = i[48622];
  assign o[48621] = i[48621];
  assign o[48620] = i[48620];
  assign o[48619] = i[48619];
  assign o[48618] = i[48618];
  assign o[48617] = i[48617];
  assign o[48616] = i[48616];
  assign o[48615] = i[48615];
  assign o[48614] = i[48614];
  assign o[48613] = i[48613];
  assign o[48612] = i[48612];
  assign o[48611] = i[48611];
  assign o[48610] = i[48610];
  assign o[48609] = i[48609];
  assign o[48608] = i[48608];
  assign o[48607] = i[48607];
  assign o[48606] = i[48606];
  assign o[48605] = i[48605];
  assign o[48604] = i[48604];
  assign o[48603] = i[48603];
  assign o[48602] = i[48602];
  assign o[48601] = i[48601];
  assign o[48600] = i[48600];
  assign o[48599] = i[48599];
  assign o[48598] = i[48598];
  assign o[48597] = i[48597];
  assign o[48596] = i[48596];
  assign o[48595] = i[48595];
  assign o[48594] = i[48594];
  assign o[48593] = i[48593];
  assign o[48592] = i[48592];
  assign o[48591] = i[48591];
  assign o[48590] = i[48590];
  assign o[48589] = i[48589];
  assign o[48588] = i[48588];
  assign o[48587] = i[48587];
  assign o[48586] = i[48586];
  assign o[48585] = i[48585];
  assign o[48584] = i[48584];
  assign o[48583] = i[48583];
  assign o[48582] = i[48582];
  assign o[48581] = i[48581];
  assign o[48580] = i[48580];
  assign o[48579] = i[48579];
  assign o[48578] = i[48578];
  assign o[48577] = i[48577];
  assign o[48576] = i[48576];
  assign o[48575] = i[48575];
  assign o[48574] = i[48574];
  assign o[48573] = i[48573];
  assign o[48572] = i[48572];
  assign o[48571] = i[48571];
  assign o[48570] = i[48570];
  assign o[48569] = i[48569];
  assign o[48568] = i[48568];
  assign o[48567] = i[48567];
  assign o[48566] = i[48566];
  assign o[48565] = i[48565];
  assign o[48564] = i[48564];
  assign o[48563] = i[48563];
  assign o[48562] = i[48562];
  assign o[48561] = i[48561];
  assign o[48560] = i[48560];
  assign o[48559] = i[48559];
  assign o[48558] = i[48558];
  assign o[48557] = i[48557];
  assign o[48556] = i[48556];
  assign o[48555] = i[48555];
  assign o[48554] = i[48554];
  assign o[48553] = i[48553];
  assign o[48552] = i[48552];
  assign o[48551] = i[48551];
  assign o[48550] = i[48550];
  assign o[48549] = i[48549];
  assign o[48548] = i[48548];
  assign o[48547] = i[48547];
  assign o[48546] = i[48546];
  assign o[48545] = i[48545];
  assign o[48544] = i[48544];
  assign o[48543] = i[48543];
  assign o[48542] = i[48542];
  assign o[48541] = i[48541];
  assign o[48540] = i[48540];
  assign o[48539] = i[48539];
  assign o[48538] = i[48538];
  assign o[48537] = i[48537];
  assign o[48536] = i[48536];
  assign o[48535] = i[48535];
  assign o[48534] = i[48534];
  assign o[48533] = i[48533];
  assign o[48532] = i[48532];
  assign o[48531] = i[48531];
  assign o[48530] = i[48530];
  assign o[48529] = i[48529];
  assign o[48528] = i[48528];
  assign o[48527] = i[48527];
  assign o[48526] = i[48526];
  assign o[48525] = i[48525];
  assign o[48524] = i[48524];
  assign o[48523] = i[48523];
  assign o[48522] = i[48522];
  assign o[48521] = i[48521];
  assign o[48520] = i[48520];
  assign o[48519] = i[48519];
  assign o[48518] = i[48518];
  assign o[48517] = i[48517];
  assign o[48516] = i[48516];
  assign o[48515] = i[48515];
  assign o[48514] = i[48514];
  assign o[48513] = i[48513];
  assign o[48512] = i[48512];
  assign o[48511] = i[48511];
  assign o[48510] = i[48510];
  assign o[48509] = i[48509];
  assign o[48508] = i[48508];
  assign o[48507] = i[48507];
  assign o[48506] = i[48506];
  assign o[48505] = i[48505];
  assign o[48504] = i[48504];
  assign o[48503] = i[48503];
  assign o[48502] = i[48502];
  assign o[48501] = i[48501];
  assign o[48500] = i[48500];
  assign o[48499] = i[48499];
  assign o[48498] = i[48498];
  assign o[48497] = i[48497];
  assign o[48496] = i[48496];
  assign o[48495] = i[48495];
  assign o[48494] = i[48494];
  assign o[48493] = i[48493];
  assign o[48492] = i[48492];
  assign o[48491] = i[48491];
  assign o[48490] = i[48490];
  assign o[48489] = i[48489];
  assign o[48488] = i[48488];
  assign o[48487] = i[48487];
  assign o[48486] = i[48486];
  assign o[48485] = i[48485];
  assign o[48484] = i[48484];
  assign o[48483] = i[48483];
  assign o[48482] = i[48482];
  assign o[48481] = i[48481];
  assign o[48480] = i[48480];
  assign o[48479] = i[48479];
  assign o[48478] = i[48478];
  assign o[48477] = i[48477];
  assign o[48476] = i[48476];
  assign o[48475] = i[48475];
  assign o[48474] = i[48474];
  assign o[48473] = i[48473];
  assign o[48472] = i[48472];
  assign o[48471] = i[48471];
  assign o[48470] = i[48470];
  assign o[48469] = i[48469];
  assign o[48468] = i[48468];
  assign o[48467] = i[48467];
  assign o[48466] = i[48466];
  assign o[48465] = i[48465];
  assign o[48464] = i[48464];
  assign o[48463] = i[48463];
  assign o[48462] = i[48462];
  assign o[48461] = i[48461];
  assign o[48460] = i[48460];
  assign o[48459] = i[48459];
  assign o[48458] = i[48458];
  assign o[48457] = i[48457];
  assign o[48456] = i[48456];
  assign o[48455] = i[48455];
  assign o[48454] = i[48454];
  assign o[48453] = i[48453];
  assign o[48452] = i[48452];
  assign o[48451] = i[48451];
  assign o[48450] = i[48450];
  assign o[48449] = i[48449];
  assign o[48448] = i[48448];
  assign o[48447] = i[48447];
  assign o[48446] = i[48446];
  assign o[48445] = i[48445];
  assign o[48444] = i[48444];
  assign o[48443] = i[48443];
  assign o[48442] = i[48442];
  assign o[48441] = i[48441];
  assign o[48440] = i[48440];
  assign o[48439] = i[48439];
  assign o[48438] = i[48438];
  assign o[48437] = i[48437];
  assign o[48436] = i[48436];
  assign o[48435] = i[48435];
  assign o[48434] = i[48434];
  assign o[48433] = i[48433];
  assign o[48432] = i[48432];
  assign o[48431] = i[48431];
  assign o[48430] = i[48430];
  assign o[48429] = i[48429];
  assign o[48428] = i[48428];
  assign o[48427] = i[48427];
  assign o[48426] = i[48426];
  assign o[48425] = i[48425];
  assign o[48424] = i[48424];
  assign o[48423] = i[48423];
  assign o[48422] = i[48422];
  assign o[48421] = i[48421];
  assign o[48420] = i[48420];
  assign o[48419] = i[48419];
  assign o[48418] = i[48418];
  assign o[48417] = i[48417];
  assign o[48416] = i[48416];
  assign o[48415] = i[48415];
  assign o[48414] = i[48414];
  assign o[48413] = i[48413];
  assign o[48412] = i[48412];
  assign o[48411] = i[48411];
  assign o[48410] = i[48410];
  assign o[48409] = i[48409];
  assign o[48408] = i[48408];
  assign o[48407] = i[48407];
  assign o[48406] = i[48406];
  assign o[48405] = i[48405];
  assign o[48404] = i[48404];
  assign o[48403] = i[48403];
  assign o[48402] = i[48402];
  assign o[48401] = i[48401];
  assign o[48400] = i[48400];
  assign o[48399] = i[48399];
  assign o[48398] = i[48398];
  assign o[48397] = i[48397];
  assign o[48396] = i[48396];
  assign o[48395] = i[48395];
  assign o[48394] = i[48394];
  assign o[48393] = i[48393];
  assign o[48392] = i[48392];
  assign o[48391] = i[48391];
  assign o[48390] = i[48390];
  assign o[48389] = i[48389];
  assign o[48388] = i[48388];
  assign o[48387] = i[48387];
  assign o[48386] = i[48386];
  assign o[48385] = i[48385];
  assign o[48384] = i[48384];
  assign o[48383] = i[48383];
  assign o[48382] = i[48382];
  assign o[48381] = i[48381];
  assign o[48380] = i[48380];
  assign o[48379] = i[48379];
  assign o[48378] = i[48378];
  assign o[48377] = i[48377];
  assign o[48376] = i[48376];
  assign o[48375] = i[48375];
  assign o[48374] = i[48374];
  assign o[48373] = i[48373];
  assign o[48372] = i[48372];
  assign o[48371] = i[48371];
  assign o[48370] = i[48370];
  assign o[48369] = i[48369];
  assign o[48368] = i[48368];
  assign o[48367] = i[48367];
  assign o[48366] = i[48366];
  assign o[48365] = i[48365];
  assign o[48364] = i[48364];
  assign o[48363] = i[48363];
  assign o[48362] = i[48362];
  assign o[48361] = i[48361];
  assign o[48360] = i[48360];
  assign o[48359] = i[48359];
  assign o[48358] = i[48358];
  assign o[48357] = i[48357];
  assign o[48356] = i[48356];
  assign o[48355] = i[48355];
  assign o[48354] = i[48354];
  assign o[48353] = i[48353];
  assign o[48352] = i[48352];
  assign o[48351] = i[48351];
  assign o[48350] = i[48350];
  assign o[48349] = i[48349];
  assign o[48348] = i[48348];
  assign o[48347] = i[48347];
  assign o[48346] = i[48346];
  assign o[48345] = i[48345];
  assign o[48344] = i[48344];
  assign o[48343] = i[48343];
  assign o[48342] = i[48342];
  assign o[48341] = i[48341];
  assign o[48340] = i[48340];
  assign o[48339] = i[48339];
  assign o[48338] = i[48338];
  assign o[48337] = i[48337];
  assign o[48336] = i[48336];
  assign o[48335] = i[48335];
  assign o[48334] = i[48334];
  assign o[48333] = i[48333];
  assign o[48332] = i[48332];
  assign o[48331] = i[48331];
  assign o[48330] = i[48330];
  assign o[48329] = i[48329];
  assign o[48328] = i[48328];
  assign o[48327] = i[48327];
  assign o[48326] = i[48326];
  assign o[48325] = i[48325];
  assign o[48324] = i[48324];
  assign o[48323] = i[48323];
  assign o[48322] = i[48322];
  assign o[48321] = i[48321];
  assign o[48320] = i[48320];
  assign o[48319] = i[48319];
  assign o[48318] = i[48318];
  assign o[48317] = i[48317];
  assign o[48316] = i[48316];
  assign o[48315] = i[48315];
  assign o[48314] = i[48314];
  assign o[48313] = i[48313];
  assign o[48312] = i[48312];
  assign o[48311] = i[48311];
  assign o[48310] = i[48310];
  assign o[48309] = i[48309];
  assign o[48308] = i[48308];
  assign o[48307] = i[48307];
  assign o[48306] = i[48306];
  assign o[48305] = i[48305];
  assign o[48304] = i[48304];
  assign o[48303] = i[48303];
  assign o[48302] = i[48302];
  assign o[48301] = i[48301];
  assign o[48300] = i[48300];
  assign o[48299] = i[48299];
  assign o[48298] = i[48298];
  assign o[48297] = i[48297];
  assign o[48296] = i[48296];
  assign o[48295] = i[48295];
  assign o[48294] = i[48294];
  assign o[48293] = i[48293];
  assign o[48292] = i[48292];
  assign o[48291] = i[48291];
  assign o[48290] = i[48290];
  assign o[48289] = i[48289];
  assign o[48288] = i[48288];
  assign o[48287] = i[48287];
  assign o[48286] = i[48286];
  assign o[48285] = i[48285];
  assign o[48284] = i[48284];
  assign o[48283] = i[48283];
  assign o[48282] = i[48282];
  assign o[48281] = i[48281];
  assign o[48280] = i[48280];
  assign o[48279] = i[48279];
  assign o[48278] = i[48278];
  assign o[48277] = i[48277];
  assign o[48276] = i[48276];
  assign o[48275] = i[48275];
  assign o[48274] = i[48274];
  assign o[48273] = i[48273];
  assign o[48272] = i[48272];
  assign o[48271] = i[48271];
  assign o[48270] = i[48270];
  assign o[48269] = i[48269];
  assign o[48268] = i[48268];
  assign o[48267] = i[48267];
  assign o[48266] = i[48266];
  assign o[48265] = i[48265];
  assign o[48264] = i[48264];
  assign o[48263] = i[48263];
  assign o[48262] = i[48262];
  assign o[48261] = i[48261];
  assign o[48260] = i[48260];
  assign o[48259] = i[48259];
  assign o[48258] = i[48258];
  assign o[48257] = i[48257];
  assign o[48256] = i[48256];
  assign o[48255] = i[48255];
  assign o[48254] = i[48254];
  assign o[48253] = i[48253];
  assign o[48252] = i[48252];
  assign o[48251] = i[48251];
  assign o[48250] = i[48250];
  assign o[48249] = i[48249];
  assign o[48248] = i[48248];
  assign o[48247] = i[48247];
  assign o[48246] = i[48246];
  assign o[48245] = i[48245];
  assign o[48244] = i[48244];
  assign o[48243] = i[48243];
  assign o[48242] = i[48242];
  assign o[48241] = i[48241];
  assign o[48240] = i[48240];
  assign o[48239] = i[48239];
  assign o[48238] = i[48238];
  assign o[48237] = i[48237];
  assign o[48236] = i[48236];
  assign o[48235] = i[48235];
  assign o[48234] = i[48234];
  assign o[48233] = i[48233];
  assign o[48232] = i[48232];
  assign o[48231] = i[48231];
  assign o[48230] = i[48230];
  assign o[48229] = i[48229];
  assign o[48228] = i[48228];
  assign o[48227] = i[48227];
  assign o[48226] = i[48226];
  assign o[48225] = i[48225];
  assign o[48224] = i[48224];
  assign o[48223] = i[48223];
  assign o[48222] = i[48222];
  assign o[48221] = i[48221];
  assign o[48220] = i[48220];
  assign o[48219] = i[48219];
  assign o[48218] = i[48218];
  assign o[48217] = i[48217];
  assign o[48216] = i[48216];
  assign o[48215] = i[48215];
  assign o[48214] = i[48214];
  assign o[48213] = i[48213];
  assign o[48212] = i[48212];
  assign o[48211] = i[48211];
  assign o[48210] = i[48210];
  assign o[48209] = i[48209];
  assign o[48208] = i[48208];
  assign o[48207] = i[48207];
  assign o[48206] = i[48206];
  assign o[48205] = i[48205];
  assign o[48204] = i[48204];
  assign o[48203] = i[48203];
  assign o[48202] = i[48202];
  assign o[48201] = i[48201];
  assign o[48200] = i[48200];
  assign o[48199] = i[48199];
  assign o[48198] = i[48198];
  assign o[48197] = i[48197];
  assign o[48196] = i[48196];
  assign o[48195] = i[48195];
  assign o[48194] = i[48194];
  assign o[48193] = i[48193];
  assign o[48192] = i[48192];
  assign o[48191] = i[48191];
  assign o[48190] = i[48190];
  assign o[48189] = i[48189];
  assign o[48188] = i[48188];
  assign o[48187] = i[48187];
  assign o[48186] = i[48186];
  assign o[48185] = i[48185];
  assign o[48184] = i[48184];
  assign o[48183] = i[48183];
  assign o[48182] = i[48182];
  assign o[48181] = i[48181];
  assign o[48180] = i[48180];
  assign o[48179] = i[48179];
  assign o[48178] = i[48178];
  assign o[48177] = i[48177];
  assign o[48176] = i[48176];
  assign o[48175] = i[48175];
  assign o[48174] = i[48174];
  assign o[48173] = i[48173];
  assign o[48172] = i[48172];
  assign o[48171] = i[48171];
  assign o[48170] = i[48170];
  assign o[48169] = i[48169];
  assign o[48168] = i[48168];
  assign o[48167] = i[48167];
  assign o[48166] = i[48166];
  assign o[48165] = i[48165];
  assign o[48164] = i[48164];
  assign o[48163] = i[48163];
  assign o[48162] = i[48162];
  assign o[48161] = i[48161];
  assign o[48160] = i[48160];
  assign o[48159] = i[48159];
  assign o[48158] = i[48158];
  assign o[48157] = i[48157];
  assign o[48156] = i[48156];
  assign o[48155] = i[48155];
  assign o[48154] = i[48154];
  assign o[48153] = i[48153];
  assign o[48152] = i[48152];
  assign o[48151] = i[48151];
  assign o[48150] = i[48150];
  assign o[48149] = i[48149];
  assign o[48148] = i[48148];
  assign o[48147] = i[48147];
  assign o[48146] = i[48146];
  assign o[48145] = i[48145];
  assign o[48144] = i[48144];
  assign o[48143] = i[48143];
  assign o[48142] = i[48142];
  assign o[48141] = i[48141];
  assign o[48140] = i[48140];
  assign o[48139] = i[48139];
  assign o[48138] = i[48138];
  assign o[48137] = i[48137];
  assign o[48136] = i[48136];
  assign o[48135] = i[48135];
  assign o[48134] = i[48134];
  assign o[48133] = i[48133];
  assign o[48132] = i[48132];
  assign o[48131] = i[48131];
  assign o[48130] = i[48130];
  assign o[48129] = i[48129];
  assign o[48128] = i[48128];
  assign o[48127] = i[48127];
  assign o[48126] = i[48126];
  assign o[48125] = i[48125];
  assign o[48124] = i[48124];
  assign o[48123] = i[48123];
  assign o[48122] = i[48122];
  assign o[48121] = i[48121];
  assign o[48120] = i[48120];
  assign o[48119] = i[48119];
  assign o[48118] = i[48118];
  assign o[48117] = i[48117];
  assign o[48116] = i[48116];
  assign o[48115] = i[48115];
  assign o[48114] = i[48114];
  assign o[48113] = i[48113];
  assign o[48112] = i[48112];
  assign o[48111] = i[48111];
  assign o[48110] = i[48110];
  assign o[48109] = i[48109];
  assign o[48108] = i[48108];
  assign o[48107] = i[48107];
  assign o[48106] = i[48106];
  assign o[48105] = i[48105];
  assign o[48104] = i[48104];
  assign o[48103] = i[48103];
  assign o[48102] = i[48102];
  assign o[48101] = i[48101];
  assign o[48100] = i[48100];
  assign o[48099] = i[48099];
  assign o[48098] = i[48098];
  assign o[48097] = i[48097];
  assign o[48096] = i[48096];
  assign o[48095] = i[48095];
  assign o[48094] = i[48094];
  assign o[48093] = i[48093];
  assign o[48092] = i[48092];
  assign o[48091] = i[48091];
  assign o[48090] = i[48090];
  assign o[48089] = i[48089];
  assign o[48088] = i[48088];
  assign o[48087] = i[48087];
  assign o[48086] = i[48086];
  assign o[48085] = i[48085];
  assign o[48084] = i[48084];
  assign o[48083] = i[48083];
  assign o[48082] = i[48082];
  assign o[48081] = i[48081];
  assign o[48080] = i[48080];
  assign o[48079] = i[48079];
  assign o[48078] = i[48078];
  assign o[48077] = i[48077];
  assign o[48076] = i[48076];
  assign o[48075] = i[48075];
  assign o[48074] = i[48074];
  assign o[48073] = i[48073];
  assign o[48072] = i[48072];
  assign o[48071] = i[48071];
  assign o[48070] = i[48070];
  assign o[48069] = i[48069];
  assign o[48068] = i[48068];
  assign o[48067] = i[48067];
  assign o[48066] = i[48066];
  assign o[48065] = i[48065];
  assign o[48064] = i[48064];
  assign o[48063] = i[48063];
  assign o[48062] = i[48062];
  assign o[48061] = i[48061];
  assign o[48060] = i[48060];
  assign o[48059] = i[48059];
  assign o[48058] = i[48058];
  assign o[48057] = i[48057];
  assign o[48056] = i[48056];
  assign o[48055] = i[48055];
  assign o[48054] = i[48054];
  assign o[48053] = i[48053];
  assign o[48052] = i[48052];
  assign o[48051] = i[48051];
  assign o[48050] = i[48050];
  assign o[48049] = i[48049];
  assign o[48048] = i[48048];
  assign o[48047] = i[48047];
  assign o[48046] = i[48046];
  assign o[48045] = i[48045];
  assign o[48044] = i[48044];
  assign o[48043] = i[48043];
  assign o[48042] = i[48042];
  assign o[48041] = i[48041];
  assign o[48040] = i[48040];
  assign o[48039] = i[48039];
  assign o[48038] = i[48038];
  assign o[48037] = i[48037];
  assign o[48036] = i[48036];
  assign o[48035] = i[48035];
  assign o[48034] = i[48034];
  assign o[48033] = i[48033];
  assign o[48032] = i[48032];
  assign o[48031] = i[48031];
  assign o[48030] = i[48030];
  assign o[48029] = i[48029];
  assign o[48028] = i[48028];
  assign o[48027] = i[48027];
  assign o[48026] = i[48026];
  assign o[48025] = i[48025];
  assign o[48024] = i[48024];
  assign o[48023] = i[48023];
  assign o[48022] = i[48022];
  assign o[48021] = i[48021];
  assign o[48020] = i[48020];
  assign o[48019] = i[48019];
  assign o[48018] = i[48018];
  assign o[48017] = i[48017];
  assign o[48016] = i[48016];
  assign o[48015] = i[48015];
  assign o[48014] = i[48014];
  assign o[48013] = i[48013];
  assign o[48012] = i[48012];
  assign o[48011] = i[48011];
  assign o[48010] = i[48010];
  assign o[48009] = i[48009];
  assign o[48008] = i[48008];
  assign o[48007] = i[48007];
  assign o[48006] = i[48006];
  assign o[48005] = i[48005];
  assign o[48004] = i[48004];
  assign o[48003] = i[48003];
  assign o[48002] = i[48002];
  assign o[48001] = i[48001];
  assign o[48000] = i[48000];
  assign o[47999] = i[47999];
  assign o[47998] = i[47998];
  assign o[47997] = i[47997];
  assign o[47996] = i[47996];
  assign o[47995] = i[47995];
  assign o[47994] = i[47994];
  assign o[47993] = i[47993];
  assign o[47992] = i[47992];
  assign o[47991] = i[47991];
  assign o[47990] = i[47990];
  assign o[47989] = i[47989];
  assign o[47988] = i[47988];
  assign o[47987] = i[47987];
  assign o[47986] = i[47986];
  assign o[47985] = i[47985];
  assign o[47984] = i[47984];
  assign o[47983] = i[47983];
  assign o[47982] = i[47982];
  assign o[47981] = i[47981];
  assign o[47980] = i[47980];
  assign o[47979] = i[47979];
  assign o[47978] = i[47978];
  assign o[47977] = i[47977];
  assign o[47976] = i[47976];
  assign o[47975] = i[47975];
  assign o[47974] = i[47974];
  assign o[47973] = i[47973];
  assign o[47972] = i[47972];
  assign o[47971] = i[47971];
  assign o[47970] = i[47970];
  assign o[47969] = i[47969];
  assign o[47968] = i[47968];
  assign o[47967] = i[47967];
  assign o[47966] = i[47966];
  assign o[47965] = i[47965];
  assign o[47964] = i[47964];
  assign o[47963] = i[47963];
  assign o[47962] = i[47962];
  assign o[47961] = i[47961];
  assign o[47960] = i[47960];
  assign o[47959] = i[47959];
  assign o[47958] = i[47958];
  assign o[47957] = i[47957];
  assign o[47956] = i[47956];
  assign o[47955] = i[47955];
  assign o[47954] = i[47954];
  assign o[47953] = i[47953];
  assign o[47952] = i[47952];
  assign o[47951] = i[47951];
  assign o[47950] = i[47950];
  assign o[47949] = i[47949];
  assign o[47948] = i[47948];
  assign o[47947] = i[47947];
  assign o[47946] = i[47946];
  assign o[47945] = i[47945];
  assign o[47944] = i[47944];
  assign o[47943] = i[47943];
  assign o[47942] = i[47942];
  assign o[47941] = i[47941];
  assign o[47940] = i[47940];
  assign o[47939] = i[47939];
  assign o[47938] = i[47938];
  assign o[47937] = i[47937];
  assign o[47936] = i[47936];
  assign o[47935] = i[47935];
  assign o[47934] = i[47934];
  assign o[47933] = i[47933];
  assign o[47932] = i[47932];
  assign o[47931] = i[47931];
  assign o[47930] = i[47930];
  assign o[47929] = i[47929];
  assign o[47928] = i[47928];
  assign o[47927] = i[47927];
  assign o[47926] = i[47926];
  assign o[47925] = i[47925];
  assign o[47924] = i[47924];
  assign o[47923] = i[47923];
  assign o[47922] = i[47922];
  assign o[47921] = i[47921];
  assign o[47920] = i[47920];
  assign o[47919] = i[47919];
  assign o[47918] = i[47918];
  assign o[47917] = i[47917];
  assign o[47916] = i[47916];
  assign o[47915] = i[47915];
  assign o[47914] = i[47914];
  assign o[47913] = i[47913];
  assign o[47912] = i[47912];
  assign o[47911] = i[47911];
  assign o[47910] = i[47910];
  assign o[47909] = i[47909];
  assign o[47908] = i[47908];
  assign o[47907] = i[47907];
  assign o[47906] = i[47906];
  assign o[47905] = i[47905];
  assign o[47904] = i[47904];
  assign o[47903] = i[47903];
  assign o[47902] = i[47902];
  assign o[47901] = i[47901];
  assign o[47900] = i[47900];
  assign o[47899] = i[47899];
  assign o[47898] = i[47898];
  assign o[47897] = i[47897];
  assign o[47896] = i[47896];
  assign o[47895] = i[47895];
  assign o[47894] = i[47894];
  assign o[47893] = i[47893];
  assign o[47892] = i[47892];
  assign o[47891] = i[47891];
  assign o[47890] = i[47890];
  assign o[47889] = i[47889];
  assign o[47888] = i[47888];
  assign o[47887] = i[47887];
  assign o[47886] = i[47886];
  assign o[47885] = i[47885];
  assign o[47884] = i[47884];
  assign o[47883] = i[47883];
  assign o[47882] = i[47882];
  assign o[47881] = i[47881];
  assign o[47880] = i[47880];
  assign o[47879] = i[47879];
  assign o[47878] = i[47878];
  assign o[47877] = i[47877];
  assign o[47876] = i[47876];
  assign o[47875] = i[47875];
  assign o[47874] = i[47874];
  assign o[47873] = i[47873];
  assign o[47872] = i[47872];
  assign o[47871] = i[47871];
  assign o[47870] = i[47870];
  assign o[47869] = i[47869];
  assign o[47868] = i[47868];
  assign o[47867] = i[47867];
  assign o[47866] = i[47866];
  assign o[47865] = i[47865];
  assign o[47864] = i[47864];
  assign o[47863] = i[47863];
  assign o[47862] = i[47862];
  assign o[47861] = i[47861];
  assign o[47860] = i[47860];
  assign o[47859] = i[47859];
  assign o[47858] = i[47858];
  assign o[47857] = i[47857];
  assign o[47856] = i[47856];
  assign o[47855] = i[47855];
  assign o[47854] = i[47854];
  assign o[47853] = i[47853];
  assign o[47852] = i[47852];
  assign o[47851] = i[47851];
  assign o[47850] = i[47850];
  assign o[47849] = i[47849];
  assign o[47848] = i[47848];
  assign o[47847] = i[47847];
  assign o[47846] = i[47846];
  assign o[47845] = i[47845];
  assign o[47844] = i[47844];
  assign o[47843] = i[47843];
  assign o[47842] = i[47842];
  assign o[47841] = i[47841];
  assign o[47840] = i[47840];
  assign o[47839] = i[47839];
  assign o[47838] = i[47838];
  assign o[47837] = i[47837];
  assign o[47836] = i[47836];
  assign o[47835] = i[47835];
  assign o[47834] = i[47834];
  assign o[47833] = i[47833];
  assign o[47832] = i[47832];
  assign o[47831] = i[47831];
  assign o[47830] = i[47830];
  assign o[47829] = i[47829];
  assign o[47828] = i[47828];
  assign o[47827] = i[47827];
  assign o[47826] = i[47826];
  assign o[47825] = i[47825];
  assign o[47824] = i[47824];
  assign o[47823] = i[47823];
  assign o[47822] = i[47822];
  assign o[47821] = i[47821];
  assign o[47820] = i[47820];
  assign o[47819] = i[47819];
  assign o[47818] = i[47818];
  assign o[47817] = i[47817];
  assign o[47816] = i[47816];
  assign o[47815] = i[47815];
  assign o[47814] = i[47814];
  assign o[47813] = i[47813];
  assign o[47812] = i[47812];
  assign o[47811] = i[47811];
  assign o[47810] = i[47810];
  assign o[47809] = i[47809];
  assign o[47808] = i[47808];
  assign o[47807] = i[47807];
  assign o[47806] = i[47806];
  assign o[47805] = i[47805];
  assign o[47804] = i[47804];
  assign o[47803] = i[47803];
  assign o[47802] = i[47802];
  assign o[47801] = i[47801];
  assign o[47800] = i[47800];
  assign o[47799] = i[47799];
  assign o[47798] = i[47798];
  assign o[47797] = i[47797];
  assign o[47796] = i[47796];
  assign o[47795] = i[47795];
  assign o[47794] = i[47794];
  assign o[47793] = i[47793];
  assign o[47792] = i[47792];
  assign o[47791] = i[47791];
  assign o[47790] = i[47790];
  assign o[47789] = i[47789];
  assign o[47788] = i[47788];
  assign o[47787] = i[47787];
  assign o[47786] = i[47786];
  assign o[47785] = i[47785];
  assign o[47784] = i[47784];
  assign o[47783] = i[47783];
  assign o[47782] = i[47782];
  assign o[47781] = i[47781];
  assign o[47780] = i[47780];
  assign o[47779] = i[47779];
  assign o[47778] = i[47778];
  assign o[47777] = i[47777];
  assign o[47776] = i[47776];
  assign o[47775] = i[47775];
  assign o[47774] = i[47774];
  assign o[47773] = i[47773];
  assign o[47772] = i[47772];
  assign o[47771] = i[47771];
  assign o[47770] = i[47770];
  assign o[47769] = i[47769];
  assign o[47768] = i[47768];
  assign o[47767] = i[47767];
  assign o[47766] = i[47766];
  assign o[47765] = i[47765];
  assign o[47764] = i[47764];
  assign o[47763] = i[47763];
  assign o[47762] = i[47762];
  assign o[47761] = i[47761];
  assign o[47760] = i[47760];
  assign o[47759] = i[47759];
  assign o[47758] = i[47758];
  assign o[47757] = i[47757];
  assign o[47756] = i[47756];
  assign o[47755] = i[47755];
  assign o[47754] = i[47754];
  assign o[47753] = i[47753];
  assign o[47752] = i[47752];
  assign o[47751] = i[47751];
  assign o[47750] = i[47750];
  assign o[47749] = i[47749];
  assign o[47748] = i[47748];
  assign o[47747] = i[47747];
  assign o[47746] = i[47746];
  assign o[47745] = i[47745];
  assign o[47744] = i[47744];
  assign o[47743] = i[47743];
  assign o[47742] = i[47742];
  assign o[47741] = i[47741];
  assign o[47740] = i[47740];
  assign o[47739] = i[47739];
  assign o[47738] = i[47738];
  assign o[47737] = i[47737];
  assign o[47736] = i[47736];
  assign o[47735] = i[47735];
  assign o[47734] = i[47734];
  assign o[47733] = i[47733];
  assign o[47732] = i[47732];
  assign o[47731] = i[47731];
  assign o[47730] = i[47730];
  assign o[47729] = i[47729];
  assign o[47728] = i[47728];
  assign o[47727] = i[47727];
  assign o[47726] = i[47726];
  assign o[47725] = i[47725];
  assign o[47724] = i[47724];
  assign o[47723] = i[47723];
  assign o[47722] = i[47722];
  assign o[47721] = i[47721];
  assign o[47720] = i[47720];
  assign o[47719] = i[47719];
  assign o[47718] = i[47718];
  assign o[47717] = i[47717];
  assign o[47716] = i[47716];
  assign o[47715] = i[47715];
  assign o[47714] = i[47714];
  assign o[47713] = i[47713];
  assign o[47712] = i[47712];
  assign o[47711] = i[47711];
  assign o[47710] = i[47710];
  assign o[47709] = i[47709];
  assign o[47708] = i[47708];
  assign o[47707] = i[47707];
  assign o[47706] = i[47706];
  assign o[47705] = i[47705];
  assign o[47704] = i[47704];
  assign o[47703] = i[47703];
  assign o[47702] = i[47702];
  assign o[47701] = i[47701];
  assign o[47700] = i[47700];
  assign o[47699] = i[47699];
  assign o[47698] = i[47698];
  assign o[47697] = i[47697];
  assign o[47696] = i[47696];
  assign o[47695] = i[47695];
  assign o[47694] = i[47694];
  assign o[47693] = i[47693];
  assign o[47692] = i[47692];
  assign o[47691] = i[47691];
  assign o[47690] = i[47690];
  assign o[47689] = i[47689];
  assign o[47688] = i[47688];
  assign o[47687] = i[47687];
  assign o[47686] = i[47686];
  assign o[47685] = i[47685];
  assign o[47684] = i[47684];
  assign o[47683] = i[47683];
  assign o[47682] = i[47682];
  assign o[47681] = i[47681];
  assign o[47680] = i[47680];
  assign o[47679] = i[47679];
  assign o[47678] = i[47678];
  assign o[47677] = i[47677];
  assign o[47676] = i[47676];
  assign o[47675] = i[47675];
  assign o[47674] = i[47674];
  assign o[47673] = i[47673];
  assign o[47672] = i[47672];
  assign o[47671] = i[47671];
  assign o[47670] = i[47670];
  assign o[47669] = i[47669];
  assign o[47668] = i[47668];
  assign o[47667] = i[47667];
  assign o[47666] = i[47666];
  assign o[47665] = i[47665];
  assign o[47664] = i[47664];
  assign o[47663] = i[47663];
  assign o[47662] = i[47662];
  assign o[47661] = i[47661];
  assign o[47660] = i[47660];
  assign o[47659] = i[47659];
  assign o[47658] = i[47658];
  assign o[47657] = i[47657];
  assign o[47656] = i[47656];
  assign o[47655] = i[47655];
  assign o[47654] = i[47654];
  assign o[47653] = i[47653];
  assign o[47652] = i[47652];
  assign o[47651] = i[47651];
  assign o[47650] = i[47650];
  assign o[47649] = i[47649];
  assign o[47648] = i[47648];
  assign o[47647] = i[47647];
  assign o[47646] = i[47646];
  assign o[47645] = i[47645];
  assign o[47644] = i[47644];
  assign o[47643] = i[47643];
  assign o[47642] = i[47642];
  assign o[47641] = i[47641];
  assign o[47640] = i[47640];
  assign o[47639] = i[47639];
  assign o[47638] = i[47638];
  assign o[47637] = i[47637];
  assign o[47636] = i[47636];
  assign o[47635] = i[47635];
  assign o[47634] = i[47634];
  assign o[47633] = i[47633];
  assign o[47632] = i[47632];
  assign o[47631] = i[47631];
  assign o[47630] = i[47630];
  assign o[47629] = i[47629];
  assign o[47628] = i[47628];
  assign o[47627] = i[47627];
  assign o[47626] = i[47626];
  assign o[47625] = i[47625];
  assign o[47624] = i[47624];
  assign o[47623] = i[47623];
  assign o[47622] = i[47622];
  assign o[47621] = i[47621];
  assign o[47620] = i[47620];
  assign o[47619] = i[47619];
  assign o[47618] = i[47618];
  assign o[47617] = i[47617];
  assign o[47616] = i[47616];
  assign o[47615] = i[47615];
  assign o[47614] = i[47614];
  assign o[47613] = i[47613];
  assign o[47612] = i[47612];
  assign o[47611] = i[47611];
  assign o[47610] = i[47610];
  assign o[47609] = i[47609];
  assign o[47608] = i[47608];
  assign o[47607] = i[47607];
  assign o[47606] = i[47606];
  assign o[47605] = i[47605];
  assign o[47604] = i[47604];
  assign o[47603] = i[47603];
  assign o[47602] = i[47602];
  assign o[47601] = i[47601];
  assign o[47600] = i[47600];
  assign o[47599] = i[47599];
  assign o[47598] = i[47598];
  assign o[47597] = i[47597];
  assign o[47596] = i[47596];
  assign o[47595] = i[47595];
  assign o[47594] = i[47594];
  assign o[47593] = i[47593];
  assign o[47592] = i[47592];
  assign o[47591] = i[47591];
  assign o[47590] = i[47590];
  assign o[47589] = i[47589];
  assign o[47588] = i[47588];
  assign o[47587] = i[47587];
  assign o[47586] = i[47586];
  assign o[47585] = i[47585];
  assign o[47584] = i[47584];
  assign o[47583] = i[47583];
  assign o[47582] = i[47582];
  assign o[47581] = i[47581];
  assign o[47580] = i[47580];
  assign o[47579] = i[47579];
  assign o[47578] = i[47578];
  assign o[47577] = i[47577];
  assign o[47576] = i[47576];
  assign o[47575] = i[47575];
  assign o[47574] = i[47574];
  assign o[47573] = i[47573];
  assign o[47572] = i[47572];
  assign o[47571] = i[47571];
  assign o[47570] = i[47570];
  assign o[47569] = i[47569];
  assign o[47568] = i[47568];
  assign o[47567] = i[47567];
  assign o[47566] = i[47566];
  assign o[47565] = i[47565];
  assign o[47564] = i[47564];
  assign o[47563] = i[47563];
  assign o[47562] = i[47562];
  assign o[47561] = i[47561];
  assign o[47560] = i[47560];
  assign o[47559] = i[47559];
  assign o[47558] = i[47558];
  assign o[47557] = i[47557];
  assign o[47556] = i[47556];
  assign o[47555] = i[47555];
  assign o[47554] = i[47554];
  assign o[47553] = i[47553];
  assign o[47552] = i[47552];
  assign o[47551] = i[47551];
  assign o[47550] = i[47550];
  assign o[47549] = i[47549];
  assign o[47548] = i[47548];
  assign o[47547] = i[47547];
  assign o[47546] = i[47546];
  assign o[47545] = i[47545];
  assign o[47544] = i[47544];
  assign o[47543] = i[47543];
  assign o[47542] = i[47542];
  assign o[47541] = i[47541];
  assign o[47540] = i[47540];
  assign o[47539] = i[47539];
  assign o[47538] = i[47538];
  assign o[47537] = i[47537];
  assign o[47536] = i[47536];
  assign o[47535] = i[47535];
  assign o[47534] = i[47534];
  assign o[47533] = i[47533];
  assign o[47532] = i[47532];
  assign o[47531] = i[47531];
  assign o[47530] = i[47530];
  assign o[47529] = i[47529];
  assign o[47528] = i[47528];
  assign o[47527] = i[47527];
  assign o[47526] = i[47526];
  assign o[47525] = i[47525];
  assign o[47524] = i[47524];
  assign o[47523] = i[47523];
  assign o[47522] = i[47522];
  assign o[47521] = i[47521];
  assign o[47520] = i[47520];
  assign o[47519] = i[47519];
  assign o[47518] = i[47518];
  assign o[47517] = i[47517];
  assign o[47516] = i[47516];
  assign o[47515] = i[47515];
  assign o[47514] = i[47514];
  assign o[47513] = i[47513];
  assign o[47512] = i[47512];
  assign o[47511] = i[47511];
  assign o[47510] = i[47510];
  assign o[47509] = i[47509];
  assign o[47508] = i[47508];
  assign o[47507] = i[47507];
  assign o[47506] = i[47506];
  assign o[47505] = i[47505];
  assign o[47504] = i[47504];
  assign o[47503] = i[47503];
  assign o[47502] = i[47502];
  assign o[47501] = i[47501];
  assign o[47500] = i[47500];
  assign o[47499] = i[47499];
  assign o[47498] = i[47498];
  assign o[47497] = i[47497];
  assign o[47496] = i[47496];
  assign o[47495] = i[47495];
  assign o[47494] = i[47494];
  assign o[47493] = i[47493];
  assign o[47492] = i[47492];
  assign o[47491] = i[47491];
  assign o[47490] = i[47490];
  assign o[47489] = i[47489];
  assign o[47488] = i[47488];
  assign o[47487] = i[47487];
  assign o[47486] = i[47486];
  assign o[47485] = i[47485];
  assign o[47484] = i[47484];
  assign o[47483] = i[47483];
  assign o[47482] = i[47482];
  assign o[47481] = i[47481];
  assign o[47480] = i[47480];
  assign o[47479] = i[47479];
  assign o[47478] = i[47478];
  assign o[47477] = i[47477];
  assign o[47476] = i[47476];
  assign o[47475] = i[47475];
  assign o[47474] = i[47474];
  assign o[47473] = i[47473];
  assign o[47472] = i[47472];
  assign o[47471] = i[47471];
  assign o[47470] = i[47470];
  assign o[47469] = i[47469];
  assign o[47468] = i[47468];
  assign o[47467] = i[47467];
  assign o[47466] = i[47466];
  assign o[47465] = i[47465];
  assign o[47464] = i[47464];
  assign o[47463] = i[47463];
  assign o[47462] = i[47462];
  assign o[47461] = i[47461];
  assign o[47460] = i[47460];
  assign o[47459] = i[47459];
  assign o[47458] = i[47458];
  assign o[47457] = i[47457];
  assign o[47456] = i[47456];
  assign o[47455] = i[47455];
  assign o[47454] = i[47454];
  assign o[47453] = i[47453];
  assign o[47452] = i[47452];
  assign o[47451] = i[47451];
  assign o[47450] = i[47450];
  assign o[47449] = i[47449];
  assign o[47448] = i[47448];
  assign o[47447] = i[47447];
  assign o[47446] = i[47446];
  assign o[47445] = i[47445];
  assign o[47444] = i[47444];
  assign o[47443] = i[47443];
  assign o[47442] = i[47442];
  assign o[47441] = i[47441];
  assign o[47440] = i[47440];
  assign o[47439] = i[47439];
  assign o[47438] = i[47438];
  assign o[47437] = i[47437];
  assign o[47436] = i[47436];
  assign o[47435] = i[47435];
  assign o[47434] = i[47434];
  assign o[47433] = i[47433];
  assign o[47432] = i[47432];
  assign o[47431] = i[47431];
  assign o[47430] = i[47430];
  assign o[47429] = i[47429];
  assign o[47428] = i[47428];
  assign o[47427] = i[47427];
  assign o[47426] = i[47426];
  assign o[47425] = i[47425];
  assign o[47424] = i[47424];
  assign o[47423] = i[47423];
  assign o[47422] = i[47422];
  assign o[47421] = i[47421];
  assign o[47420] = i[47420];
  assign o[47419] = i[47419];
  assign o[47418] = i[47418];
  assign o[47417] = i[47417];
  assign o[47416] = i[47416];
  assign o[47415] = i[47415];
  assign o[47414] = i[47414];
  assign o[47413] = i[47413];
  assign o[47412] = i[47412];
  assign o[47411] = i[47411];
  assign o[47410] = i[47410];
  assign o[47409] = i[47409];
  assign o[47408] = i[47408];
  assign o[47407] = i[47407];
  assign o[47406] = i[47406];
  assign o[47405] = i[47405];
  assign o[47404] = i[47404];
  assign o[47403] = i[47403];
  assign o[47402] = i[47402];
  assign o[47401] = i[47401];
  assign o[47400] = i[47400];
  assign o[47399] = i[47399];
  assign o[47398] = i[47398];
  assign o[47397] = i[47397];
  assign o[47396] = i[47396];
  assign o[47395] = i[47395];
  assign o[47394] = i[47394];
  assign o[47393] = i[47393];
  assign o[47392] = i[47392];
  assign o[47391] = i[47391];
  assign o[47390] = i[47390];
  assign o[47389] = i[47389];
  assign o[47388] = i[47388];
  assign o[47387] = i[47387];
  assign o[47386] = i[47386];
  assign o[47385] = i[47385];
  assign o[47384] = i[47384];
  assign o[47383] = i[47383];
  assign o[47382] = i[47382];
  assign o[47381] = i[47381];
  assign o[47380] = i[47380];
  assign o[47379] = i[47379];
  assign o[47378] = i[47378];
  assign o[47377] = i[47377];
  assign o[47376] = i[47376];
  assign o[47375] = i[47375];
  assign o[47374] = i[47374];
  assign o[47373] = i[47373];
  assign o[47372] = i[47372];
  assign o[47371] = i[47371];
  assign o[47370] = i[47370];
  assign o[47369] = i[47369];
  assign o[47368] = i[47368];
  assign o[47367] = i[47367];
  assign o[47366] = i[47366];
  assign o[47365] = i[47365];
  assign o[47364] = i[47364];
  assign o[47363] = i[47363];
  assign o[47362] = i[47362];
  assign o[47361] = i[47361];
  assign o[47360] = i[47360];
  assign o[47359] = i[47359];
  assign o[47358] = i[47358];
  assign o[47357] = i[47357];
  assign o[47356] = i[47356];
  assign o[47355] = i[47355];
  assign o[47354] = i[47354];
  assign o[47353] = i[47353];
  assign o[47352] = i[47352];
  assign o[47351] = i[47351];
  assign o[47350] = i[47350];
  assign o[47349] = i[47349];
  assign o[47348] = i[47348];
  assign o[47347] = i[47347];
  assign o[47346] = i[47346];
  assign o[47345] = i[47345];
  assign o[47344] = i[47344];
  assign o[47343] = i[47343];
  assign o[47342] = i[47342];
  assign o[47341] = i[47341];
  assign o[47340] = i[47340];
  assign o[47339] = i[47339];
  assign o[47338] = i[47338];
  assign o[47337] = i[47337];
  assign o[47336] = i[47336];
  assign o[47335] = i[47335];
  assign o[47334] = i[47334];
  assign o[47333] = i[47333];
  assign o[47332] = i[47332];
  assign o[47331] = i[47331];
  assign o[47330] = i[47330];
  assign o[47329] = i[47329];
  assign o[47328] = i[47328];
  assign o[47327] = i[47327];
  assign o[47326] = i[47326];
  assign o[47325] = i[47325];
  assign o[47324] = i[47324];
  assign o[47323] = i[47323];
  assign o[47322] = i[47322];
  assign o[47321] = i[47321];
  assign o[47320] = i[47320];
  assign o[47319] = i[47319];
  assign o[47318] = i[47318];
  assign o[47317] = i[47317];
  assign o[47316] = i[47316];
  assign o[47315] = i[47315];
  assign o[47314] = i[47314];
  assign o[47313] = i[47313];
  assign o[47312] = i[47312];
  assign o[47311] = i[47311];
  assign o[47310] = i[47310];
  assign o[47309] = i[47309];
  assign o[47308] = i[47308];
  assign o[47307] = i[47307];
  assign o[47306] = i[47306];
  assign o[47305] = i[47305];
  assign o[47304] = i[47304];
  assign o[47303] = i[47303];
  assign o[47302] = i[47302];
  assign o[47301] = i[47301];
  assign o[47300] = i[47300];
  assign o[47299] = i[47299];
  assign o[47298] = i[47298];
  assign o[47297] = i[47297];
  assign o[47296] = i[47296];
  assign o[47295] = i[47295];
  assign o[47294] = i[47294];
  assign o[47293] = i[47293];
  assign o[47292] = i[47292];
  assign o[47291] = i[47291];
  assign o[47290] = i[47290];
  assign o[47289] = i[47289];
  assign o[47288] = i[47288];
  assign o[47287] = i[47287];
  assign o[47286] = i[47286];
  assign o[47285] = i[47285];
  assign o[47284] = i[47284];
  assign o[47283] = i[47283];
  assign o[47282] = i[47282];
  assign o[47281] = i[47281];
  assign o[47280] = i[47280];
  assign o[47279] = i[47279];
  assign o[47278] = i[47278];
  assign o[47277] = i[47277];
  assign o[47276] = i[47276];
  assign o[47275] = i[47275];
  assign o[47274] = i[47274];
  assign o[47273] = i[47273];
  assign o[47272] = i[47272];
  assign o[47271] = i[47271];
  assign o[47270] = i[47270];
  assign o[47269] = i[47269];
  assign o[47268] = i[47268];
  assign o[47267] = i[47267];
  assign o[47266] = i[47266];
  assign o[47265] = i[47265];
  assign o[47264] = i[47264];
  assign o[47263] = i[47263];
  assign o[47262] = i[47262];
  assign o[47261] = i[47261];
  assign o[47260] = i[47260];
  assign o[47259] = i[47259];
  assign o[47258] = i[47258];
  assign o[47257] = i[47257];
  assign o[47256] = i[47256];
  assign o[47255] = i[47255];
  assign o[47254] = i[47254];
  assign o[47253] = i[47253];
  assign o[47252] = i[47252];
  assign o[47251] = i[47251];
  assign o[47250] = i[47250];
  assign o[47249] = i[47249];
  assign o[47248] = i[47248];
  assign o[47247] = i[47247];
  assign o[47246] = i[47246];
  assign o[47245] = i[47245];
  assign o[47244] = i[47244];
  assign o[47243] = i[47243];
  assign o[47242] = i[47242];
  assign o[47241] = i[47241];
  assign o[47240] = i[47240];
  assign o[47239] = i[47239];
  assign o[47238] = i[47238];
  assign o[47237] = i[47237];
  assign o[47236] = i[47236];
  assign o[47235] = i[47235];
  assign o[47234] = i[47234];
  assign o[47233] = i[47233];
  assign o[47232] = i[47232];
  assign o[47231] = i[47231];
  assign o[47230] = i[47230];
  assign o[47229] = i[47229];
  assign o[47228] = i[47228];
  assign o[47227] = i[47227];
  assign o[47226] = i[47226];
  assign o[47225] = i[47225];
  assign o[47224] = i[47224];
  assign o[47223] = i[47223];
  assign o[47222] = i[47222];
  assign o[47221] = i[47221];
  assign o[47220] = i[47220];
  assign o[47219] = i[47219];
  assign o[47218] = i[47218];
  assign o[47217] = i[47217];
  assign o[47216] = i[47216];
  assign o[47215] = i[47215];
  assign o[47214] = i[47214];
  assign o[47213] = i[47213];
  assign o[47212] = i[47212];
  assign o[47211] = i[47211];
  assign o[47210] = i[47210];
  assign o[47209] = i[47209];
  assign o[47208] = i[47208];
  assign o[47207] = i[47207];
  assign o[47206] = i[47206];
  assign o[47205] = i[47205];
  assign o[47204] = i[47204];
  assign o[47203] = i[47203];
  assign o[47202] = i[47202];
  assign o[47201] = i[47201];
  assign o[47200] = i[47200];
  assign o[47199] = i[47199];
  assign o[47198] = i[47198];
  assign o[47197] = i[47197];
  assign o[47196] = i[47196];
  assign o[47195] = i[47195];
  assign o[47194] = i[47194];
  assign o[47193] = i[47193];
  assign o[47192] = i[47192];
  assign o[47191] = i[47191];
  assign o[47190] = i[47190];
  assign o[47189] = i[47189];
  assign o[47188] = i[47188];
  assign o[47187] = i[47187];
  assign o[47186] = i[47186];
  assign o[47185] = i[47185];
  assign o[47184] = i[47184];
  assign o[47183] = i[47183];
  assign o[47182] = i[47182];
  assign o[47181] = i[47181];
  assign o[47180] = i[47180];
  assign o[47179] = i[47179];
  assign o[47178] = i[47178];
  assign o[47177] = i[47177];
  assign o[47176] = i[47176];
  assign o[47175] = i[47175];
  assign o[47174] = i[47174];
  assign o[47173] = i[47173];
  assign o[47172] = i[47172];
  assign o[47171] = i[47171];
  assign o[47170] = i[47170];
  assign o[47169] = i[47169];
  assign o[47168] = i[47168];
  assign o[47167] = i[47167];
  assign o[47166] = i[47166];
  assign o[47165] = i[47165];
  assign o[47164] = i[47164];
  assign o[47163] = i[47163];
  assign o[47162] = i[47162];
  assign o[47161] = i[47161];
  assign o[47160] = i[47160];
  assign o[47159] = i[47159];
  assign o[47158] = i[47158];
  assign o[47157] = i[47157];
  assign o[47156] = i[47156];
  assign o[47155] = i[47155];
  assign o[47154] = i[47154];
  assign o[47153] = i[47153];
  assign o[47152] = i[47152];
  assign o[47151] = i[47151];
  assign o[47150] = i[47150];
  assign o[47149] = i[47149];
  assign o[47148] = i[47148];
  assign o[47147] = i[47147];
  assign o[47146] = i[47146];
  assign o[47145] = i[47145];
  assign o[47144] = i[47144];
  assign o[47143] = i[47143];
  assign o[47142] = i[47142];
  assign o[47141] = i[47141];
  assign o[47140] = i[47140];
  assign o[47139] = i[47139];
  assign o[47138] = i[47138];
  assign o[47137] = i[47137];
  assign o[47136] = i[47136];
  assign o[47135] = i[47135];
  assign o[47134] = i[47134];
  assign o[47133] = i[47133];
  assign o[47132] = i[47132];
  assign o[47131] = i[47131];
  assign o[47130] = i[47130];
  assign o[47129] = i[47129];
  assign o[47128] = i[47128];
  assign o[47127] = i[47127];
  assign o[47126] = i[47126];
  assign o[47125] = i[47125];
  assign o[47124] = i[47124];
  assign o[47123] = i[47123];
  assign o[47122] = i[47122];
  assign o[47121] = i[47121];
  assign o[47120] = i[47120];
  assign o[47119] = i[47119];
  assign o[47118] = i[47118];
  assign o[47117] = i[47117];
  assign o[47116] = i[47116];
  assign o[47115] = i[47115];
  assign o[47114] = i[47114];
  assign o[47113] = i[47113];
  assign o[47112] = i[47112];
  assign o[47111] = i[47111];
  assign o[47110] = i[47110];
  assign o[47109] = i[47109];
  assign o[47108] = i[47108];
  assign o[47107] = i[47107];
  assign o[47106] = i[47106];
  assign o[47105] = i[47105];
  assign o[47104] = i[47104];
  assign o[47103] = i[47103];
  assign o[47102] = i[47102];
  assign o[47101] = i[47101];
  assign o[47100] = i[47100];
  assign o[47099] = i[47099];
  assign o[47098] = i[47098];
  assign o[47097] = i[47097];
  assign o[47096] = i[47096];
  assign o[47095] = i[47095];
  assign o[47094] = i[47094];
  assign o[47093] = i[47093];
  assign o[47092] = i[47092];
  assign o[47091] = i[47091];
  assign o[47090] = i[47090];
  assign o[47089] = i[47089];
  assign o[47088] = i[47088];
  assign o[47087] = i[47087];
  assign o[47086] = i[47086];
  assign o[47085] = i[47085];
  assign o[47084] = i[47084];
  assign o[47083] = i[47083];
  assign o[47082] = i[47082];
  assign o[47081] = i[47081];
  assign o[47080] = i[47080];
  assign o[47079] = i[47079];
  assign o[47078] = i[47078];
  assign o[47077] = i[47077];
  assign o[47076] = i[47076];
  assign o[47075] = i[47075];
  assign o[47074] = i[47074];
  assign o[47073] = i[47073];
  assign o[47072] = i[47072];
  assign o[47071] = i[47071];
  assign o[47070] = i[47070];
  assign o[47069] = i[47069];
  assign o[47068] = i[47068];
  assign o[47067] = i[47067];
  assign o[47066] = i[47066];
  assign o[47065] = i[47065];
  assign o[47064] = i[47064];
  assign o[47063] = i[47063];
  assign o[47062] = i[47062];
  assign o[47061] = i[47061];
  assign o[47060] = i[47060];
  assign o[47059] = i[47059];
  assign o[47058] = i[47058];
  assign o[47057] = i[47057];
  assign o[47056] = i[47056];
  assign o[47055] = i[47055];
  assign o[47054] = i[47054];
  assign o[47053] = i[47053];
  assign o[47052] = i[47052];
  assign o[47051] = i[47051];
  assign o[47050] = i[47050];
  assign o[47049] = i[47049];
  assign o[47048] = i[47048];
  assign o[47047] = i[47047];
  assign o[47046] = i[47046];
  assign o[47045] = i[47045];
  assign o[47044] = i[47044];
  assign o[47043] = i[47043];
  assign o[47042] = i[47042];
  assign o[47041] = i[47041];
  assign o[47040] = i[47040];
  assign o[47039] = i[47039];
  assign o[47038] = i[47038];
  assign o[47037] = i[47037];
  assign o[47036] = i[47036];
  assign o[47035] = i[47035];
  assign o[47034] = i[47034];
  assign o[47033] = i[47033];
  assign o[47032] = i[47032];
  assign o[47031] = i[47031];
  assign o[47030] = i[47030];
  assign o[47029] = i[47029];
  assign o[47028] = i[47028];
  assign o[47027] = i[47027];
  assign o[47026] = i[47026];
  assign o[47025] = i[47025];
  assign o[47024] = i[47024];
  assign o[47023] = i[47023];
  assign o[47022] = i[47022];
  assign o[47021] = i[47021];
  assign o[47020] = i[47020];
  assign o[47019] = i[47019];
  assign o[47018] = i[47018];
  assign o[47017] = i[47017];
  assign o[47016] = i[47016];
  assign o[47015] = i[47015];
  assign o[47014] = i[47014];
  assign o[47013] = i[47013];
  assign o[47012] = i[47012];
  assign o[47011] = i[47011];
  assign o[47010] = i[47010];
  assign o[47009] = i[47009];
  assign o[47008] = i[47008];
  assign o[47007] = i[47007];
  assign o[47006] = i[47006];
  assign o[47005] = i[47005];
  assign o[47004] = i[47004];
  assign o[47003] = i[47003];
  assign o[47002] = i[47002];
  assign o[47001] = i[47001];
  assign o[47000] = i[47000];
  assign o[46999] = i[46999];
  assign o[46998] = i[46998];
  assign o[46997] = i[46997];
  assign o[46996] = i[46996];
  assign o[46995] = i[46995];
  assign o[46994] = i[46994];
  assign o[46993] = i[46993];
  assign o[46992] = i[46992];
  assign o[46991] = i[46991];
  assign o[46990] = i[46990];
  assign o[46989] = i[46989];
  assign o[46988] = i[46988];
  assign o[46987] = i[46987];
  assign o[46986] = i[46986];
  assign o[46985] = i[46985];
  assign o[46984] = i[46984];
  assign o[46983] = i[46983];
  assign o[46982] = i[46982];
  assign o[46981] = i[46981];
  assign o[46980] = i[46980];
  assign o[46979] = i[46979];
  assign o[46978] = i[46978];
  assign o[46977] = i[46977];
  assign o[46976] = i[46976];
  assign o[46975] = i[46975];
  assign o[46974] = i[46974];
  assign o[46973] = i[46973];
  assign o[46972] = i[46972];
  assign o[46971] = i[46971];
  assign o[46970] = i[46970];
  assign o[46969] = i[46969];
  assign o[46968] = i[46968];
  assign o[46967] = i[46967];
  assign o[46966] = i[46966];
  assign o[46965] = i[46965];
  assign o[46964] = i[46964];
  assign o[46963] = i[46963];
  assign o[46962] = i[46962];
  assign o[46961] = i[46961];
  assign o[46960] = i[46960];
  assign o[46959] = i[46959];
  assign o[46958] = i[46958];
  assign o[46957] = i[46957];
  assign o[46956] = i[46956];
  assign o[46955] = i[46955];
  assign o[46954] = i[46954];
  assign o[46953] = i[46953];
  assign o[46952] = i[46952];
  assign o[46951] = i[46951];
  assign o[46950] = i[46950];
  assign o[46949] = i[46949];
  assign o[46948] = i[46948];
  assign o[46947] = i[46947];
  assign o[46946] = i[46946];
  assign o[46945] = i[46945];
  assign o[46944] = i[46944];
  assign o[46943] = i[46943];
  assign o[46942] = i[46942];
  assign o[46941] = i[46941];
  assign o[46940] = i[46940];
  assign o[46939] = i[46939];
  assign o[46938] = i[46938];
  assign o[46937] = i[46937];
  assign o[46936] = i[46936];
  assign o[46935] = i[46935];
  assign o[46934] = i[46934];
  assign o[46933] = i[46933];
  assign o[46932] = i[46932];
  assign o[46931] = i[46931];
  assign o[46930] = i[46930];
  assign o[46929] = i[46929];
  assign o[46928] = i[46928];
  assign o[46927] = i[46927];
  assign o[46926] = i[46926];
  assign o[46925] = i[46925];
  assign o[46924] = i[46924];
  assign o[46923] = i[46923];
  assign o[46922] = i[46922];
  assign o[46921] = i[46921];
  assign o[46920] = i[46920];
  assign o[46919] = i[46919];
  assign o[46918] = i[46918];
  assign o[46917] = i[46917];
  assign o[46916] = i[46916];
  assign o[46915] = i[46915];
  assign o[46914] = i[46914];
  assign o[46913] = i[46913];
  assign o[46912] = i[46912];
  assign o[46911] = i[46911];
  assign o[46910] = i[46910];
  assign o[46909] = i[46909];
  assign o[46908] = i[46908];
  assign o[46907] = i[46907];
  assign o[46906] = i[46906];
  assign o[46905] = i[46905];
  assign o[46904] = i[46904];
  assign o[46903] = i[46903];
  assign o[46902] = i[46902];
  assign o[46901] = i[46901];
  assign o[46900] = i[46900];
  assign o[46899] = i[46899];
  assign o[46898] = i[46898];
  assign o[46897] = i[46897];
  assign o[46896] = i[46896];
  assign o[46895] = i[46895];
  assign o[46894] = i[46894];
  assign o[46893] = i[46893];
  assign o[46892] = i[46892];
  assign o[46891] = i[46891];
  assign o[46890] = i[46890];
  assign o[46889] = i[46889];
  assign o[46888] = i[46888];
  assign o[46887] = i[46887];
  assign o[46886] = i[46886];
  assign o[46885] = i[46885];
  assign o[46884] = i[46884];
  assign o[46883] = i[46883];
  assign o[46882] = i[46882];
  assign o[46881] = i[46881];
  assign o[46880] = i[46880];
  assign o[46879] = i[46879];
  assign o[46878] = i[46878];
  assign o[46877] = i[46877];
  assign o[46876] = i[46876];
  assign o[46875] = i[46875];
  assign o[46874] = i[46874];
  assign o[46873] = i[46873];
  assign o[46872] = i[46872];
  assign o[46871] = i[46871];
  assign o[46870] = i[46870];
  assign o[46869] = i[46869];
  assign o[46868] = i[46868];
  assign o[46867] = i[46867];
  assign o[46866] = i[46866];
  assign o[46865] = i[46865];
  assign o[46864] = i[46864];
  assign o[46863] = i[46863];
  assign o[46862] = i[46862];
  assign o[46861] = i[46861];
  assign o[46860] = i[46860];
  assign o[46859] = i[46859];
  assign o[46858] = i[46858];
  assign o[46857] = i[46857];
  assign o[46856] = i[46856];
  assign o[46855] = i[46855];
  assign o[46854] = i[46854];
  assign o[46853] = i[46853];
  assign o[46852] = i[46852];
  assign o[46851] = i[46851];
  assign o[46850] = i[46850];
  assign o[46849] = i[46849];
  assign o[46848] = i[46848];
  assign o[46847] = i[46847];
  assign o[46846] = i[46846];
  assign o[46845] = i[46845];
  assign o[46844] = i[46844];
  assign o[46843] = i[46843];
  assign o[46842] = i[46842];
  assign o[46841] = i[46841];
  assign o[46840] = i[46840];
  assign o[46839] = i[46839];
  assign o[46838] = i[46838];
  assign o[46837] = i[46837];
  assign o[46836] = i[46836];
  assign o[46835] = i[46835];
  assign o[46834] = i[46834];
  assign o[46833] = i[46833];
  assign o[46832] = i[46832];
  assign o[46831] = i[46831];
  assign o[46830] = i[46830];
  assign o[46829] = i[46829];
  assign o[46828] = i[46828];
  assign o[46827] = i[46827];
  assign o[46826] = i[46826];
  assign o[46825] = i[46825];
  assign o[46824] = i[46824];
  assign o[46823] = i[46823];
  assign o[46822] = i[46822];
  assign o[46821] = i[46821];
  assign o[46820] = i[46820];
  assign o[46819] = i[46819];
  assign o[46818] = i[46818];
  assign o[46817] = i[46817];
  assign o[46816] = i[46816];
  assign o[46815] = i[46815];
  assign o[46814] = i[46814];
  assign o[46813] = i[46813];
  assign o[46812] = i[46812];
  assign o[46811] = i[46811];
  assign o[46810] = i[46810];
  assign o[46809] = i[46809];
  assign o[46808] = i[46808];
  assign o[46807] = i[46807];
  assign o[46806] = i[46806];
  assign o[46805] = i[46805];
  assign o[46804] = i[46804];
  assign o[46803] = i[46803];
  assign o[46802] = i[46802];
  assign o[46801] = i[46801];
  assign o[46800] = i[46800];
  assign o[46799] = i[46799];
  assign o[46798] = i[46798];
  assign o[46797] = i[46797];
  assign o[46796] = i[46796];
  assign o[46795] = i[46795];
  assign o[46794] = i[46794];
  assign o[46793] = i[46793];
  assign o[46792] = i[46792];
  assign o[46791] = i[46791];
  assign o[46790] = i[46790];
  assign o[46789] = i[46789];
  assign o[46788] = i[46788];
  assign o[46787] = i[46787];
  assign o[46786] = i[46786];
  assign o[46785] = i[46785];
  assign o[46784] = i[46784];
  assign o[46783] = i[46783];
  assign o[46782] = i[46782];
  assign o[46781] = i[46781];
  assign o[46780] = i[46780];
  assign o[46779] = i[46779];
  assign o[46778] = i[46778];
  assign o[46777] = i[46777];
  assign o[46776] = i[46776];
  assign o[46775] = i[46775];
  assign o[46774] = i[46774];
  assign o[46773] = i[46773];
  assign o[46772] = i[46772];
  assign o[46771] = i[46771];
  assign o[46770] = i[46770];
  assign o[46769] = i[46769];
  assign o[46768] = i[46768];
  assign o[46767] = i[46767];
  assign o[46766] = i[46766];
  assign o[46765] = i[46765];
  assign o[46764] = i[46764];
  assign o[46763] = i[46763];
  assign o[46762] = i[46762];
  assign o[46761] = i[46761];
  assign o[46760] = i[46760];
  assign o[46759] = i[46759];
  assign o[46758] = i[46758];
  assign o[46757] = i[46757];
  assign o[46756] = i[46756];
  assign o[46755] = i[46755];
  assign o[46754] = i[46754];
  assign o[46753] = i[46753];
  assign o[46752] = i[46752];
  assign o[46751] = i[46751];
  assign o[46750] = i[46750];
  assign o[46749] = i[46749];
  assign o[46748] = i[46748];
  assign o[46747] = i[46747];
  assign o[46746] = i[46746];
  assign o[46745] = i[46745];
  assign o[46744] = i[46744];
  assign o[46743] = i[46743];
  assign o[46742] = i[46742];
  assign o[46741] = i[46741];
  assign o[46740] = i[46740];
  assign o[46739] = i[46739];
  assign o[46738] = i[46738];
  assign o[46737] = i[46737];
  assign o[46736] = i[46736];
  assign o[46735] = i[46735];
  assign o[46734] = i[46734];
  assign o[46733] = i[46733];
  assign o[46732] = i[46732];
  assign o[46731] = i[46731];
  assign o[46730] = i[46730];
  assign o[46729] = i[46729];
  assign o[46728] = i[46728];
  assign o[46727] = i[46727];
  assign o[46726] = i[46726];
  assign o[46725] = i[46725];
  assign o[46724] = i[46724];
  assign o[46723] = i[46723];
  assign o[46722] = i[46722];
  assign o[46721] = i[46721];
  assign o[46720] = i[46720];
  assign o[46719] = i[46719];
  assign o[46718] = i[46718];
  assign o[46717] = i[46717];
  assign o[46716] = i[46716];
  assign o[46715] = i[46715];
  assign o[46714] = i[46714];
  assign o[46713] = i[46713];
  assign o[46712] = i[46712];
  assign o[46711] = i[46711];
  assign o[46710] = i[46710];
  assign o[46709] = i[46709];
  assign o[46708] = i[46708];
  assign o[46707] = i[46707];
  assign o[46706] = i[46706];
  assign o[46705] = i[46705];
  assign o[46704] = i[46704];
  assign o[46703] = i[46703];
  assign o[46702] = i[46702];
  assign o[46701] = i[46701];
  assign o[46700] = i[46700];
  assign o[46699] = i[46699];
  assign o[46698] = i[46698];
  assign o[46697] = i[46697];
  assign o[46696] = i[46696];
  assign o[46695] = i[46695];
  assign o[46694] = i[46694];
  assign o[46693] = i[46693];
  assign o[46692] = i[46692];
  assign o[46691] = i[46691];
  assign o[46690] = i[46690];
  assign o[46689] = i[46689];
  assign o[46688] = i[46688];
  assign o[46687] = i[46687];
  assign o[46686] = i[46686];
  assign o[46685] = i[46685];
  assign o[46684] = i[46684];
  assign o[46683] = i[46683];
  assign o[46682] = i[46682];
  assign o[46681] = i[46681];
  assign o[46680] = i[46680];
  assign o[46679] = i[46679];
  assign o[46678] = i[46678];
  assign o[46677] = i[46677];
  assign o[46676] = i[46676];
  assign o[46675] = i[46675];
  assign o[46674] = i[46674];
  assign o[46673] = i[46673];
  assign o[46672] = i[46672];
  assign o[46671] = i[46671];
  assign o[46670] = i[46670];
  assign o[46669] = i[46669];
  assign o[46668] = i[46668];
  assign o[46667] = i[46667];
  assign o[46666] = i[46666];
  assign o[46665] = i[46665];
  assign o[46664] = i[46664];
  assign o[46663] = i[46663];
  assign o[46662] = i[46662];
  assign o[46661] = i[46661];
  assign o[46660] = i[46660];
  assign o[46659] = i[46659];
  assign o[46658] = i[46658];
  assign o[46657] = i[46657];
  assign o[46656] = i[46656];
  assign o[46655] = i[46655];
  assign o[46654] = i[46654];
  assign o[46653] = i[46653];
  assign o[46652] = i[46652];
  assign o[46651] = i[46651];
  assign o[46650] = i[46650];
  assign o[46649] = i[46649];
  assign o[46648] = i[46648];
  assign o[46647] = i[46647];
  assign o[46646] = i[46646];
  assign o[46645] = i[46645];
  assign o[46644] = i[46644];
  assign o[46643] = i[46643];
  assign o[46642] = i[46642];
  assign o[46641] = i[46641];
  assign o[46640] = i[46640];
  assign o[46639] = i[46639];
  assign o[46638] = i[46638];
  assign o[46637] = i[46637];
  assign o[46636] = i[46636];
  assign o[46635] = i[46635];
  assign o[46634] = i[46634];
  assign o[46633] = i[46633];
  assign o[46632] = i[46632];
  assign o[46631] = i[46631];
  assign o[46630] = i[46630];
  assign o[46629] = i[46629];
  assign o[46628] = i[46628];
  assign o[46627] = i[46627];
  assign o[46626] = i[46626];
  assign o[46625] = i[46625];
  assign o[46624] = i[46624];
  assign o[46623] = i[46623];
  assign o[46622] = i[46622];
  assign o[46621] = i[46621];
  assign o[46620] = i[46620];
  assign o[46619] = i[46619];
  assign o[46618] = i[46618];
  assign o[46617] = i[46617];
  assign o[46616] = i[46616];
  assign o[46615] = i[46615];
  assign o[46614] = i[46614];
  assign o[46613] = i[46613];
  assign o[46612] = i[46612];
  assign o[46611] = i[46611];
  assign o[46610] = i[46610];
  assign o[46609] = i[46609];
  assign o[46608] = i[46608];
  assign o[46607] = i[46607];
  assign o[46606] = i[46606];
  assign o[46605] = i[46605];
  assign o[46604] = i[46604];
  assign o[46603] = i[46603];
  assign o[46602] = i[46602];
  assign o[46601] = i[46601];
  assign o[46600] = i[46600];
  assign o[46599] = i[46599];
  assign o[46598] = i[46598];
  assign o[46597] = i[46597];
  assign o[46596] = i[46596];
  assign o[46595] = i[46595];
  assign o[46594] = i[46594];
  assign o[46593] = i[46593];
  assign o[46592] = i[46592];
  assign o[46591] = i[46591];
  assign o[46590] = i[46590];
  assign o[46589] = i[46589];
  assign o[46588] = i[46588];
  assign o[46587] = i[46587];
  assign o[46586] = i[46586];
  assign o[46585] = i[46585];
  assign o[46584] = i[46584];
  assign o[46583] = i[46583];
  assign o[46582] = i[46582];
  assign o[46581] = i[46581];
  assign o[46580] = i[46580];
  assign o[46579] = i[46579];
  assign o[46578] = i[46578];
  assign o[46577] = i[46577];
  assign o[46576] = i[46576];
  assign o[46575] = i[46575];
  assign o[46574] = i[46574];
  assign o[46573] = i[46573];
  assign o[46572] = i[46572];
  assign o[46571] = i[46571];
  assign o[46570] = i[46570];
  assign o[46569] = i[46569];
  assign o[46568] = i[46568];
  assign o[46567] = i[46567];
  assign o[46566] = i[46566];
  assign o[46565] = i[46565];
  assign o[46564] = i[46564];
  assign o[46563] = i[46563];
  assign o[46562] = i[46562];
  assign o[46561] = i[46561];
  assign o[46560] = i[46560];
  assign o[46559] = i[46559];
  assign o[46558] = i[46558];
  assign o[46557] = i[46557];
  assign o[46556] = i[46556];
  assign o[46555] = i[46555];
  assign o[46554] = i[46554];
  assign o[46553] = i[46553];
  assign o[46552] = i[46552];
  assign o[46551] = i[46551];
  assign o[46550] = i[46550];
  assign o[46549] = i[46549];
  assign o[46548] = i[46548];
  assign o[46547] = i[46547];
  assign o[46546] = i[46546];
  assign o[46545] = i[46545];
  assign o[46544] = i[46544];
  assign o[46543] = i[46543];
  assign o[46542] = i[46542];
  assign o[46541] = i[46541];
  assign o[46540] = i[46540];
  assign o[46539] = i[46539];
  assign o[46538] = i[46538];
  assign o[46537] = i[46537];
  assign o[46536] = i[46536];
  assign o[46535] = i[46535];
  assign o[46534] = i[46534];
  assign o[46533] = i[46533];
  assign o[46532] = i[46532];
  assign o[46531] = i[46531];
  assign o[46530] = i[46530];
  assign o[46529] = i[46529];
  assign o[46528] = i[46528];
  assign o[46527] = i[46527];
  assign o[46526] = i[46526];
  assign o[46525] = i[46525];
  assign o[46524] = i[46524];
  assign o[46523] = i[46523];
  assign o[46522] = i[46522];
  assign o[46521] = i[46521];
  assign o[46520] = i[46520];
  assign o[46519] = i[46519];
  assign o[46518] = i[46518];
  assign o[46517] = i[46517];
  assign o[46516] = i[46516];
  assign o[46515] = i[46515];
  assign o[46514] = i[46514];
  assign o[46513] = i[46513];
  assign o[46512] = i[46512];
  assign o[46511] = i[46511];
  assign o[46510] = i[46510];
  assign o[46509] = i[46509];
  assign o[46508] = i[46508];
  assign o[46507] = i[46507];
  assign o[46506] = i[46506];
  assign o[46505] = i[46505];
  assign o[46504] = i[46504];
  assign o[46503] = i[46503];
  assign o[46502] = i[46502];
  assign o[46501] = i[46501];
  assign o[46500] = i[46500];
  assign o[46499] = i[46499];
  assign o[46498] = i[46498];
  assign o[46497] = i[46497];
  assign o[46496] = i[46496];
  assign o[46495] = i[46495];
  assign o[46494] = i[46494];
  assign o[46493] = i[46493];
  assign o[46492] = i[46492];
  assign o[46491] = i[46491];
  assign o[46490] = i[46490];
  assign o[46489] = i[46489];
  assign o[46488] = i[46488];
  assign o[46487] = i[46487];
  assign o[46486] = i[46486];
  assign o[46485] = i[46485];
  assign o[46484] = i[46484];
  assign o[46483] = i[46483];
  assign o[46482] = i[46482];
  assign o[46481] = i[46481];
  assign o[46480] = i[46480];
  assign o[46479] = i[46479];
  assign o[46478] = i[46478];
  assign o[46477] = i[46477];
  assign o[46476] = i[46476];
  assign o[46475] = i[46475];
  assign o[46474] = i[46474];
  assign o[46473] = i[46473];
  assign o[46472] = i[46472];
  assign o[46471] = i[46471];
  assign o[46470] = i[46470];
  assign o[46469] = i[46469];
  assign o[46468] = i[46468];
  assign o[46467] = i[46467];
  assign o[46466] = i[46466];
  assign o[46465] = i[46465];
  assign o[46464] = i[46464];
  assign o[46463] = i[46463];
  assign o[46462] = i[46462];
  assign o[46461] = i[46461];
  assign o[46460] = i[46460];
  assign o[46459] = i[46459];
  assign o[46458] = i[46458];
  assign o[46457] = i[46457];
  assign o[46456] = i[46456];
  assign o[46455] = i[46455];
  assign o[46454] = i[46454];
  assign o[46453] = i[46453];
  assign o[46452] = i[46452];
  assign o[46451] = i[46451];
  assign o[46450] = i[46450];
  assign o[46449] = i[46449];
  assign o[46448] = i[46448];
  assign o[46447] = i[46447];
  assign o[46446] = i[46446];
  assign o[46445] = i[46445];
  assign o[46444] = i[46444];
  assign o[46443] = i[46443];
  assign o[46442] = i[46442];
  assign o[46441] = i[46441];
  assign o[46440] = i[46440];
  assign o[46439] = i[46439];
  assign o[46438] = i[46438];
  assign o[46437] = i[46437];
  assign o[46436] = i[46436];
  assign o[46435] = i[46435];
  assign o[46434] = i[46434];
  assign o[46433] = i[46433];
  assign o[46432] = i[46432];
  assign o[46431] = i[46431];
  assign o[46430] = i[46430];
  assign o[46429] = i[46429];
  assign o[46428] = i[46428];
  assign o[46427] = i[46427];
  assign o[46426] = i[46426];
  assign o[46425] = i[46425];
  assign o[46424] = i[46424];
  assign o[46423] = i[46423];
  assign o[46422] = i[46422];
  assign o[46421] = i[46421];
  assign o[46420] = i[46420];
  assign o[46419] = i[46419];
  assign o[46418] = i[46418];
  assign o[46417] = i[46417];
  assign o[46416] = i[46416];
  assign o[46415] = i[46415];
  assign o[46414] = i[46414];
  assign o[46413] = i[46413];
  assign o[46412] = i[46412];
  assign o[46411] = i[46411];
  assign o[46410] = i[46410];
  assign o[46409] = i[46409];
  assign o[46408] = i[46408];
  assign o[46407] = i[46407];
  assign o[46406] = i[46406];
  assign o[46405] = i[46405];
  assign o[46404] = i[46404];
  assign o[46403] = i[46403];
  assign o[46402] = i[46402];
  assign o[46401] = i[46401];
  assign o[46400] = i[46400];
  assign o[46399] = i[46399];
  assign o[46398] = i[46398];
  assign o[46397] = i[46397];
  assign o[46396] = i[46396];
  assign o[46395] = i[46395];
  assign o[46394] = i[46394];
  assign o[46393] = i[46393];
  assign o[46392] = i[46392];
  assign o[46391] = i[46391];
  assign o[46390] = i[46390];
  assign o[46389] = i[46389];
  assign o[46388] = i[46388];
  assign o[46387] = i[46387];
  assign o[46386] = i[46386];
  assign o[46385] = i[46385];
  assign o[46384] = i[46384];
  assign o[46383] = i[46383];
  assign o[46382] = i[46382];
  assign o[46381] = i[46381];
  assign o[46380] = i[46380];
  assign o[46379] = i[46379];
  assign o[46378] = i[46378];
  assign o[46377] = i[46377];
  assign o[46376] = i[46376];
  assign o[46375] = i[46375];
  assign o[46374] = i[46374];
  assign o[46373] = i[46373];
  assign o[46372] = i[46372];
  assign o[46371] = i[46371];
  assign o[46370] = i[46370];
  assign o[46369] = i[46369];
  assign o[46368] = i[46368];
  assign o[46367] = i[46367];
  assign o[46366] = i[46366];
  assign o[46365] = i[46365];
  assign o[46364] = i[46364];
  assign o[46363] = i[46363];
  assign o[46362] = i[46362];
  assign o[46361] = i[46361];
  assign o[46360] = i[46360];
  assign o[46359] = i[46359];
  assign o[46358] = i[46358];
  assign o[46357] = i[46357];
  assign o[46356] = i[46356];
  assign o[46355] = i[46355];
  assign o[46354] = i[46354];
  assign o[46353] = i[46353];
  assign o[46352] = i[46352];
  assign o[46351] = i[46351];
  assign o[46350] = i[46350];
  assign o[46349] = i[46349];
  assign o[46348] = i[46348];
  assign o[46347] = i[46347];
  assign o[46346] = i[46346];
  assign o[46345] = i[46345];
  assign o[46344] = i[46344];
  assign o[46343] = i[46343];
  assign o[46342] = i[46342];
  assign o[46341] = i[46341];
  assign o[46340] = i[46340];
  assign o[46339] = i[46339];
  assign o[46338] = i[46338];
  assign o[46337] = i[46337];
  assign o[46336] = i[46336];
  assign o[46335] = i[46335];
  assign o[46334] = i[46334];
  assign o[46333] = i[46333];
  assign o[46332] = i[46332];
  assign o[46331] = i[46331];
  assign o[46330] = i[46330];
  assign o[46329] = i[46329];
  assign o[46328] = i[46328];
  assign o[46327] = i[46327];
  assign o[46326] = i[46326];
  assign o[46325] = i[46325];
  assign o[46324] = i[46324];
  assign o[46323] = i[46323];
  assign o[46322] = i[46322];
  assign o[46321] = i[46321];
  assign o[46320] = i[46320];
  assign o[46319] = i[46319];
  assign o[46318] = i[46318];
  assign o[46317] = i[46317];
  assign o[46316] = i[46316];
  assign o[46315] = i[46315];
  assign o[46314] = i[46314];
  assign o[46313] = i[46313];
  assign o[46312] = i[46312];
  assign o[46311] = i[46311];
  assign o[46310] = i[46310];
  assign o[46309] = i[46309];
  assign o[46308] = i[46308];
  assign o[46307] = i[46307];
  assign o[46306] = i[46306];
  assign o[46305] = i[46305];
  assign o[46304] = i[46304];
  assign o[46303] = i[46303];
  assign o[46302] = i[46302];
  assign o[46301] = i[46301];
  assign o[46300] = i[46300];
  assign o[46299] = i[46299];
  assign o[46298] = i[46298];
  assign o[46297] = i[46297];
  assign o[46296] = i[46296];
  assign o[46295] = i[46295];
  assign o[46294] = i[46294];
  assign o[46293] = i[46293];
  assign o[46292] = i[46292];
  assign o[46291] = i[46291];
  assign o[46290] = i[46290];
  assign o[46289] = i[46289];
  assign o[46288] = i[46288];
  assign o[46287] = i[46287];
  assign o[46286] = i[46286];
  assign o[46285] = i[46285];
  assign o[46284] = i[46284];
  assign o[46283] = i[46283];
  assign o[46282] = i[46282];
  assign o[46281] = i[46281];
  assign o[46280] = i[46280];
  assign o[46279] = i[46279];
  assign o[46278] = i[46278];
  assign o[46277] = i[46277];
  assign o[46276] = i[46276];
  assign o[46275] = i[46275];
  assign o[46274] = i[46274];
  assign o[46273] = i[46273];
  assign o[46272] = i[46272];
  assign o[46271] = i[46271];
  assign o[46270] = i[46270];
  assign o[46269] = i[46269];
  assign o[46268] = i[46268];
  assign o[46267] = i[46267];
  assign o[46266] = i[46266];
  assign o[46265] = i[46265];
  assign o[46264] = i[46264];
  assign o[46263] = i[46263];
  assign o[46262] = i[46262];
  assign o[46261] = i[46261];
  assign o[46260] = i[46260];
  assign o[46259] = i[46259];
  assign o[46258] = i[46258];
  assign o[46257] = i[46257];
  assign o[46256] = i[46256];
  assign o[46255] = i[46255];
  assign o[46254] = i[46254];
  assign o[46253] = i[46253];
  assign o[46252] = i[46252];
  assign o[46251] = i[46251];
  assign o[46250] = i[46250];
  assign o[46249] = i[46249];
  assign o[46248] = i[46248];
  assign o[46247] = i[46247];
  assign o[46246] = i[46246];
  assign o[46245] = i[46245];
  assign o[46244] = i[46244];
  assign o[46243] = i[46243];
  assign o[46242] = i[46242];
  assign o[46241] = i[46241];
  assign o[46240] = i[46240];
  assign o[46239] = i[46239];
  assign o[46238] = i[46238];
  assign o[46237] = i[46237];
  assign o[46236] = i[46236];
  assign o[46235] = i[46235];
  assign o[46234] = i[46234];
  assign o[46233] = i[46233];
  assign o[46232] = i[46232];
  assign o[46231] = i[46231];
  assign o[46230] = i[46230];
  assign o[46229] = i[46229];
  assign o[46228] = i[46228];
  assign o[46227] = i[46227];
  assign o[46226] = i[46226];
  assign o[46225] = i[46225];
  assign o[46224] = i[46224];
  assign o[46223] = i[46223];
  assign o[46222] = i[46222];
  assign o[46221] = i[46221];
  assign o[46220] = i[46220];
  assign o[46219] = i[46219];
  assign o[46218] = i[46218];
  assign o[46217] = i[46217];
  assign o[46216] = i[46216];
  assign o[46215] = i[46215];
  assign o[46214] = i[46214];
  assign o[46213] = i[46213];
  assign o[46212] = i[46212];
  assign o[46211] = i[46211];
  assign o[46210] = i[46210];
  assign o[46209] = i[46209];
  assign o[46208] = i[46208];
  assign o[46207] = i[46207];
  assign o[46206] = i[46206];
  assign o[46205] = i[46205];
  assign o[46204] = i[46204];
  assign o[46203] = i[46203];
  assign o[46202] = i[46202];
  assign o[46201] = i[46201];
  assign o[46200] = i[46200];
  assign o[46199] = i[46199];
  assign o[46198] = i[46198];
  assign o[46197] = i[46197];
  assign o[46196] = i[46196];
  assign o[46195] = i[46195];
  assign o[46194] = i[46194];
  assign o[46193] = i[46193];
  assign o[46192] = i[46192];
  assign o[46191] = i[46191];
  assign o[46190] = i[46190];
  assign o[46189] = i[46189];
  assign o[46188] = i[46188];
  assign o[46187] = i[46187];
  assign o[46186] = i[46186];
  assign o[46185] = i[46185];
  assign o[46184] = i[46184];
  assign o[46183] = i[46183];
  assign o[46182] = i[46182];
  assign o[46181] = i[46181];
  assign o[46180] = i[46180];
  assign o[46179] = i[46179];
  assign o[46178] = i[46178];
  assign o[46177] = i[46177];
  assign o[46176] = i[46176];
  assign o[46175] = i[46175];
  assign o[46174] = i[46174];
  assign o[46173] = i[46173];
  assign o[46172] = i[46172];
  assign o[46171] = i[46171];
  assign o[46170] = i[46170];
  assign o[46169] = i[46169];
  assign o[46168] = i[46168];
  assign o[46167] = i[46167];
  assign o[46166] = i[46166];
  assign o[46165] = i[46165];
  assign o[46164] = i[46164];
  assign o[46163] = i[46163];
  assign o[46162] = i[46162];
  assign o[46161] = i[46161];
  assign o[46160] = i[46160];
  assign o[46159] = i[46159];
  assign o[46158] = i[46158];
  assign o[46157] = i[46157];
  assign o[46156] = i[46156];
  assign o[46155] = i[46155];
  assign o[46154] = i[46154];
  assign o[46153] = i[46153];
  assign o[46152] = i[46152];
  assign o[46151] = i[46151];
  assign o[46150] = i[46150];
  assign o[46149] = i[46149];
  assign o[46148] = i[46148];
  assign o[46147] = i[46147];
  assign o[46146] = i[46146];
  assign o[46145] = i[46145];
  assign o[46144] = i[46144];
  assign o[46143] = i[46143];
  assign o[46142] = i[46142];
  assign o[46141] = i[46141];
  assign o[46140] = i[46140];
  assign o[46139] = i[46139];
  assign o[46138] = i[46138];
  assign o[46137] = i[46137];
  assign o[46136] = i[46136];
  assign o[46135] = i[46135];
  assign o[46134] = i[46134];
  assign o[46133] = i[46133];
  assign o[46132] = i[46132];
  assign o[46131] = i[46131];
  assign o[46130] = i[46130];
  assign o[46129] = i[46129];
  assign o[46128] = i[46128];
  assign o[46127] = i[46127];
  assign o[46126] = i[46126];
  assign o[46125] = i[46125];
  assign o[46124] = i[46124];
  assign o[46123] = i[46123];
  assign o[46122] = i[46122];
  assign o[46121] = i[46121];
  assign o[46120] = i[46120];
  assign o[46119] = i[46119];
  assign o[46118] = i[46118];
  assign o[46117] = i[46117];
  assign o[46116] = i[46116];
  assign o[46115] = i[46115];
  assign o[46114] = i[46114];
  assign o[46113] = i[46113];
  assign o[46112] = i[46112];
  assign o[46111] = i[46111];
  assign o[46110] = i[46110];
  assign o[46109] = i[46109];
  assign o[46108] = i[46108];
  assign o[46107] = i[46107];
  assign o[46106] = i[46106];
  assign o[46105] = i[46105];
  assign o[46104] = i[46104];
  assign o[46103] = i[46103];
  assign o[46102] = i[46102];
  assign o[46101] = i[46101];
  assign o[46100] = i[46100];
  assign o[46099] = i[46099];
  assign o[46098] = i[46098];
  assign o[46097] = i[46097];
  assign o[46096] = i[46096];
  assign o[46095] = i[46095];
  assign o[46094] = i[46094];
  assign o[46093] = i[46093];
  assign o[46092] = i[46092];
  assign o[46091] = i[46091];
  assign o[46090] = i[46090];
  assign o[46089] = i[46089];
  assign o[46088] = i[46088];
  assign o[46087] = i[46087];
  assign o[46086] = i[46086];
  assign o[46085] = i[46085];
  assign o[46084] = i[46084];
  assign o[46083] = i[46083];
  assign o[46082] = i[46082];
  assign o[46081] = i[46081];
  assign o[46080] = i[46080];
  assign o[46079] = i[46079];
  assign o[46078] = i[46078];
  assign o[46077] = i[46077];
  assign o[46076] = i[46076];
  assign o[46075] = i[46075];
  assign o[46074] = i[46074];
  assign o[46073] = i[46073];
  assign o[46072] = i[46072];
  assign o[46071] = i[46071];
  assign o[46070] = i[46070];
  assign o[46069] = i[46069];
  assign o[46068] = i[46068];
  assign o[46067] = i[46067];
  assign o[46066] = i[46066];
  assign o[46065] = i[46065];
  assign o[46064] = i[46064];
  assign o[46063] = i[46063];
  assign o[46062] = i[46062];
  assign o[46061] = i[46061];
  assign o[46060] = i[46060];
  assign o[46059] = i[46059];
  assign o[46058] = i[46058];
  assign o[46057] = i[46057];
  assign o[46056] = i[46056];
  assign o[46055] = i[46055];
  assign o[46054] = i[46054];
  assign o[46053] = i[46053];
  assign o[46052] = i[46052];
  assign o[46051] = i[46051];
  assign o[46050] = i[46050];
  assign o[46049] = i[46049];
  assign o[46048] = i[46048];
  assign o[46047] = i[46047];
  assign o[46046] = i[46046];
  assign o[46045] = i[46045];
  assign o[46044] = i[46044];
  assign o[46043] = i[46043];
  assign o[46042] = i[46042];
  assign o[46041] = i[46041];
  assign o[46040] = i[46040];
  assign o[46039] = i[46039];
  assign o[46038] = i[46038];
  assign o[46037] = i[46037];
  assign o[46036] = i[46036];
  assign o[46035] = i[46035];
  assign o[46034] = i[46034];
  assign o[46033] = i[46033];
  assign o[46032] = i[46032];
  assign o[46031] = i[46031];
  assign o[46030] = i[46030];
  assign o[46029] = i[46029];
  assign o[46028] = i[46028];
  assign o[46027] = i[46027];
  assign o[46026] = i[46026];
  assign o[46025] = i[46025];
  assign o[46024] = i[46024];
  assign o[46023] = i[46023];
  assign o[46022] = i[46022];
  assign o[46021] = i[46021];
  assign o[46020] = i[46020];
  assign o[46019] = i[46019];
  assign o[46018] = i[46018];
  assign o[46017] = i[46017];
  assign o[46016] = i[46016];
  assign o[46015] = i[46015];
  assign o[46014] = i[46014];
  assign o[46013] = i[46013];
  assign o[46012] = i[46012];
  assign o[46011] = i[46011];
  assign o[46010] = i[46010];
  assign o[46009] = i[46009];
  assign o[46008] = i[46008];
  assign o[46007] = i[46007];
  assign o[46006] = i[46006];
  assign o[46005] = i[46005];
  assign o[46004] = i[46004];
  assign o[46003] = i[46003];
  assign o[46002] = i[46002];
  assign o[46001] = i[46001];
  assign o[46000] = i[46000];
  assign o[45999] = i[45999];
  assign o[45998] = i[45998];
  assign o[45997] = i[45997];
  assign o[45996] = i[45996];
  assign o[45995] = i[45995];
  assign o[45994] = i[45994];
  assign o[45993] = i[45993];
  assign o[45992] = i[45992];
  assign o[45991] = i[45991];
  assign o[45990] = i[45990];
  assign o[45989] = i[45989];
  assign o[45988] = i[45988];
  assign o[45987] = i[45987];
  assign o[45986] = i[45986];
  assign o[45985] = i[45985];
  assign o[45984] = i[45984];
  assign o[45983] = i[45983];
  assign o[45982] = i[45982];
  assign o[45981] = i[45981];
  assign o[45980] = i[45980];
  assign o[45979] = i[45979];
  assign o[45978] = i[45978];
  assign o[45977] = i[45977];
  assign o[45976] = i[45976];
  assign o[45975] = i[45975];
  assign o[45974] = i[45974];
  assign o[45973] = i[45973];
  assign o[45972] = i[45972];
  assign o[45971] = i[45971];
  assign o[45970] = i[45970];
  assign o[45969] = i[45969];
  assign o[45968] = i[45968];
  assign o[45967] = i[45967];
  assign o[45966] = i[45966];
  assign o[45965] = i[45965];
  assign o[45964] = i[45964];
  assign o[45963] = i[45963];
  assign o[45962] = i[45962];
  assign o[45961] = i[45961];
  assign o[45960] = i[45960];
  assign o[45959] = i[45959];
  assign o[45958] = i[45958];
  assign o[45957] = i[45957];
  assign o[45956] = i[45956];
  assign o[45955] = i[45955];
  assign o[45954] = i[45954];
  assign o[45953] = i[45953];
  assign o[45952] = i[45952];
  assign o[45951] = i[45951];
  assign o[45950] = i[45950];
  assign o[45949] = i[45949];
  assign o[45948] = i[45948];
  assign o[45947] = i[45947];
  assign o[45946] = i[45946];
  assign o[45945] = i[45945];
  assign o[45944] = i[45944];
  assign o[45943] = i[45943];
  assign o[45942] = i[45942];
  assign o[45941] = i[45941];
  assign o[45940] = i[45940];
  assign o[45939] = i[45939];
  assign o[45938] = i[45938];
  assign o[45937] = i[45937];
  assign o[45936] = i[45936];
  assign o[45935] = i[45935];
  assign o[45934] = i[45934];
  assign o[45933] = i[45933];
  assign o[45932] = i[45932];
  assign o[45931] = i[45931];
  assign o[45930] = i[45930];
  assign o[45929] = i[45929];
  assign o[45928] = i[45928];
  assign o[45927] = i[45927];
  assign o[45926] = i[45926];
  assign o[45925] = i[45925];
  assign o[45924] = i[45924];
  assign o[45923] = i[45923];
  assign o[45922] = i[45922];
  assign o[45921] = i[45921];
  assign o[45920] = i[45920];
  assign o[45919] = i[45919];
  assign o[45918] = i[45918];
  assign o[45917] = i[45917];
  assign o[45916] = i[45916];
  assign o[45915] = i[45915];
  assign o[45914] = i[45914];
  assign o[45913] = i[45913];
  assign o[45912] = i[45912];
  assign o[45911] = i[45911];
  assign o[45910] = i[45910];
  assign o[45909] = i[45909];
  assign o[45908] = i[45908];
  assign o[45907] = i[45907];
  assign o[45906] = i[45906];
  assign o[45905] = i[45905];
  assign o[45904] = i[45904];
  assign o[45903] = i[45903];
  assign o[45902] = i[45902];
  assign o[45901] = i[45901];
  assign o[45900] = i[45900];
  assign o[45899] = i[45899];
  assign o[45898] = i[45898];
  assign o[45897] = i[45897];
  assign o[45896] = i[45896];
  assign o[45895] = i[45895];
  assign o[45894] = i[45894];
  assign o[45893] = i[45893];
  assign o[45892] = i[45892];
  assign o[45891] = i[45891];
  assign o[45890] = i[45890];
  assign o[45889] = i[45889];
  assign o[45888] = i[45888];
  assign o[45887] = i[45887];
  assign o[45886] = i[45886];
  assign o[45885] = i[45885];
  assign o[45884] = i[45884];
  assign o[45883] = i[45883];
  assign o[45882] = i[45882];
  assign o[45881] = i[45881];
  assign o[45880] = i[45880];
  assign o[45879] = i[45879];
  assign o[45878] = i[45878];
  assign o[45877] = i[45877];
  assign o[45876] = i[45876];
  assign o[45875] = i[45875];
  assign o[45874] = i[45874];
  assign o[45873] = i[45873];
  assign o[45872] = i[45872];
  assign o[45871] = i[45871];
  assign o[45870] = i[45870];
  assign o[45869] = i[45869];
  assign o[45868] = i[45868];
  assign o[45867] = i[45867];
  assign o[45866] = i[45866];
  assign o[45865] = i[45865];
  assign o[45864] = i[45864];
  assign o[45863] = i[45863];
  assign o[45862] = i[45862];
  assign o[45861] = i[45861];
  assign o[45860] = i[45860];
  assign o[45859] = i[45859];
  assign o[45858] = i[45858];
  assign o[45857] = i[45857];
  assign o[45856] = i[45856];
  assign o[45855] = i[45855];
  assign o[45854] = i[45854];
  assign o[45853] = i[45853];
  assign o[45852] = i[45852];
  assign o[45851] = i[45851];
  assign o[45850] = i[45850];
  assign o[45849] = i[45849];
  assign o[45848] = i[45848];
  assign o[45847] = i[45847];
  assign o[45846] = i[45846];
  assign o[45845] = i[45845];
  assign o[45844] = i[45844];
  assign o[45843] = i[45843];
  assign o[45842] = i[45842];
  assign o[45841] = i[45841];
  assign o[45840] = i[45840];
  assign o[45839] = i[45839];
  assign o[45838] = i[45838];
  assign o[45837] = i[45837];
  assign o[45836] = i[45836];
  assign o[45835] = i[45835];
  assign o[45834] = i[45834];
  assign o[45833] = i[45833];
  assign o[45832] = i[45832];
  assign o[45831] = i[45831];
  assign o[45830] = i[45830];
  assign o[45829] = i[45829];
  assign o[45828] = i[45828];
  assign o[45827] = i[45827];
  assign o[45826] = i[45826];
  assign o[45825] = i[45825];
  assign o[45824] = i[45824];
  assign o[45823] = i[45823];
  assign o[45822] = i[45822];
  assign o[45821] = i[45821];
  assign o[45820] = i[45820];
  assign o[45819] = i[45819];
  assign o[45818] = i[45818];
  assign o[45817] = i[45817];
  assign o[45816] = i[45816];
  assign o[45815] = i[45815];
  assign o[45814] = i[45814];
  assign o[45813] = i[45813];
  assign o[45812] = i[45812];
  assign o[45811] = i[45811];
  assign o[45810] = i[45810];
  assign o[45809] = i[45809];
  assign o[45808] = i[45808];
  assign o[45807] = i[45807];
  assign o[45806] = i[45806];
  assign o[45805] = i[45805];
  assign o[45804] = i[45804];
  assign o[45803] = i[45803];
  assign o[45802] = i[45802];
  assign o[45801] = i[45801];
  assign o[45800] = i[45800];
  assign o[45799] = i[45799];
  assign o[45798] = i[45798];
  assign o[45797] = i[45797];
  assign o[45796] = i[45796];
  assign o[45795] = i[45795];
  assign o[45794] = i[45794];
  assign o[45793] = i[45793];
  assign o[45792] = i[45792];
  assign o[45791] = i[45791];
  assign o[45790] = i[45790];
  assign o[45789] = i[45789];
  assign o[45788] = i[45788];
  assign o[45787] = i[45787];
  assign o[45786] = i[45786];
  assign o[45785] = i[45785];
  assign o[45784] = i[45784];
  assign o[45783] = i[45783];
  assign o[45782] = i[45782];
  assign o[45781] = i[45781];
  assign o[45780] = i[45780];
  assign o[45779] = i[45779];
  assign o[45778] = i[45778];
  assign o[45777] = i[45777];
  assign o[45776] = i[45776];
  assign o[45775] = i[45775];
  assign o[45774] = i[45774];
  assign o[45773] = i[45773];
  assign o[45772] = i[45772];
  assign o[45771] = i[45771];
  assign o[45770] = i[45770];
  assign o[45769] = i[45769];
  assign o[45768] = i[45768];
  assign o[45767] = i[45767];
  assign o[45766] = i[45766];
  assign o[45765] = i[45765];
  assign o[45764] = i[45764];
  assign o[45763] = i[45763];
  assign o[45762] = i[45762];
  assign o[45761] = i[45761];
  assign o[45760] = i[45760];
  assign o[45759] = i[45759];
  assign o[45758] = i[45758];
  assign o[45757] = i[45757];
  assign o[45756] = i[45756];
  assign o[45755] = i[45755];
  assign o[45754] = i[45754];
  assign o[45753] = i[45753];
  assign o[45752] = i[45752];
  assign o[45751] = i[45751];
  assign o[45750] = i[45750];
  assign o[45749] = i[45749];
  assign o[45748] = i[45748];
  assign o[45747] = i[45747];
  assign o[45746] = i[45746];
  assign o[45745] = i[45745];
  assign o[45744] = i[45744];
  assign o[45743] = i[45743];
  assign o[45742] = i[45742];
  assign o[45741] = i[45741];
  assign o[45740] = i[45740];
  assign o[45739] = i[45739];
  assign o[45738] = i[45738];
  assign o[45737] = i[45737];
  assign o[45736] = i[45736];
  assign o[45735] = i[45735];
  assign o[45734] = i[45734];
  assign o[45733] = i[45733];
  assign o[45732] = i[45732];
  assign o[45731] = i[45731];
  assign o[45730] = i[45730];
  assign o[45729] = i[45729];
  assign o[45728] = i[45728];
  assign o[45727] = i[45727];
  assign o[45726] = i[45726];
  assign o[45725] = i[45725];
  assign o[45724] = i[45724];
  assign o[45723] = i[45723];
  assign o[45722] = i[45722];
  assign o[45721] = i[45721];
  assign o[45720] = i[45720];
  assign o[45719] = i[45719];
  assign o[45718] = i[45718];
  assign o[45717] = i[45717];
  assign o[45716] = i[45716];
  assign o[45715] = i[45715];
  assign o[45714] = i[45714];
  assign o[45713] = i[45713];
  assign o[45712] = i[45712];
  assign o[45711] = i[45711];
  assign o[45710] = i[45710];
  assign o[45709] = i[45709];
  assign o[45708] = i[45708];
  assign o[45707] = i[45707];
  assign o[45706] = i[45706];
  assign o[45705] = i[45705];
  assign o[45704] = i[45704];
  assign o[45703] = i[45703];
  assign o[45702] = i[45702];
  assign o[45701] = i[45701];
  assign o[45700] = i[45700];
  assign o[45699] = i[45699];
  assign o[45698] = i[45698];
  assign o[45697] = i[45697];
  assign o[45696] = i[45696];
  assign o[45695] = i[45695];
  assign o[45694] = i[45694];
  assign o[45693] = i[45693];
  assign o[45692] = i[45692];
  assign o[45691] = i[45691];
  assign o[45690] = i[45690];
  assign o[45689] = i[45689];
  assign o[45688] = i[45688];
  assign o[45687] = i[45687];
  assign o[45686] = i[45686];
  assign o[45685] = i[45685];
  assign o[45684] = i[45684];
  assign o[45683] = i[45683];
  assign o[45682] = i[45682];
  assign o[45681] = i[45681];
  assign o[45680] = i[45680];
  assign o[45679] = i[45679];
  assign o[45678] = i[45678];
  assign o[45677] = i[45677];
  assign o[45676] = i[45676];
  assign o[45675] = i[45675];
  assign o[45674] = i[45674];
  assign o[45673] = i[45673];
  assign o[45672] = i[45672];
  assign o[45671] = i[45671];
  assign o[45670] = i[45670];
  assign o[45669] = i[45669];
  assign o[45668] = i[45668];
  assign o[45667] = i[45667];
  assign o[45666] = i[45666];
  assign o[45665] = i[45665];
  assign o[45664] = i[45664];
  assign o[45663] = i[45663];
  assign o[45662] = i[45662];
  assign o[45661] = i[45661];
  assign o[45660] = i[45660];
  assign o[45659] = i[45659];
  assign o[45658] = i[45658];
  assign o[45657] = i[45657];
  assign o[45656] = i[45656];
  assign o[45655] = i[45655];
  assign o[45654] = i[45654];
  assign o[45653] = i[45653];
  assign o[45652] = i[45652];
  assign o[45651] = i[45651];
  assign o[45650] = i[45650];
  assign o[45649] = i[45649];
  assign o[45648] = i[45648];
  assign o[45647] = i[45647];
  assign o[45646] = i[45646];
  assign o[45645] = i[45645];
  assign o[45644] = i[45644];
  assign o[45643] = i[45643];
  assign o[45642] = i[45642];
  assign o[45641] = i[45641];
  assign o[45640] = i[45640];
  assign o[45639] = i[45639];
  assign o[45638] = i[45638];
  assign o[45637] = i[45637];
  assign o[45636] = i[45636];
  assign o[45635] = i[45635];
  assign o[45634] = i[45634];
  assign o[45633] = i[45633];
  assign o[45632] = i[45632];
  assign o[45631] = i[45631];
  assign o[45630] = i[45630];
  assign o[45629] = i[45629];
  assign o[45628] = i[45628];
  assign o[45627] = i[45627];
  assign o[45626] = i[45626];
  assign o[45625] = i[45625];
  assign o[45624] = i[45624];
  assign o[45623] = i[45623];
  assign o[45622] = i[45622];
  assign o[45621] = i[45621];
  assign o[45620] = i[45620];
  assign o[45619] = i[45619];
  assign o[45618] = i[45618];
  assign o[45617] = i[45617];
  assign o[45616] = i[45616];
  assign o[45615] = i[45615];
  assign o[45614] = i[45614];
  assign o[45613] = i[45613];
  assign o[45612] = i[45612];
  assign o[45611] = i[45611];
  assign o[45610] = i[45610];
  assign o[45609] = i[45609];
  assign o[45608] = i[45608];
  assign o[45607] = i[45607];
  assign o[45606] = i[45606];
  assign o[45605] = i[45605];
  assign o[45604] = i[45604];
  assign o[45603] = i[45603];
  assign o[45602] = i[45602];
  assign o[45601] = i[45601];
  assign o[45600] = i[45600];
  assign o[45599] = i[45599];
  assign o[45598] = i[45598];
  assign o[45597] = i[45597];
  assign o[45596] = i[45596];
  assign o[45595] = i[45595];
  assign o[45594] = i[45594];
  assign o[45593] = i[45593];
  assign o[45592] = i[45592];
  assign o[45591] = i[45591];
  assign o[45590] = i[45590];
  assign o[45589] = i[45589];
  assign o[45588] = i[45588];
  assign o[45587] = i[45587];
  assign o[45586] = i[45586];
  assign o[45585] = i[45585];
  assign o[45584] = i[45584];
  assign o[45583] = i[45583];
  assign o[45582] = i[45582];
  assign o[45581] = i[45581];
  assign o[45580] = i[45580];
  assign o[45579] = i[45579];
  assign o[45578] = i[45578];
  assign o[45577] = i[45577];
  assign o[45576] = i[45576];
  assign o[45575] = i[45575];
  assign o[45574] = i[45574];
  assign o[45573] = i[45573];
  assign o[45572] = i[45572];
  assign o[45571] = i[45571];
  assign o[45570] = i[45570];
  assign o[45569] = i[45569];
  assign o[45568] = i[45568];
  assign o[45567] = i[45567];
  assign o[45566] = i[45566];
  assign o[45565] = i[45565];
  assign o[45564] = i[45564];
  assign o[45563] = i[45563];
  assign o[45562] = i[45562];
  assign o[45561] = i[45561];
  assign o[45560] = i[45560];
  assign o[45559] = i[45559];
  assign o[45558] = i[45558];
  assign o[45557] = i[45557];
  assign o[45556] = i[45556];
  assign o[45555] = i[45555];
  assign o[45554] = i[45554];
  assign o[45553] = i[45553];
  assign o[45552] = i[45552];
  assign o[45551] = i[45551];
  assign o[45550] = i[45550];
  assign o[45549] = i[45549];
  assign o[45548] = i[45548];
  assign o[45547] = i[45547];
  assign o[45546] = i[45546];
  assign o[45545] = i[45545];
  assign o[45544] = i[45544];
  assign o[45543] = i[45543];
  assign o[45542] = i[45542];
  assign o[45541] = i[45541];
  assign o[45540] = i[45540];
  assign o[45539] = i[45539];
  assign o[45538] = i[45538];
  assign o[45537] = i[45537];
  assign o[45536] = i[45536];
  assign o[45535] = i[45535];
  assign o[45534] = i[45534];
  assign o[45533] = i[45533];
  assign o[45532] = i[45532];
  assign o[45531] = i[45531];
  assign o[45530] = i[45530];
  assign o[45529] = i[45529];
  assign o[45528] = i[45528];
  assign o[45527] = i[45527];
  assign o[45526] = i[45526];
  assign o[45525] = i[45525];
  assign o[45524] = i[45524];
  assign o[45523] = i[45523];
  assign o[45522] = i[45522];
  assign o[45521] = i[45521];
  assign o[45520] = i[45520];
  assign o[45519] = i[45519];
  assign o[45518] = i[45518];
  assign o[45517] = i[45517];
  assign o[45516] = i[45516];
  assign o[45515] = i[45515];
  assign o[45514] = i[45514];
  assign o[45513] = i[45513];
  assign o[45512] = i[45512];
  assign o[45511] = i[45511];
  assign o[45510] = i[45510];
  assign o[45509] = i[45509];
  assign o[45508] = i[45508];
  assign o[45507] = i[45507];
  assign o[45506] = i[45506];
  assign o[45505] = i[45505];
  assign o[45504] = i[45504];
  assign o[45503] = i[45503];
  assign o[45502] = i[45502];
  assign o[45501] = i[45501];
  assign o[45500] = i[45500];
  assign o[45499] = i[45499];
  assign o[45498] = i[45498];
  assign o[45497] = i[45497];
  assign o[45496] = i[45496];
  assign o[45495] = i[45495];
  assign o[45494] = i[45494];
  assign o[45493] = i[45493];
  assign o[45492] = i[45492];
  assign o[45491] = i[45491];
  assign o[45490] = i[45490];
  assign o[45489] = i[45489];
  assign o[45488] = i[45488];
  assign o[45487] = i[45487];
  assign o[45486] = i[45486];
  assign o[45485] = i[45485];
  assign o[45484] = i[45484];
  assign o[45483] = i[45483];
  assign o[45482] = i[45482];
  assign o[45481] = i[45481];
  assign o[45480] = i[45480];
  assign o[45479] = i[45479];
  assign o[45478] = i[45478];
  assign o[45477] = i[45477];
  assign o[45476] = i[45476];
  assign o[45475] = i[45475];
  assign o[45474] = i[45474];
  assign o[45473] = i[45473];
  assign o[45472] = i[45472];
  assign o[45471] = i[45471];
  assign o[45470] = i[45470];
  assign o[45469] = i[45469];
  assign o[45468] = i[45468];
  assign o[45467] = i[45467];
  assign o[45466] = i[45466];
  assign o[45465] = i[45465];
  assign o[45464] = i[45464];
  assign o[45463] = i[45463];
  assign o[45462] = i[45462];
  assign o[45461] = i[45461];
  assign o[45460] = i[45460];
  assign o[45459] = i[45459];
  assign o[45458] = i[45458];
  assign o[45457] = i[45457];
  assign o[45456] = i[45456];
  assign o[45455] = i[45455];
  assign o[45454] = i[45454];
  assign o[45453] = i[45453];
  assign o[45452] = i[45452];
  assign o[45451] = i[45451];
  assign o[45450] = i[45450];
  assign o[45449] = i[45449];
  assign o[45448] = i[45448];
  assign o[45447] = i[45447];
  assign o[45446] = i[45446];
  assign o[45445] = i[45445];
  assign o[45444] = i[45444];
  assign o[45443] = i[45443];
  assign o[45442] = i[45442];
  assign o[45441] = i[45441];
  assign o[45440] = i[45440];
  assign o[45439] = i[45439];
  assign o[45438] = i[45438];
  assign o[45437] = i[45437];
  assign o[45436] = i[45436];
  assign o[45435] = i[45435];
  assign o[45434] = i[45434];
  assign o[45433] = i[45433];
  assign o[45432] = i[45432];
  assign o[45431] = i[45431];
  assign o[45430] = i[45430];
  assign o[45429] = i[45429];
  assign o[45428] = i[45428];
  assign o[45427] = i[45427];
  assign o[45426] = i[45426];
  assign o[45425] = i[45425];
  assign o[45424] = i[45424];
  assign o[45423] = i[45423];
  assign o[45422] = i[45422];
  assign o[45421] = i[45421];
  assign o[45420] = i[45420];
  assign o[45419] = i[45419];
  assign o[45418] = i[45418];
  assign o[45417] = i[45417];
  assign o[45416] = i[45416];
  assign o[45415] = i[45415];
  assign o[45414] = i[45414];
  assign o[45413] = i[45413];
  assign o[45412] = i[45412];
  assign o[45411] = i[45411];
  assign o[45410] = i[45410];
  assign o[45409] = i[45409];
  assign o[45408] = i[45408];
  assign o[45407] = i[45407];
  assign o[45406] = i[45406];
  assign o[45405] = i[45405];
  assign o[45404] = i[45404];
  assign o[45403] = i[45403];
  assign o[45402] = i[45402];
  assign o[45401] = i[45401];
  assign o[45400] = i[45400];
  assign o[45399] = i[45399];
  assign o[45398] = i[45398];
  assign o[45397] = i[45397];
  assign o[45396] = i[45396];
  assign o[45395] = i[45395];
  assign o[45394] = i[45394];
  assign o[45393] = i[45393];
  assign o[45392] = i[45392];
  assign o[45391] = i[45391];
  assign o[45390] = i[45390];
  assign o[45389] = i[45389];
  assign o[45388] = i[45388];
  assign o[45387] = i[45387];
  assign o[45386] = i[45386];
  assign o[45385] = i[45385];
  assign o[45384] = i[45384];
  assign o[45383] = i[45383];
  assign o[45382] = i[45382];
  assign o[45381] = i[45381];
  assign o[45380] = i[45380];
  assign o[45379] = i[45379];
  assign o[45378] = i[45378];
  assign o[45377] = i[45377];
  assign o[45376] = i[45376];
  assign o[45375] = i[45375];
  assign o[45374] = i[45374];
  assign o[45373] = i[45373];
  assign o[45372] = i[45372];
  assign o[45371] = i[45371];
  assign o[45370] = i[45370];
  assign o[45369] = i[45369];
  assign o[45368] = i[45368];
  assign o[45367] = i[45367];
  assign o[45366] = i[45366];
  assign o[45365] = i[45365];
  assign o[45364] = i[45364];
  assign o[45363] = i[45363];
  assign o[45362] = i[45362];
  assign o[45361] = i[45361];
  assign o[45360] = i[45360];
  assign o[45359] = i[45359];
  assign o[45358] = i[45358];
  assign o[45357] = i[45357];
  assign o[45356] = i[45356];
  assign o[45355] = i[45355];
  assign o[45354] = i[45354];
  assign o[45353] = i[45353];
  assign o[45352] = i[45352];
  assign o[45351] = i[45351];
  assign o[45350] = i[45350];
  assign o[45349] = i[45349];
  assign o[45348] = i[45348];
  assign o[45347] = i[45347];
  assign o[45346] = i[45346];
  assign o[45345] = i[45345];
  assign o[45344] = i[45344];
  assign o[45343] = i[45343];
  assign o[45342] = i[45342];
  assign o[45341] = i[45341];
  assign o[45340] = i[45340];
  assign o[45339] = i[45339];
  assign o[45338] = i[45338];
  assign o[45337] = i[45337];
  assign o[45336] = i[45336];
  assign o[45335] = i[45335];
  assign o[45334] = i[45334];
  assign o[45333] = i[45333];
  assign o[45332] = i[45332];
  assign o[45331] = i[45331];
  assign o[45330] = i[45330];
  assign o[45329] = i[45329];
  assign o[45328] = i[45328];
  assign o[45327] = i[45327];
  assign o[45326] = i[45326];
  assign o[45325] = i[45325];
  assign o[45324] = i[45324];
  assign o[45323] = i[45323];
  assign o[45322] = i[45322];
  assign o[45321] = i[45321];
  assign o[45320] = i[45320];
  assign o[45319] = i[45319];
  assign o[45318] = i[45318];
  assign o[45317] = i[45317];
  assign o[45316] = i[45316];
  assign o[45315] = i[45315];
  assign o[45314] = i[45314];
  assign o[45313] = i[45313];
  assign o[45312] = i[45312];
  assign o[45311] = i[45311];
  assign o[45310] = i[45310];
  assign o[45309] = i[45309];
  assign o[45308] = i[45308];
  assign o[45307] = i[45307];
  assign o[45306] = i[45306];
  assign o[45305] = i[45305];
  assign o[45304] = i[45304];
  assign o[45303] = i[45303];
  assign o[45302] = i[45302];
  assign o[45301] = i[45301];
  assign o[45300] = i[45300];
  assign o[45299] = i[45299];
  assign o[45298] = i[45298];
  assign o[45297] = i[45297];
  assign o[45296] = i[45296];
  assign o[45295] = i[45295];
  assign o[45294] = i[45294];
  assign o[45293] = i[45293];
  assign o[45292] = i[45292];
  assign o[45291] = i[45291];
  assign o[45290] = i[45290];
  assign o[45289] = i[45289];
  assign o[45288] = i[45288];
  assign o[45287] = i[45287];
  assign o[45286] = i[45286];
  assign o[45285] = i[45285];
  assign o[45284] = i[45284];
  assign o[45283] = i[45283];
  assign o[45282] = i[45282];
  assign o[45281] = i[45281];
  assign o[45280] = i[45280];
  assign o[45279] = i[45279];
  assign o[45278] = i[45278];
  assign o[45277] = i[45277];
  assign o[45276] = i[45276];
  assign o[45275] = i[45275];
  assign o[45274] = i[45274];
  assign o[45273] = i[45273];
  assign o[45272] = i[45272];
  assign o[45271] = i[45271];
  assign o[45270] = i[45270];
  assign o[45269] = i[45269];
  assign o[45268] = i[45268];
  assign o[45267] = i[45267];
  assign o[45266] = i[45266];
  assign o[45265] = i[45265];
  assign o[45264] = i[45264];
  assign o[45263] = i[45263];
  assign o[45262] = i[45262];
  assign o[45261] = i[45261];
  assign o[45260] = i[45260];
  assign o[45259] = i[45259];
  assign o[45258] = i[45258];
  assign o[45257] = i[45257];
  assign o[45256] = i[45256];
  assign o[45255] = i[45255];
  assign o[45254] = i[45254];
  assign o[45253] = i[45253];
  assign o[45252] = i[45252];
  assign o[45251] = i[45251];
  assign o[45250] = i[45250];
  assign o[45249] = i[45249];
  assign o[45248] = i[45248];
  assign o[45247] = i[45247];
  assign o[45246] = i[45246];
  assign o[45245] = i[45245];
  assign o[45244] = i[45244];
  assign o[45243] = i[45243];
  assign o[45242] = i[45242];
  assign o[45241] = i[45241];
  assign o[45240] = i[45240];
  assign o[45239] = i[45239];
  assign o[45238] = i[45238];
  assign o[45237] = i[45237];
  assign o[45236] = i[45236];
  assign o[45235] = i[45235];
  assign o[45234] = i[45234];
  assign o[45233] = i[45233];
  assign o[45232] = i[45232];
  assign o[45231] = i[45231];
  assign o[45230] = i[45230];
  assign o[45229] = i[45229];
  assign o[45228] = i[45228];
  assign o[45227] = i[45227];
  assign o[45226] = i[45226];
  assign o[45225] = i[45225];
  assign o[45224] = i[45224];
  assign o[45223] = i[45223];
  assign o[45222] = i[45222];
  assign o[45221] = i[45221];
  assign o[45220] = i[45220];
  assign o[45219] = i[45219];
  assign o[45218] = i[45218];
  assign o[45217] = i[45217];
  assign o[45216] = i[45216];
  assign o[45215] = i[45215];
  assign o[45214] = i[45214];
  assign o[45213] = i[45213];
  assign o[45212] = i[45212];
  assign o[45211] = i[45211];
  assign o[45210] = i[45210];
  assign o[45209] = i[45209];
  assign o[45208] = i[45208];
  assign o[45207] = i[45207];
  assign o[45206] = i[45206];
  assign o[45205] = i[45205];
  assign o[45204] = i[45204];
  assign o[45203] = i[45203];
  assign o[45202] = i[45202];
  assign o[45201] = i[45201];
  assign o[45200] = i[45200];
  assign o[45199] = i[45199];
  assign o[45198] = i[45198];
  assign o[45197] = i[45197];
  assign o[45196] = i[45196];
  assign o[45195] = i[45195];
  assign o[45194] = i[45194];
  assign o[45193] = i[45193];
  assign o[45192] = i[45192];
  assign o[45191] = i[45191];
  assign o[45190] = i[45190];
  assign o[45189] = i[45189];
  assign o[45188] = i[45188];
  assign o[45187] = i[45187];
  assign o[45186] = i[45186];
  assign o[45185] = i[45185];
  assign o[45184] = i[45184];
  assign o[45183] = i[45183];
  assign o[45182] = i[45182];
  assign o[45181] = i[45181];
  assign o[45180] = i[45180];
  assign o[45179] = i[45179];
  assign o[45178] = i[45178];
  assign o[45177] = i[45177];
  assign o[45176] = i[45176];
  assign o[45175] = i[45175];
  assign o[45174] = i[45174];
  assign o[45173] = i[45173];
  assign o[45172] = i[45172];
  assign o[45171] = i[45171];
  assign o[45170] = i[45170];
  assign o[45169] = i[45169];
  assign o[45168] = i[45168];
  assign o[45167] = i[45167];
  assign o[45166] = i[45166];
  assign o[45165] = i[45165];
  assign o[45164] = i[45164];
  assign o[45163] = i[45163];
  assign o[45162] = i[45162];
  assign o[45161] = i[45161];
  assign o[45160] = i[45160];
  assign o[45159] = i[45159];
  assign o[45158] = i[45158];
  assign o[45157] = i[45157];
  assign o[45156] = i[45156];
  assign o[45155] = i[45155];
  assign o[45154] = i[45154];
  assign o[45153] = i[45153];
  assign o[45152] = i[45152];
  assign o[45151] = i[45151];
  assign o[45150] = i[45150];
  assign o[45149] = i[45149];
  assign o[45148] = i[45148];
  assign o[45147] = i[45147];
  assign o[45146] = i[45146];
  assign o[45145] = i[45145];
  assign o[45144] = i[45144];
  assign o[45143] = i[45143];
  assign o[45142] = i[45142];
  assign o[45141] = i[45141];
  assign o[45140] = i[45140];
  assign o[45139] = i[45139];
  assign o[45138] = i[45138];
  assign o[45137] = i[45137];
  assign o[45136] = i[45136];
  assign o[45135] = i[45135];
  assign o[45134] = i[45134];
  assign o[45133] = i[45133];
  assign o[45132] = i[45132];
  assign o[45131] = i[45131];
  assign o[45130] = i[45130];
  assign o[45129] = i[45129];
  assign o[45128] = i[45128];
  assign o[45127] = i[45127];
  assign o[45126] = i[45126];
  assign o[45125] = i[45125];
  assign o[45124] = i[45124];
  assign o[45123] = i[45123];
  assign o[45122] = i[45122];
  assign o[45121] = i[45121];
  assign o[45120] = i[45120];
  assign o[45119] = i[45119];
  assign o[45118] = i[45118];
  assign o[45117] = i[45117];
  assign o[45116] = i[45116];
  assign o[45115] = i[45115];
  assign o[45114] = i[45114];
  assign o[45113] = i[45113];
  assign o[45112] = i[45112];
  assign o[45111] = i[45111];
  assign o[45110] = i[45110];
  assign o[45109] = i[45109];
  assign o[45108] = i[45108];
  assign o[45107] = i[45107];
  assign o[45106] = i[45106];
  assign o[45105] = i[45105];
  assign o[45104] = i[45104];
  assign o[45103] = i[45103];
  assign o[45102] = i[45102];
  assign o[45101] = i[45101];
  assign o[45100] = i[45100];
  assign o[45099] = i[45099];
  assign o[45098] = i[45098];
  assign o[45097] = i[45097];
  assign o[45096] = i[45096];
  assign o[45095] = i[45095];
  assign o[45094] = i[45094];
  assign o[45093] = i[45093];
  assign o[45092] = i[45092];
  assign o[45091] = i[45091];
  assign o[45090] = i[45090];
  assign o[45089] = i[45089];
  assign o[45088] = i[45088];
  assign o[45087] = i[45087];
  assign o[45086] = i[45086];
  assign o[45085] = i[45085];
  assign o[45084] = i[45084];
  assign o[45083] = i[45083];
  assign o[45082] = i[45082];
  assign o[45081] = i[45081];
  assign o[45080] = i[45080];
  assign o[45079] = i[45079];
  assign o[45078] = i[45078];
  assign o[45077] = i[45077];
  assign o[45076] = i[45076];
  assign o[45075] = i[45075];
  assign o[45074] = i[45074];
  assign o[45073] = i[45073];
  assign o[45072] = i[45072];
  assign o[45071] = i[45071];
  assign o[45070] = i[45070];
  assign o[45069] = i[45069];
  assign o[45068] = i[45068];
  assign o[45067] = i[45067];
  assign o[45066] = i[45066];
  assign o[45065] = i[45065];
  assign o[45064] = i[45064];
  assign o[45063] = i[45063];
  assign o[45062] = i[45062];
  assign o[45061] = i[45061];
  assign o[45060] = i[45060];
  assign o[45059] = i[45059];
  assign o[45058] = i[45058];
  assign o[45057] = i[45057];
  assign o[45056] = i[45056];
  assign o[45055] = i[45055];
  assign o[45054] = i[45054];
  assign o[45053] = i[45053];
  assign o[45052] = i[45052];
  assign o[45051] = i[45051];
  assign o[45050] = i[45050];
  assign o[45049] = i[45049];
  assign o[45048] = i[45048];
  assign o[45047] = i[45047];
  assign o[45046] = i[45046];
  assign o[45045] = i[45045];
  assign o[45044] = i[45044];
  assign o[45043] = i[45043];
  assign o[45042] = i[45042];
  assign o[45041] = i[45041];
  assign o[45040] = i[45040];
  assign o[45039] = i[45039];
  assign o[45038] = i[45038];
  assign o[45037] = i[45037];
  assign o[45036] = i[45036];
  assign o[45035] = i[45035];
  assign o[45034] = i[45034];
  assign o[45033] = i[45033];
  assign o[45032] = i[45032];
  assign o[45031] = i[45031];
  assign o[45030] = i[45030];
  assign o[45029] = i[45029];
  assign o[45028] = i[45028];
  assign o[45027] = i[45027];
  assign o[45026] = i[45026];
  assign o[45025] = i[45025];
  assign o[45024] = i[45024];
  assign o[45023] = i[45023];
  assign o[45022] = i[45022];
  assign o[45021] = i[45021];
  assign o[45020] = i[45020];
  assign o[45019] = i[45019];
  assign o[45018] = i[45018];
  assign o[45017] = i[45017];
  assign o[45016] = i[45016];
  assign o[45015] = i[45015];
  assign o[45014] = i[45014];
  assign o[45013] = i[45013];
  assign o[45012] = i[45012];
  assign o[45011] = i[45011];
  assign o[45010] = i[45010];
  assign o[45009] = i[45009];
  assign o[45008] = i[45008];
  assign o[45007] = i[45007];
  assign o[45006] = i[45006];
  assign o[45005] = i[45005];
  assign o[45004] = i[45004];
  assign o[45003] = i[45003];
  assign o[45002] = i[45002];
  assign o[45001] = i[45001];
  assign o[45000] = i[45000];
  assign o[44999] = i[44999];
  assign o[44998] = i[44998];
  assign o[44997] = i[44997];
  assign o[44996] = i[44996];
  assign o[44995] = i[44995];
  assign o[44994] = i[44994];
  assign o[44993] = i[44993];
  assign o[44992] = i[44992];
  assign o[44991] = i[44991];
  assign o[44990] = i[44990];
  assign o[44989] = i[44989];
  assign o[44988] = i[44988];
  assign o[44987] = i[44987];
  assign o[44986] = i[44986];
  assign o[44985] = i[44985];
  assign o[44984] = i[44984];
  assign o[44983] = i[44983];
  assign o[44982] = i[44982];
  assign o[44981] = i[44981];
  assign o[44980] = i[44980];
  assign o[44979] = i[44979];
  assign o[44978] = i[44978];
  assign o[44977] = i[44977];
  assign o[44976] = i[44976];
  assign o[44975] = i[44975];
  assign o[44974] = i[44974];
  assign o[44973] = i[44973];
  assign o[44972] = i[44972];
  assign o[44971] = i[44971];
  assign o[44970] = i[44970];
  assign o[44969] = i[44969];
  assign o[44968] = i[44968];
  assign o[44967] = i[44967];
  assign o[44966] = i[44966];
  assign o[44965] = i[44965];
  assign o[44964] = i[44964];
  assign o[44963] = i[44963];
  assign o[44962] = i[44962];
  assign o[44961] = i[44961];
  assign o[44960] = i[44960];
  assign o[44959] = i[44959];
  assign o[44958] = i[44958];
  assign o[44957] = i[44957];
  assign o[44956] = i[44956];
  assign o[44955] = i[44955];
  assign o[44954] = i[44954];
  assign o[44953] = i[44953];
  assign o[44952] = i[44952];
  assign o[44951] = i[44951];
  assign o[44950] = i[44950];
  assign o[44949] = i[44949];
  assign o[44948] = i[44948];
  assign o[44947] = i[44947];
  assign o[44946] = i[44946];
  assign o[44945] = i[44945];
  assign o[44944] = i[44944];
  assign o[44943] = i[44943];
  assign o[44942] = i[44942];
  assign o[44941] = i[44941];
  assign o[44940] = i[44940];
  assign o[44939] = i[44939];
  assign o[44938] = i[44938];
  assign o[44937] = i[44937];
  assign o[44936] = i[44936];
  assign o[44935] = i[44935];
  assign o[44934] = i[44934];
  assign o[44933] = i[44933];
  assign o[44932] = i[44932];
  assign o[44931] = i[44931];
  assign o[44930] = i[44930];
  assign o[44929] = i[44929];
  assign o[44928] = i[44928];
  assign o[44927] = i[44927];
  assign o[44926] = i[44926];
  assign o[44925] = i[44925];
  assign o[44924] = i[44924];
  assign o[44923] = i[44923];
  assign o[44922] = i[44922];
  assign o[44921] = i[44921];
  assign o[44920] = i[44920];
  assign o[44919] = i[44919];
  assign o[44918] = i[44918];
  assign o[44917] = i[44917];
  assign o[44916] = i[44916];
  assign o[44915] = i[44915];
  assign o[44914] = i[44914];
  assign o[44913] = i[44913];
  assign o[44912] = i[44912];
  assign o[44911] = i[44911];
  assign o[44910] = i[44910];
  assign o[44909] = i[44909];
  assign o[44908] = i[44908];
  assign o[44907] = i[44907];
  assign o[44906] = i[44906];
  assign o[44905] = i[44905];
  assign o[44904] = i[44904];
  assign o[44903] = i[44903];
  assign o[44902] = i[44902];
  assign o[44901] = i[44901];
  assign o[44900] = i[44900];
  assign o[44899] = i[44899];
  assign o[44898] = i[44898];
  assign o[44897] = i[44897];
  assign o[44896] = i[44896];
  assign o[44895] = i[44895];
  assign o[44894] = i[44894];
  assign o[44893] = i[44893];
  assign o[44892] = i[44892];
  assign o[44891] = i[44891];
  assign o[44890] = i[44890];
  assign o[44889] = i[44889];
  assign o[44888] = i[44888];
  assign o[44887] = i[44887];
  assign o[44886] = i[44886];
  assign o[44885] = i[44885];
  assign o[44884] = i[44884];
  assign o[44883] = i[44883];
  assign o[44882] = i[44882];
  assign o[44881] = i[44881];
  assign o[44880] = i[44880];
  assign o[44879] = i[44879];
  assign o[44878] = i[44878];
  assign o[44877] = i[44877];
  assign o[44876] = i[44876];
  assign o[44875] = i[44875];
  assign o[44874] = i[44874];
  assign o[44873] = i[44873];
  assign o[44872] = i[44872];
  assign o[44871] = i[44871];
  assign o[44870] = i[44870];
  assign o[44869] = i[44869];
  assign o[44868] = i[44868];
  assign o[44867] = i[44867];
  assign o[44866] = i[44866];
  assign o[44865] = i[44865];
  assign o[44864] = i[44864];
  assign o[44863] = i[44863];
  assign o[44862] = i[44862];
  assign o[44861] = i[44861];
  assign o[44860] = i[44860];
  assign o[44859] = i[44859];
  assign o[44858] = i[44858];
  assign o[44857] = i[44857];
  assign o[44856] = i[44856];
  assign o[44855] = i[44855];
  assign o[44854] = i[44854];
  assign o[44853] = i[44853];
  assign o[44852] = i[44852];
  assign o[44851] = i[44851];
  assign o[44850] = i[44850];
  assign o[44849] = i[44849];
  assign o[44848] = i[44848];
  assign o[44847] = i[44847];
  assign o[44846] = i[44846];
  assign o[44845] = i[44845];
  assign o[44844] = i[44844];
  assign o[44843] = i[44843];
  assign o[44842] = i[44842];
  assign o[44841] = i[44841];
  assign o[44840] = i[44840];
  assign o[44839] = i[44839];
  assign o[44838] = i[44838];
  assign o[44837] = i[44837];
  assign o[44836] = i[44836];
  assign o[44835] = i[44835];
  assign o[44834] = i[44834];
  assign o[44833] = i[44833];
  assign o[44832] = i[44832];
  assign o[44831] = i[44831];
  assign o[44830] = i[44830];
  assign o[44829] = i[44829];
  assign o[44828] = i[44828];
  assign o[44827] = i[44827];
  assign o[44826] = i[44826];
  assign o[44825] = i[44825];
  assign o[44824] = i[44824];
  assign o[44823] = i[44823];
  assign o[44822] = i[44822];
  assign o[44821] = i[44821];
  assign o[44820] = i[44820];
  assign o[44819] = i[44819];
  assign o[44818] = i[44818];
  assign o[44817] = i[44817];
  assign o[44816] = i[44816];
  assign o[44815] = i[44815];
  assign o[44814] = i[44814];
  assign o[44813] = i[44813];
  assign o[44812] = i[44812];
  assign o[44811] = i[44811];
  assign o[44810] = i[44810];
  assign o[44809] = i[44809];
  assign o[44808] = i[44808];
  assign o[44807] = i[44807];
  assign o[44806] = i[44806];
  assign o[44805] = i[44805];
  assign o[44804] = i[44804];
  assign o[44803] = i[44803];
  assign o[44802] = i[44802];
  assign o[44801] = i[44801];
  assign o[44800] = i[44800];
  assign o[44799] = i[44799];
  assign o[44798] = i[44798];
  assign o[44797] = i[44797];
  assign o[44796] = i[44796];
  assign o[44795] = i[44795];
  assign o[44794] = i[44794];
  assign o[44793] = i[44793];
  assign o[44792] = i[44792];
  assign o[44791] = i[44791];
  assign o[44790] = i[44790];
  assign o[44789] = i[44789];
  assign o[44788] = i[44788];
  assign o[44787] = i[44787];
  assign o[44786] = i[44786];
  assign o[44785] = i[44785];
  assign o[44784] = i[44784];
  assign o[44783] = i[44783];
  assign o[44782] = i[44782];
  assign o[44781] = i[44781];
  assign o[44780] = i[44780];
  assign o[44779] = i[44779];
  assign o[44778] = i[44778];
  assign o[44777] = i[44777];
  assign o[44776] = i[44776];
  assign o[44775] = i[44775];
  assign o[44774] = i[44774];
  assign o[44773] = i[44773];
  assign o[44772] = i[44772];
  assign o[44771] = i[44771];
  assign o[44770] = i[44770];
  assign o[44769] = i[44769];
  assign o[44768] = i[44768];
  assign o[44767] = i[44767];
  assign o[44766] = i[44766];
  assign o[44765] = i[44765];
  assign o[44764] = i[44764];
  assign o[44763] = i[44763];
  assign o[44762] = i[44762];
  assign o[44761] = i[44761];
  assign o[44760] = i[44760];
  assign o[44759] = i[44759];
  assign o[44758] = i[44758];
  assign o[44757] = i[44757];
  assign o[44756] = i[44756];
  assign o[44755] = i[44755];
  assign o[44754] = i[44754];
  assign o[44753] = i[44753];
  assign o[44752] = i[44752];
  assign o[44751] = i[44751];
  assign o[44750] = i[44750];
  assign o[44749] = i[44749];
  assign o[44748] = i[44748];
  assign o[44747] = i[44747];
  assign o[44746] = i[44746];
  assign o[44745] = i[44745];
  assign o[44744] = i[44744];
  assign o[44743] = i[44743];
  assign o[44742] = i[44742];
  assign o[44741] = i[44741];
  assign o[44740] = i[44740];
  assign o[44739] = i[44739];
  assign o[44738] = i[44738];
  assign o[44737] = i[44737];
  assign o[44736] = i[44736];
  assign o[44735] = i[44735];
  assign o[44734] = i[44734];
  assign o[44733] = i[44733];
  assign o[44732] = i[44732];
  assign o[44731] = i[44731];
  assign o[44730] = i[44730];
  assign o[44729] = i[44729];
  assign o[44728] = i[44728];
  assign o[44727] = i[44727];
  assign o[44726] = i[44726];
  assign o[44725] = i[44725];
  assign o[44724] = i[44724];
  assign o[44723] = i[44723];
  assign o[44722] = i[44722];
  assign o[44721] = i[44721];
  assign o[44720] = i[44720];
  assign o[44719] = i[44719];
  assign o[44718] = i[44718];
  assign o[44717] = i[44717];
  assign o[44716] = i[44716];
  assign o[44715] = i[44715];
  assign o[44714] = i[44714];
  assign o[44713] = i[44713];
  assign o[44712] = i[44712];
  assign o[44711] = i[44711];
  assign o[44710] = i[44710];
  assign o[44709] = i[44709];
  assign o[44708] = i[44708];
  assign o[44707] = i[44707];
  assign o[44706] = i[44706];
  assign o[44705] = i[44705];
  assign o[44704] = i[44704];
  assign o[44703] = i[44703];
  assign o[44702] = i[44702];
  assign o[44701] = i[44701];
  assign o[44700] = i[44700];
  assign o[44699] = i[44699];
  assign o[44698] = i[44698];
  assign o[44697] = i[44697];
  assign o[44696] = i[44696];
  assign o[44695] = i[44695];
  assign o[44694] = i[44694];
  assign o[44693] = i[44693];
  assign o[44692] = i[44692];
  assign o[44691] = i[44691];
  assign o[44690] = i[44690];
  assign o[44689] = i[44689];
  assign o[44688] = i[44688];
  assign o[44687] = i[44687];
  assign o[44686] = i[44686];
  assign o[44685] = i[44685];
  assign o[44684] = i[44684];
  assign o[44683] = i[44683];
  assign o[44682] = i[44682];
  assign o[44681] = i[44681];
  assign o[44680] = i[44680];
  assign o[44679] = i[44679];
  assign o[44678] = i[44678];
  assign o[44677] = i[44677];
  assign o[44676] = i[44676];
  assign o[44675] = i[44675];
  assign o[44674] = i[44674];
  assign o[44673] = i[44673];
  assign o[44672] = i[44672];
  assign o[44671] = i[44671];
  assign o[44670] = i[44670];
  assign o[44669] = i[44669];
  assign o[44668] = i[44668];
  assign o[44667] = i[44667];
  assign o[44666] = i[44666];
  assign o[44665] = i[44665];
  assign o[44664] = i[44664];
  assign o[44663] = i[44663];
  assign o[44662] = i[44662];
  assign o[44661] = i[44661];
  assign o[44660] = i[44660];
  assign o[44659] = i[44659];
  assign o[44658] = i[44658];
  assign o[44657] = i[44657];
  assign o[44656] = i[44656];
  assign o[44655] = i[44655];
  assign o[44654] = i[44654];
  assign o[44653] = i[44653];
  assign o[44652] = i[44652];
  assign o[44651] = i[44651];
  assign o[44650] = i[44650];
  assign o[44649] = i[44649];
  assign o[44648] = i[44648];
  assign o[44647] = i[44647];
  assign o[44646] = i[44646];
  assign o[44645] = i[44645];
  assign o[44644] = i[44644];
  assign o[44643] = i[44643];
  assign o[44642] = i[44642];
  assign o[44641] = i[44641];
  assign o[44640] = i[44640];
  assign o[44639] = i[44639];
  assign o[44638] = i[44638];
  assign o[44637] = i[44637];
  assign o[44636] = i[44636];
  assign o[44635] = i[44635];
  assign o[44634] = i[44634];
  assign o[44633] = i[44633];
  assign o[44632] = i[44632];
  assign o[44631] = i[44631];
  assign o[44630] = i[44630];
  assign o[44629] = i[44629];
  assign o[44628] = i[44628];
  assign o[44627] = i[44627];
  assign o[44626] = i[44626];
  assign o[44625] = i[44625];
  assign o[44624] = i[44624];
  assign o[44623] = i[44623];
  assign o[44622] = i[44622];
  assign o[44621] = i[44621];
  assign o[44620] = i[44620];
  assign o[44619] = i[44619];
  assign o[44618] = i[44618];
  assign o[44617] = i[44617];
  assign o[44616] = i[44616];
  assign o[44615] = i[44615];
  assign o[44614] = i[44614];
  assign o[44613] = i[44613];
  assign o[44612] = i[44612];
  assign o[44611] = i[44611];
  assign o[44610] = i[44610];
  assign o[44609] = i[44609];
  assign o[44608] = i[44608];
  assign o[44607] = i[44607];
  assign o[44606] = i[44606];
  assign o[44605] = i[44605];
  assign o[44604] = i[44604];
  assign o[44603] = i[44603];
  assign o[44602] = i[44602];
  assign o[44601] = i[44601];
  assign o[44600] = i[44600];
  assign o[44599] = i[44599];
  assign o[44598] = i[44598];
  assign o[44597] = i[44597];
  assign o[44596] = i[44596];
  assign o[44595] = i[44595];
  assign o[44594] = i[44594];
  assign o[44593] = i[44593];
  assign o[44592] = i[44592];
  assign o[44591] = i[44591];
  assign o[44590] = i[44590];
  assign o[44589] = i[44589];
  assign o[44588] = i[44588];
  assign o[44587] = i[44587];
  assign o[44586] = i[44586];
  assign o[44585] = i[44585];
  assign o[44584] = i[44584];
  assign o[44583] = i[44583];
  assign o[44582] = i[44582];
  assign o[44581] = i[44581];
  assign o[44580] = i[44580];
  assign o[44579] = i[44579];
  assign o[44578] = i[44578];
  assign o[44577] = i[44577];
  assign o[44576] = i[44576];
  assign o[44575] = i[44575];
  assign o[44574] = i[44574];
  assign o[44573] = i[44573];
  assign o[44572] = i[44572];
  assign o[44571] = i[44571];
  assign o[44570] = i[44570];
  assign o[44569] = i[44569];
  assign o[44568] = i[44568];
  assign o[44567] = i[44567];
  assign o[44566] = i[44566];
  assign o[44565] = i[44565];
  assign o[44564] = i[44564];
  assign o[44563] = i[44563];
  assign o[44562] = i[44562];
  assign o[44561] = i[44561];
  assign o[44560] = i[44560];
  assign o[44559] = i[44559];
  assign o[44558] = i[44558];
  assign o[44557] = i[44557];
  assign o[44556] = i[44556];
  assign o[44555] = i[44555];
  assign o[44554] = i[44554];
  assign o[44553] = i[44553];
  assign o[44552] = i[44552];
  assign o[44551] = i[44551];
  assign o[44550] = i[44550];
  assign o[44549] = i[44549];
  assign o[44548] = i[44548];
  assign o[44547] = i[44547];
  assign o[44546] = i[44546];
  assign o[44545] = i[44545];
  assign o[44544] = i[44544];
  assign o[44543] = i[44543];
  assign o[44542] = i[44542];
  assign o[44541] = i[44541];
  assign o[44540] = i[44540];
  assign o[44539] = i[44539];
  assign o[44538] = i[44538];
  assign o[44537] = i[44537];
  assign o[44536] = i[44536];
  assign o[44535] = i[44535];
  assign o[44534] = i[44534];
  assign o[44533] = i[44533];
  assign o[44532] = i[44532];
  assign o[44531] = i[44531];
  assign o[44530] = i[44530];
  assign o[44529] = i[44529];
  assign o[44528] = i[44528];
  assign o[44527] = i[44527];
  assign o[44526] = i[44526];
  assign o[44525] = i[44525];
  assign o[44524] = i[44524];
  assign o[44523] = i[44523];
  assign o[44522] = i[44522];
  assign o[44521] = i[44521];
  assign o[44520] = i[44520];
  assign o[44519] = i[44519];
  assign o[44518] = i[44518];
  assign o[44517] = i[44517];
  assign o[44516] = i[44516];
  assign o[44515] = i[44515];
  assign o[44514] = i[44514];
  assign o[44513] = i[44513];
  assign o[44512] = i[44512];
  assign o[44511] = i[44511];
  assign o[44510] = i[44510];
  assign o[44509] = i[44509];
  assign o[44508] = i[44508];
  assign o[44507] = i[44507];
  assign o[44506] = i[44506];
  assign o[44505] = i[44505];
  assign o[44504] = i[44504];
  assign o[44503] = i[44503];
  assign o[44502] = i[44502];
  assign o[44501] = i[44501];
  assign o[44500] = i[44500];
  assign o[44499] = i[44499];
  assign o[44498] = i[44498];
  assign o[44497] = i[44497];
  assign o[44496] = i[44496];
  assign o[44495] = i[44495];
  assign o[44494] = i[44494];
  assign o[44493] = i[44493];
  assign o[44492] = i[44492];
  assign o[44491] = i[44491];
  assign o[44490] = i[44490];
  assign o[44489] = i[44489];
  assign o[44488] = i[44488];
  assign o[44487] = i[44487];
  assign o[44486] = i[44486];
  assign o[44485] = i[44485];
  assign o[44484] = i[44484];
  assign o[44483] = i[44483];
  assign o[44482] = i[44482];
  assign o[44481] = i[44481];
  assign o[44480] = i[44480];
  assign o[44479] = i[44479];
  assign o[44478] = i[44478];
  assign o[44477] = i[44477];
  assign o[44476] = i[44476];
  assign o[44475] = i[44475];
  assign o[44474] = i[44474];
  assign o[44473] = i[44473];
  assign o[44472] = i[44472];
  assign o[44471] = i[44471];
  assign o[44470] = i[44470];
  assign o[44469] = i[44469];
  assign o[44468] = i[44468];
  assign o[44467] = i[44467];
  assign o[44466] = i[44466];
  assign o[44465] = i[44465];
  assign o[44464] = i[44464];
  assign o[44463] = i[44463];
  assign o[44462] = i[44462];
  assign o[44461] = i[44461];
  assign o[44460] = i[44460];
  assign o[44459] = i[44459];
  assign o[44458] = i[44458];
  assign o[44457] = i[44457];
  assign o[44456] = i[44456];
  assign o[44455] = i[44455];
  assign o[44454] = i[44454];
  assign o[44453] = i[44453];
  assign o[44452] = i[44452];
  assign o[44451] = i[44451];
  assign o[44450] = i[44450];
  assign o[44449] = i[44449];
  assign o[44448] = i[44448];
  assign o[44447] = i[44447];
  assign o[44446] = i[44446];
  assign o[44445] = i[44445];
  assign o[44444] = i[44444];
  assign o[44443] = i[44443];
  assign o[44442] = i[44442];
  assign o[44441] = i[44441];
  assign o[44440] = i[44440];
  assign o[44439] = i[44439];
  assign o[44438] = i[44438];
  assign o[44437] = i[44437];
  assign o[44436] = i[44436];
  assign o[44435] = i[44435];
  assign o[44434] = i[44434];
  assign o[44433] = i[44433];
  assign o[44432] = i[44432];
  assign o[44431] = i[44431];
  assign o[44430] = i[44430];
  assign o[44429] = i[44429];
  assign o[44428] = i[44428];
  assign o[44427] = i[44427];
  assign o[44426] = i[44426];
  assign o[44425] = i[44425];
  assign o[44424] = i[44424];
  assign o[44423] = i[44423];
  assign o[44422] = i[44422];
  assign o[44421] = i[44421];
  assign o[44420] = i[44420];
  assign o[44419] = i[44419];
  assign o[44418] = i[44418];
  assign o[44417] = i[44417];
  assign o[44416] = i[44416];
  assign o[44415] = i[44415];
  assign o[44414] = i[44414];
  assign o[44413] = i[44413];
  assign o[44412] = i[44412];
  assign o[44411] = i[44411];
  assign o[44410] = i[44410];
  assign o[44409] = i[44409];
  assign o[44408] = i[44408];
  assign o[44407] = i[44407];
  assign o[44406] = i[44406];
  assign o[44405] = i[44405];
  assign o[44404] = i[44404];
  assign o[44403] = i[44403];
  assign o[44402] = i[44402];
  assign o[44401] = i[44401];
  assign o[44400] = i[44400];
  assign o[44399] = i[44399];
  assign o[44398] = i[44398];
  assign o[44397] = i[44397];
  assign o[44396] = i[44396];
  assign o[44395] = i[44395];
  assign o[44394] = i[44394];
  assign o[44393] = i[44393];
  assign o[44392] = i[44392];
  assign o[44391] = i[44391];
  assign o[44390] = i[44390];
  assign o[44389] = i[44389];
  assign o[44388] = i[44388];
  assign o[44387] = i[44387];
  assign o[44386] = i[44386];
  assign o[44385] = i[44385];
  assign o[44384] = i[44384];
  assign o[44383] = i[44383];
  assign o[44382] = i[44382];
  assign o[44381] = i[44381];
  assign o[44380] = i[44380];
  assign o[44379] = i[44379];
  assign o[44378] = i[44378];
  assign o[44377] = i[44377];
  assign o[44376] = i[44376];
  assign o[44375] = i[44375];
  assign o[44374] = i[44374];
  assign o[44373] = i[44373];
  assign o[44372] = i[44372];
  assign o[44371] = i[44371];
  assign o[44370] = i[44370];
  assign o[44369] = i[44369];
  assign o[44368] = i[44368];
  assign o[44367] = i[44367];
  assign o[44366] = i[44366];
  assign o[44365] = i[44365];
  assign o[44364] = i[44364];
  assign o[44363] = i[44363];
  assign o[44362] = i[44362];
  assign o[44361] = i[44361];
  assign o[44360] = i[44360];
  assign o[44359] = i[44359];
  assign o[44358] = i[44358];
  assign o[44357] = i[44357];
  assign o[44356] = i[44356];
  assign o[44355] = i[44355];
  assign o[44354] = i[44354];
  assign o[44353] = i[44353];
  assign o[44352] = i[44352];
  assign o[44351] = i[44351];
  assign o[44350] = i[44350];
  assign o[44349] = i[44349];
  assign o[44348] = i[44348];
  assign o[44347] = i[44347];
  assign o[44346] = i[44346];
  assign o[44345] = i[44345];
  assign o[44344] = i[44344];
  assign o[44343] = i[44343];
  assign o[44342] = i[44342];
  assign o[44341] = i[44341];
  assign o[44340] = i[44340];
  assign o[44339] = i[44339];
  assign o[44338] = i[44338];
  assign o[44337] = i[44337];
  assign o[44336] = i[44336];
  assign o[44335] = i[44335];
  assign o[44334] = i[44334];
  assign o[44333] = i[44333];
  assign o[44332] = i[44332];
  assign o[44331] = i[44331];
  assign o[44330] = i[44330];
  assign o[44329] = i[44329];
  assign o[44328] = i[44328];
  assign o[44327] = i[44327];
  assign o[44326] = i[44326];
  assign o[44325] = i[44325];
  assign o[44324] = i[44324];
  assign o[44323] = i[44323];
  assign o[44322] = i[44322];
  assign o[44321] = i[44321];
  assign o[44320] = i[44320];
  assign o[44319] = i[44319];
  assign o[44318] = i[44318];
  assign o[44317] = i[44317];
  assign o[44316] = i[44316];
  assign o[44315] = i[44315];
  assign o[44314] = i[44314];
  assign o[44313] = i[44313];
  assign o[44312] = i[44312];
  assign o[44311] = i[44311];
  assign o[44310] = i[44310];
  assign o[44309] = i[44309];
  assign o[44308] = i[44308];
  assign o[44307] = i[44307];
  assign o[44306] = i[44306];
  assign o[44305] = i[44305];
  assign o[44304] = i[44304];
  assign o[44303] = i[44303];
  assign o[44302] = i[44302];
  assign o[44301] = i[44301];
  assign o[44300] = i[44300];
  assign o[44299] = i[44299];
  assign o[44298] = i[44298];
  assign o[44297] = i[44297];
  assign o[44296] = i[44296];
  assign o[44295] = i[44295];
  assign o[44294] = i[44294];
  assign o[44293] = i[44293];
  assign o[44292] = i[44292];
  assign o[44291] = i[44291];
  assign o[44290] = i[44290];
  assign o[44289] = i[44289];
  assign o[44288] = i[44288];
  assign o[44287] = i[44287];
  assign o[44286] = i[44286];
  assign o[44285] = i[44285];
  assign o[44284] = i[44284];
  assign o[44283] = i[44283];
  assign o[44282] = i[44282];
  assign o[44281] = i[44281];
  assign o[44280] = i[44280];
  assign o[44279] = i[44279];
  assign o[44278] = i[44278];
  assign o[44277] = i[44277];
  assign o[44276] = i[44276];
  assign o[44275] = i[44275];
  assign o[44274] = i[44274];
  assign o[44273] = i[44273];
  assign o[44272] = i[44272];
  assign o[44271] = i[44271];
  assign o[44270] = i[44270];
  assign o[44269] = i[44269];
  assign o[44268] = i[44268];
  assign o[44267] = i[44267];
  assign o[44266] = i[44266];
  assign o[44265] = i[44265];
  assign o[44264] = i[44264];
  assign o[44263] = i[44263];
  assign o[44262] = i[44262];
  assign o[44261] = i[44261];
  assign o[44260] = i[44260];
  assign o[44259] = i[44259];
  assign o[44258] = i[44258];
  assign o[44257] = i[44257];
  assign o[44256] = i[44256];
  assign o[44255] = i[44255];
  assign o[44254] = i[44254];
  assign o[44253] = i[44253];
  assign o[44252] = i[44252];
  assign o[44251] = i[44251];
  assign o[44250] = i[44250];
  assign o[44249] = i[44249];
  assign o[44248] = i[44248];
  assign o[44247] = i[44247];
  assign o[44246] = i[44246];
  assign o[44245] = i[44245];
  assign o[44244] = i[44244];
  assign o[44243] = i[44243];
  assign o[44242] = i[44242];
  assign o[44241] = i[44241];
  assign o[44240] = i[44240];
  assign o[44239] = i[44239];
  assign o[44238] = i[44238];
  assign o[44237] = i[44237];
  assign o[44236] = i[44236];
  assign o[44235] = i[44235];
  assign o[44234] = i[44234];
  assign o[44233] = i[44233];
  assign o[44232] = i[44232];
  assign o[44231] = i[44231];
  assign o[44230] = i[44230];
  assign o[44229] = i[44229];
  assign o[44228] = i[44228];
  assign o[44227] = i[44227];
  assign o[44226] = i[44226];
  assign o[44225] = i[44225];
  assign o[44224] = i[44224];
  assign o[44223] = i[44223];
  assign o[44222] = i[44222];
  assign o[44221] = i[44221];
  assign o[44220] = i[44220];
  assign o[44219] = i[44219];
  assign o[44218] = i[44218];
  assign o[44217] = i[44217];
  assign o[44216] = i[44216];
  assign o[44215] = i[44215];
  assign o[44214] = i[44214];
  assign o[44213] = i[44213];
  assign o[44212] = i[44212];
  assign o[44211] = i[44211];
  assign o[44210] = i[44210];
  assign o[44209] = i[44209];
  assign o[44208] = i[44208];
  assign o[44207] = i[44207];
  assign o[44206] = i[44206];
  assign o[44205] = i[44205];
  assign o[44204] = i[44204];
  assign o[44203] = i[44203];
  assign o[44202] = i[44202];
  assign o[44201] = i[44201];
  assign o[44200] = i[44200];
  assign o[44199] = i[44199];
  assign o[44198] = i[44198];
  assign o[44197] = i[44197];
  assign o[44196] = i[44196];
  assign o[44195] = i[44195];
  assign o[44194] = i[44194];
  assign o[44193] = i[44193];
  assign o[44192] = i[44192];
  assign o[44191] = i[44191];
  assign o[44190] = i[44190];
  assign o[44189] = i[44189];
  assign o[44188] = i[44188];
  assign o[44187] = i[44187];
  assign o[44186] = i[44186];
  assign o[44185] = i[44185];
  assign o[44184] = i[44184];
  assign o[44183] = i[44183];
  assign o[44182] = i[44182];
  assign o[44181] = i[44181];
  assign o[44180] = i[44180];
  assign o[44179] = i[44179];
  assign o[44178] = i[44178];
  assign o[44177] = i[44177];
  assign o[44176] = i[44176];
  assign o[44175] = i[44175];
  assign o[44174] = i[44174];
  assign o[44173] = i[44173];
  assign o[44172] = i[44172];
  assign o[44171] = i[44171];
  assign o[44170] = i[44170];
  assign o[44169] = i[44169];
  assign o[44168] = i[44168];
  assign o[44167] = i[44167];
  assign o[44166] = i[44166];
  assign o[44165] = i[44165];
  assign o[44164] = i[44164];
  assign o[44163] = i[44163];
  assign o[44162] = i[44162];
  assign o[44161] = i[44161];
  assign o[44160] = i[44160];
  assign o[44159] = i[44159];
  assign o[44158] = i[44158];
  assign o[44157] = i[44157];
  assign o[44156] = i[44156];
  assign o[44155] = i[44155];
  assign o[44154] = i[44154];
  assign o[44153] = i[44153];
  assign o[44152] = i[44152];
  assign o[44151] = i[44151];
  assign o[44150] = i[44150];
  assign o[44149] = i[44149];
  assign o[44148] = i[44148];
  assign o[44147] = i[44147];
  assign o[44146] = i[44146];
  assign o[44145] = i[44145];
  assign o[44144] = i[44144];
  assign o[44143] = i[44143];
  assign o[44142] = i[44142];
  assign o[44141] = i[44141];
  assign o[44140] = i[44140];
  assign o[44139] = i[44139];
  assign o[44138] = i[44138];
  assign o[44137] = i[44137];
  assign o[44136] = i[44136];
  assign o[44135] = i[44135];
  assign o[44134] = i[44134];
  assign o[44133] = i[44133];
  assign o[44132] = i[44132];
  assign o[44131] = i[44131];
  assign o[44130] = i[44130];
  assign o[44129] = i[44129];
  assign o[44128] = i[44128];
  assign o[44127] = i[44127];
  assign o[44126] = i[44126];
  assign o[44125] = i[44125];
  assign o[44124] = i[44124];
  assign o[44123] = i[44123];
  assign o[44122] = i[44122];
  assign o[44121] = i[44121];
  assign o[44120] = i[44120];
  assign o[44119] = i[44119];
  assign o[44118] = i[44118];
  assign o[44117] = i[44117];
  assign o[44116] = i[44116];
  assign o[44115] = i[44115];
  assign o[44114] = i[44114];
  assign o[44113] = i[44113];
  assign o[44112] = i[44112];
  assign o[44111] = i[44111];
  assign o[44110] = i[44110];
  assign o[44109] = i[44109];
  assign o[44108] = i[44108];
  assign o[44107] = i[44107];
  assign o[44106] = i[44106];
  assign o[44105] = i[44105];
  assign o[44104] = i[44104];
  assign o[44103] = i[44103];
  assign o[44102] = i[44102];
  assign o[44101] = i[44101];
  assign o[44100] = i[44100];
  assign o[44099] = i[44099];
  assign o[44098] = i[44098];
  assign o[44097] = i[44097];
  assign o[44096] = i[44096];
  assign o[44095] = i[44095];
  assign o[44094] = i[44094];
  assign o[44093] = i[44093];
  assign o[44092] = i[44092];
  assign o[44091] = i[44091];
  assign o[44090] = i[44090];
  assign o[44089] = i[44089];
  assign o[44088] = i[44088];
  assign o[44087] = i[44087];
  assign o[44086] = i[44086];
  assign o[44085] = i[44085];
  assign o[44084] = i[44084];
  assign o[44083] = i[44083];
  assign o[44082] = i[44082];
  assign o[44081] = i[44081];
  assign o[44080] = i[44080];
  assign o[44079] = i[44079];
  assign o[44078] = i[44078];
  assign o[44077] = i[44077];
  assign o[44076] = i[44076];
  assign o[44075] = i[44075];
  assign o[44074] = i[44074];
  assign o[44073] = i[44073];
  assign o[44072] = i[44072];
  assign o[44071] = i[44071];
  assign o[44070] = i[44070];
  assign o[44069] = i[44069];
  assign o[44068] = i[44068];
  assign o[44067] = i[44067];
  assign o[44066] = i[44066];
  assign o[44065] = i[44065];
  assign o[44064] = i[44064];
  assign o[44063] = i[44063];
  assign o[44062] = i[44062];
  assign o[44061] = i[44061];
  assign o[44060] = i[44060];
  assign o[44059] = i[44059];
  assign o[44058] = i[44058];
  assign o[44057] = i[44057];
  assign o[44056] = i[44056];
  assign o[44055] = i[44055];
  assign o[44054] = i[44054];
  assign o[44053] = i[44053];
  assign o[44052] = i[44052];
  assign o[44051] = i[44051];
  assign o[44050] = i[44050];
  assign o[44049] = i[44049];
  assign o[44048] = i[44048];
  assign o[44047] = i[44047];
  assign o[44046] = i[44046];
  assign o[44045] = i[44045];
  assign o[44044] = i[44044];
  assign o[44043] = i[44043];
  assign o[44042] = i[44042];
  assign o[44041] = i[44041];
  assign o[44040] = i[44040];
  assign o[44039] = i[44039];
  assign o[44038] = i[44038];
  assign o[44037] = i[44037];
  assign o[44036] = i[44036];
  assign o[44035] = i[44035];
  assign o[44034] = i[44034];
  assign o[44033] = i[44033];
  assign o[44032] = i[44032];
  assign o[44031] = i[44031];
  assign o[44030] = i[44030];
  assign o[44029] = i[44029];
  assign o[44028] = i[44028];
  assign o[44027] = i[44027];
  assign o[44026] = i[44026];
  assign o[44025] = i[44025];
  assign o[44024] = i[44024];
  assign o[44023] = i[44023];
  assign o[44022] = i[44022];
  assign o[44021] = i[44021];
  assign o[44020] = i[44020];
  assign o[44019] = i[44019];
  assign o[44018] = i[44018];
  assign o[44017] = i[44017];
  assign o[44016] = i[44016];
  assign o[44015] = i[44015];
  assign o[44014] = i[44014];
  assign o[44013] = i[44013];
  assign o[44012] = i[44012];
  assign o[44011] = i[44011];
  assign o[44010] = i[44010];
  assign o[44009] = i[44009];
  assign o[44008] = i[44008];
  assign o[44007] = i[44007];
  assign o[44006] = i[44006];
  assign o[44005] = i[44005];
  assign o[44004] = i[44004];
  assign o[44003] = i[44003];
  assign o[44002] = i[44002];
  assign o[44001] = i[44001];
  assign o[44000] = i[44000];
  assign o[43999] = i[43999];
  assign o[43998] = i[43998];
  assign o[43997] = i[43997];
  assign o[43996] = i[43996];
  assign o[43995] = i[43995];
  assign o[43994] = i[43994];
  assign o[43993] = i[43993];
  assign o[43992] = i[43992];
  assign o[43991] = i[43991];
  assign o[43990] = i[43990];
  assign o[43989] = i[43989];
  assign o[43988] = i[43988];
  assign o[43987] = i[43987];
  assign o[43986] = i[43986];
  assign o[43985] = i[43985];
  assign o[43984] = i[43984];
  assign o[43983] = i[43983];
  assign o[43982] = i[43982];
  assign o[43981] = i[43981];
  assign o[43980] = i[43980];
  assign o[43979] = i[43979];
  assign o[43978] = i[43978];
  assign o[43977] = i[43977];
  assign o[43976] = i[43976];
  assign o[43975] = i[43975];
  assign o[43974] = i[43974];
  assign o[43973] = i[43973];
  assign o[43972] = i[43972];
  assign o[43971] = i[43971];
  assign o[43970] = i[43970];
  assign o[43969] = i[43969];
  assign o[43968] = i[43968];
  assign o[43967] = i[43967];
  assign o[43966] = i[43966];
  assign o[43965] = i[43965];
  assign o[43964] = i[43964];
  assign o[43963] = i[43963];
  assign o[43962] = i[43962];
  assign o[43961] = i[43961];
  assign o[43960] = i[43960];
  assign o[43959] = i[43959];
  assign o[43958] = i[43958];
  assign o[43957] = i[43957];
  assign o[43956] = i[43956];
  assign o[43955] = i[43955];
  assign o[43954] = i[43954];
  assign o[43953] = i[43953];
  assign o[43952] = i[43952];
  assign o[43951] = i[43951];
  assign o[43950] = i[43950];
  assign o[43949] = i[43949];
  assign o[43948] = i[43948];
  assign o[43947] = i[43947];
  assign o[43946] = i[43946];
  assign o[43945] = i[43945];
  assign o[43944] = i[43944];
  assign o[43943] = i[43943];
  assign o[43942] = i[43942];
  assign o[43941] = i[43941];
  assign o[43940] = i[43940];
  assign o[43939] = i[43939];
  assign o[43938] = i[43938];
  assign o[43937] = i[43937];
  assign o[43936] = i[43936];
  assign o[43935] = i[43935];
  assign o[43934] = i[43934];
  assign o[43933] = i[43933];
  assign o[43932] = i[43932];
  assign o[43931] = i[43931];
  assign o[43930] = i[43930];
  assign o[43929] = i[43929];
  assign o[43928] = i[43928];
  assign o[43927] = i[43927];
  assign o[43926] = i[43926];
  assign o[43925] = i[43925];
  assign o[43924] = i[43924];
  assign o[43923] = i[43923];
  assign o[43922] = i[43922];
  assign o[43921] = i[43921];
  assign o[43920] = i[43920];
  assign o[43919] = i[43919];
  assign o[43918] = i[43918];
  assign o[43917] = i[43917];
  assign o[43916] = i[43916];
  assign o[43915] = i[43915];
  assign o[43914] = i[43914];
  assign o[43913] = i[43913];
  assign o[43912] = i[43912];
  assign o[43911] = i[43911];
  assign o[43910] = i[43910];
  assign o[43909] = i[43909];
  assign o[43908] = i[43908];
  assign o[43907] = i[43907];
  assign o[43906] = i[43906];
  assign o[43905] = i[43905];
  assign o[43904] = i[43904];
  assign o[43903] = i[43903];
  assign o[43902] = i[43902];
  assign o[43901] = i[43901];
  assign o[43900] = i[43900];
  assign o[43899] = i[43899];
  assign o[43898] = i[43898];
  assign o[43897] = i[43897];
  assign o[43896] = i[43896];
  assign o[43895] = i[43895];
  assign o[43894] = i[43894];
  assign o[43893] = i[43893];
  assign o[43892] = i[43892];
  assign o[43891] = i[43891];
  assign o[43890] = i[43890];
  assign o[43889] = i[43889];
  assign o[43888] = i[43888];
  assign o[43887] = i[43887];
  assign o[43886] = i[43886];
  assign o[43885] = i[43885];
  assign o[43884] = i[43884];
  assign o[43883] = i[43883];
  assign o[43882] = i[43882];
  assign o[43881] = i[43881];
  assign o[43880] = i[43880];
  assign o[43879] = i[43879];
  assign o[43878] = i[43878];
  assign o[43877] = i[43877];
  assign o[43876] = i[43876];
  assign o[43875] = i[43875];
  assign o[43874] = i[43874];
  assign o[43873] = i[43873];
  assign o[43872] = i[43872];
  assign o[43871] = i[43871];
  assign o[43870] = i[43870];
  assign o[43869] = i[43869];
  assign o[43868] = i[43868];
  assign o[43867] = i[43867];
  assign o[43866] = i[43866];
  assign o[43865] = i[43865];
  assign o[43864] = i[43864];
  assign o[43863] = i[43863];
  assign o[43862] = i[43862];
  assign o[43861] = i[43861];
  assign o[43860] = i[43860];
  assign o[43859] = i[43859];
  assign o[43858] = i[43858];
  assign o[43857] = i[43857];
  assign o[43856] = i[43856];
  assign o[43855] = i[43855];
  assign o[43854] = i[43854];
  assign o[43853] = i[43853];
  assign o[43852] = i[43852];
  assign o[43851] = i[43851];
  assign o[43850] = i[43850];
  assign o[43849] = i[43849];
  assign o[43848] = i[43848];
  assign o[43847] = i[43847];
  assign o[43846] = i[43846];
  assign o[43845] = i[43845];
  assign o[43844] = i[43844];
  assign o[43843] = i[43843];
  assign o[43842] = i[43842];
  assign o[43841] = i[43841];
  assign o[43840] = i[43840];
  assign o[43839] = i[43839];
  assign o[43838] = i[43838];
  assign o[43837] = i[43837];
  assign o[43836] = i[43836];
  assign o[43835] = i[43835];
  assign o[43834] = i[43834];
  assign o[43833] = i[43833];
  assign o[43832] = i[43832];
  assign o[43831] = i[43831];
  assign o[43830] = i[43830];
  assign o[43829] = i[43829];
  assign o[43828] = i[43828];
  assign o[43827] = i[43827];
  assign o[43826] = i[43826];
  assign o[43825] = i[43825];
  assign o[43824] = i[43824];
  assign o[43823] = i[43823];
  assign o[43822] = i[43822];
  assign o[43821] = i[43821];
  assign o[43820] = i[43820];
  assign o[43819] = i[43819];
  assign o[43818] = i[43818];
  assign o[43817] = i[43817];
  assign o[43816] = i[43816];
  assign o[43815] = i[43815];
  assign o[43814] = i[43814];
  assign o[43813] = i[43813];
  assign o[43812] = i[43812];
  assign o[43811] = i[43811];
  assign o[43810] = i[43810];
  assign o[43809] = i[43809];
  assign o[43808] = i[43808];
  assign o[43807] = i[43807];
  assign o[43806] = i[43806];
  assign o[43805] = i[43805];
  assign o[43804] = i[43804];
  assign o[43803] = i[43803];
  assign o[43802] = i[43802];
  assign o[43801] = i[43801];
  assign o[43800] = i[43800];
  assign o[43799] = i[43799];
  assign o[43798] = i[43798];
  assign o[43797] = i[43797];
  assign o[43796] = i[43796];
  assign o[43795] = i[43795];
  assign o[43794] = i[43794];
  assign o[43793] = i[43793];
  assign o[43792] = i[43792];
  assign o[43791] = i[43791];
  assign o[43790] = i[43790];
  assign o[43789] = i[43789];
  assign o[43788] = i[43788];
  assign o[43787] = i[43787];
  assign o[43786] = i[43786];
  assign o[43785] = i[43785];
  assign o[43784] = i[43784];
  assign o[43783] = i[43783];
  assign o[43782] = i[43782];
  assign o[43781] = i[43781];
  assign o[43780] = i[43780];
  assign o[43779] = i[43779];
  assign o[43778] = i[43778];
  assign o[43777] = i[43777];
  assign o[43776] = i[43776];
  assign o[43775] = i[43775];
  assign o[43774] = i[43774];
  assign o[43773] = i[43773];
  assign o[43772] = i[43772];
  assign o[43771] = i[43771];
  assign o[43770] = i[43770];
  assign o[43769] = i[43769];
  assign o[43768] = i[43768];
  assign o[43767] = i[43767];
  assign o[43766] = i[43766];
  assign o[43765] = i[43765];
  assign o[43764] = i[43764];
  assign o[43763] = i[43763];
  assign o[43762] = i[43762];
  assign o[43761] = i[43761];
  assign o[43760] = i[43760];
  assign o[43759] = i[43759];
  assign o[43758] = i[43758];
  assign o[43757] = i[43757];
  assign o[43756] = i[43756];
  assign o[43755] = i[43755];
  assign o[43754] = i[43754];
  assign o[43753] = i[43753];
  assign o[43752] = i[43752];
  assign o[43751] = i[43751];
  assign o[43750] = i[43750];
  assign o[43749] = i[43749];
  assign o[43748] = i[43748];
  assign o[43747] = i[43747];
  assign o[43746] = i[43746];
  assign o[43745] = i[43745];
  assign o[43744] = i[43744];
  assign o[43743] = i[43743];
  assign o[43742] = i[43742];
  assign o[43741] = i[43741];
  assign o[43740] = i[43740];
  assign o[43739] = i[43739];
  assign o[43738] = i[43738];
  assign o[43737] = i[43737];
  assign o[43736] = i[43736];
  assign o[43735] = i[43735];
  assign o[43734] = i[43734];
  assign o[43733] = i[43733];
  assign o[43732] = i[43732];
  assign o[43731] = i[43731];
  assign o[43730] = i[43730];
  assign o[43729] = i[43729];
  assign o[43728] = i[43728];
  assign o[43727] = i[43727];
  assign o[43726] = i[43726];
  assign o[43725] = i[43725];
  assign o[43724] = i[43724];
  assign o[43723] = i[43723];
  assign o[43722] = i[43722];
  assign o[43721] = i[43721];
  assign o[43720] = i[43720];
  assign o[43719] = i[43719];
  assign o[43718] = i[43718];
  assign o[43717] = i[43717];
  assign o[43716] = i[43716];
  assign o[43715] = i[43715];
  assign o[43714] = i[43714];
  assign o[43713] = i[43713];
  assign o[43712] = i[43712];
  assign o[43711] = i[43711];
  assign o[43710] = i[43710];
  assign o[43709] = i[43709];
  assign o[43708] = i[43708];
  assign o[43707] = i[43707];
  assign o[43706] = i[43706];
  assign o[43705] = i[43705];
  assign o[43704] = i[43704];
  assign o[43703] = i[43703];
  assign o[43702] = i[43702];
  assign o[43701] = i[43701];
  assign o[43700] = i[43700];
  assign o[43699] = i[43699];
  assign o[43698] = i[43698];
  assign o[43697] = i[43697];
  assign o[43696] = i[43696];
  assign o[43695] = i[43695];
  assign o[43694] = i[43694];
  assign o[43693] = i[43693];
  assign o[43692] = i[43692];
  assign o[43691] = i[43691];
  assign o[43690] = i[43690];
  assign o[43689] = i[43689];
  assign o[43688] = i[43688];
  assign o[43687] = i[43687];
  assign o[43686] = i[43686];
  assign o[43685] = i[43685];
  assign o[43684] = i[43684];
  assign o[43683] = i[43683];
  assign o[43682] = i[43682];
  assign o[43681] = i[43681];
  assign o[43680] = i[43680];
  assign o[43679] = i[43679];
  assign o[43678] = i[43678];
  assign o[43677] = i[43677];
  assign o[43676] = i[43676];
  assign o[43675] = i[43675];
  assign o[43674] = i[43674];
  assign o[43673] = i[43673];
  assign o[43672] = i[43672];
  assign o[43671] = i[43671];
  assign o[43670] = i[43670];
  assign o[43669] = i[43669];
  assign o[43668] = i[43668];
  assign o[43667] = i[43667];
  assign o[43666] = i[43666];
  assign o[43665] = i[43665];
  assign o[43664] = i[43664];
  assign o[43663] = i[43663];
  assign o[43662] = i[43662];
  assign o[43661] = i[43661];
  assign o[43660] = i[43660];
  assign o[43659] = i[43659];
  assign o[43658] = i[43658];
  assign o[43657] = i[43657];
  assign o[43656] = i[43656];
  assign o[43655] = i[43655];
  assign o[43654] = i[43654];
  assign o[43653] = i[43653];
  assign o[43652] = i[43652];
  assign o[43651] = i[43651];
  assign o[43650] = i[43650];
  assign o[43649] = i[43649];
  assign o[43648] = i[43648];
  assign o[43647] = i[43647];
  assign o[43646] = i[43646];
  assign o[43645] = i[43645];
  assign o[43644] = i[43644];
  assign o[43643] = i[43643];
  assign o[43642] = i[43642];
  assign o[43641] = i[43641];
  assign o[43640] = i[43640];
  assign o[43639] = i[43639];
  assign o[43638] = i[43638];
  assign o[43637] = i[43637];
  assign o[43636] = i[43636];
  assign o[43635] = i[43635];
  assign o[43634] = i[43634];
  assign o[43633] = i[43633];
  assign o[43632] = i[43632];
  assign o[43631] = i[43631];
  assign o[43630] = i[43630];
  assign o[43629] = i[43629];
  assign o[43628] = i[43628];
  assign o[43627] = i[43627];
  assign o[43626] = i[43626];
  assign o[43625] = i[43625];
  assign o[43624] = i[43624];
  assign o[43623] = i[43623];
  assign o[43622] = i[43622];
  assign o[43621] = i[43621];
  assign o[43620] = i[43620];
  assign o[43619] = i[43619];
  assign o[43618] = i[43618];
  assign o[43617] = i[43617];
  assign o[43616] = i[43616];
  assign o[43615] = i[43615];
  assign o[43614] = i[43614];
  assign o[43613] = i[43613];
  assign o[43612] = i[43612];
  assign o[43611] = i[43611];
  assign o[43610] = i[43610];
  assign o[43609] = i[43609];
  assign o[43608] = i[43608];
  assign o[43607] = i[43607];
  assign o[43606] = i[43606];
  assign o[43605] = i[43605];
  assign o[43604] = i[43604];
  assign o[43603] = i[43603];
  assign o[43602] = i[43602];
  assign o[43601] = i[43601];
  assign o[43600] = i[43600];
  assign o[43599] = i[43599];
  assign o[43598] = i[43598];
  assign o[43597] = i[43597];
  assign o[43596] = i[43596];
  assign o[43595] = i[43595];
  assign o[43594] = i[43594];
  assign o[43593] = i[43593];
  assign o[43592] = i[43592];
  assign o[43591] = i[43591];
  assign o[43590] = i[43590];
  assign o[43589] = i[43589];
  assign o[43588] = i[43588];
  assign o[43587] = i[43587];
  assign o[43586] = i[43586];
  assign o[43585] = i[43585];
  assign o[43584] = i[43584];
  assign o[43583] = i[43583];
  assign o[43582] = i[43582];
  assign o[43581] = i[43581];
  assign o[43580] = i[43580];
  assign o[43579] = i[43579];
  assign o[43578] = i[43578];
  assign o[43577] = i[43577];
  assign o[43576] = i[43576];
  assign o[43575] = i[43575];
  assign o[43574] = i[43574];
  assign o[43573] = i[43573];
  assign o[43572] = i[43572];
  assign o[43571] = i[43571];
  assign o[43570] = i[43570];
  assign o[43569] = i[43569];
  assign o[43568] = i[43568];
  assign o[43567] = i[43567];
  assign o[43566] = i[43566];
  assign o[43565] = i[43565];
  assign o[43564] = i[43564];
  assign o[43563] = i[43563];
  assign o[43562] = i[43562];
  assign o[43561] = i[43561];
  assign o[43560] = i[43560];
  assign o[43559] = i[43559];
  assign o[43558] = i[43558];
  assign o[43557] = i[43557];
  assign o[43556] = i[43556];
  assign o[43555] = i[43555];
  assign o[43554] = i[43554];
  assign o[43553] = i[43553];
  assign o[43552] = i[43552];
  assign o[43551] = i[43551];
  assign o[43550] = i[43550];
  assign o[43549] = i[43549];
  assign o[43548] = i[43548];
  assign o[43547] = i[43547];
  assign o[43546] = i[43546];
  assign o[43545] = i[43545];
  assign o[43544] = i[43544];
  assign o[43543] = i[43543];
  assign o[43542] = i[43542];
  assign o[43541] = i[43541];
  assign o[43540] = i[43540];
  assign o[43539] = i[43539];
  assign o[43538] = i[43538];
  assign o[43537] = i[43537];
  assign o[43536] = i[43536];
  assign o[43535] = i[43535];
  assign o[43534] = i[43534];
  assign o[43533] = i[43533];
  assign o[43532] = i[43532];
  assign o[43531] = i[43531];
  assign o[43530] = i[43530];
  assign o[43529] = i[43529];
  assign o[43528] = i[43528];
  assign o[43527] = i[43527];
  assign o[43526] = i[43526];
  assign o[43525] = i[43525];
  assign o[43524] = i[43524];
  assign o[43523] = i[43523];
  assign o[43522] = i[43522];
  assign o[43521] = i[43521];
  assign o[43520] = i[43520];
  assign o[43519] = i[43519];
  assign o[43518] = i[43518];
  assign o[43517] = i[43517];
  assign o[43516] = i[43516];
  assign o[43515] = i[43515];
  assign o[43514] = i[43514];
  assign o[43513] = i[43513];
  assign o[43512] = i[43512];
  assign o[43511] = i[43511];
  assign o[43510] = i[43510];
  assign o[43509] = i[43509];
  assign o[43508] = i[43508];
  assign o[43507] = i[43507];
  assign o[43506] = i[43506];
  assign o[43505] = i[43505];
  assign o[43504] = i[43504];
  assign o[43503] = i[43503];
  assign o[43502] = i[43502];
  assign o[43501] = i[43501];
  assign o[43500] = i[43500];
  assign o[43499] = i[43499];
  assign o[43498] = i[43498];
  assign o[43497] = i[43497];
  assign o[43496] = i[43496];
  assign o[43495] = i[43495];
  assign o[43494] = i[43494];
  assign o[43493] = i[43493];
  assign o[43492] = i[43492];
  assign o[43491] = i[43491];
  assign o[43490] = i[43490];
  assign o[43489] = i[43489];
  assign o[43488] = i[43488];
  assign o[43487] = i[43487];
  assign o[43486] = i[43486];
  assign o[43485] = i[43485];
  assign o[43484] = i[43484];
  assign o[43483] = i[43483];
  assign o[43482] = i[43482];
  assign o[43481] = i[43481];
  assign o[43480] = i[43480];
  assign o[43479] = i[43479];
  assign o[43478] = i[43478];
  assign o[43477] = i[43477];
  assign o[43476] = i[43476];
  assign o[43475] = i[43475];
  assign o[43474] = i[43474];
  assign o[43473] = i[43473];
  assign o[43472] = i[43472];
  assign o[43471] = i[43471];
  assign o[43470] = i[43470];
  assign o[43469] = i[43469];
  assign o[43468] = i[43468];
  assign o[43467] = i[43467];
  assign o[43466] = i[43466];
  assign o[43465] = i[43465];
  assign o[43464] = i[43464];
  assign o[43463] = i[43463];
  assign o[43462] = i[43462];
  assign o[43461] = i[43461];
  assign o[43460] = i[43460];
  assign o[43459] = i[43459];
  assign o[43458] = i[43458];
  assign o[43457] = i[43457];
  assign o[43456] = i[43456];
  assign o[43455] = i[43455];
  assign o[43454] = i[43454];
  assign o[43453] = i[43453];
  assign o[43452] = i[43452];
  assign o[43451] = i[43451];
  assign o[43450] = i[43450];
  assign o[43449] = i[43449];
  assign o[43448] = i[43448];
  assign o[43447] = i[43447];
  assign o[43446] = i[43446];
  assign o[43445] = i[43445];
  assign o[43444] = i[43444];
  assign o[43443] = i[43443];
  assign o[43442] = i[43442];
  assign o[43441] = i[43441];
  assign o[43440] = i[43440];
  assign o[43439] = i[43439];
  assign o[43438] = i[43438];
  assign o[43437] = i[43437];
  assign o[43436] = i[43436];
  assign o[43435] = i[43435];
  assign o[43434] = i[43434];
  assign o[43433] = i[43433];
  assign o[43432] = i[43432];
  assign o[43431] = i[43431];
  assign o[43430] = i[43430];
  assign o[43429] = i[43429];
  assign o[43428] = i[43428];
  assign o[43427] = i[43427];
  assign o[43426] = i[43426];
  assign o[43425] = i[43425];
  assign o[43424] = i[43424];
  assign o[43423] = i[43423];
  assign o[43422] = i[43422];
  assign o[43421] = i[43421];
  assign o[43420] = i[43420];
  assign o[43419] = i[43419];
  assign o[43418] = i[43418];
  assign o[43417] = i[43417];
  assign o[43416] = i[43416];
  assign o[43415] = i[43415];
  assign o[43414] = i[43414];
  assign o[43413] = i[43413];
  assign o[43412] = i[43412];
  assign o[43411] = i[43411];
  assign o[43410] = i[43410];
  assign o[43409] = i[43409];
  assign o[43408] = i[43408];
  assign o[43407] = i[43407];
  assign o[43406] = i[43406];
  assign o[43405] = i[43405];
  assign o[43404] = i[43404];
  assign o[43403] = i[43403];
  assign o[43402] = i[43402];
  assign o[43401] = i[43401];
  assign o[43400] = i[43400];
  assign o[43399] = i[43399];
  assign o[43398] = i[43398];
  assign o[43397] = i[43397];
  assign o[43396] = i[43396];
  assign o[43395] = i[43395];
  assign o[43394] = i[43394];
  assign o[43393] = i[43393];
  assign o[43392] = i[43392];
  assign o[43391] = i[43391];
  assign o[43390] = i[43390];
  assign o[43389] = i[43389];
  assign o[43388] = i[43388];
  assign o[43387] = i[43387];
  assign o[43386] = i[43386];
  assign o[43385] = i[43385];
  assign o[43384] = i[43384];
  assign o[43383] = i[43383];
  assign o[43382] = i[43382];
  assign o[43381] = i[43381];
  assign o[43380] = i[43380];
  assign o[43379] = i[43379];
  assign o[43378] = i[43378];
  assign o[43377] = i[43377];
  assign o[43376] = i[43376];
  assign o[43375] = i[43375];
  assign o[43374] = i[43374];
  assign o[43373] = i[43373];
  assign o[43372] = i[43372];
  assign o[43371] = i[43371];
  assign o[43370] = i[43370];
  assign o[43369] = i[43369];
  assign o[43368] = i[43368];
  assign o[43367] = i[43367];
  assign o[43366] = i[43366];
  assign o[43365] = i[43365];
  assign o[43364] = i[43364];
  assign o[43363] = i[43363];
  assign o[43362] = i[43362];
  assign o[43361] = i[43361];
  assign o[43360] = i[43360];
  assign o[43359] = i[43359];
  assign o[43358] = i[43358];
  assign o[43357] = i[43357];
  assign o[43356] = i[43356];
  assign o[43355] = i[43355];
  assign o[43354] = i[43354];
  assign o[43353] = i[43353];
  assign o[43352] = i[43352];
  assign o[43351] = i[43351];
  assign o[43350] = i[43350];
  assign o[43349] = i[43349];
  assign o[43348] = i[43348];
  assign o[43347] = i[43347];
  assign o[43346] = i[43346];
  assign o[43345] = i[43345];
  assign o[43344] = i[43344];
  assign o[43343] = i[43343];
  assign o[43342] = i[43342];
  assign o[43341] = i[43341];
  assign o[43340] = i[43340];
  assign o[43339] = i[43339];
  assign o[43338] = i[43338];
  assign o[43337] = i[43337];
  assign o[43336] = i[43336];
  assign o[43335] = i[43335];
  assign o[43334] = i[43334];
  assign o[43333] = i[43333];
  assign o[43332] = i[43332];
  assign o[43331] = i[43331];
  assign o[43330] = i[43330];
  assign o[43329] = i[43329];
  assign o[43328] = i[43328];
  assign o[43327] = i[43327];
  assign o[43326] = i[43326];
  assign o[43325] = i[43325];
  assign o[43324] = i[43324];
  assign o[43323] = i[43323];
  assign o[43322] = i[43322];
  assign o[43321] = i[43321];
  assign o[43320] = i[43320];
  assign o[43319] = i[43319];
  assign o[43318] = i[43318];
  assign o[43317] = i[43317];
  assign o[43316] = i[43316];
  assign o[43315] = i[43315];
  assign o[43314] = i[43314];
  assign o[43313] = i[43313];
  assign o[43312] = i[43312];
  assign o[43311] = i[43311];
  assign o[43310] = i[43310];
  assign o[43309] = i[43309];
  assign o[43308] = i[43308];
  assign o[43307] = i[43307];
  assign o[43306] = i[43306];
  assign o[43305] = i[43305];
  assign o[43304] = i[43304];
  assign o[43303] = i[43303];
  assign o[43302] = i[43302];
  assign o[43301] = i[43301];
  assign o[43300] = i[43300];
  assign o[43299] = i[43299];
  assign o[43298] = i[43298];
  assign o[43297] = i[43297];
  assign o[43296] = i[43296];
  assign o[43295] = i[43295];
  assign o[43294] = i[43294];
  assign o[43293] = i[43293];
  assign o[43292] = i[43292];
  assign o[43291] = i[43291];
  assign o[43290] = i[43290];
  assign o[43289] = i[43289];
  assign o[43288] = i[43288];
  assign o[43287] = i[43287];
  assign o[43286] = i[43286];
  assign o[43285] = i[43285];
  assign o[43284] = i[43284];
  assign o[43283] = i[43283];
  assign o[43282] = i[43282];
  assign o[43281] = i[43281];
  assign o[43280] = i[43280];
  assign o[43279] = i[43279];
  assign o[43278] = i[43278];
  assign o[43277] = i[43277];
  assign o[43276] = i[43276];
  assign o[43275] = i[43275];
  assign o[43274] = i[43274];
  assign o[43273] = i[43273];
  assign o[43272] = i[43272];
  assign o[43271] = i[43271];
  assign o[43270] = i[43270];
  assign o[43269] = i[43269];
  assign o[43268] = i[43268];
  assign o[43267] = i[43267];
  assign o[43266] = i[43266];
  assign o[43265] = i[43265];
  assign o[43264] = i[43264];
  assign o[43263] = i[43263];
  assign o[43262] = i[43262];
  assign o[43261] = i[43261];
  assign o[43260] = i[43260];
  assign o[43259] = i[43259];
  assign o[43258] = i[43258];
  assign o[43257] = i[43257];
  assign o[43256] = i[43256];
  assign o[43255] = i[43255];
  assign o[43254] = i[43254];
  assign o[43253] = i[43253];
  assign o[43252] = i[43252];
  assign o[43251] = i[43251];
  assign o[43250] = i[43250];
  assign o[43249] = i[43249];
  assign o[43248] = i[43248];
  assign o[43247] = i[43247];
  assign o[43246] = i[43246];
  assign o[43245] = i[43245];
  assign o[43244] = i[43244];
  assign o[43243] = i[43243];
  assign o[43242] = i[43242];
  assign o[43241] = i[43241];
  assign o[43240] = i[43240];
  assign o[43239] = i[43239];
  assign o[43238] = i[43238];
  assign o[43237] = i[43237];
  assign o[43236] = i[43236];
  assign o[43235] = i[43235];
  assign o[43234] = i[43234];
  assign o[43233] = i[43233];
  assign o[43232] = i[43232];
  assign o[43231] = i[43231];
  assign o[43230] = i[43230];
  assign o[43229] = i[43229];
  assign o[43228] = i[43228];
  assign o[43227] = i[43227];
  assign o[43226] = i[43226];
  assign o[43225] = i[43225];
  assign o[43224] = i[43224];
  assign o[43223] = i[43223];
  assign o[43222] = i[43222];
  assign o[43221] = i[43221];
  assign o[43220] = i[43220];
  assign o[43219] = i[43219];
  assign o[43218] = i[43218];
  assign o[43217] = i[43217];
  assign o[43216] = i[43216];
  assign o[43215] = i[43215];
  assign o[43214] = i[43214];
  assign o[43213] = i[43213];
  assign o[43212] = i[43212];
  assign o[43211] = i[43211];
  assign o[43210] = i[43210];
  assign o[43209] = i[43209];
  assign o[43208] = i[43208];
  assign o[43207] = i[43207];
  assign o[43206] = i[43206];
  assign o[43205] = i[43205];
  assign o[43204] = i[43204];
  assign o[43203] = i[43203];
  assign o[43202] = i[43202];
  assign o[43201] = i[43201];
  assign o[43200] = i[43200];
  assign o[43199] = i[43199];
  assign o[43198] = i[43198];
  assign o[43197] = i[43197];
  assign o[43196] = i[43196];
  assign o[43195] = i[43195];
  assign o[43194] = i[43194];
  assign o[43193] = i[43193];
  assign o[43192] = i[43192];
  assign o[43191] = i[43191];
  assign o[43190] = i[43190];
  assign o[43189] = i[43189];
  assign o[43188] = i[43188];
  assign o[43187] = i[43187];
  assign o[43186] = i[43186];
  assign o[43185] = i[43185];
  assign o[43184] = i[43184];
  assign o[43183] = i[43183];
  assign o[43182] = i[43182];
  assign o[43181] = i[43181];
  assign o[43180] = i[43180];
  assign o[43179] = i[43179];
  assign o[43178] = i[43178];
  assign o[43177] = i[43177];
  assign o[43176] = i[43176];
  assign o[43175] = i[43175];
  assign o[43174] = i[43174];
  assign o[43173] = i[43173];
  assign o[43172] = i[43172];
  assign o[43171] = i[43171];
  assign o[43170] = i[43170];
  assign o[43169] = i[43169];
  assign o[43168] = i[43168];
  assign o[43167] = i[43167];
  assign o[43166] = i[43166];
  assign o[43165] = i[43165];
  assign o[43164] = i[43164];
  assign o[43163] = i[43163];
  assign o[43162] = i[43162];
  assign o[43161] = i[43161];
  assign o[43160] = i[43160];
  assign o[43159] = i[43159];
  assign o[43158] = i[43158];
  assign o[43157] = i[43157];
  assign o[43156] = i[43156];
  assign o[43155] = i[43155];
  assign o[43154] = i[43154];
  assign o[43153] = i[43153];
  assign o[43152] = i[43152];
  assign o[43151] = i[43151];
  assign o[43150] = i[43150];
  assign o[43149] = i[43149];
  assign o[43148] = i[43148];
  assign o[43147] = i[43147];
  assign o[43146] = i[43146];
  assign o[43145] = i[43145];
  assign o[43144] = i[43144];
  assign o[43143] = i[43143];
  assign o[43142] = i[43142];
  assign o[43141] = i[43141];
  assign o[43140] = i[43140];
  assign o[43139] = i[43139];
  assign o[43138] = i[43138];
  assign o[43137] = i[43137];
  assign o[43136] = i[43136];
  assign o[43135] = i[43135];
  assign o[43134] = i[43134];
  assign o[43133] = i[43133];
  assign o[43132] = i[43132];
  assign o[43131] = i[43131];
  assign o[43130] = i[43130];
  assign o[43129] = i[43129];
  assign o[43128] = i[43128];
  assign o[43127] = i[43127];
  assign o[43126] = i[43126];
  assign o[43125] = i[43125];
  assign o[43124] = i[43124];
  assign o[43123] = i[43123];
  assign o[43122] = i[43122];
  assign o[43121] = i[43121];
  assign o[43120] = i[43120];
  assign o[43119] = i[43119];
  assign o[43118] = i[43118];
  assign o[43117] = i[43117];
  assign o[43116] = i[43116];
  assign o[43115] = i[43115];
  assign o[43114] = i[43114];
  assign o[43113] = i[43113];
  assign o[43112] = i[43112];
  assign o[43111] = i[43111];
  assign o[43110] = i[43110];
  assign o[43109] = i[43109];
  assign o[43108] = i[43108];
  assign o[43107] = i[43107];
  assign o[43106] = i[43106];
  assign o[43105] = i[43105];
  assign o[43104] = i[43104];
  assign o[43103] = i[43103];
  assign o[43102] = i[43102];
  assign o[43101] = i[43101];
  assign o[43100] = i[43100];
  assign o[43099] = i[43099];
  assign o[43098] = i[43098];
  assign o[43097] = i[43097];
  assign o[43096] = i[43096];
  assign o[43095] = i[43095];
  assign o[43094] = i[43094];
  assign o[43093] = i[43093];
  assign o[43092] = i[43092];
  assign o[43091] = i[43091];
  assign o[43090] = i[43090];
  assign o[43089] = i[43089];
  assign o[43088] = i[43088];
  assign o[43087] = i[43087];
  assign o[43086] = i[43086];
  assign o[43085] = i[43085];
  assign o[43084] = i[43084];
  assign o[43083] = i[43083];
  assign o[43082] = i[43082];
  assign o[43081] = i[43081];
  assign o[43080] = i[43080];
  assign o[43079] = i[43079];
  assign o[43078] = i[43078];
  assign o[43077] = i[43077];
  assign o[43076] = i[43076];
  assign o[43075] = i[43075];
  assign o[43074] = i[43074];
  assign o[43073] = i[43073];
  assign o[43072] = i[43072];
  assign o[43071] = i[43071];
  assign o[43070] = i[43070];
  assign o[43069] = i[43069];
  assign o[43068] = i[43068];
  assign o[43067] = i[43067];
  assign o[43066] = i[43066];
  assign o[43065] = i[43065];
  assign o[43064] = i[43064];
  assign o[43063] = i[43063];
  assign o[43062] = i[43062];
  assign o[43061] = i[43061];
  assign o[43060] = i[43060];
  assign o[43059] = i[43059];
  assign o[43058] = i[43058];
  assign o[43057] = i[43057];
  assign o[43056] = i[43056];
  assign o[43055] = i[43055];
  assign o[43054] = i[43054];
  assign o[43053] = i[43053];
  assign o[43052] = i[43052];
  assign o[43051] = i[43051];
  assign o[43050] = i[43050];
  assign o[43049] = i[43049];
  assign o[43048] = i[43048];
  assign o[43047] = i[43047];
  assign o[43046] = i[43046];
  assign o[43045] = i[43045];
  assign o[43044] = i[43044];
  assign o[43043] = i[43043];
  assign o[43042] = i[43042];
  assign o[43041] = i[43041];
  assign o[43040] = i[43040];
  assign o[43039] = i[43039];
  assign o[43038] = i[43038];
  assign o[43037] = i[43037];
  assign o[43036] = i[43036];
  assign o[43035] = i[43035];
  assign o[43034] = i[43034];
  assign o[43033] = i[43033];
  assign o[43032] = i[43032];
  assign o[43031] = i[43031];
  assign o[43030] = i[43030];
  assign o[43029] = i[43029];
  assign o[43028] = i[43028];
  assign o[43027] = i[43027];
  assign o[43026] = i[43026];
  assign o[43025] = i[43025];
  assign o[43024] = i[43024];
  assign o[43023] = i[43023];
  assign o[43022] = i[43022];
  assign o[43021] = i[43021];
  assign o[43020] = i[43020];
  assign o[43019] = i[43019];
  assign o[43018] = i[43018];
  assign o[43017] = i[43017];
  assign o[43016] = i[43016];
  assign o[43015] = i[43015];
  assign o[43014] = i[43014];
  assign o[43013] = i[43013];
  assign o[43012] = i[43012];
  assign o[43011] = i[43011];
  assign o[43010] = i[43010];
  assign o[43009] = i[43009];
  assign o[43008] = i[43008];
  assign o[43007] = i[43007];
  assign o[43006] = i[43006];
  assign o[43005] = i[43005];
  assign o[43004] = i[43004];
  assign o[43003] = i[43003];
  assign o[43002] = i[43002];
  assign o[43001] = i[43001];
  assign o[43000] = i[43000];
  assign o[42999] = i[42999];
  assign o[42998] = i[42998];
  assign o[42997] = i[42997];
  assign o[42996] = i[42996];
  assign o[42995] = i[42995];
  assign o[42994] = i[42994];
  assign o[42993] = i[42993];
  assign o[42992] = i[42992];
  assign o[42991] = i[42991];
  assign o[42990] = i[42990];
  assign o[42989] = i[42989];
  assign o[42988] = i[42988];
  assign o[42987] = i[42987];
  assign o[42986] = i[42986];
  assign o[42985] = i[42985];
  assign o[42984] = i[42984];
  assign o[42983] = i[42983];
  assign o[42982] = i[42982];
  assign o[42981] = i[42981];
  assign o[42980] = i[42980];
  assign o[42979] = i[42979];
  assign o[42978] = i[42978];
  assign o[42977] = i[42977];
  assign o[42976] = i[42976];
  assign o[42975] = i[42975];
  assign o[42974] = i[42974];
  assign o[42973] = i[42973];
  assign o[42972] = i[42972];
  assign o[42971] = i[42971];
  assign o[42970] = i[42970];
  assign o[42969] = i[42969];
  assign o[42968] = i[42968];
  assign o[42967] = i[42967];
  assign o[42966] = i[42966];
  assign o[42965] = i[42965];
  assign o[42964] = i[42964];
  assign o[42963] = i[42963];
  assign o[42962] = i[42962];
  assign o[42961] = i[42961];
  assign o[42960] = i[42960];
  assign o[42959] = i[42959];
  assign o[42958] = i[42958];
  assign o[42957] = i[42957];
  assign o[42956] = i[42956];
  assign o[42955] = i[42955];
  assign o[42954] = i[42954];
  assign o[42953] = i[42953];
  assign o[42952] = i[42952];
  assign o[42951] = i[42951];
  assign o[42950] = i[42950];
  assign o[42949] = i[42949];
  assign o[42948] = i[42948];
  assign o[42947] = i[42947];
  assign o[42946] = i[42946];
  assign o[42945] = i[42945];
  assign o[42944] = i[42944];
  assign o[42943] = i[42943];
  assign o[42942] = i[42942];
  assign o[42941] = i[42941];
  assign o[42940] = i[42940];
  assign o[42939] = i[42939];
  assign o[42938] = i[42938];
  assign o[42937] = i[42937];
  assign o[42936] = i[42936];
  assign o[42935] = i[42935];
  assign o[42934] = i[42934];
  assign o[42933] = i[42933];
  assign o[42932] = i[42932];
  assign o[42931] = i[42931];
  assign o[42930] = i[42930];
  assign o[42929] = i[42929];
  assign o[42928] = i[42928];
  assign o[42927] = i[42927];
  assign o[42926] = i[42926];
  assign o[42925] = i[42925];
  assign o[42924] = i[42924];
  assign o[42923] = i[42923];
  assign o[42922] = i[42922];
  assign o[42921] = i[42921];
  assign o[42920] = i[42920];
  assign o[42919] = i[42919];
  assign o[42918] = i[42918];
  assign o[42917] = i[42917];
  assign o[42916] = i[42916];
  assign o[42915] = i[42915];
  assign o[42914] = i[42914];
  assign o[42913] = i[42913];
  assign o[42912] = i[42912];
  assign o[42911] = i[42911];
  assign o[42910] = i[42910];
  assign o[42909] = i[42909];
  assign o[42908] = i[42908];
  assign o[42907] = i[42907];
  assign o[42906] = i[42906];
  assign o[42905] = i[42905];
  assign o[42904] = i[42904];
  assign o[42903] = i[42903];
  assign o[42902] = i[42902];
  assign o[42901] = i[42901];
  assign o[42900] = i[42900];
  assign o[42899] = i[42899];
  assign o[42898] = i[42898];
  assign o[42897] = i[42897];
  assign o[42896] = i[42896];
  assign o[42895] = i[42895];
  assign o[42894] = i[42894];
  assign o[42893] = i[42893];
  assign o[42892] = i[42892];
  assign o[42891] = i[42891];
  assign o[42890] = i[42890];
  assign o[42889] = i[42889];
  assign o[42888] = i[42888];
  assign o[42887] = i[42887];
  assign o[42886] = i[42886];
  assign o[42885] = i[42885];
  assign o[42884] = i[42884];
  assign o[42883] = i[42883];
  assign o[42882] = i[42882];
  assign o[42881] = i[42881];
  assign o[42880] = i[42880];
  assign o[42879] = i[42879];
  assign o[42878] = i[42878];
  assign o[42877] = i[42877];
  assign o[42876] = i[42876];
  assign o[42875] = i[42875];
  assign o[42874] = i[42874];
  assign o[42873] = i[42873];
  assign o[42872] = i[42872];
  assign o[42871] = i[42871];
  assign o[42870] = i[42870];
  assign o[42869] = i[42869];
  assign o[42868] = i[42868];
  assign o[42867] = i[42867];
  assign o[42866] = i[42866];
  assign o[42865] = i[42865];
  assign o[42864] = i[42864];
  assign o[42863] = i[42863];
  assign o[42862] = i[42862];
  assign o[42861] = i[42861];
  assign o[42860] = i[42860];
  assign o[42859] = i[42859];
  assign o[42858] = i[42858];
  assign o[42857] = i[42857];
  assign o[42856] = i[42856];
  assign o[42855] = i[42855];
  assign o[42854] = i[42854];
  assign o[42853] = i[42853];
  assign o[42852] = i[42852];
  assign o[42851] = i[42851];
  assign o[42850] = i[42850];
  assign o[42849] = i[42849];
  assign o[42848] = i[42848];
  assign o[42847] = i[42847];
  assign o[42846] = i[42846];
  assign o[42845] = i[42845];
  assign o[42844] = i[42844];
  assign o[42843] = i[42843];
  assign o[42842] = i[42842];
  assign o[42841] = i[42841];
  assign o[42840] = i[42840];
  assign o[42839] = i[42839];
  assign o[42838] = i[42838];
  assign o[42837] = i[42837];
  assign o[42836] = i[42836];
  assign o[42835] = i[42835];
  assign o[42834] = i[42834];
  assign o[42833] = i[42833];
  assign o[42832] = i[42832];
  assign o[42831] = i[42831];
  assign o[42830] = i[42830];
  assign o[42829] = i[42829];
  assign o[42828] = i[42828];
  assign o[42827] = i[42827];
  assign o[42826] = i[42826];
  assign o[42825] = i[42825];
  assign o[42824] = i[42824];
  assign o[42823] = i[42823];
  assign o[42822] = i[42822];
  assign o[42821] = i[42821];
  assign o[42820] = i[42820];
  assign o[42819] = i[42819];
  assign o[42818] = i[42818];
  assign o[42817] = i[42817];
  assign o[42816] = i[42816];
  assign o[42815] = i[42815];
  assign o[42814] = i[42814];
  assign o[42813] = i[42813];
  assign o[42812] = i[42812];
  assign o[42811] = i[42811];
  assign o[42810] = i[42810];
  assign o[42809] = i[42809];
  assign o[42808] = i[42808];
  assign o[42807] = i[42807];
  assign o[42806] = i[42806];
  assign o[42805] = i[42805];
  assign o[42804] = i[42804];
  assign o[42803] = i[42803];
  assign o[42802] = i[42802];
  assign o[42801] = i[42801];
  assign o[42800] = i[42800];
  assign o[42799] = i[42799];
  assign o[42798] = i[42798];
  assign o[42797] = i[42797];
  assign o[42796] = i[42796];
  assign o[42795] = i[42795];
  assign o[42794] = i[42794];
  assign o[42793] = i[42793];
  assign o[42792] = i[42792];
  assign o[42791] = i[42791];
  assign o[42790] = i[42790];
  assign o[42789] = i[42789];
  assign o[42788] = i[42788];
  assign o[42787] = i[42787];
  assign o[42786] = i[42786];
  assign o[42785] = i[42785];
  assign o[42784] = i[42784];
  assign o[42783] = i[42783];
  assign o[42782] = i[42782];
  assign o[42781] = i[42781];
  assign o[42780] = i[42780];
  assign o[42779] = i[42779];
  assign o[42778] = i[42778];
  assign o[42777] = i[42777];
  assign o[42776] = i[42776];
  assign o[42775] = i[42775];
  assign o[42774] = i[42774];
  assign o[42773] = i[42773];
  assign o[42772] = i[42772];
  assign o[42771] = i[42771];
  assign o[42770] = i[42770];
  assign o[42769] = i[42769];
  assign o[42768] = i[42768];
  assign o[42767] = i[42767];
  assign o[42766] = i[42766];
  assign o[42765] = i[42765];
  assign o[42764] = i[42764];
  assign o[42763] = i[42763];
  assign o[42762] = i[42762];
  assign o[42761] = i[42761];
  assign o[42760] = i[42760];
  assign o[42759] = i[42759];
  assign o[42758] = i[42758];
  assign o[42757] = i[42757];
  assign o[42756] = i[42756];
  assign o[42755] = i[42755];
  assign o[42754] = i[42754];
  assign o[42753] = i[42753];
  assign o[42752] = i[42752];
  assign o[42751] = i[42751];
  assign o[42750] = i[42750];
  assign o[42749] = i[42749];
  assign o[42748] = i[42748];
  assign o[42747] = i[42747];
  assign o[42746] = i[42746];
  assign o[42745] = i[42745];
  assign o[42744] = i[42744];
  assign o[42743] = i[42743];
  assign o[42742] = i[42742];
  assign o[42741] = i[42741];
  assign o[42740] = i[42740];
  assign o[42739] = i[42739];
  assign o[42738] = i[42738];
  assign o[42737] = i[42737];
  assign o[42736] = i[42736];
  assign o[42735] = i[42735];
  assign o[42734] = i[42734];
  assign o[42733] = i[42733];
  assign o[42732] = i[42732];
  assign o[42731] = i[42731];
  assign o[42730] = i[42730];
  assign o[42729] = i[42729];
  assign o[42728] = i[42728];
  assign o[42727] = i[42727];
  assign o[42726] = i[42726];
  assign o[42725] = i[42725];
  assign o[42724] = i[42724];
  assign o[42723] = i[42723];
  assign o[42722] = i[42722];
  assign o[42721] = i[42721];
  assign o[42720] = i[42720];
  assign o[42719] = i[42719];
  assign o[42718] = i[42718];
  assign o[42717] = i[42717];
  assign o[42716] = i[42716];
  assign o[42715] = i[42715];
  assign o[42714] = i[42714];
  assign o[42713] = i[42713];
  assign o[42712] = i[42712];
  assign o[42711] = i[42711];
  assign o[42710] = i[42710];
  assign o[42709] = i[42709];
  assign o[42708] = i[42708];
  assign o[42707] = i[42707];
  assign o[42706] = i[42706];
  assign o[42705] = i[42705];
  assign o[42704] = i[42704];
  assign o[42703] = i[42703];
  assign o[42702] = i[42702];
  assign o[42701] = i[42701];
  assign o[42700] = i[42700];
  assign o[42699] = i[42699];
  assign o[42698] = i[42698];
  assign o[42697] = i[42697];
  assign o[42696] = i[42696];
  assign o[42695] = i[42695];
  assign o[42694] = i[42694];
  assign o[42693] = i[42693];
  assign o[42692] = i[42692];
  assign o[42691] = i[42691];
  assign o[42690] = i[42690];
  assign o[42689] = i[42689];
  assign o[42688] = i[42688];
  assign o[42687] = i[42687];
  assign o[42686] = i[42686];
  assign o[42685] = i[42685];
  assign o[42684] = i[42684];
  assign o[42683] = i[42683];
  assign o[42682] = i[42682];
  assign o[42681] = i[42681];
  assign o[42680] = i[42680];
  assign o[42679] = i[42679];
  assign o[42678] = i[42678];
  assign o[42677] = i[42677];
  assign o[42676] = i[42676];
  assign o[42675] = i[42675];
  assign o[42674] = i[42674];
  assign o[42673] = i[42673];
  assign o[42672] = i[42672];
  assign o[42671] = i[42671];
  assign o[42670] = i[42670];
  assign o[42669] = i[42669];
  assign o[42668] = i[42668];
  assign o[42667] = i[42667];
  assign o[42666] = i[42666];
  assign o[42665] = i[42665];
  assign o[42664] = i[42664];
  assign o[42663] = i[42663];
  assign o[42662] = i[42662];
  assign o[42661] = i[42661];
  assign o[42660] = i[42660];
  assign o[42659] = i[42659];
  assign o[42658] = i[42658];
  assign o[42657] = i[42657];
  assign o[42656] = i[42656];
  assign o[42655] = i[42655];
  assign o[42654] = i[42654];
  assign o[42653] = i[42653];
  assign o[42652] = i[42652];
  assign o[42651] = i[42651];
  assign o[42650] = i[42650];
  assign o[42649] = i[42649];
  assign o[42648] = i[42648];
  assign o[42647] = i[42647];
  assign o[42646] = i[42646];
  assign o[42645] = i[42645];
  assign o[42644] = i[42644];
  assign o[42643] = i[42643];
  assign o[42642] = i[42642];
  assign o[42641] = i[42641];
  assign o[42640] = i[42640];
  assign o[42639] = i[42639];
  assign o[42638] = i[42638];
  assign o[42637] = i[42637];
  assign o[42636] = i[42636];
  assign o[42635] = i[42635];
  assign o[42634] = i[42634];
  assign o[42633] = i[42633];
  assign o[42632] = i[42632];
  assign o[42631] = i[42631];
  assign o[42630] = i[42630];
  assign o[42629] = i[42629];
  assign o[42628] = i[42628];
  assign o[42627] = i[42627];
  assign o[42626] = i[42626];
  assign o[42625] = i[42625];
  assign o[42624] = i[42624];
  assign o[42623] = i[42623];
  assign o[42622] = i[42622];
  assign o[42621] = i[42621];
  assign o[42620] = i[42620];
  assign o[42619] = i[42619];
  assign o[42618] = i[42618];
  assign o[42617] = i[42617];
  assign o[42616] = i[42616];
  assign o[42615] = i[42615];
  assign o[42614] = i[42614];
  assign o[42613] = i[42613];
  assign o[42612] = i[42612];
  assign o[42611] = i[42611];
  assign o[42610] = i[42610];
  assign o[42609] = i[42609];
  assign o[42608] = i[42608];
  assign o[42607] = i[42607];
  assign o[42606] = i[42606];
  assign o[42605] = i[42605];
  assign o[42604] = i[42604];
  assign o[42603] = i[42603];
  assign o[42602] = i[42602];
  assign o[42601] = i[42601];
  assign o[42600] = i[42600];
  assign o[42599] = i[42599];
  assign o[42598] = i[42598];
  assign o[42597] = i[42597];
  assign o[42596] = i[42596];
  assign o[42595] = i[42595];
  assign o[42594] = i[42594];
  assign o[42593] = i[42593];
  assign o[42592] = i[42592];
  assign o[42591] = i[42591];
  assign o[42590] = i[42590];
  assign o[42589] = i[42589];
  assign o[42588] = i[42588];
  assign o[42587] = i[42587];
  assign o[42586] = i[42586];
  assign o[42585] = i[42585];
  assign o[42584] = i[42584];
  assign o[42583] = i[42583];
  assign o[42582] = i[42582];
  assign o[42581] = i[42581];
  assign o[42580] = i[42580];
  assign o[42579] = i[42579];
  assign o[42578] = i[42578];
  assign o[42577] = i[42577];
  assign o[42576] = i[42576];
  assign o[42575] = i[42575];
  assign o[42574] = i[42574];
  assign o[42573] = i[42573];
  assign o[42572] = i[42572];
  assign o[42571] = i[42571];
  assign o[42570] = i[42570];
  assign o[42569] = i[42569];
  assign o[42568] = i[42568];
  assign o[42567] = i[42567];
  assign o[42566] = i[42566];
  assign o[42565] = i[42565];
  assign o[42564] = i[42564];
  assign o[42563] = i[42563];
  assign o[42562] = i[42562];
  assign o[42561] = i[42561];
  assign o[42560] = i[42560];
  assign o[42559] = i[42559];
  assign o[42558] = i[42558];
  assign o[42557] = i[42557];
  assign o[42556] = i[42556];
  assign o[42555] = i[42555];
  assign o[42554] = i[42554];
  assign o[42553] = i[42553];
  assign o[42552] = i[42552];
  assign o[42551] = i[42551];
  assign o[42550] = i[42550];
  assign o[42549] = i[42549];
  assign o[42548] = i[42548];
  assign o[42547] = i[42547];
  assign o[42546] = i[42546];
  assign o[42545] = i[42545];
  assign o[42544] = i[42544];
  assign o[42543] = i[42543];
  assign o[42542] = i[42542];
  assign o[42541] = i[42541];
  assign o[42540] = i[42540];
  assign o[42539] = i[42539];
  assign o[42538] = i[42538];
  assign o[42537] = i[42537];
  assign o[42536] = i[42536];
  assign o[42535] = i[42535];
  assign o[42534] = i[42534];
  assign o[42533] = i[42533];
  assign o[42532] = i[42532];
  assign o[42531] = i[42531];
  assign o[42530] = i[42530];
  assign o[42529] = i[42529];
  assign o[42528] = i[42528];
  assign o[42527] = i[42527];
  assign o[42526] = i[42526];
  assign o[42525] = i[42525];
  assign o[42524] = i[42524];
  assign o[42523] = i[42523];
  assign o[42522] = i[42522];
  assign o[42521] = i[42521];
  assign o[42520] = i[42520];
  assign o[42519] = i[42519];
  assign o[42518] = i[42518];
  assign o[42517] = i[42517];
  assign o[42516] = i[42516];
  assign o[42515] = i[42515];
  assign o[42514] = i[42514];
  assign o[42513] = i[42513];
  assign o[42512] = i[42512];
  assign o[42511] = i[42511];
  assign o[42510] = i[42510];
  assign o[42509] = i[42509];
  assign o[42508] = i[42508];
  assign o[42507] = i[42507];
  assign o[42506] = i[42506];
  assign o[42505] = i[42505];
  assign o[42504] = i[42504];
  assign o[42503] = i[42503];
  assign o[42502] = i[42502];
  assign o[42501] = i[42501];
  assign o[42500] = i[42500];
  assign o[42499] = i[42499];
  assign o[42498] = i[42498];
  assign o[42497] = i[42497];
  assign o[42496] = i[42496];
  assign o[42495] = i[42495];
  assign o[42494] = i[42494];
  assign o[42493] = i[42493];
  assign o[42492] = i[42492];
  assign o[42491] = i[42491];
  assign o[42490] = i[42490];
  assign o[42489] = i[42489];
  assign o[42488] = i[42488];
  assign o[42487] = i[42487];
  assign o[42486] = i[42486];
  assign o[42485] = i[42485];
  assign o[42484] = i[42484];
  assign o[42483] = i[42483];
  assign o[42482] = i[42482];
  assign o[42481] = i[42481];
  assign o[42480] = i[42480];
  assign o[42479] = i[42479];
  assign o[42478] = i[42478];
  assign o[42477] = i[42477];
  assign o[42476] = i[42476];
  assign o[42475] = i[42475];
  assign o[42474] = i[42474];
  assign o[42473] = i[42473];
  assign o[42472] = i[42472];
  assign o[42471] = i[42471];
  assign o[42470] = i[42470];
  assign o[42469] = i[42469];
  assign o[42468] = i[42468];
  assign o[42467] = i[42467];
  assign o[42466] = i[42466];
  assign o[42465] = i[42465];
  assign o[42464] = i[42464];
  assign o[42463] = i[42463];
  assign o[42462] = i[42462];
  assign o[42461] = i[42461];
  assign o[42460] = i[42460];
  assign o[42459] = i[42459];
  assign o[42458] = i[42458];
  assign o[42457] = i[42457];
  assign o[42456] = i[42456];
  assign o[42455] = i[42455];
  assign o[42454] = i[42454];
  assign o[42453] = i[42453];
  assign o[42452] = i[42452];
  assign o[42451] = i[42451];
  assign o[42450] = i[42450];
  assign o[42449] = i[42449];
  assign o[42448] = i[42448];
  assign o[42447] = i[42447];
  assign o[42446] = i[42446];
  assign o[42445] = i[42445];
  assign o[42444] = i[42444];
  assign o[42443] = i[42443];
  assign o[42442] = i[42442];
  assign o[42441] = i[42441];
  assign o[42440] = i[42440];
  assign o[42439] = i[42439];
  assign o[42438] = i[42438];
  assign o[42437] = i[42437];
  assign o[42436] = i[42436];
  assign o[42435] = i[42435];
  assign o[42434] = i[42434];
  assign o[42433] = i[42433];
  assign o[42432] = i[42432];
  assign o[42431] = i[42431];
  assign o[42430] = i[42430];
  assign o[42429] = i[42429];
  assign o[42428] = i[42428];
  assign o[42427] = i[42427];
  assign o[42426] = i[42426];
  assign o[42425] = i[42425];
  assign o[42424] = i[42424];
  assign o[42423] = i[42423];
  assign o[42422] = i[42422];
  assign o[42421] = i[42421];
  assign o[42420] = i[42420];
  assign o[42419] = i[42419];
  assign o[42418] = i[42418];
  assign o[42417] = i[42417];
  assign o[42416] = i[42416];
  assign o[42415] = i[42415];
  assign o[42414] = i[42414];
  assign o[42413] = i[42413];
  assign o[42412] = i[42412];
  assign o[42411] = i[42411];
  assign o[42410] = i[42410];
  assign o[42409] = i[42409];
  assign o[42408] = i[42408];
  assign o[42407] = i[42407];
  assign o[42406] = i[42406];
  assign o[42405] = i[42405];
  assign o[42404] = i[42404];
  assign o[42403] = i[42403];
  assign o[42402] = i[42402];
  assign o[42401] = i[42401];
  assign o[42400] = i[42400];
  assign o[42399] = i[42399];
  assign o[42398] = i[42398];
  assign o[42397] = i[42397];
  assign o[42396] = i[42396];
  assign o[42395] = i[42395];
  assign o[42394] = i[42394];
  assign o[42393] = i[42393];
  assign o[42392] = i[42392];
  assign o[42391] = i[42391];
  assign o[42390] = i[42390];
  assign o[42389] = i[42389];
  assign o[42388] = i[42388];
  assign o[42387] = i[42387];
  assign o[42386] = i[42386];
  assign o[42385] = i[42385];
  assign o[42384] = i[42384];
  assign o[42383] = i[42383];
  assign o[42382] = i[42382];
  assign o[42381] = i[42381];
  assign o[42380] = i[42380];
  assign o[42379] = i[42379];
  assign o[42378] = i[42378];
  assign o[42377] = i[42377];
  assign o[42376] = i[42376];
  assign o[42375] = i[42375];
  assign o[42374] = i[42374];
  assign o[42373] = i[42373];
  assign o[42372] = i[42372];
  assign o[42371] = i[42371];
  assign o[42370] = i[42370];
  assign o[42369] = i[42369];
  assign o[42368] = i[42368];
  assign o[42367] = i[42367];
  assign o[42366] = i[42366];
  assign o[42365] = i[42365];
  assign o[42364] = i[42364];
  assign o[42363] = i[42363];
  assign o[42362] = i[42362];
  assign o[42361] = i[42361];
  assign o[42360] = i[42360];
  assign o[42359] = i[42359];
  assign o[42358] = i[42358];
  assign o[42357] = i[42357];
  assign o[42356] = i[42356];
  assign o[42355] = i[42355];
  assign o[42354] = i[42354];
  assign o[42353] = i[42353];
  assign o[42352] = i[42352];
  assign o[42351] = i[42351];
  assign o[42350] = i[42350];
  assign o[42349] = i[42349];
  assign o[42348] = i[42348];
  assign o[42347] = i[42347];
  assign o[42346] = i[42346];
  assign o[42345] = i[42345];
  assign o[42344] = i[42344];
  assign o[42343] = i[42343];
  assign o[42342] = i[42342];
  assign o[42341] = i[42341];
  assign o[42340] = i[42340];
  assign o[42339] = i[42339];
  assign o[42338] = i[42338];
  assign o[42337] = i[42337];
  assign o[42336] = i[42336];
  assign o[42335] = i[42335];
  assign o[42334] = i[42334];
  assign o[42333] = i[42333];
  assign o[42332] = i[42332];
  assign o[42331] = i[42331];
  assign o[42330] = i[42330];
  assign o[42329] = i[42329];
  assign o[42328] = i[42328];
  assign o[42327] = i[42327];
  assign o[42326] = i[42326];
  assign o[42325] = i[42325];
  assign o[42324] = i[42324];
  assign o[42323] = i[42323];
  assign o[42322] = i[42322];
  assign o[42321] = i[42321];
  assign o[42320] = i[42320];
  assign o[42319] = i[42319];
  assign o[42318] = i[42318];
  assign o[42317] = i[42317];
  assign o[42316] = i[42316];
  assign o[42315] = i[42315];
  assign o[42314] = i[42314];
  assign o[42313] = i[42313];
  assign o[42312] = i[42312];
  assign o[42311] = i[42311];
  assign o[42310] = i[42310];
  assign o[42309] = i[42309];
  assign o[42308] = i[42308];
  assign o[42307] = i[42307];
  assign o[42306] = i[42306];
  assign o[42305] = i[42305];
  assign o[42304] = i[42304];
  assign o[42303] = i[42303];
  assign o[42302] = i[42302];
  assign o[42301] = i[42301];
  assign o[42300] = i[42300];
  assign o[42299] = i[42299];
  assign o[42298] = i[42298];
  assign o[42297] = i[42297];
  assign o[42296] = i[42296];
  assign o[42295] = i[42295];
  assign o[42294] = i[42294];
  assign o[42293] = i[42293];
  assign o[42292] = i[42292];
  assign o[42291] = i[42291];
  assign o[42290] = i[42290];
  assign o[42289] = i[42289];
  assign o[42288] = i[42288];
  assign o[42287] = i[42287];
  assign o[42286] = i[42286];
  assign o[42285] = i[42285];
  assign o[42284] = i[42284];
  assign o[42283] = i[42283];
  assign o[42282] = i[42282];
  assign o[42281] = i[42281];
  assign o[42280] = i[42280];
  assign o[42279] = i[42279];
  assign o[42278] = i[42278];
  assign o[42277] = i[42277];
  assign o[42276] = i[42276];
  assign o[42275] = i[42275];
  assign o[42274] = i[42274];
  assign o[42273] = i[42273];
  assign o[42272] = i[42272];
  assign o[42271] = i[42271];
  assign o[42270] = i[42270];
  assign o[42269] = i[42269];
  assign o[42268] = i[42268];
  assign o[42267] = i[42267];
  assign o[42266] = i[42266];
  assign o[42265] = i[42265];
  assign o[42264] = i[42264];
  assign o[42263] = i[42263];
  assign o[42262] = i[42262];
  assign o[42261] = i[42261];
  assign o[42260] = i[42260];
  assign o[42259] = i[42259];
  assign o[42258] = i[42258];
  assign o[42257] = i[42257];
  assign o[42256] = i[42256];
  assign o[42255] = i[42255];
  assign o[42254] = i[42254];
  assign o[42253] = i[42253];
  assign o[42252] = i[42252];
  assign o[42251] = i[42251];
  assign o[42250] = i[42250];
  assign o[42249] = i[42249];
  assign o[42248] = i[42248];
  assign o[42247] = i[42247];
  assign o[42246] = i[42246];
  assign o[42245] = i[42245];
  assign o[42244] = i[42244];
  assign o[42243] = i[42243];
  assign o[42242] = i[42242];
  assign o[42241] = i[42241];
  assign o[42240] = i[42240];
  assign o[42239] = i[42239];
  assign o[42238] = i[42238];
  assign o[42237] = i[42237];
  assign o[42236] = i[42236];
  assign o[42235] = i[42235];
  assign o[42234] = i[42234];
  assign o[42233] = i[42233];
  assign o[42232] = i[42232];
  assign o[42231] = i[42231];
  assign o[42230] = i[42230];
  assign o[42229] = i[42229];
  assign o[42228] = i[42228];
  assign o[42227] = i[42227];
  assign o[42226] = i[42226];
  assign o[42225] = i[42225];
  assign o[42224] = i[42224];
  assign o[42223] = i[42223];
  assign o[42222] = i[42222];
  assign o[42221] = i[42221];
  assign o[42220] = i[42220];
  assign o[42219] = i[42219];
  assign o[42218] = i[42218];
  assign o[42217] = i[42217];
  assign o[42216] = i[42216];
  assign o[42215] = i[42215];
  assign o[42214] = i[42214];
  assign o[42213] = i[42213];
  assign o[42212] = i[42212];
  assign o[42211] = i[42211];
  assign o[42210] = i[42210];
  assign o[42209] = i[42209];
  assign o[42208] = i[42208];
  assign o[42207] = i[42207];
  assign o[42206] = i[42206];
  assign o[42205] = i[42205];
  assign o[42204] = i[42204];
  assign o[42203] = i[42203];
  assign o[42202] = i[42202];
  assign o[42201] = i[42201];
  assign o[42200] = i[42200];
  assign o[42199] = i[42199];
  assign o[42198] = i[42198];
  assign o[42197] = i[42197];
  assign o[42196] = i[42196];
  assign o[42195] = i[42195];
  assign o[42194] = i[42194];
  assign o[42193] = i[42193];
  assign o[42192] = i[42192];
  assign o[42191] = i[42191];
  assign o[42190] = i[42190];
  assign o[42189] = i[42189];
  assign o[42188] = i[42188];
  assign o[42187] = i[42187];
  assign o[42186] = i[42186];
  assign o[42185] = i[42185];
  assign o[42184] = i[42184];
  assign o[42183] = i[42183];
  assign o[42182] = i[42182];
  assign o[42181] = i[42181];
  assign o[42180] = i[42180];
  assign o[42179] = i[42179];
  assign o[42178] = i[42178];
  assign o[42177] = i[42177];
  assign o[42176] = i[42176];
  assign o[42175] = i[42175];
  assign o[42174] = i[42174];
  assign o[42173] = i[42173];
  assign o[42172] = i[42172];
  assign o[42171] = i[42171];
  assign o[42170] = i[42170];
  assign o[42169] = i[42169];
  assign o[42168] = i[42168];
  assign o[42167] = i[42167];
  assign o[42166] = i[42166];
  assign o[42165] = i[42165];
  assign o[42164] = i[42164];
  assign o[42163] = i[42163];
  assign o[42162] = i[42162];
  assign o[42161] = i[42161];
  assign o[42160] = i[42160];
  assign o[42159] = i[42159];
  assign o[42158] = i[42158];
  assign o[42157] = i[42157];
  assign o[42156] = i[42156];
  assign o[42155] = i[42155];
  assign o[42154] = i[42154];
  assign o[42153] = i[42153];
  assign o[42152] = i[42152];
  assign o[42151] = i[42151];
  assign o[42150] = i[42150];
  assign o[42149] = i[42149];
  assign o[42148] = i[42148];
  assign o[42147] = i[42147];
  assign o[42146] = i[42146];
  assign o[42145] = i[42145];
  assign o[42144] = i[42144];
  assign o[42143] = i[42143];
  assign o[42142] = i[42142];
  assign o[42141] = i[42141];
  assign o[42140] = i[42140];
  assign o[42139] = i[42139];
  assign o[42138] = i[42138];
  assign o[42137] = i[42137];
  assign o[42136] = i[42136];
  assign o[42135] = i[42135];
  assign o[42134] = i[42134];
  assign o[42133] = i[42133];
  assign o[42132] = i[42132];
  assign o[42131] = i[42131];
  assign o[42130] = i[42130];
  assign o[42129] = i[42129];
  assign o[42128] = i[42128];
  assign o[42127] = i[42127];
  assign o[42126] = i[42126];
  assign o[42125] = i[42125];
  assign o[42124] = i[42124];
  assign o[42123] = i[42123];
  assign o[42122] = i[42122];
  assign o[42121] = i[42121];
  assign o[42120] = i[42120];
  assign o[42119] = i[42119];
  assign o[42118] = i[42118];
  assign o[42117] = i[42117];
  assign o[42116] = i[42116];
  assign o[42115] = i[42115];
  assign o[42114] = i[42114];
  assign o[42113] = i[42113];
  assign o[42112] = i[42112];
  assign o[42111] = i[42111];
  assign o[42110] = i[42110];
  assign o[42109] = i[42109];
  assign o[42108] = i[42108];
  assign o[42107] = i[42107];
  assign o[42106] = i[42106];
  assign o[42105] = i[42105];
  assign o[42104] = i[42104];
  assign o[42103] = i[42103];
  assign o[42102] = i[42102];
  assign o[42101] = i[42101];
  assign o[42100] = i[42100];
  assign o[42099] = i[42099];
  assign o[42098] = i[42098];
  assign o[42097] = i[42097];
  assign o[42096] = i[42096];
  assign o[42095] = i[42095];
  assign o[42094] = i[42094];
  assign o[42093] = i[42093];
  assign o[42092] = i[42092];
  assign o[42091] = i[42091];
  assign o[42090] = i[42090];
  assign o[42089] = i[42089];
  assign o[42088] = i[42088];
  assign o[42087] = i[42087];
  assign o[42086] = i[42086];
  assign o[42085] = i[42085];
  assign o[42084] = i[42084];
  assign o[42083] = i[42083];
  assign o[42082] = i[42082];
  assign o[42081] = i[42081];
  assign o[42080] = i[42080];
  assign o[42079] = i[42079];
  assign o[42078] = i[42078];
  assign o[42077] = i[42077];
  assign o[42076] = i[42076];
  assign o[42075] = i[42075];
  assign o[42074] = i[42074];
  assign o[42073] = i[42073];
  assign o[42072] = i[42072];
  assign o[42071] = i[42071];
  assign o[42070] = i[42070];
  assign o[42069] = i[42069];
  assign o[42068] = i[42068];
  assign o[42067] = i[42067];
  assign o[42066] = i[42066];
  assign o[42065] = i[42065];
  assign o[42064] = i[42064];
  assign o[42063] = i[42063];
  assign o[42062] = i[42062];
  assign o[42061] = i[42061];
  assign o[42060] = i[42060];
  assign o[42059] = i[42059];
  assign o[42058] = i[42058];
  assign o[42057] = i[42057];
  assign o[42056] = i[42056];
  assign o[42055] = i[42055];
  assign o[42054] = i[42054];
  assign o[42053] = i[42053];
  assign o[42052] = i[42052];
  assign o[42051] = i[42051];
  assign o[42050] = i[42050];
  assign o[42049] = i[42049];
  assign o[42048] = i[42048];
  assign o[42047] = i[42047];
  assign o[42046] = i[42046];
  assign o[42045] = i[42045];
  assign o[42044] = i[42044];
  assign o[42043] = i[42043];
  assign o[42042] = i[42042];
  assign o[42041] = i[42041];
  assign o[42040] = i[42040];
  assign o[42039] = i[42039];
  assign o[42038] = i[42038];
  assign o[42037] = i[42037];
  assign o[42036] = i[42036];
  assign o[42035] = i[42035];
  assign o[42034] = i[42034];
  assign o[42033] = i[42033];
  assign o[42032] = i[42032];
  assign o[42031] = i[42031];
  assign o[42030] = i[42030];
  assign o[42029] = i[42029];
  assign o[42028] = i[42028];
  assign o[42027] = i[42027];
  assign o[42026] = i[42026];
  assign o[42025] = i[42025];
  assign o[42024] = i[42024];
  assign o[42023] = i[42023];
  assign o[42022] = i[42022];
  assign o[42021] = i[42021];
  assign o[42020] = i[42020];
  assign o[42019] = i[42019];
  assign o[42018] = i[42018];
  assign o[42017] = i[42017];
  assign o[42016] = i[42016];
  assign o[42015] = i[42015];
  assign o[42014] = i[42014];
  assign o[42013] = i[42013];
  assign o[42012] = i[42012];
  assign o[42011] = i[42011];
  assign o[42010] = i[42010];
  assign o[42009] = i[42009];
  assign o[42008] = i[42008];
  assign o[42007] = i[42007];
  assign o[42006] = i[42006];
  assign o[42005] = i[42005];
  assign o[42004] = i[42004];
  assign o[42003] = i[42003];
  assign o[42002] = i[42002];
  assign o[42001] = i[42001];
  assign o[42000] = i[42000];
  assign o[41999] = i[41999];
  assign o[41998] = i[41998];
  assign o[41997] = i[41997];
  assign o[41996] = i[41996];
  assign o[41995] = i[41995];
  assign o[41994] = i[41994];
  assign o[41993] = i[41993];
  assign o[41992] = i[41992];
  assign o[41991] = i[41991];
  assign o[41990] = i[41990];
  assign o[41989] = i[41989];
  assign o[41988] = i[41988];
  assign o[41987] = i[41987];
  assign o[41986] = i[41986];
  assign o[41985] = i[41985];
  assign o[41984] = i[41984];
  assign o[41983] = i[41983];
  assign o[41982] = i[41982];
  assign o[41981] = i[41981];
  assign o[41980] = i[41980];
  assign o[41979] = i[41979];
  assign o[41978] = i[41978];
  assign o[41977] = i[41977];
  assign o[41976] = i[41976];
  assign o[41975] = i[41975];
  assign o[41974] = i[41974];
  assign o[41973] = i[41973];
  assign o[41972] = i[41972];
  assign o[41971] = i[41971];
  assign o[41970] = i[41970];
  assign o[41969] = i[41969];
  assign o[41968] = i[41968];
  assign o[41967] = i[41967];
  assign o[41966] = i[41966];
  assign o[41965] = i[41965];
  assign o[41964] = i[41964];
  assign o[41963] = i[41963];
  assign o[41962] = i[41962];
  assign o[41961] = i[41961];
  assign o[41960] = i[41960];
  assign o[41959] = i[41959];
  assign o[41958] = i[41958];
  assign o[41957] = i[41957];
  assign o[41956] = i[41956];
  assign o[41955] = i[41955];
  assign o[41954] = i[41954];
  assign o[41953] = i[41953];
  assign o[41952] = i[41952];
  assign o[41951] = i[41951];
  assign o[41950] = i[41950];
  assign o[41949] = i[41949];
  assign o[41948] = i[41948];
  assign o[41947] = i[41947];
  assign o[41946] = i[41946];
  assign o[41945] = i[41945];
  assign o[41944] = i[41944];
  assign o[41943] = i[41943];
  assign o[41942] = i[41942];
  assign o[41941] = i[41941];
  assign o[41940] = i[41940];
  assign o[41939] = i[41939];
  assign o[41938] = i[41938];
  assign o[41937] = i[41937];
  assign o[41936] = i[41936];
  assign o[41935] = i[41935];
  assign o[41934] = i[41934];
  assign o[41933] = i[41933];
  assign o[41932] = i[41932];
  assign o[41931] = i[41931];
  assign o[41930] = i[41930];
  assign o[41929] = i[41929];
  assign o[41928] = i[41928];
  assign o[41927] = i[41927];
  assign o[41926] = i[41926];
  assign o[41925] = i[41925];
  assign o[41924] = i[41924];
  assign o[41923] = i[41923];
  assign o[41922] = i[41922];
  assign o[41921] = i[41921];
  assign o[41920] = i[41920];
  assign o[41919] = i[41919];
  assign o[41918] = i[41918];
  assign o[41917] = i[41917];
  assign o[41916] = i[41916];
  assign o[41915] = i[41915];
  assign o[41914] = i[41914];
  assign o[41913] = i[41913];
  assign o[41912] = i[41912];
  assign o[41911] = i[41911];
  assign o[41910] = i[41910];
  assign o[41909] = i[41909];
  assign o[41908] = i[41908];
  assign o[41907] = i[41907];
  assign o[41906] = i[41906];
  assign o[41905] = i[41905];
  assign o[41904] = i[41904];
  assign o[41903] = i[41903];
  assign o[41902] = i[41902];
  assign o[41901] = i[41901];
  assign o[41900] = i[41900];
  assign o[41899] = i[41899];
  assign o[41898] = i[41898];
  assign o[41897] = i[41897];
  assign o[41896] = i[41896];
  assign o[41895] = i[41895];
  assign o[41894] = i[41894];
  assign o[41893] = i[41893];
  assign o[41892] = i[41892];
  assign o[41891] = i[41891];
  assign o[41890] = i[41890];
  assign o[41889] = i[41889];
  assign o[41888] = i[41888];
  assign o[41887] = i[41887];
  assign o[41886] = i[41886];
  assign o[41885] = i[41885];
  assign o[41884] = i[41884];
  assign o[41883] = i[41883];
  assign o[41882] = i[41882];
  assign o[41881] = i[41881];
  assign o[41880] = i[41880];
  assign o[41879] = i[41879];
  assign o[41878] = i[41878];
  assign o[41877] = i[41877];
  assign o[41876] = i[41876];
  assign o[41875] = i[41875];
  assign o[41874] = i[41874];
  assign o[41873] = i[41873];
  assign o[41872] = i[41872];
  assign o[41871] = i[41871];
  assign o[41870] = i[41870];
  assign o[41869] = i[41869];
  assign o[41868] = i[41868];
  assign o[41867] = i[41867];
  assign o[41866] = i[41866];
  assign o[41865] = i[41865];
  assign o[41864] = i[41864];
  assign o[41863] = i[41863];
  assign o[41862] = i[41862];
  assign o[41861] = i[41861];
  assign o[41860] = i[41860];
  assign o[41859] = i[41859];
  assign o[41858] = i[41858];
  assign o[41857] = i[41857];
  assign o[41856] = i[41856];
  assign o[41855] = i[41855];
  assign o[41854] = i[41854];
  assign o[41853] = i[41853];
  assign o[41852] = i[41852];
  assign o[41851] = i[41851];
  assign o[41850] = i[41850];
  assign o[41849] = i[41849];
  assign o[41848] = i[41848];
  assign o[41847] = i[41847];
  assign o[41846] = i[41846];
  assign o[41845] = i[41845];
  assign o[41844] = i[41844];
  assign o[41843] = i[41843];
  assign o[41842] = i[41842];
  assign o[41841] = i[41841];
  assign o[41840] = i[41840];
  assign o[41839] = i[41839];
  assign o[41838] = i[41838];
  assign o[41837] = i[41837];
  assign o[41836] = i[41836];
  assign o[41835] = i[41835];
  assign o[41834] = i[41834];
  assign o[41833] = i[41833];
  assign o[41832] = i[41832];
  assign o[41831] = i[41831];
  assign o[41830] = i[41830];
  assign o[41829] = i[41829];
  assign o[41828] = i[41828];
  assign o[41827] = i[41827];
  assign o[41826] = i[41826];
  assign o[41825] = i[41825];
  assign o[41824] = i[41824];
  assign o[41823] = i[41823];
  assign o[41822] = i[41822];
  assign o[41821] = i[41821];
  assign o[41820] = i[41820];
  assign o[41819] = i[41819];
  assign o[41818] = i[41818];
  assign o[41817] = i[41817];
  assign o[41816] = i[41816];
  assign o[41815] = i[41815];
  assign o[41814] = i[41814];
  assign o[41813] = i[41813];
  assign o[41812] = i[41812];
  assign o[41811] = i[41811];
  assign o[41810] = i[41810];
  assign o[41809] = i[41809];
  assign o[41808] = i[41808];
  assign o[41807] = i[41807];
  assign o[41806] = i[41806];
  assign o[41805] = i[41805];
  assign o[41804] = i[41804];
  assign o[41803] = i[41803];
  assign o[41802] = i[41802];
  assign o[41801] = i[41801];
  assign o[41800] = i[41800];
  assign o[41799] = i[41799];
  assign o[41798] = i[41798];
  assign o[41797] = i[41797];
  assign o[41796] = i[41796];
  assign o[41795] = i[41795];
  assign o[41794] = i[41794];
  assign o[41793] = i[41793];
  assign o[41792] = i[41792];
  assign o[41791] = i[41791];
  assign o[41790] = i[41790];
  assign o[41789] = i[41789];
  assign o[41788] = i[41788];
  assign o[41787] = i[41787];
  assign o[41786] = i[41786];
  assign o[41785] = i[41785];
  assign o[41784] = i[41784];
  assign o[41783] = i[41783];
  assign o[41782] = i[41782];
  assign o[41781] = i[41781];
  assign o[41780] = i[41780];
  assign o[41779] = i[41779];
  assign o[41778] = i[41778];
  assign o[41777] = i[41777];
  assign o[41776] = i[41776];
  assign o[41775] = i[41775];
  assign o[41774] = i[41774];
  assign o[41773] = i[41773];
  assign o[41772] = i[41772];
  assign o[41771] = i[41771];
  assign o[41770] = i[41770];
  assign o[41769] = i[41769];
  assign o[41768] = i[41768];
  assign o[41767] = i[41767];
  assign o[41766] = i[41766];
  assign o[41765] = i[41765];
  assign o[41764] = i[41764];
  assign o[41763] = i[41763];
  assign o[41762] = i[41762];
  assign o[41761] = i[41761];
  assign o[41760] = i[41760];
  assign o[41759] = i[41759];
  assign o[41758] = i[41758];
  assign o[41757] = i[41757];
  assign o[41756] = i[41756];
  assign o[41755] = i[41755];
  assign o[41754] = i[41754];
  assign o[41753] = i[41753];
  assign o[41752] = i[41752];
  assign o[41751] = i[41751];
  assign o[41750] = i[41750];
  assign o[41749] = i[41749];
  assign o[41748] = i[41748];
  assign o[41747] = i[41747];
  assign o[41746] = i[41746];
  assign o[41745] = i[41745];
  assign o[41744] = i[41744];
  assign o[41743] = i[41743];
  assign o[41742] = i[41742];
  assign o[41741] = i[41741];
  assign o[41740] = i[41740];
  assign o[41739] = i[41739];
  assign o[41738] = i[41738];
  assign o[41737] = i[41737];
  assign o[41736] = i[41736];
  assign o[41735] = i[41735];
  assign o[41734] = i[41734];
  assign o[41733] = i[41733];
  assign o[41732] = i[41732];
  assign o[41731] = i[41731];
  assign o[41730] = i[41730];
  assign o[41729] = i[41729];
  assign o[41728] = i[41728];
  assign o[41727] = i[41727];
  assign o[41726] = i[41726];
  assign o[41725] = i[41725];
  assign o[41724] = i[41724];
  assign o[41723] = i[41723];
  assign o[41722] = i[41722];
  assign o[41721] = i[41721];
  assign o[41720] = i[41720];
  assign o[41719] = i[41719];
  assign o[41718] = i[41718];
  assign o[41717] = i[41717];
  assign o[41716] = i[41716];
  assign o[41715] = i[41715];
  assign o[41714] = i[41714];
  assign o[41713] = i[41713];
  assign o[41712] = i[41712];
  assign o[41711] = i[41711];
  assign o[41710] = i[41710];
  assign o[41709] = i[41709];
  assign o[41708] = i[41708];
  assign o[41707] = i[41707];
  assign o[41706] = i[41706];
  assign o[41705] = i[41705];
  assign o[41704] = i[41704];
  assign o[41703] = i[41703];
  assign o[41702] = i[41702];
  assign o[41701] = i[41701];
  assign o[41700] = i[41700];
  assign o[41699] = i[41699];
  assign o[41698] = i[41698];
  assign o[41697] = i[41697];
  assign o[41696] = i[41696];
  assign o[41695] = i[41695];
  assign o[41694] = i[41694];
  assign o[41693] = i[41693];
  assign o[41692] = i[41692];
  assign o[41691] = i[41691];
  assign o[41690] = i[41690];
  assign o[41689] = i[41689];
  assign o[41688] = i[41688];
  assign o[41687] = i[41687];
  assign o[41686] = i[41686];
  assign o[41685] = i[41685];
  assign o[41684] = i[41684];
  assign o[41683] = i[41683];
  assign o[41682] = i[41682];
  assign o[41681] = i[41681];
  assign o[41680] = i[41680];
  assign o[41679] = i[41679];
  assign o[41678] = i[41678];
  assign o[41677] = i[41677];
  assign o[41676] = i[41676];
  assign o[41675] = i[41675];
  assign o[41674] = i[41674];
  assign o[41673] = i[41673];
  assign o[41672] = i[41672];
  assign o[41671] = i[41671];
  assign o[41670] = i[41670];
  assign o[41669] = i[41669];
  assign o[41668] = i[41668];
  assign o[41667] = i[41667];
  assign o[41666] = i[41666];
  assign o[41665] = i[41665];
  assign o[41664] = i[41664];
  assign o[41663] = i[41663];
  assign o[41662] = i[41662];
  assign o[41661] = i[41661];
  assign o[41660] = i[41660];
  assign o[41659] = i[41659];
  assign o[41658] = i[41658];
  assign o[41657] = i[41657];
  assign o[41656] = i[41656];
  assign o[41655] = i[41655];
  assign o[41654] = i[41654];
  assign o[41653] = i[41653];
  assign o[41652] = i[41652];
  assign o[41651] = i[41651];
  assign o[41650] = i[41650];
  assign o[41649] = i[41649];
  assign o[41648] = i[41648];
  assign o[41647] = i[41647];
  assign o[41646] = i[41646];
  assign o[41645] = i[41645];
  assign o[41644] = i[41644];
  assign o[41643] = i[41643];
  assign o[41642] = i[41642];
  assign o[41641] = i[41641];
  assign o[41640] = i[41640];
  assign o[41639] = i[41639];
  assign o[41638] = i[41638];
  assign o[41637] = i[41637];
  assign o[41636] = i[41636];
  assign o[41635] = i[41635];
  assign o[41634] = i[41634];
  assign o[41633] = i[41633];
  assign o[41632] = i[41632];
  assign o[41631] = i[41631];
  assign o[41630] = i[41630];
  assign o[41629] = i[41629];
  assign o[41628] = i[41628];
  assign o[41627] = i[41627];
  assign o[41626] = i[41626];
  assign o[41625] = i[41625];
  assign o[41624] = i[41624];
  assign o[41623] = i[41623];
  assign o[41622] = i[41622];
  assign o[41621] = i[41621];
  assign o[41620] = i[41620];
  assign o[41619] = i[41619];
  assign o[41618] = i[41618];
  assign o[41617] = i[41617];
  assign o[41616] = i[41616];
  assign o[41615] = i[41615];
  assign o[41614] = i[41614];
  assign o[41613] = i[41613];
  assign o[41612] = i[41612];
  assign o[41611] = i[41611];
  assign o[41610] = i[41610];
  assign o[41609] = i[41609];
  assign o[41608] = i[41608];
  assign o[41607] = i[41607];
  assign o[41606] = i[41606];
  assign o[41605] = i[41605];
  assign o[41604] = i[41604];
  assign o[41603] = i[41603];
  assign o[41602] = i[41602];
  assign o[41601] = i[41601];
  assign o[41600] = i[41600];
  assign o[41599] = i[41599];
  assign o[41598] = i[41598];
  assign o[41597] = i[41597];
  assign o[41596] = i[41596];
  assign o[41595] = i[41595];
  assign o[41594] = i[41594];
  assign o[41593] = i[41593];
  assign o[41592] = i[41592];
  assign o[41591] = i[41591];
  assign o[41590] = i[41590];
  assign o[41589] = i[41589];
  assign o[41588] = i[41588];
  assign o[41587] = i[41587];
  assign o[41586] = i[41586];
  assign o[41585] = i[41585];
  assign o[41584] = i[41584];
  assign o[41583] = i[41583];
  assign o[41582] = i[41582];
  assign o[41581] = i[41581];
  assign o[41580] = i[41580];
  assign o[41579] = i[41579];
  assign o[41578] = i[41578];
  assign o[41577] = i[41577];
  assign o[41576] = i[41576];
  assign o[41575] = i[41575];
  assign o[41574] = i[41574];
  assign o[41573] = i[41573];
  assign o[41572] = i[41572];
  assign o[41571] = i[41571];
  assign o[41570] = i[41570];
  assign o[41569] = i[41569];
  assign o[41568] = i[41568];
  assign o[41567] = i[41567];
  assign o[41566] = i[41566];
  assign o[41565] = i[41565];
  assign o[41564] = i[41564];
  assign o[41563] = i[41563];
  assign o[41562] = i[41562];
  assign o[41561] = i[41561];
  assign o[41560] = i[41560];
  assign o[41559] = i[41559];
  assign o[41558] = i[41558];
  assign o[41557] = i[41557];
  assign o[41556] = i[41556];
  assign o[41555] = i[41555];
  assign o[41554] = i[41554];
  assign o[41553] = i[41553];
  assign o[41552] = i[41552];
  assign o[41551] = i[41551];
  assign o[41550] = i[41550];
  assign o[41549] = i[41549];
  assign o[41548] = i[41548];
  assign o[41547] = i[41547];
  assign o[41546] = i[41546];
  assign o[41545] = i[41545];
  assign o[41544] = i[41544];
  assign o[41543] = i[41543];
  assign o[41542] = i[41542];
  assign o[41541] = i[41541];
  assign o[41540] = i[41540];
  assign o[41539] = i[41539];
  assign o[41538] = i[41538];
  assign o[41537] = i[41537];
  assign o[41536] = i[41536];
  assign o[41535] = i[41535];
  assign o[41534] = i[41534];
  assign o[41533] = i[41533];
  assign o[41532] = i[41532];
  assign o[41531] = i[41531];
  assign o[41530] = i[41530];
  assign o[41529] = i[41529];
  assign o[41528] = i[41528];
  assign o[41527] = i[41527];
  assign o[41526] = i[41526];
  assign o[41525] = i[41525];
  assign o[41524] = i[41524];
  assign o[41523] = i[41523];
  assign o[41522] = i[41522];
  assign o[41521] = i[41521];
  assign o[41520] = i[41520];
  assign o[41519] = i[41519];
  assign o[41518] = i[41518];
  assign o[41517] = i[41517];
  assign o[41516] = i[41516];
  assign o[41515] = i[41515];
  assign o[41514] = i[41514];
  assign o[41513] = i[41513];
  assign o[41512] = i[41512];
  assign o[41511] = i[41511];
  assign o[41510] = i[41510];
  assign o[41509] = i[41509];
  assign o[41508] = i[41508];
  assign o[41507] = i[41507];
  assign o[41506] = i[41506];
  assign o[41505] = i[41505];
  assign o[41504] = i[41504];
  assign o[41503] = i[41503];
  assign o[41502] = i[41502];
  assign o[41501] = i[41501];
  assign o[41500] = i[41500];
  assign o[41499] = i[41499];
  assign o[41498] = i[41498];
  assign o[41497] = i[41497];
  assign o[41496] = i[41496];
  assign o[41495] = i[41495];
  assign o[41494] = i[41494];
  assign o[41493] = i[41493];
  assign o[41492] = i[41492];
  assign o[41491] = i[41491];
  assign o[41490] = i[41490];
  assign o[41489] = i[41489];
  assign o[41488] = i[41488];
  assign o[41487] = i[41487];
  assign o[41486] = i[41486];
  assign o[41485] = i[41485];
  assign o[41484] = i[41484];
  assign o[41483] = i[41483];
  assign o[41482] = i[41482];
  assign o[41481] = i[41481];
  assign o[41480] = i[41480];
  assign o[41479] = i[41479];
  assign o[41478] = i[41478];
  assign o[41477] = i[41477];
  assign o[41476] = i[41476];
  assign o[41475] = i[41475];
  assign o[41474] = i[41474];
  assign o[41473] = i[41473];
  assign o[41472] = i[41472];
  assign o[41471] = i[41471];
  assign o[41470] = i[41470];
  assign o[41469] = i[41469];
  assign o[41468] = i[41468];
  assign o[41467] = i[41467];
  assign o[41466] = i[41466];
  assign o[41465] = i[41465];
  assign o[41464] = i[41464];
  assign o[41463] = i[41463];
  assign o[41462] = i[41462];
  assign o[41461] = i[41461];
  assign o[41460] = i[41460];
  assign o[41459] = i[41459];
  assign o[41458] = i[41458];
  assign o[41457] = i[41457];
  assign o[41456] = i[41456];
  assign o[41455] = i[41455];
  assign o[41454] = i[41454];
  assign o[41453] = i[41453];
  assign o[41452] = i[41452];
  assign o[41451] = i[41451];
  assign o[41450] = i[41450];
  assign o[41449] = i[41449];
  assign o[41448] = i[41448];
  assign o[41447] = i[41447];
  assign o[41446] = i[41446];
  assign o[41445] = i[41445];
  assign o[41444] = i[41444];
  assign o[41443] = i[41443];
  assign o[41442] = i[41442];
  assign o[41441] = i[41441];
  assign o[41440] = i[41440];
  assign o[41439] = i[41439];
  assign o[41438] = i[41438];
  assign o[41437] = i[41437];
  assign o[41436] = i[41436];
  assign o[41435] = i[41435];
  assign o[41434] = i[41434];
  assign o[41433] = i[41433];
  assign o[41432] = i[41432];
  assign o[41431] = i[41431];
  assign o[41430] = i[41430];
  assign o[41429] = i[41429];
  assign o[41428] = i[41428];
  assign o[41427] = i[41427];
  assign o[41426] = i[41426];
  assign o[41425] = i[41425];
  assign o[41424] = i[41424];
  assign o[41423] = i[41423];
  assign o[41422] = i[41422];
  assign o[41421] = i[41421];
  assign o[41420] = i[41420];
  assign o[41419] = i[41419];
  assign o[41418] = i[41418];
  assign o[41417] = i[41417];
  assign o[41416] = i[41416];
  assign o[41415] = i[41415];
  assign o[41414] = i[41414];
  assign o[41413] = i[41413];
  assign o[41412] = i[41412];
  assign o[41411] = i[41411];
  assign o[41410] = i[41410];
  assign o[41409] = i[41409];
  assign o[41408] = i[41408];
  assign o[41407] = i[41407];
  assign o[41406] = i[41406];
  assign o[41405] = i[41405];
  assign o[41404] = i[41404];
  assign o[41403] = i[41403];
  assign o[41402] = i[41402];
  assign o[41401] = i[41401];
  assign o[41400] = i[41400];
  assign o[41399] = i[41399];
  assign o[41398] = i[41398];
  assign o[41397] = i[41397];
  assign o[41396] = i[41396];
  assign o[41395] = i[41395];
  assign o[41394] = i[41394];
  assign o[41393] = i[41393];
  assign o[41392] = i[41392];
  assign o[41391] = i[41391];
  assign o[41390] = i[41390];
  assign o[41389] = i[41389];
  assign o[41388] = i[41388];
  assign o[41387] = i[41387];
  assign o[41386] = i[41386];
  assign o[41385] = i[41385];
  assign o[41384] = i[41384];
  assign o[41383] = i[41383];
  assign o[41382] = i[41382];
  assign o[41381] = i[41381];
  assign o[41380] = i[41380];
  assign o[41379] = i[41379];
  assign o[41378] = i[41378];
  assign o[41377] = i[41377];
  assign o[41376] = i[41376];
  assign o[41375] = i[41375];
  assign o[41374] = i[41374];
  assign o[41373] = i[41373];
  assign o[41372] = i[41372];
  assign o[41371] = i[41371];
  assign o[41370] = i[41370];
  assign o[41369] = i[41369];
  assign o[41368] = i[41368];
  assign o[41367] = i[41367];
  assign o[41366] = i[41366];
  assign o[41365] = i[41365];
  assign o[41364] = i[41364];
  assign o[41363] = i[41363];
  assign o[41362] = i[41362];
  assign o[41361] = i[41361];
  assign o[41360] = i[41360];
  assign o[41359] = i[41359];
  assign o[41358] = i[41358];
  assign o[41357] = i[41357];
  assign o[41356] = i[41356];
  assign o[41355] = i[41355];
  assign o[41354] = i[41354];
  assign o[41353] = i[41353];
  assign o[41352] = i[41352];
  assign o[41351] = i[41351];
  assign o[41350] = i[41350];
  assign o[41349] = i[41349];
  assign o[41348] = i[41348];
  assign o[41347] = i[41347];
  assign o[41346] = i[41346];
  assign o[41345] = i[41345];
  assign o[41344] = i[41344];
  assign o[41343] = i[41343];
  assign o[41342] = i[41342];
  assign o[41341] = i[41341];
  assign o[41340] = i[41340];
  assign o[41339] = i[41339];
  assign o[41338] = i[41338];
  assign o[41337] = i[41337];
  assign o[41336] = i[41336];
  assign o[41335] = i[41335];
  assign o[41334] = i[41334];
  assign o[41333] = i[41333];
  assign o[41332] = i[41332];
  assign o[41331] = i[41331];
  assign o[41330] = i[41330];
  assign o[41329] = i[41329];
  assign o[41328] = i[41328];
  assign o[41327] = i[41327];
  assign o[41326] = i[41326];
  assign o[41325] = i[41325];
  assign o[41324] = i[41324];
  assign o[41323] = i[41323];
  assign o[41322] = i[41322];
  assign o[41321] = i[41321];
  assign o[41320] = i[41320];
  assign o[41319] = i[41319];
  assign o[41318] = i[41318];
  assign o[41317] = i[41317];
  assign o[41316] = i[41316];
  assign o[41315] = i[41315];
  assign o[41314] = i[41314];
  assign o[41313] = i[41313];
  assign o[41312] = i[41312];
  assign o[41311] = i[41311];
  assign o[41310] = i[41310];
  assign o[41309] = i[41309];
  assign o[41308] = i[41308];
  assign o[41307] = i[41307];
  assign o[41306] = i[41306];
  assign o[41305] = i[41305];
  assign o[41304] = i[41304];
  assign o[41303] = i[41303];
  assign o[41302] = i[41302];
  assign o[41301] = i[41301];
  assign o[41300] = i[41300];
  assign o[41299] = i[41299];
  assign o[41298] = i[41298];
  assign o[41297] = i[41297];
  assign o[41296] = i[41296];
  assign o[41295] = i[41295];
  assign o[41294] = i[41294];
  assign o[41293] = i[41293];
  assign o[41292] = i[41292];
  assign o[41291] = i[41291];
  assign o[41290] = i[41290];
  assign o[41289] = i[41289];
  assign o[41288] = i[41288];
  assign o[41287] = i[41287];
  assign o[41286] = i[41286];
  assign o[41285] = i[41285];
  assign o[41284] = i[41284];
  assign o[41283] = i[41283];
  assign o[41282] = i[41282];
  assign o[41281] = i[41281];
  assign o[41280] = i[41280];
  assign o[41279] = i[41279];
  assign o[41278] = i[41278];
  assign o[41277] = i[41277];
  assign o[41276] = i[41276];
  assign o[41275] = i[41275];
  assign o[41274] = i[41274];
  assign o[41273] = i[41273];
  assign o[41272] = i[41272];
  assign o[41271] = i[41271];
  assign o[41270] = i[41270];
  assign o[41269] = i[41269];
  assign o[41268] = i[41268];
  assign o[41267] = i[41267];
  assign o[41266] = i[41266];
  assign o[41265] = i[41265];
  assign o[41264] = i[41264];
  assign o[41263] = i[41263];
  assign o[41262] = i[41262];
  assign o[41261] = i[41261];
  assign o[41260] = i[41260];
  assign o[41259] = i[41259];
  assign o[41258] = i[41258];
  assign o[41257] = i[41257];
  assign o[41256] = i[41256];
  assign o[41255] = i[41255];
  assign o[41254] = i[41254];
  assign o[41253] = i[41253];
  assign o[41252] = i[41252];
  assign o[41251] = i[41251];
  assign o[41250] = i[41250];
  assign o[41249] = i[41249];
  assign o[41248] = i[41248];
  assign o[41247] = i[41247];
  assign o[41246] = i[41246];
  assign o[41245] = i[41245];
  assign o[41244] = i[41244];
  assign o[41243] = i[41243];
  assign o[41242] = i[41242];
  assign o[41241] = i[41241];
  assign o[41240] = i[41240];
  assign o[41239] = i[41239];
  assign o[41238] = i[41238];
  assign o[41237] = i[41237];
  assign o[41236] = i[41236];
  assign o[41235] = i[41235];
  assign o[41234] = i[41234];
  assign o[41233] = i[41233];
  assign o[41232] = i[41232];
  assign o[41231] = i[41231];
  assign o[41230] = i[41230];
  assign o[41229] = i[41229];
  assign o[41228] = i[41228];
  assign o[41227] = i[41227];
  assign o[41226] = i[41226];
  assign o[41225] = i[41225];
  assign o[41224] = i[41224];
  assign o[41223] = i[41223];
  assign o[41222] = i[41222];
  assign o[41221] = i[41221];
  assign o[41220] = i[41220];
  assign o[41219] = i[41219];
  assign o[41218] = i[41218];
  assign o[41217] = i[41217];
  assign o[41216] = i[41216];
  assign o[41215] = i[41215];
  assign o[41214] = i[41214];
  assign o[41213] = i[41213];
  assign o[41212] = i[41212];
  assign o[41211] = i[41211];
  assign o[41210] = i[41210];
  assign o[41209] = i[41209];
  assign o[41208] = i[41208];
  assign o[41207] = i[41207];
  assign o[41206] = i[41206];
  assign o[41205] = i[41205];
  assign o[41204] = i[41204];
  assign o[41203] = i[41203];
  assign o[41202] = i[41202];
  assign o[41201] = i[41201];
  assign o[41200] = i[41200];
  assign o[41199] = i[41199];
  assign o[41198] = i[41198];
  assign o[41197] = i[41197];
  assign o[41196] = i[41196];
  assign o[41195] = i[41195];
  assign o[41194] = i[41194];
  assign o[41193] = i[41193];
  assign o[41192] = i[41192];
  assign o[41191] = i[41191];
  assign o[41190] = i[41190];
  assign o[41189] = i[41189];
  assign o[41188] = i[41188];
  assign o[41187] = i[41187];
  assign o[41186] = i[41186];
  assign o[41185] = i[41185];
  assign o[41184] = i[41184];
  assign o[41183] = i[41183];
  assign o[41182] = i[41182];
  assign o[41181] = i[41181];
  assign o[41180] = i[41180];
  assign o[41179] = i[41179];
  assign o[41178] = i[41178];
  assign o[41177] = i[41177];
  assign o[41176] = i[41176];
  assign o[41175] = i[41175];
  assign o[41174] = i[41174];
  assign o[41173] = i[41173];
  assign o[41172] = i[41172];
  assign o[41171] = i[41171];
  assign o[41170] = i[41170];
  assign o[41169] = i[41169];
  assign o[41168] = i[41168];
  assign o[41167] = i[41167];
  assign o[41166] = i[41166];
  assign o[41165] = i[41165];
  assign o[41164] = i[41164];
  assign o[41163] = i[41163];
  assign o[41162] = i[41162];
  assign o[41161] = i[41161];
  assign o[41160] = i[41160];
  assign o[41159] = i[41159];
  assign o[41158] = i[41158];
  assign o[41157] = i[41157];
  assign o[41156] = i[41156];
  assign o[41155] = i[41155];
  assign o[41154] = i[41154];
  assign o[41153] = i[41153];
  assign o[41152] = i[41152];
  assign o[41151] = i[41151];
  assign o[41150] = i[41150];
  assign o[41149] = i[41149];
  assign o[41148] = i[41148];
  assign o[41147] = i[41147];
  assign o[41146] = i[41146];
  assign o[41145] = i[41145];
  assign o[41144] = i[41144];
  assign o[41143] = i[41143];
  assign o[41142] = i[41142];
  assign o[41141] = i[41141];
  assign o[41140] = i[41140];
  assign o[41139] = i[41139];
  assign o[41138] = i[41138];
  assign o[41137] = i[41137];
  assign o[41136] = i[41136];
  assign o[41135] = i[41135];
  assign o[41134] = i[41134];
  assign o[41133] = i[41133];
  assign o[41132] = i[41132];
  assign o[41131] = i[41131];
  assign o[41130] = i[41130];
  assign o[41129] = i[41129];
  assign o[41128] = i[41128];
  assign o[41127] = i[41127];
  assign o[41126] = i[41126];
  assign o[41125] = i[41125];
  assign o[41124] = i[41124];
  assign o[41123] = i[41123];
  assign o[41122] = i[41122];
  assign o[41121] = i[41121];
  assign o[41120] = i[41120];
  assign o[41119] = i[41119];
  assign o[41118] = i[41118];
  assign o[41117] = i[41117];
  assign o[41116] = i[41116];
  assign o[41115] = i[41115];
  assign o[41114] = i[41114];
  assign o[41113] = i[41113];
  assign o[41112] = i[41112];
  assign o[41111] = i[41111];
  assign o[41110] = i[41110];
  assign o[41109] = i[41109];
  assign o[41108] = i[41108];
  assign o[41107] = i[41107];
  assign o[41106] = i[41106];
  assign o[41105] = i[41105];
  assign o[41104] = i[41104];
  assign o[41103] = i[41103];
  assign o[41102] = i[41102];
  assign o[41101] = i[41101];
  assign o[41100] = i[41100];
  assign o[41099] = i[41099];
  assign o[41098] = i[41098];
  assign o[41097] = i[41097];
  assign o[41096] = i[41096];
  assign o[41095] = i[41095];
  assign o[41094] = i[41094];
  assign o[41093] = i[41093];
  assign o[41092] = i[41092];
  assign o[41091] = i[41091];
  assign o[41090] = i[41090];
  assign o[41089] = i[41089];
  assign o[41088] = i[41088];
  assign o[41087] = i[41087];
  assign o[41086] = i[41086];
  assign o[41085] = i[41085];
  assign o[41084] = i[41084];
  assign o[41083] = i[41083];
  assign o[41082] = i[41082];
  assign o[41081] = i[41081];
  assign o[41080] = i[41080];
  assign o[41079] = i[41079];
  assign o[41078] = i[41078];
  assign o[41077] = i[41077];
  assign o[41076] = i[41076];
  assign o[41075] = i[41075];
  assign o[41074] = i[41074];
  assign o[41073] = i[41073];
  assign o[41072] = i[41072];
  assign o[41071] = i[41071];
  assign o[41070] = i[41070];
  assign o[41069] = i[41069];
  assign o[41068] = i[41068];
  assign o[41067] = i[41067];
  assign o[41066] = i[41066];
  assign o[41065] = i[41065];
  assign o[41064] = i[41064];
  assign o[41063] = i[41063];
  assign o[41062] = i[41062];
  assign o[41061] = i[41061];
  assign o[41060] = i[41060];
  assign o[41059] = i[41059];
  assign o[41058] = i[41058];
  assign o[41057] = i[41057];
  assign o[41056] = i[41056];
  assign o[41055] = i[41055];
  assign o[41054] = i[41054];
  assign o[41053] = i[41053];
  assign o[41052] = i[41052];
  assign o[41051] = i[41051];
  assign o[41050] = i[41050];
  assign o[41049] = i[41049];
  assign o[41048] = i[41048];
  assign o[41047] = i[41047];
  assign o[41046] = i[41046];
  assign o[41045] = i[41045];
  assign o[41044] = i[41044];
  assign o[41043] = i[41043];
  assign o[41042] = i[41042];
  assign o[41041] = i[41041];
  assign o[41040] = i[41040];
  assign o[41039] = i[41039];
  assign o[41038] = i[41038];
  assign o[41037] = i[41037];
  assign o[41036] = i[41036];
  assign o[41035] = i[41035];
  assign o[41034] = i[41034];
  assign o[41033] = i[41033];
  assign o[41032] = i[41032];
  assign o[41031] = i[41031];
  assign o[41030] = i[41030];
  assign o[41029] = i[41029];
  assign o[41028] = i[41028];
  assign o[41027] = i[41027];
  assign o[41026] = i[41026];
  assign o[41025] = i[41025];
  assign o[41024] = i[41024];
  assign o[41023] = i[41023];
  assign o[41022] = i[41022];
  assign o[41021] = i[41021];
  assign o[41020] = i[41020];
  assign o[41019] = i[41019];
  assign o[41018] = i[41018];
  assign o[41017] = i[41017];
  assign o[41016] = i[41016];
  assign o[41015] = i[41015];
  assign o[41014] = i[41014];
  assign o[41013] = i[41013];
  assign o[41012] = i[41012];
  assign o[41011] = i[41011];
  assign o[41010] = i[41010];
  assign o[41009] = i[41009];
  assign o[41008] = i[41008];
  assign o[41007] = i[41007];
  assign o[41006] = i[41006];
  assign o[41005] = i[41005];
  assign o[41004] = i[41004];
  assign o[41003] = i[41003];
  assign o[41002] = i[41002];
  assign o[41001] = i[41001];
  assign o[41000] = i[41000];
  assign o[40999] = i[40999];
  assign o[40998] = i[40998];
  assign o[40997] = i[40997];
  assign o[40996] = i[40996];
  assign o[40995] = i[40995];
  assign o[40994] = i[40994];
  assign o[40993] = i[40993];
  assign o[40992] = i[40992];
  assign o[40991] = i[40991];
  assign o[40990] = i[40990];
  assign o[40989] = i[40989];
  assign o[40988] = i[40988];
  assign o[40987] = i[40987];
  assign o[40986] = i[40986];
  assign o[40985] = i[40985];
  assign o[40984] = i[40984];
  assign o[40983] = i[40983];
  assign o[40982] = i[40982];
  assign o[40981] = i[40981];
  assign o[40980] = i[40980];
  assign o[40979] = i[40979];
  assign o[40978] = i[40978];
  assign o[40977] = i[40977];
  assign o[40976] = i[40976];
  assign o[40975] = i[40975];
  assign o[40974] = i[40974];
  assign o[40973] = i[40973];
  assign o[40972] = i[40972];
  assign o[40971] = i[40971];
  assign o[40970] = i[40970];
  assign o[40969] = i[40969];
  assign o[40968] = i[40968];
  assign o[40967] = i[40967];
  assign o[40966] = i[40966];
  assign o[40965] = i[40965];
  assign o[40964] = i[40964];
  assign o[40963] = i[40963];
  assign o[40962] = i[40962];
  assign o[40961] = i[40961];
  assign o[40960] = i[40960];
  assign o[40959] = i[40959];
  assign o[40958] = i[40958];
  assign o[40957] = i[40957];
  assign o[40956] = i[40956];
  assign o[40955] = i[40955];
  assign o[40954] = i[40954];
  assign o[40953] = i[40953];
  assign o[40952] = i[40952];
  assign o[40951] = i[40951];
  assign o[40950] = i[40950];
  assign o[40949] = i[40949];
  assign o[40948] = i[40948];
  assign o[40947] = i[40947];
  assign o[40946] = i[40946];
  assign o[40945] = i[40945];
  assign o[40944] = i[40944];
  assign o[40943] = i[40943];
  assign o[40942] = i[40942];
  assign o[40941] = i[40941];
  assign o[40940] = i[40940];
  assign o[40939] = i[40939];
  assign o[40938] = i[40938];
  assign o[40937] = i[40937];
  assign o[40936] = i[40936];
  assign o[40935] = i[40935];
  assign o[40934] = i[40934];
  assign o[40933] = i[40933];
  assign o[40932] = i[40932];
  assign o[40931] = i[40931];
  assign o[40930] = i[40930];
  assign o[40929] = i[40929];
  assign o[40928] = i[40928];
  assign o[40927] = i[40927];
  assign o[40926] = i[40926];
  assign o[40925] = i[40925];
  assign o[40924] = i[40924];
  assign o[40923] = i[40923];
  assign o[40922] = i[40922];
  assign o[40921] = i[40921];
  assign o[40920] = i[40920];
  assign o[40919] = i[40919];
  assign o[40918] = i[40918];
  assign o[40917] = i[40917];
  assign o[40916] = i[40916];
  assign o[40915] = i[40915];
  assign o[40914] = i[40914];
  assign o[40913] = i[40913];
  assign o[40912] = i[40912];
  assign o[40911] = i[40911];
  assign o[40910] = i[40910];
  assign o[40909] = i[40909];
  assign o[40908] = i[40908];
  assign o[40907] = i[40907];
  assign o[40906] = i[40906];
  assign o[40905] = i[40905];
  assign o[40904] = i[40904];
  assign o[40903] = i[40903];
  assign o[40902] = i[40902];
  assign o[40901] = i[40901];
  assign o[40900] = i[40900];
  assign o[40899] = i[40899];
  assign o[40898] = i[40898];
  assign o[40897] = i[40897];
  assign o[40896] = i[40896];
  assign o[40895] = i[40895];
  assign o[40894] = i[40894];
  assign o[40893] = i[40893];
  assign o[40892] = i[40892];
  assign o[40891] = i[40891];
  assign o[40890] = i[40890];
  assign o[40889] = i[40889];
  assign o[40888] = i[40888];
  assign o[40887] = i[40887];
  assign o[40886] = i[40886];
  assign o[40885] = i[40885];
  assign o[40884] = i[40884];
  assign o[40883] = i[40883];
  assign o[40882] = i[40882];
  assign o[40881] = i[40881];
  assign o[40880] = i[40880];
  assign o[40879] = i[40879];
  assign o[40878] = i[40878];
  assign o[40877] = i[40877];
  assign o[40876] = i[40876];
  assign o[40875] = i[40875];
  assign o[40874] = i[40874];
  assign o[40873] = i[40873];
  assign o[40872] = i[40872];
  assign o[40871] = i[40871];
  assign o[40870] = i[40870];
  assign o[40869] = i[40869];
  assign o[40868] = i[40868];
  assign o[40867] = i[40867];
  assign o[40866] = i[40866];
  assign o[40865] = i[40865];
  assign o[40864] = i[40864];
  assign o[40863] = i[40863];
  assign o[40862] = i[40862];
  assign o[40861] = i[40861];
  assign o[40860] = i[40860];
  assign o[40859] = i[40859];
  assign o[40858] = i[40858];
  assign o[40857] = i[40857];
  assign o[40856] = i[40856];
  assign o[40855] = i[40855];
  assign o[40854] = i[40854];
  assign o[40853] = i[40853];
  assign o[40852] = i[40852];
  assign o[40851] = i[40851];
  assign o[40850] = i[40850];
  assign o[40849] = i[40849];
  assign o[40848] = i[40848];
  assign o[40847] = i[40847];
  assign o[40846] = i[40846];
  assign o[40845] = i[40845];
  assign o[40844] = i[40844];
  assign o[40843] = i[40843];
  assign o[40842] = i[40842];
  assign o[40841] = i[40841];
  assign o[40840] = i[40840];
  assign o[40839] = i[40839];
  assign o[40838] = i[40838];
  assign o[40837] = i[40837];
  assign o[40836] = i[40836];
  assign o[40835] = i[40835];
  assign o[40834] = i[40834];
  assign o[40833] = i[40833];
  assign o[40832] = i[40832];
  assign o[40831] = i[40831];
  assign o[40830] = i[40830];
  assign o[40829] = i[40829];
  assign o[40828] = i[40828];
  assign o[40827] = i[40827];
  assign o[40826] = i[40826];
  assign o[40825] = i[40825];
  assign o[40824] = i[40824];
  assign o[40823] = i[40823];
  assign o[40822] = i[40822];
  assign o[40821] = i[40821];
  assign o[40820] = i[40820];
  assign o[40819] = i[40819];
  assign o[40818] = i[40818];
  assign o[40817] = i[40817];
  assign o[40816] = i[40816];
  assign o[40815] = i[40815];
  assign o[40814] = i[40814];
  assign o[40813] = i[40813];
  assign o[40812] = i[40812];
  assign o[40811] = i[40811];
  assign o[40810] = i[40810];
  assign o[40809] = i[40809];
  assign o[40808] = i[40808];
  assign o[40807] = i[40807];
  assign o[40806] = i[40806];
  assign o[40805] = i[40805];
  assign o[40804] = i[40804];
  assign o[40803] = i[40803];
  assign o[40802] = i[40802];
  assign o[40801] = i[40801];
  assign o[40800] = i[40800];
  assign o[40799] = i[40799];
  assign o[40798] = i[40798];
  assign o[40797] = i[40797];
  assign o[40796] = i[40796];
  assign o[40795] = i[40795];
  assign o[40794] = i[40794];
  assign o[40793] = i[40793];
  assign o[40792] = i[40792];
  assign o[40791] = i[40791];
  assign o[40790] = i[40790];
  assign o[40789] = i[40789];
  assign o[40788] = i[40788];
  assign o[40787] = i[40787];
  assign o[40786] = i[40786];
  assign o[40785] = i[40785];
  assign o[40784] = i[40784];
  assign o[40783] = i[40783];
  assign o[40782] = i[40782];
  assign o[40781] = i[40781];
  assign o[40780] = i[40780];
  assign o[40779] = i[40779];
  assign o[40778] = i[40778];
  assign o[40777] = i[40777];
  assign o[40776] = i[40776];
  assign o[40775] = i[40775];
  assign o[40774] = i[40774];
  assign o[40773] = i[40773];
  assign o[40772] = i[40772];
  assign o[40771] = i[40771];
  assign o[40770] = i[40770];
  assign o[40769] = i[40769];
  assign o[40768] = i[40768];
  assign o[40767] = i[40767];
  assign o[40766] = i[40766];
  assign o[40765] = i[40765];
  assign o[40764] = i[40764];
  assign o[40763] = i[40763];
  assign o[40762] = i[40762];
  assign o[40761] = i[40761];
  assign o[40760] = i[40760];
  assign o[40759] = i[40759];
  assign o[40758] = i[40758];
  assign o[40757] = i[40757];
  assign o[40756] = i[40756];
  assign o[40755] = i[40755];
  assign o[40754] = i[40754];
  assign o[40753] = i[40753];
  assign o[40752] = i[40752];
  assign o[40751] = i[40751];
  assign o[40750] = i[40750];
  assign o[40749] = i[40749];
  assign o[40748] = i[40748];
  assign o[40747] = i[40747];
  assign o[40746] = i[40746];
  assign o[40745] = i[40745];
  assign o[40744] = i[40744];
  assign o[40743] = i[40743];
  assign o[40742] = i[40742];
  assign o[40741] = i[40741];
  assign o[40740] = i[40740];
  assign o[40739] = i[40739];
  assign o[40738] = i[40738];
  assign o[40737] = i[40737];
  assign o[40736] = i[40736];
  assign o[40735] = i[40735];
  assign o[40734] = i[40734];
  assign o[40733] = i[40733];
  assign o[40732] = i[40732];
  assign o[40731] = i[40731];
  assign o[40730] = i[40730];
  assign o[40729] = i[40729];
  assign o[40728] = i[40728];
  assign o[40727] = i[40727];
  assign o[40726] = i[40726];
  assign o[40725] = i[40725];
  assign o[40724] = i[40724];
  assign o[40723] = i[40723];
  assign o[40722] = i[40722];
  assign o[40721] = i[40721];
  assign o[40720] = i[40720];
  assign o[40719] = i[40719];
  assign o[40718] = i[40718];
  assign o[40717] = i[40717];
  assign o[40716] = i[40716];
  assign o[40715] = i[40715];
  assign o[40714] = i[40714];
  assign o[40713] = i[40713];
  assign o[40712] = i[40712];
  assign o[40711] = i[40711];
  assign o[40710] = i[40710];
  assign o[40709] = i[40709];
  assign o[40708] = i[40708];
  assign o[40707] = i[40707];
  assign o[40706] = i[40706];
  assign o[40705] = i[40705];
  assign o[40704] = i[40704];
  assign o[40703] = i[40703];
  assign o[40702] = i[40702];
  assign o[40701] = i[40701];
  assign o[40700] = i[40700];
  assign o[40699] = i[40699];
  assign o[40698] = i[40698];
  assign o[40697] = i[40697];
  assign o[40696] = i[40696];
  assign o[40695] = i[40695];
  assign o[40694] = i[40694];
  assign o[40693] = i[40693];
  assign o[40692] = i[40692];
  assign o[40691] = i[40691];
  assign o[40690] = i[40690];
  assign o[40689] = i[40689];
  assign o[40688] = i[40688];
  assign o[40687] = i[40687];
  assign o[40686] = i[40686];
  assign o[40685] = i[40685];
  assign o[40684] = i[40684];
  assign o[40683] = i[40683];
  assign o[40682] = i[40682];
  assign o[40681] = i[40681];
  assign o[40680] = i[40680];
  assign o[40679] = i[40679];
  assign o[40678] = i[40678];
  assign o[40677] = i[40677];
  assign o[40676] = i[40676];
  assign o[40675] = i[40675];
  assign o[40674] = i[40674];
  assign o[40673] = i[40673];
  assign o[40672] = i[40672];
  assign o[40671] = i[40671];
  assign o[40670] = i[40670];
  assign o[40669] = i[40669];
  assign o[40668] = i[40668];
  assign o[40667] = i[40667];
  assign o[40666] = i[40666];
  assign o[40665] = i[40665];
  assign o[40664] = i[40664];
  assign o[40663] = i[40663];
  assign o[40662] = i[40662];
  assign o[40661] = i[40661];
  assign o[40660] = i[40660];
  assign o[40659] = i[40659];
  assign o[40658] = i[40658];
  assign o[40657] = i[40657];
  assign o[40656] = i[40656];
  assign o[40655] = i[40655];
  assign o[40654] = i[40654];
  assign o[40653] = i[40653];
  assign o[40652] = i[40652];
  assign o[40651] = i[40651];
  assign o[40650] = i[40650];
  assign o[40649] = i[40649];
  assign o[40648] = i[40648];
  assign o[40647] = i[40647];
  assign o[40646] = i[40646];
  assign o[40645] = i[40645];
  assign o[40644] = i[40644];
  assign o[40643] = i[40643];
  assign o[40642] = i[40642];
  assign o[40641] = i[40641];
  assign o[40640] = i[40640];
  assign o[40639] = i[40639];
  assign o[40638] = i[40638];
  assign o[40637] = i[40637];
  assign o[40636] = i[40636];
  assign o[40635] = i[40635];
  assign o[40634] = i[40634];
  assign o[40633] = i[40633];
  assign o[40632] = i[40632];
  assign o[40631] = i[40631];
  assign o[40630] = i[40630];
  assign o[40629] = i[40629];
  assign o[40628] = i[40628];
  assign o[40627] = i[40627];
  assign o[40626] = i[40626];
  assign o[40625] = i[40625];
  assign o[40624] = i[40624];
  assign o[40623] = i[40623];
  assign o[40622] = i[40622];
  assign o[40621] = i[40621];
  assign o[40620] = i[40620];
  assign o[40619] = i[40619];
  assign o[40618] = i[40618];
  assign o[40617] = i[40617];
  assign o[40616] = i[40616];
  assign o[40615] = i[40615];
  assign o[40614] = i[40614];
  assign o[40613] = i[40613];
  assign o[40612] = i[40612];
  assign o[40611] = i[40611];
  assign o[40610] = i[40610];
  assign o[40609] = i[40609];
  assign o[40608] = i[40608];
  assign o[40607] = i[40607];
  assign o[40606] = i[40606];
  assign o[40605] = i[40605];
  assign o[40604] = i[40604];
  assign o[40603] = i[40603];
  assign o[40602] = i[40602];
  assign o[40601] = i[40601];
  assign o[40600] = i[40600];
  assign o[40599] = i[40599];
  assign o[40598] = i[40598];
  assign o[40597] = i[40597];
  assign o[40596] = i[40596];
  assign o[40595] = i[40595];
  assign o[40594] = i[40594];
  assign o[40593] = i[40593];
  assign o[40592] = i[40592];
  assign o[40591] = i[40591];
  assign o[40590] = i[40590];
  assign o[40589] = i[40589];
  assign o[40588] = i[40588];
  assign o[40587] = i[40587];
  assign o[40586] = i[40586];
  assign o[40585] = i[40585];
  assign o[40584] = i[40584];
  assign o[40583] = i[40583];
  assign o[40582] = i[40582];
  assign o[40581] = i[40581];
  assign o[40580] = i[40580];
  assign o[40579] = i[40579];
  assign o[40578] = i[40578];
  assign o[40577] = i[40577];
  assign o[40576] = i[40576];
  assign o[40575] = i[40575];
  assign o[40574] = i[40574];
  assign o[40573] = i[40573];
  assign o[40572] = i[40572];
  assign o[40571] = i[40571];
  assign o[40570] = i[40570];
  assign o[40569] = i[40569];
  assign o[40568] = i[40568];
  assign o[40567] = i[40567];
  assign o[40566] = i[40566];
  assign o[40565] = i[40565];
  assign o[40564] = i[40564];
  assign o[40563] = i[40563];
  assign o[40562] = i[40562];
  assign o[40561] = i[40561];
  assign o[40560] = i[40560];
  assign o[40559] = i[40559];
  assign o[40558] = i[40558];
  assign o[40557] = i[40557];
  assign o[40556] = i[40556];
  assign o[40555] = i[40555];
  assign o[40554] = i[40554];
  assign o[40553] = i[40553];
  assign o[40552] = i[40552];
  assign o[40551] = i[40551];
  assign o[40550] = i[40550];
  assign o[40549] = i[40549];
  assign o[40548] = i[40548];
  assign o[40547] = i[40547];
  assign o[40546] = i[40546];
  assign o[40545] = i[40545];
  assign o[40544] = i[40544];
  assign o[40543] = i[40543];
  assign o[40542] = i[40542];
  assign o[40541] = i[40541];
  assign o[40540] = i[40540];
  assign o[40539] = i[40539];
  assign o[40538] = i[40538];
  assign o[40537] = i[40537];
  assign o[40536] = i[40536];
  assign o[40535] = i[40535];
  assign o[40534] = i[40534];
  assign o[40533] = i[40533];
  assign o[40532] = i[40532];
  assign o[40531] = i[40531];
  assign o[40530] = i[40530];
  assign o[40529] = i[40529];
  assign o[40528] = i[40528];
  assign o[40527] = i[40527];
  assign o[40526] = i[40526];
  assign o[40525] = i[40525];
  assign o[40524] = i[40524];
  assign o[40523] = i[40523];
  assign o[40522] = i[40522];
  assign o[40521] = i[40521];
  assign o[40520] = i[40520];
  assign o[40519] = i[40519];
  assign o[40518] = i[40518];
  assign o[40517] = i[40517];
  assign o[40516] = i[40516];
  assign o[40515] = i[40515];
  assign o[40514] = i[40514];
  assign o[40513] = i[40513];
  assign o[40512] = i[40512];
  assign o[40511] = i[40511];
  assign o[40510] = i[40510];
  assign o[40509] = i[40509];
  assign o[40508] = i[40508];
  assign o[40507] = i[40507];
  assign o[40506] = i[40506];
  assign o[40505] = i[40505];
  assign o[40504] = i[40504];
  assign o[40503] = i[40503];
  assign o[40502] = i[40502];
  assign o[40501] = i[40501];
  assign o[40500] = i[40500];
  assign o[40499] = i[40499];
  assign o[40498] = i[40498];
  assign o[40497] = i[40497];
  assign o[40496] = i[40496];
  assign o[40495] = i[40495];
  assign o[40494] = i[40494];
  assign o[40493] = i[40493];
  assign o[40492] = i[40492];
  assign o[40491] = i[40491];
  assign o[40490] = i[40490];
  assign o[40489] = i[40489];
  assign o[40488] = i[40488];
  assign o[40487] = i[40487];
  assign o[40486] = i[40486];
  assign o[40485] = i[40485];
  assign o[40484] = i[40484];
  assign o[40483] = i[40483];
  assign o[40482] = i[40482];
  assign o[40481] = i[40481];
  assign o[40480] = i[40480];
  assign o[40479] = i[40479];
  assign o[40478] = i[40478];
  assign o[40477] = i[40477];
  assign o[40476] = i[40476];
  assign o[40475] = i[40475];
  assign o[40474] = i[40474];
  assign o[40473] = i[40473];
  assign o[40472] = i[40472];
  assign o[40471] = i[40471];
  assign o[40470] = i[40470];
  assign o[40469] = i[40469];
  assign o[40468] = i[40468];
  assign o[40467] = i[40467];
  assign o[40466] = i[40466];
  assign o[40465] = i[40465];
  assign o[40464] = i[40464];
  assign o[40463] = i[40463];
  assign o[40462] = i[40462];
  assign o[40461] = i[40461];
  assign o[40460] = i[40460];
  assign o[40459] = i[40459];
  assign o[40458] = i[40458];
  assign o[40457] = i[40457];
  assign o[40456] = i[40456];
  assign o[40455] = i[40455];
  assign o[40454] = i[40454];
  assign o[40453] = i[40453];
  assign o[40452] = i[40452];
  assign o[40451] = i[40451];
  assign o[40450] = i[40450];
  assign o[40449] = i[40449];
  assign o[40448] = i[40448];
  assign o[40447] = i[40447];
  assign o[40446] = i[40446];
  assign o[40445] = i[40445];
  assign o[40444] = i[40444];
  assign o[40443] = i[40443];
  assign o[40442] = i[40442];
  assign o[40441] = i[40441];
  assign o[40440] = i[40440];
  assign o[40439] = i[40439];
  assign o[40438] = i[40438];
  assign o[40437] = i[40437];
  assign o[40436] = i[40436];
  assign o[40435] = i[40435];
  assign o[40434] = i[40434];
  assign o[40433] = i[40433];
  assign o[40432] = i[40432];
  assign o[40431] = i[40431];
  assign o[40430] = i[40430];
  assign o[40429] = i[40429];
  assign o[40428] = i[40428];
  assign o[40427] = i[40427];
  assign o[40426] = i[40426];
  assign o[40425] = i[40425];
  assign o[40424] = i[40424];
  assign o[40423] = i[40423];
  assign o[40422] = i[40422];
  assign o[40421] = i[40421];
  assign o[40420] = i[40420];
  assign o[40419] = i[40419];
  assign o[40418] = i[40418];
  assign o[40417] = i[40417];
  assign o[40416] = i[40416];
  assign o[40415] = i[40415];
  assign o[40414] = i[40414];
  assign o[40413] = i[40413];
  assign o[40412] = i[40412];
  assign o[40411] = i[40411];
  assign o[40410] = i[40410];
  assign o[40409] = i[40409];
  assign o[40408] = i[40408];
  assign o[40407] = i[40407];
  assign o[40406] = i[40406];
  assign o[40405] = i[40405];
  assign o[40404] = i[40404];
  assign o[40403] = i[40403];
  assign o[40402] = i[40402];
  assign o[40401] = i[40401];
  assign o[40400] = i[40400];
  assign o[40399] = i[40399];
  assign o[40398] = i[40398];
  assign o[40397] = i[40397];
  assign o[40396] = i[40396];
  assign o[40395] = i[40395];
  assign o[40394] = i[40394];
  assign o[40393] = i[40393];
  assign o[40392] = i[40392];
  assign o[40391] = i[40391];
  assign o[40390] = i[40390];
  assign o[40389] = i[40389];
  assign o[40388] = i[40388];
  assign o[40387] = i[40387];
  assign o[40386] = i[40386];
  assign o[40385] = i[40385];
  assign o[40384] = i[40384];
  assign o[40383] = i[40383];
  assign o[40382] = i[40382];
  assign o[40381] = i[40381];
  assign o[40380] = i[40380];
  assign o[40379] = i[40379];
  assign o[40378] = i[40378];
  assign o[40377] = i[40377];
  assign o[40376] = i[40376];
  assign o[40375] = i[40375];
  assign o[40374] = i[40374];
  assign o[40373] = i[40373];
  assign o[40372] = i[40372];
  assign o[40371] = i[40371];
  assign o[40370] = i[40370];
  assign o[40369] = i[40369];
  assign o[40368] = i[40368];
  assign o[40367] = i[40367];
  assign o[40366] = i[40366];
  assign o[40365] = i[40365];
  assign o[40364] = i[40364];
  assign o[40363] = i[40363];
  assign o[40362] = i[40362];
  assign o[40361] = i[40361];
  assign o[40360] = i[40360];
  assign o[40359] = i[40359];
  assign o[40358] = i[40358];
  assign o[40357] = i[40357];
  assign o[40356] = i[40356];
  assign o[40355] = i[40355];
  assign o[40354] = i[40354];
  assign o[40353] = i[40353];
  assign o[40352] = i[40352];
  assign o[40351] = i[40351];
  assign o[40350] = i[40350];
  assign o[40349] = i[40349];
  assign o[40348] = i[40348];
  assign o[40347] = i[40347];
  assign o[40346] = i[40346];
  assign o[40345] = i[40345];
  assign o[40344] = i[40344];
  assign o[40343] = i[40343];
  assign o[40342] = i[40342];
  assign o[40341] = i[40341];
  assign o[40340] = i[40340];
  assign o[40339] = i[40339];
  assign o[40338] = i[40338];
  assign o[40337] = i[40337];
  assign o[40336] = i[40336];
  assign o[40335] = i[40335];
  assign o[40334] = i[40334];
  assign o[40333] = i[40333];
  assign o[40332] = i[40332];
  assign o[40331] = i[40331];
  assign o[40330] = i[40330];
  assign o[40329] = i[40329];
  assign o[40328] = i[40328];
  assign o[40327] = i[40327];
  assign o[40326] = i[40326];
  assign o[40325] = i[40325];
  assign o[40324] = i[40324];
  assign o[40323] = i[40323];
  assign o[40322] = i[40322];
  assign o[40321] = i[40321];
  assign o[40320] = i[40320];
  assign o[40319] = i[40319];
  assign o[40318] = i[40318];
  assign o[40317] = i[40317];
  assign o[40316] = i[40316];
  assign o[40315] = i[40315];
  assign o[40314] = i[40314];
  assign o[40313] = i[40313];
  assign o[40312] = i[40312];
  assign o[40311] = i[40311];
  assign o[40310] = i[40310];
  assign o[40309] = i[40309];
  assign o[40308] = i[40308];
  assign o[40307] = i[40307];
  assign o[40306] = i[40306];
  assign o[40305] = i[40305];
  assign o[40304] = i[40304];
  assign o[40303] = i[40303];
  assign o[40302] = i[40302];
  assign o[40301] = i[40301];
  assign o[40300] = i[40300];
  assign o[40299] = i[40299];
  assign o[40298] = i[40298];
  assign o[40297] = i[40297];
  assign o[40296] = i[40296];
  assign o[40295] = i[40295];
  assign o[40294] = i[40294];
  assign o[40293] = i[40293];
  assign o[40292] = i[40292];
  assign o[40291] = i[40291];
  assign o[40290] = i[40290];
  assign o[40289] = i[40289];
  assign o[40288] = i[40288];
  assign o[40287] = i[40287];
  assign o[40286] = i[40286];
  assign o[40285] = i[40285];
  assign o[40284] = i[40284];
  assign o[40283] = i[40283];
  assign o[40282] = i[40282];
  assign o[40281] = i[40281];
  assign o[40280] = i[40280];
  assign o[40279] = i[40279];
  assign o[40278] = i[40278];
  assign o[40277] = i[40277];
  assign o[40276] = i[40276];
  assign o[40275] = i[40275];
  assign o[40274] = i[40274];
  assign o[40273] = i[40273];
  assign o[40272] = i[40272];
  assign o[40271] = i[40271];
  assign o[40270] = i[40270];
  assign o[40269] = i[40269];
  assign o[40268] = i[40268];
  assign o[40267] = i[40267];
  assign o[40266] = i[40266];
  assign o[40265] = i[40265];
  assign o[40264] = i[40264];
  assign o[40263] = i[40263];
  assign o[40262] = i[40262];
  assign o[40261] = i[40261];
  assign o[40260] = i[40260];
  assign o[40259] = i[40259];
  assign o[40258] = i[40258];
  assign o[40257] = i[40257];
  assign o[40256] = i[40256];
  assign o[40255] = i[40255];
  assign o[40254] = i[40254];
  assign o[40253] = i[40253];
  assign o[40252] = i[40252];
  assign o[40251] = i[40251];
  assign o[40250] = i[40250];
  assign o[40249] = i[40249];
  assign o[40248] = i[40248];
  assign o[40247] = i[40247];
  assign o[40246] = i[40246];
  assign o[40245] = i[40245];
  assign o[40244] = i[40244];
  assign o[40243] = i[40243];
  assign o[40242] = i[40242];
  assign o[40241] = i[40241];
  assign o[40240] = i[40240];
  assign o[40239] = i[40239];
  assign o[40238] = i[40238];
  assign o[40237] = i[40237];
  assign o[40236] = i[40236];
  assign o[40235] = i[40235];
  assign o[40234] = i[40234];
  assign o[40233] = i[40233];
  assign o[40232] = i[40232];
  assign o[40231] = i[40231];
  assign o[40230] = i[40230];
  assign o[40229] = i[40229];
  assign o[40228] = i[40228];
  assign o[40227] = i[40227];
  assign o[40226] = i[40226];
  assign o[40225] = i[40225];
  assign o[40224] = i[40224];
  assign o[40223] = i[40223];
  assign o[40222] = i[40222];
  assign o[40221] = i[40221];
  assign o[40220] = i[40220];
  assign o[40219] = i[40219];
  assign o[40218] = i[40218];
  assign o[40217] = i[40217];
  assign o[40216] = i[40216];
  assign o[40215] = i[40215];
  assign o[40214] = i[40214];
  assign o[40213] = i[40213];
  assign o[40212] = i[40212];
  assign o[40211] = i[40211];
  assign o[40210] = i[40210];
  assign o[40209] = i[40209];
  assign o[40208] = i[40208];
  assign o[40207] = i[40207];
  assign o[40206] = i[40206];
  assign o[40205] = i[40205];
  assign o[40204] = i[40204];
  assign o[40203] = i[40203];
  assign o[40202] = i[40202];
  assign o[40201] = i[40201];
  assign o[40200] = i[40200];
  assign o[40199] = i[40199];
  assign o[40198] = i[40198];
  assign o[40197] = i[40197];
  assign o[40196] = i[40196];
  assign o[40195] = i[40195];
  assign o[40194] = i[40194];
  assign o[40193] = i[40193];
  assign o[40192] = i[40192];
  assign o[40191] = i[40191];
  assign o[40190] = i[40190];
  assign o[40189] = i[40189];
  assign o[40188] = i[40188];
  assign o[40187] = i[40187];
  assign o[40186] = i[40186];
  assign o[40185] = i[40185];
  assign o[40184] = i[40184];
  assign o[40183] = i[40183];
  assign o[40182] = i[40182];
  assign o[40181] = i[40181];
  assign o[40180] = i[40180];
  assign o[40179] = i[40179];
  assign o[40178] = i[40178];
  assign o[40177] = i[40177];
  assign o[40176] = i[40176];
  assign o[40175] = i[40175];
  assign o[40174] = i[40174];
  assign o[40173] = i[40173];
  assign o[40172] = i[40172];
  assign o[40171] = i[40171];
  assign o[40170] = i[40170];
  assign o[40169] = i[40169];
  assign o[40168] = i[40168];
  assign o[40167] = i[40167];
  assign o[40166] = i[40166];
  assign o[40165] = i[40165];
  assign o[40164] = i[40164];
  assign o[40163] = i[40163];
  assign o[40162] = i[40162];
  assign o[40161] = i[40161];
  assign o[40160] = i[40160];
  assign o[40159] = i[40159];
  assign o[40158] = i[40158];
  assign o[40157] = i[40157];
  assign o[40156] = i[40156];
  assign o[40155] = i[40155];
  assign o[40154] = i[40154];
  assign o[40153] = i[40153];
  assign o[40152] = i[40152];
  assign o[40151] = i[40151];
  assign o[40150] = i[40150];
  assign o[40149] = i[40149];
  assign o[40148] = i[40148];
  assign o[40147] = i[40147];
  assign o[40146] = i[40146];
  assign o[40145] = i[40145];
  assign o[40144] = i[40144];
  assign o[40143] = i[40143];
  assign o[40142] = i[40142];
  assign o[40141] = i[40141];
  assign o[40140] = i[40140];
  assign o[40139] = i[40139];
  assign o[40138] = i[40138];
  assign o[40137] = i[40137];
  assign o[40136] = i[40136];
  assign o[40135] = i[40135];
  assign o[40134] = i[40134];
  assign o[40133] = i[40133];
  assign o[40132] = i[40132];
  assign o[40131] = i[40131];
  assign o[40130] = i[40130];
  assign o[40129] = i[40129];
  assign o[40128] = i[40128];
  assign o[40127] = i[40127];
  assign o[40126] = i[40126];
  assign o[40125] = i[40125];
  assign o[40124] = i[40124];
  assign o[40123] = i[40123];
  assign o[40122] = i[40122];
  assign o[40121] = i[40121];
  assign o[40120] = i[40120];
  assign o[40119] = i[40119];
  assign o[40118] = i[40118];
  assign o[40117] = i[40117];
  assign o[40116] = i[40116];
  assign o[40115] = i[40115];
  assign o[40114] = i[40114];
  assign o[40113] = i[40113];
  assign o[40112] = i[40112];
  assign o[40111] = i[40111];
  assign o[40110] = i[40110];
  assign o[40109] = i[40109];
  assign o[40108] = i[40108];
  assign o[40107] = i[40107];
  assign o[40106] = i[40106];
  assign o[40105] = i[40105];
  assign o[40104] = i[40104];
  assign o[40103] = i[40103];
  assign o[40102] = i[40102];
  assign o[40101] = i[40101];
  assign o[40100] = i[40100];
  assign o[40099] = i[40099];
  assign o[40098] = i[40098];
  assign o[40097] = i[40097];
  assign o[40096] = i[40096];
  assign o[40095] = i[40095];
  assign o[40094] = i[40094];
  assign o[40093] = i[40093];
  assign o[40092] = i[40092];
  assign o[40091] = i[40091];
  assign o[40090] = i[40090];
  assign o[40089] = i[40089];
  assign o[40088] = i[40088];
  assign o[40087] = i[40087];
  assign o[40086] = i[40086];
  assign o[40085] = i[40085];
  assign o[40084] = i[40084];
  assign o[40083] = i[40083];
  assign o[40082] = i[40082];
  assign o[40081] = i[40081];
  assign o[40080] = i[40080];
  assign o[40079] = i[40079];
  assign o[40078] = i[40078];
  assign o[40077] = i[40077];
  assign o[40076] = i[40076];
  assign o[40075] = i[40075];
  assign o[40074] = i[40074];
  assign o[40073] = i[40073];
  assign o[40072] = i[40072];
  assign o[40071] = i[40071];
  assign o[40070] = i[40070];
  assign o[40069] = i[40069];
  assign o[40068] = i[40068];
  assign o[40067] = i[40067];
  assign o[40066] = i[40066];
  assign o[40065] = i[40065];
  assign o[40064] = i[40064];
  assign o[40063] = i[40063];
  assign o[40062] = i[40062];
  assign o[40061] = i[40061];
  assign o[40060] = i[40060];
  assign o[40059] = i[40059];
  assign o[40058] = i[40058];
  assign o[40057] = i[40057];
  assign o[40056] = i[40056];
  assign o[40055] = i[40055];
  assign o[40054] = i[40054];
  assign o[40053] = i[40053];
  assign o[40052] = i[40052];
  assign o[40051] = i[40051];
  assign o[40050] = i[40050];
  assign o[40049] = i[40049];
  assign o[40048] = i[40048];
  assign o[40047] = i[40047];
  assign o[40046] = i[40046];
  assign o[40045] = i[40045];
  assign o[40044] = i[40044];
  assign o[40043] = i[40043];
  assign o[40042] = i[40042];
  assign o[40041] = i[40041];
  assign o[40040] = i[40040];
  assign o[40039] = i[40039];
  assign o[40038] = i[40038];
  assign o[40037] = i[40037];
  assign o[40036] = i[40036];
  assign o[40035] = i[40035];
  assign o[40034] = i[40034];
  assign o[40033] = i[40033];
  assign o[40032] = i[40032];
  assign o[40031] = i[40031];
  assign o[40030] = i[40030];
  assign o[40029] = i[40029];
  assign o[40028] = i[40028];
  assign o[40027] = i[40027];
  assign o[40026] = i[40026];
  assign o[40025] = i[40025];
  assign o[40024] = i[40024];
  assign o[40023] = i[40023];
  assign o[40022] = i[40022];
  assign o[40021] = i[40021];
  assign o[40020] = i[40020];
  assign o[40019] = i[40019];
  assign o[40018] = i[40018];
  assign o[40017] = i[40017];
  assign o[40016] = i[40016];
  assign o[40015] = i[40015];
  assign o[40014] = i[40014];
  assign o[40013] = i[40013];
  assign o[40012] = i[40012];
  assign o[40011] = i[40011];
  assign o[40010] = i[40010];
  assign o[40009] = i[40009];
  assign o[40008] = i[40008];
  assign o[40007] = i[40007];
  assign o[40006] = i[40006];
  assign o[40005] = i[40005];
  assign o[40004] = i[40004];
  assign o[40003] = i[40003];
  assign o[40002] = i[40002];
  assign o[40001] = i[40001];
  assign o[40000] = i[40000];
  assign o[39999] = i[39999];
  assign o[39998] = i[39998];
  assign o[39997] = i[39997];
  assign o[39996] = i[39996];
  assign o[39995] = i[39995];
  assign o[39994] = i[39994];
  assign o[39993] = i[39993];
  assign o[39992] = i[39992];
  assign o[39991] = i[39991];
  assign o[39990] = i[39990];
  assign o[39989] = i[39989];
  assign o[39988] = i[39988];
  assign o[39987] = i[39987];
  assign o[39986] = i[39986];
  assign o[39985] = i[39985];
  assign o[39984] = i[39984];
  assign o[39983] = i[39983];
  assign o[39982] = i[39982];
  assign o[39981] = i[39981];
  assign o[39980] = i[39980];
  assign o[39979] = i[39979];
  assign o[39978] = i[39978];
  assign o[39977] = i[39977];
  assign o[39976] = i[39976];
  assign o[39975] = i[39975];
  assign o[39974] = i[39974];
  assign o[39973] = i[39973];
  assign o[39972] = i[39972];
  assign o[39971] = i[39971];
  assign o[39970] = i[39970];
  assign o[39969] = i[39969];
  assign o[39968] = i[39968];
  assign o[39967] = i[39967];
  assign o[39966] = i[39966];
  assign o[39965] = i[39965];
  assign o[39964] = i[39964];
  assign o[39963] = i[39963];
  assign o[39962] = i[39962];
  assign o[39961] = i[39961];
  assign o[39960] = i[39960];
  assign o[39959] = i[39959];
  assign o[39958] = i[39958];
  assign o[39957] = i[39957];
  assign o[39956] = i[39956];
  assign o[39955] = i[39955];
  assign o[39954] = i[39954];
  assign o[39953] = i[39953];
  assign o[39952] = i[39952];
  assign o[39951] = i[39951];
  assign o[39950] = i[39950];
  assign o[39949] = i[39949];
  assign o[39948] = i[39948];
  assign o[39947] = i[39947];
  assign o[39946] = i[39946];
  assign o[39945] = i[39945];
  assign o[39944] = i[39944];
  assign o[39943] = i[39943];
  assign o[39942] = i[39942];
  assign o[39941] = i[39941];
  assign o[39940] = i[39940];
  assign o[39939] = i[39939];
  assign o[39938] = i[39938];
  assign o[39937] = i[39937];
  assign o[39936] = i[39936];
  assign o[39935] = i[39935];
  assign o[39934] = i[39934];
  assign o[39933] = i[39933];
  assign o[39932] = i[39932];
  assign o[39931] = i[39931];
  assign o[39930] = i[39930];
  assign o[39929] = i[39929];
  assign o[39928] = i[39928];
  assign o[39927] = i[39927];
  assign o[39926] = i[39926];
  assign o[39925] = i[39925];
  assign o[39924] = i[39924];
  assign o[39923] = i[39923];
  assign o[39922] = i[39922];
  assign o[39921] = i[39921];
  assign o[39920] = i[39920];
  assign o[39919] = i[39919];
  assign o[39918] = i[39918];
  assign o[39917] = i[39917];
  assign o[39916] = i[39916];
  assign o[39915] = i[39915];
  assign o[39914] = i[39914];
  assign o[39913] = i[39913];
  assign o[39912] = i[39912];
  assign o[39911] = i[39911];
  assign o[39910] = i[39910];
  assign o[39909] = i[39909];
  assign o[39908] = i[39908];
  assign o[39907] = i[39907];
  assign o[39906] = i[39906];
  assign o[39905] = i[39905];
  assign o[39904] = i[39904];
  assign o[39903] = i[39903];
  assign o[39902] = i[39902];
  assign o[39901] = i[39901];
  assign o[39900] = i[39900];
  assign o[39899] = i[39899];
  assign o[39898] = i[39898];
  assign o[39897] = i[39897];
  assign o[39896] = i[39896];
  assign o[39895] = i[39895];
  assign o[39894] = i[39894];
  assign o[39893] = i[39893];
  assign o[39892] = i[39892];
  assign o[39891] = i[39891];
  assign o[39890] = i[39890];
  assign o[39889] = i[39889];
  assign o[39888] = i[39888];
  assign o[39887] = i[39887];
  assign o[39886] = i[39886];
  assign o[39885] = i[39885];
  assign o[39884] = i[39884];
  assign o[39883] = i[39883];
  assign o[39882] = i[39882];
  assign o[39881] = i[39881];
  assign o[39880] = i[39880];
  assign o[39879] = i[39879];
  assign o[39878] = i[39878];
  assign o[39877] = i[39877];
  assign o[39876] = i[39876];
  assign o[39875] = i[39875];
  assign o[39874] = i[39874];
  assign o[39873] = i[39873];
  assign o[39872] = i[39872];
  assign o[39871] = i[39871];
  assign o[39870] = i[39870];
  assign o[39869] = i[39869];
  assign o[39868] = i[39868];
  assign o[39867] = i[39867];
  assign o[39866] = i[39866];
  assign o[39865] = i[39865];
  assign o[39864] = i[39864];
  assign o[39863] = i[39863];
  assign o[39862] = i[39862];
  assign o[39861] = i[39861];
  assign o[39860] = i[39860];
  assign o[39859] = i[39859];
  assign o[39858] = i[39858];
  assign o[39857] = i[39857];
  assign o[39856] = i[39856];
  assign o[39855] = i[39855];
  assign o[39854] = i[39854];
  assign o[39853] = i[39853];
  assign o[39852] = i[39852];
  assign o[39851] = i[39851];
  assign o[39850] = i[39850];
  assign o[39849] = i[39849];
  assign o[39848] = i[39848];
  assign o[39847] = i[39847];
  assign o[39846] = i[39846];
  assign o[39845] = i[39845];
  assign o[39844] = i[39844];
  assign o[39843] = i[39843];
  assign o[39842] = i[39842];
  assign o[39841] = i[39841];
  assign o[39840] = i[39840];
  assign o[39839] = i[39839];
  assign o[39838] = i[39838];
  assign o[39837] = i[39837];
  assign o[39836] = i[39836];
  assign o[39835] = i[39835];
  assign o[39834] = i[39834];
  assign o[39833] = i[39833];
  assign o[39832] = i[39832];
  assign o[39831] = i[39831];
  assign o[39830] = i[39830];
  assign o[39829] = i[39829];
  assign o[39828] = i[39828];
  assign o[39827] = i[39827];
  assign o[39826] = i[39826];
  assign o[39825] = i[39825];
  assign o[39824] = i[39824];
  assign o[39823] = i[39823];
  assign o[39822] = i[39822];
  assign o[39821] = i[39821];
  assign o[39820] = i[39820];
  assign o[39819] = i[39819];
  assign o[39818] = i[39818];
  assign o[39817] = i[39817];
  assign o[39816] = i[39816];
  assign o[39815] = i[39815];
  assign o[39814] = i[39814];
  assign o[39813] = i[39813];
  assign o[39812] = i[39812];
  assign o[39811] = i[39811];
  assign o[39810] = i[39810];
  assign o[39809] = i[39809];
  assign o[39808] = i[39808];
  assign o[39807] = i[39807];
  assign o[39806] = i[39806];
  assign o[39805] = i[39805];
  assign o[39804] = i[39804];
  assign o[39803] = i[39803];
  assign o[39802] = i[39802];
  assign o[39801] = i[39801];
  assign o[39800] = i[39800];
  assign o[39799] = i[39799];
  assign o[39798] = i[39798];
  assign o[39797] = i[39797];
  assign o[39796] = i[39796];
  assign o[39795] = i[39795];
  assign o[39794] = i[39794];
  assign o[39793] = i[39793];
  assign o[39792] = i[39792];
  assign o[39791] = i[39791];
  assign o[39790] = i[39790];
  assign o[39789] = i[39789];
  assign o[39788] = i[39788];
  assign o[39787] = i[39787];
  assign o[39786] = i[39786];
  assign o[39785] = i[39785];
  assign o[39784] = i[39784];
  assign o[39783] = i[39783];
  assign o[39782] = i[39782];
  assign o[39781] = i[39781];
  assign o[39780] = i[39780];
  assign o[39779] = i[39779];
  assign o[39778] = i[39778];
  assign o[39777] = i[39777];
  assign o[39776] = i[39776];
  assign o[39775] = i[39775];
  assign o[39774] = i[39774];
  assign o[39773] = i[39773];
  assign o[39772] = i[39772];
  assign o[39771] = i[39771];
  assign o[39770] = i[39770];
  assign o[39769] = i[39769];
  assign o[39768] = i[39768];
  assign o[39767] = i[39767];
  assign o[39766] = i[39766];
  assign o[39765] = i[39765];
  assign o[39764] = i[39764];
  assign o[39763] = i[39763];
  assign o[39762] = i[39762];
  assign o[39761] = i[39761];
  assign o[39760] = i[39760];
  assign o[39759] = i[39759];
  assign o[39758] = i[39758];
  assign o[39757] = i[39757];
  assign o[39756] = i[39756];
  assign o[39755] = i[39755];
  assign o[39754] = i[39754];
  assign o[39753] = i[39753];
  assign o[39752] = i[39752];
  assign o[39751] = i[39751];
  assign o[39750] = i[39750];
  assign o[39749] = i[39749];
  assign o[39748] = i[39748];
  assign o[39747] = i[39747];
  assign o[39746] = i[39746];
  assign o[39745] = i[39745];
  assign o[39744] = i[39744];
  assign o[39743] = i[39743];
  assign o[39742] = i[39742];
  assign o[39741] = i[39741];
  assign o[39740] = i[39740];
  assign o[39739] = i[39739];
  assign o[39738] = i[39738];
  assign o[39737] = i[39737];
  assign o[39736] = i[39736];
  assign o[39735] = i[39735];
  assign o[39734] = i[39734];
  assign o[39733] = i[39733];
  assign o[39732] = i[39732];
  assign o[39731] = i[39731];
  assign o[39730] = i[39730];
  assign o[39729] = i[39729];
  assign o[39728] = i[39728];
  assign o[39727] = i[39727];
  assign o[39726] = i[39726];
  assign o[39725] = i[39725];
  assign o[39724] = i[39724];
  assign o[39723] = i[39723];
  assign o[39722] = i[39722];
  assign o[39721] = i[39721];
  assign o[39720] = i[39720];
  assign o[39719] = i[39719];
  assign o[39718] = i[39718];
  assign o[39717] = i[39717];
  assign o[39716] = i[39716];
  assign o[39715] = i[39715];
  assign o[39714] = i[39714];
  assign o[39713] = i[39713];
  assign o[39712] = i[39712];
  assign o[39711] = i[39711];
  assign o[39710] = i[39710];
  assign o[39709] = i[39709];
  assign o[39708] = i[39708];
  assign o[39707] = i[39707];
  assign o[39706] = i[39706];
  assign o[39705] = i[39705];
  assign o[39704] = i[39704];
  assign o[39703] = i[39703];
  assign o[39702] = i[39702];
  assign o[39701] = i[39701];
  assign o[39700] = i[39700];
  assign o[39699] = i[39699];
  assign o[39698] = i[39698];
  assign o[39697] = i[39697];
  assign o[39696] = i[39696];
  assign o[39695] = i[39695];
  assign o[39694] = i[39694];
  assign o[39693] = i[39693];
  assign o[39692] = i[39692];
  assign o[39691] = i[39691];
  assign o[39690] = i[39690];
  assign o[39689] = i[39689];
  assign o[39688] = i[39688];
  assign o[39687] = i[39687];
  assign o[39686] = i[39686];
  assign o[39685] = i[39685];
  assign o[39684] = i[39684];
  assign o[39683] = i[39683];
  assign o[39682] = i[39682];
  assign o[39681] = i[39681];
  assign o[39680] = i[39680];
  assign o[39679] = i[39679];
  assign o[39678] = i[39678];
  assign o[39677] = i[39677];
  assign o[39676] = i[39676];
  assign o[39675] = i[39675];
  assign o[39674] = i[39674];
  assign o[39673] = i[39673];
  assign o[39672] = i[39672];
  assign o[39671] = i[39671];
  assign o[39670] = i[39670];
  assign o[39669] = i[39669];
  assign o[39668] = i[39668];
  assign o[39667] = i[39667];
  assign o[39666] = i[39666];
  assign o[39665] = i[39665];
  assign o[39664] = i[39664];
  assign o[39663] = i[39663];
  assign o[39662] = i[39662];
  assign o[39661] = i[39661];
  assign o[39660] = i[39660];
  assign o[39659] = i[39659];
  assign o[39658] = i[39658];
  assign o[39657] = i[39657];
  assign o[39656] = i[39656];
  assign o[39655] = i[39655];
  assign o[39654] = i[39654];
  assign o[39653] = i[39653];
  assign o[39652] = i[39652];
  assign o[39651] = i[39651];
  assign o[39650] = i[39650];
  assign o[39649] = i[39649];
  assign o[39648] = i[39648];
  assign o[39647] = i[39647];
  assign o[39646] = i[39646];
  assign o[39645] = i[39645];
  assign o[39644] = i[39644];
  assign o[39643] = i[39643];
  assign o[39642] = i[39642];
  assign o[39641] = i[39641];
  assign o[39640] = i[39640];
  assign o[39639] = i[39639];
  assign o[39638] = i[39638];
  assign o[39637] = i[39637];
  assign o[39636] = i[39636];
  assign o[39635] = i[39635];
  assign o[39634] = i[39634];
  assign o[39633] = i[39633];
  assign o[39632] = i[39632];
  assign o[39631] = i[39631];
  assign o[39630] = i[39630];
  assign o[39629] = i[39629];
  assign o[39628] = i[39628];
  assign o[39627] = i[39627];
  assign o[39626] = i[39626];
  assign o[39625] = i[39625];
  assign o[39624] = i[39624];
  assign o[39623] = i[39623];
  assign o[39622] = i[39622];
  assign o[39621] = i[39621];
  assign o[39620] = i[39620];
  assign o[39619] = i[39619];
  assign o[39618] = i[39618];
  assign o[39617] = i[39617];
  assign o[39616] = i[39616];
  assign o[39615] = i[39615];
  assign o[39614] = i[39614];
  assign o[39613] = i[39613];
  assign o[39612] = i[39612];
  assign o[39611] = i[39611];
  assign o[39610] = i[39610];
  assign o[39609] = i[39609];
  assign o[39608] = i[39608];
  assign o[39607] = i[39607];
  assign o[39606] = i[39606];
  assign o[39605] = i[39605];
  assign o[39604] = i[39604];
  assign o[39603] = i[39603];
  assign o[39602] = i[39602];
  assign o[39601] = i[39601];
  assign o[39600] = i[39600];
  assign o[39599] = i[39599];
  assign o[39598] = i[39598];
  assign o[39597] = i[39597];
  assign o[39596] = i[39596];
  assign o[39595] = i[39595];
  assign o[39594] = i[39594];
  assign o[39593] = i[39593];
  assign o[39592] = i[39592];
  assign o[39591] = i[39591];
  assign o[39590] = i[39590];
  assign o[39589] = i[39589];
  assign o[39588] = i[39588];
  assign o[39587] = i[39587];
  assign o[39586] = i[39586];
  assign o[39585] = i[39585];
  assign o[39584] = i[39584];
  assign o[39583] = i[39583];
  assign o[39582] = i[39582];
  assign o[39581] = i[39581];
  assign o[39580] = i[39580];
  assign o[39579] = i[39579];
  assign o[39578] = i[39578];
  assign o[39577] = i[39577];
  assign o[39576] = i[39576];
  assign o[39575] = i[39575];
  assign o[39574] = i[39574];
  assign o[39573] = i[39573];
  assign o[39572] = i[39572];
  assign o[39571] = i[39571];
  assign o[39570] = i[39570];
  assign o[39569] = i[39569];
  assign o[39568] = i[39568];
  assign o[39567] = i[39567];
  assign o[39566] = i[39566];
  assign o[39565] = i[39565];
  assign o[39564] = i[39564];
  assign o[39563] = i[39563];
  assign o[39562] = i[39562];
  assign o[39561] = i[39561];
  assign o[39560] = i[39560];
  assign o[39559] = i[39559];
  assign o[39558] = i[39558];
  assign o[39557] = i[39557];
  assign o[39556] = i[39556];
  assign o[39555] = i[39555];
  assign o[39554] = i[39554];
  assign o[39553] = i[39553];
  assign o[39552] = i[39552];
  assign o[39551] = i[39551];
  assign o[39550] = i[39550];
  assign o[39549] = i[39549];
  assign o[39548] = i[39548];
  assign o[39547] = i[39547];
  assign o[39546] = i[39546];
  assign o[39545] = i[39545];
  assign o[39544] = i[39544];
  assign o[39543] = i[39543];
  assign o[39542] = i[39542];
  assign o[39541] = i[39541];
  assign o[39540] = i[39540];
  assign o[39539] = i[39539];
  assign o[39538] = i[39538];
  assign o[39537] = i[39537];
  assign o[39536] = i[39536];
  assign o[39535] = i[39535];
  assign o[39534] = i[39534];
  assign o[39533] = i[39533];
  assign o[39532] = i[39532];
  assign o[39531] = i[39531];
  assign o[39530] = i[39530];
  assign o[39529] = i[39529];
  assign o[39528] = i[39528];
  assign o[39527] = i[39527];
  assign o[39526] = i[39526];
  assign o[39525] = i[39525];
  assign o[39524] = i[39524];
  assign o[39523] = i[39523];
  assign o[39522] = i[39522];
  assign o[39521] = i[39521];
  assign o[39520] = i[39520];
  assign o[39519] = i[39519];
  assign o[39518] = i[39518];
  assign o[39517] = i[39517];
  assign o[39516] = i[39516];
  assign o[39515] = i[39515];
  assign o[39514] = i[39514];
  assign o[39513] = i[39513];
  assign o[39512] = i[39512];
  assign o[39511] = i[39511];
  assign o[39510] = i[39510];
  assign o[39509] = i[39509];
  assign o[39508] = i[39508];
  assign o[39507] = i[39507];
  assign o[39506] = i[39506];
  assign o[39505] = i[39505];
  assign o[39504] = i[39504];
  assign o[39503] = i[39503];
  assign o[39502] = i[39502];
  assign o[39501] = i[39501];
  assign o[39500] = i[39500];
  assign o[39499] = i[39499];
  assign o[39498] = i[39498];
  assign o[39497] = i[39497];
  assign o[39496] = i[39496];
  assign o[39495] = i[39495];
  assign o[39494] = i[39494];
  assign o[39493] = i[39493];
  assign o[39492] = i[39492];
  assign o[39491] = i[39491];
  assign o[39490] = i[39490];
  assign o[39489] = i[39489];
  assign o[39488] = i[39488];
  assign o[39487] = i[39487];
  assign o[39486] = i[39486];
  assign o[39485] = i[39485];
  assign o[39484] = i[39484];
  assign o[39483] = i[39483];
  assign o[39482] = i[39482];
  assign o[39481] = i[39481];
  assign o[39480] = i[39480];
  assign o[39479] = i[39479];
  assign o[39478] = i[39478];
  assign o[39477] = i[39477];
  assign o[39476] = i[39476];
  assign o[39475] = i[39475];
  assign o[39474] = i[39474];
  assign o[39473] = i[39473];
  assign o[39472] = i[39472];
  assign o[39471] = i[39471];
  assign o[39470] = i[39470];
  assign o[39469] = i[39469];
  assign o[39468] = i[39468];
  assign o[39467] = i[39467];
  assign o[39466] = i[39466];
  assign o[39465] = i[39465];
  assign o[39464] = i[39464];
  assign o[39463] = i[39463];
  assign o[39462] = i[39462];
  assign o[39461] = i[39461];
  assign o[39460] = i[39460];
  assign o[39459] = i[39459];
  assign o[39458] = i[39458];
  assign o[39457] = i[39457];
  assign o[39456] = i[39456];
  assign o[39455] = i[39455];
  assign o[39454] = i[39454];
  assign o[39453] = i[39453];
  assign o[39452] = i[39452];
  assign o[39451] = i[39451];
  assign o[39450] = i[39450];
  assign o[39449] = i[39449];
  assign o[39448] = i[39448];
  assign o[39447] = i[39447];
  assign o[39446] = i[39446];
  assign o[39445] = i[39445];
  assign o[39444] = i[39444];
  assign o[39443] = i[39443];
  assign o[39442] = i[39442];
  assign o[39441] = i[39441];
  assign o[39440] = i[39440];
  assign o[39439] = i[39439];
  assign o[39438] = i[39438];
  assign o[39437] = i[39437];
  assign o[39436] = i[39436];
  assign o[39435] = i[39435];
  assign o[39434] = i[39434];
  assign o[39433] = i[39433];
  assign o[39432] = i[39432];
  assign o[39431] = i[39431];
  assign o[39430] = i[39430];
  assign o[39429] = i[39429];
  assign o[39428] = i[39428];
  assign o[39427] = i[39427];
  assign o[39426] = i[39426];
  assign o[39425] = i[39425];
  assign o[39424] = i[39424];
  assign o[39423] = i[39423];
  assign o[39422] = i[39422];
  assign o[39421] = i[39421];
  assign o[39420] = i[39420];
  assign o[39419] = i[39419];
  assign o[39418] = i[39418];
  assign o[39417] = i[39417];
  assign o[39416] = i[39416];
  assign o[39415] = i[39415];
  assign o[39414] = i[39414];
  assign o[39413] = i[39413];
  assign o[39412] = i[39412];
  assign o[39411] = i[39411];
  assign o[39410] = i[39410];
  assign o[39409] = i[39409];
  assign o[39408] = i[39408];
  assign o[39407] = i[39407];
  assign o[39406] = i[39406];
  assign o[39405] = i[39405];
  assign o[39404] = i[39404];
  assign o[39403] = i[39403];
  assign o[39402] = i[39402];
  assign o[39401] = i[39401];
  assign o[39400] = i[39400];
  assign o[39399] = i[39399];
  assign o[39398] = i[39398];
  assign o[39397] = i[39397];
  assign o[39396] = i[39396];
  assign o[39395] = i[39395];
  assign o[39394] = i[39394];
  assign o[39393] = i[39393];
  assign o[39392] = i[39392];
  assign o[39391] = i[39391];
  assign o[39390] = i[39390];
  assign o[39389] = i[39389];
  assign o[39388] = i[39388];
  assign o[39387] = i[39387];
  assign o[39386] = i[39386];
  assign o[39385] = i[39385];
  assign o[39384] = i[39384];
  assign o[39383] = i[39383];
  assign o[39382] = i[39382];
  assign o[39381] = i[39381];
  assign o[39380] = i[39380];
  assign o[39379] = i[39379];
  assign o[39378] = i[39378];
  assign o[39377] = i[39377];
  assign o[39376] = i[39376];
  assign o[39375] = i[39375];
  assign o[39374] = i[39374];
  assign o[39373] = i[39373];
  assign o[39372] = i[39372];
  assign o[39371] = i[39371];
  assign o[39370] = i[39370];
  assign o[39369] = i[39369];
  assign o[39368] = i[39368];
  assign o[39367] = i[39367];
  assign o[39366] = i[39366];
  assign o[39365] = i[39365];
  assign o[39364] = i[39364];
  assign o[39363] = i[39363];
  assign o[39362] = i[39362];
  assign o[39361] = i[39361];
  assign o[39360] = i[39360];
  assign o[39359] = i[39359];
  assign o[39358] = i[39358];
  assign o[39357] = i[39357];
  assign o[39356] = i[39356];
  assign o[39355] = i[39355];
  assign o[39354] = i[39354];
  assign o[39353] = i[39353];
  assign o[39352] = i[39352];
  assign o[39351] = i[39351];
  assign o[39350] = i[39350];
  assign o[39349] = i[39349];
  assign o[39348] = i[39348];
  assign o[39347] = i[39347];
  assign o[39346] = i[39346];
  assign o[39345] = i[39345];
  assign o[39344] = i[39344];
  assign o[39343] = i[39343];
  assign o[39342] = i[39342];
  assign o[39341] = i[39341];
  assign o[39340] = i[39340];
  assign o[39339] = i[39339];
  assign o[39338] = i[39338];
  assign o[39337] = i[39337];
  assign o[39336] = i[39336];
  assign o[39335] = i[39335];
  assign o[39334] = i[39334];
  assign o[39333] = i[39333];
  assign o[39332] = i[39332];
  assign o[39331] = i[39331];
  assign o[39330] = i[39330];
  assign o[39329] = i[39329];
  assign o[39328] = i[39328];
  assign o[39327] = i[39327];
  assign o[39326] = i[39326];
  assign o[39325] = i[39325];
  assign o[39324] = i[39324];
  assign o[39323] = i[39323];
  assign o[39322] = i[39322];
  assign o[39321] = i[39321];
  assign o[39320] = i[39320];
  assign o[39319] = i[39319];
  assign o[39318] = i[39318];
  assign o[39317] = i[39317];
  assign o[39316] = i[39316];
  assign o[39315] = i[39315];
  assign o[39314] = i[39314];
  assign o[39313] = i[39313];
  assign o[39312] = i[39312];
  assign o[39311] = i[39311];
  assign o[39310] = i[39310];
  assign o[39309] = i[39309];
  assign o[39308] = i[39308];
  assign o[39307] = i[39307];
  assign o[39306] = i[39306];
  assign o[39305] = i[39305];
  assign o[39304] = i[39304];
  assign o[39303] = i[39303];
  assign o[39302] = i[39302];
  assign o[39301] = i[39301];
  assign o[39300] = i[39300];
  assign o[39299] = i[39299];
  assign o[39298] = i[39298];
  assign o[39297] = i[39297];
  assign o[39296] = i[39296];
  assign o[39295] = i[39295];
  assign o[39294] = i[39294];
  assign o[39293] = i[39293];
  assign o[39292] = i[39292];
  assign o[39291] = i[39291];
  assign o[39290] = i[39290];
  assign o[39289] = i[39289];
  assign o[39288] = i[39288];
  assign o[39287] = i[39287];
  assign o[39286] = i[39286];
  assign o[39285] = i[39285];
  assign o[39284] = i[39284];
  assign o[39283] = i[39283];
  assign o[39282] = i[39282];
  assign o[39281] = i[39281];
  assign o[39280] = i[39280];
  assign o[39279] = i[39279];
  assign o[39278] = i[39278];
  assign o[39277] = i[39277];
  assign o[39276] = i[39276];
  assign o[39275] = i[39275];
  assign o[39274] = i[39274];
  assign o[39273] = i[39273];
  assign o[39272] = i[39272];
  assign o[39271] = i[39271];
  assign o[39270] = i[39270];
  assign o[39269] = i[39269];
  assign o[39268] = i[39268];
  assign o[39267] = i[39267];
  assign o[39266] = i[39266];
  assign o[39265] = i[39265];
  assign o[39264] = i[39264];
  assign o[39263] = i[39263];
  assign o[39262] = i[39262];
  assign o[39261] = i[39261];
  assign o[39260] = i[39260];
  assign o[39259] = i[39259];
  assign o[39258] = i[39258];
  assign o[39257] = i[39257];
  assign o[39256] = i[39256];
  assign o[39255] = i[39255];
  assign o[39254] = i[39254];
  assign o[39253] = i[39253];
  assign o[39252] = i[39252];
  assign o[39251] = i[39251];
  assign o[39250] = i[39250];
  assign o[39249] = i[39249];
  assign o[39248] = i[39248];
  assign o[39247] = i[39247];
  assign o[39246] = i[39246];
  assign o[39245] = i[39245];
  assign o[39244] = i[39244];
  assign o[39243] = i[39243];
  assign o[39242] = i[39242];
  assign o[39241] = i[39241];
  assign o[39240] = i[39240];
  assign o[39239] = i[39239];
  assign o[39238] = i[39238];
  assign o[39237] = i[39237];
  assign o[39236] = i[39236];
  assign o[39235] = i[39235];
  assign o[39234] = i[39234];
  assign o[39233] = i[39233];
  assign o[39232] = i[39232];
  assign o[39231] = i[39231];
  assign o[39230] = i[39230];
  assign o[39229] = i[39229];
  assign o[39228] = i[39228];
  assign o[39227] = i[39227];
  assign o[39226] = i[39226];
  assign o[39225] = i[39225];
  assign o[39224] = i[39224];
  assign o[39223] = i[39223];
  assign o[39222] = i[39222];
  assign o[39221] = i[39221];
  assign o[39220] = i[39220];
  assign o[39219] = i[39219];
  assign o[39218] = i[39218];
  assign o[39217] = i[39217];
  assign o[39216] = i[39216];
  assign o[39215] = i[39215];
  assign o[39214] = i[39214];
  assign o[39213] = i[39213];
  assign o[39212] = i[39212];
  assign o[39211] = i[39211];
  assign o[39210] = i[39210];
  assign o[39209] = i[39209];
  assign o[39208] = i[39208];
  assign o[39207] = i[39207];
  assign o[39206] = i[39206];
  assign o[39205] = i[39205];
  assign o[39204] = i[39204];
  assign o[39203] = i[39203];
  assign o[39202] = i[39202];
  assign o[39201] = i[39201];
  assign o[39200] = i[39200];
  assign o[39199] = i[39199];
  assign o[39198] = i[39198];
  assign o[39197] = i[39197];
  assign o[39196] = i[39196];
  assign o[39195] = i[39195];
  assign o[39194] = i[39194];
  assign o[39193] = i[39193];
  assign o[39192] = i[39192];
  assign o[39191] = i[39191];
  assign o[39190] = i[39190];
  assign o[39189] = i[39189];
  assign o[39188] = i[39188];
  assign o[39187] = i[39187];
  assign o[39186] = i[39186];
  assign o[39185] = i[39185];
  assign o[39184] = i[39184];
  assign o[39183] = i[39183];
  assign o[39182] = i[39182];
  assign o[39181] = i[39181];
  assign o[39180] = i[39180];
  assign o[39179] = i[39179];
  assign o[39178] = i[39178];
  assign o[39177] = i[39177];
  assign o[39176] = i[39176];
  assign o[39175] = i[39175];
  assign o[39174] = i[39174];
  assign o[39173] = i[39173];
  assign o[39172] = i[39172];
  assign o[39171] = i[39171];
  assign o[39170] = i[39170];
  assign o[39169] = i[39169];
  assign o[39168] = i[39168];
  assign o[39167] = i[39167];
  assign o[39166] = i[39166];
  assign o[39165] = i[39165];
  assign o[39164] = i[39164];
  assign o[39163] = i[39163];
  assign o[39162] = i[39162];
  assign o[39161] = i[39161];
  assign o[39160] = i[39160];
  assign o[39159] = i[39159];
  assign o[39158] = i[39158];
  assign o[39157] = i[39157];
  assign o[39156] = i[39156];
  assign o[39155] = i[39155];
  assign o[39154] = i[39154];
  assign o[39153] = i[39153];
  assign o[39152] = i[39152];
  assign o[39151] = i[39151];
  assign o[39150] = i[39150];
  assign o[39149] = i[39149];
  assign o[39148] = i[39148];
  assign o[39147] = i[39147];
  assign o[39146] = i[39146];
  assign o[39145] = i[39145];
  assign o[39144] = i[39144];
  assign o[39143] = i[39143];
  assign o[39142] = i[39142];
  assign o[39141] = i[39141];
  assign o[39140] = i[39140];
  assign o[39139] = i[39139];
  assign o[39138] = i[39138];
  assign o[39137] = i[39137];
  assign o[39136] = i[39136];
  assign o[39135] = i[39135];
  assign o[39134] = i[39134];
  assign o[39133] = i[39133];
  assign o[39132] = i[39132];
  assign o[39131] = i[39131];
  assign o[39130] = i[39130];
  assign o[39129] = i[39129];
  assign o[39128] = i[39128];
  assign o[39127] = i[39127];
  assign o[39126] = i[39126];
  assign o[39125] = i[39125];
  assign o[39124] = i[39124];
  assign o[39123] = i[39123];
  assign o[39122] = i[39122];
  assign o[39121] = i[39121];
  assign o[39120] = i[39120];
  assign o[39119] = i[39119];
  assign o[39118] = i[39118];
  assign o[39117] = i[39117];
  assign o[39116] = i[39116];
  assign o[39115] = i[39115];
  assign o[39114] = i[39114];
  assign o[39113] = i[39113];
  assign o[39112] = i[39112];
  assign o[39111] = i[39111];
  assign o[39110] = i[39110];
  assign o[39109] = i[39109];
  assign o[39108] = i[39108];
  assign o[39107] = i[39107];
  assign o[39106] = i[39106];
  assign o[39105] = i[39105];
  assign o[39104] = i[39104];
  assign o[39103] = i[39103];
  assign o[39102] = i[39102];
  assign o[39101] = i[39101];
  assign o[39100] = i[39100];
  assign o[39099] = i[39099];
  assign o[39098] = i[39098];
  assign o[39097] = i[39097];
  assign o[39096] = i[39096];
  assign o[39095] = i[39095];
  assign o[39094] = i[39094];
  assign o[39093] = i[39093];
  assign o[39092] = i[39092];
  assign o[39091] = i[39091];
  assign o[39090] = i[39090];
  assign o[39089] = i[39089];
  assign o[39088] = i[39088];
  assign o[39087] = i[39087];
  assign o[39086] = i[39086];
  assign o[39085] = i[39085];
  assign o[39084] = i[39084];
  assign o[39083] = i[39083];
  assign o[39082] = i[39082];
  assign o[39081] = i[39081];
  assign o[39080] = i[39080];
  assign o[39079] = i[39079];
  assign o[39078] = i[39078];
  assign o[39077] = i[39077];
  assign o[39076] = i[39076];
  assign o[39075] = i[39075];
  assign o[39074] = i[39074];
  assign o[39073] = i[39073];
  assign o[39072] = i[39072];
  assign o[39071] = i[39071];
  assign o[39070] = i[39070];
  assign o[39069] = i[39069];
  assign o[39068] = i[39068];
  assign o[39067] = i[39067];
  assign o[39066] = i[39066];
  assign o[39065] = i[39065];
  assign o[39064] = i[39064];
  assign o[39063] = i[39063];
  assign o[39062] = i[39062];
  assign o[39061] = i[39061];
  assign o[39060] = i[39060];
  assign o[39059] = i[39059];
  assign o[39058] = i[39058];
  assign o[39057] = i[39057];
  assign o[39056] = i[39056];
  assign o[39055] = i[39055];
  assign o[39054] = i[39054];
  assign o[39053] = i[39053];
  assign o[39052] = i[39052];
  assign o[39051] = i[39051];
  assign o[39050] = i[39050];
  assign o[39049] = i[39049];
  assign o[39048] = i[39048];
  assign o[39047] = i[39047];
  assign o[39046] = i[39046];
  assign o[39045] = i[39045];
  assign o[39044] = i[39044];
  assign o[39043] = i[39043];
  assign o[39042] = i[39042];
  assign o[39041] = i[39041];
  assign o[39040] = i[39040];
  assign o[39039] = i[39039];
  assign o[39038] = i[39038];
  assign o[39037] = i[39037];
  assign o[39036] = i[39036];
  assign o[39035] = i[39035];
  assign o[39034] = i[39034];
  assign o[39033] = i[39033];
  assign o[39032] = i[39032];
  assign o[39031] = i[39031];
  assign o[39030] = i[39030];
  assign o[39029] = i[39029];
  assign o[39028] = i[39028];
  assign o[39027] = i[39027];
  assign o[39026] = i[39026];
  assign o[39025] = i[39025];
  assign o[39024] = i[39024];
  assign o[39023] = i[39023];
  assign o[39022] = i[39022];
  assign o[39021] = i[39021];
  assign o[39020] = i[39020];
  assign o[39019] = i[39019];
  assign o[39018] = i[39018];
  assign o[39017] = i[39017];
  assign o[39016] = i[39016];
  assign o[39015] = i[39015];
  assign o[39014] = i[39014];
  assign o[39013] = i[39013];
  assign o[39012] = i[39012];
  assign o[39011] = i[39011];
  assign o[39010] = i[39010];
  assign o[39009] = i[39009];
  assign o[39008] = i[39008];
  assign o[39007] = i[39007];
  assign o[39006] = i[39006];
  assign o[39005] = i[39005];
  assign o[39004] = i[39004];
  assign o[39003] = i[39003];
  assign o[39002] = i[39002];
  assign o[39001] = i[39001];
  assign o[39000] = i[39000];
  assign o[38999] = i[38999];
  assign o[38998] = i[38998];
  assign o[38997] = i[38997];
  assign o[38996] = i[38996];
  assign o[38995] = i[38995];
  assign o[38994] = i[38994];
  assign o[38993] = i[38993];
  assign o[38992] = i[38992];
  assign o[38991] = i[38991];
  assign o[38990] = i[38990];
  assign o[38989] = i[38989];
  assign o[38988] = i[38988];
  assign o[38987] = i[38987];
  assign o[38986] = i[38986];
  assign o[38985] = i[38985];
  assign o[38984] = i[38984];
  assign o[38983] = i[38983];
  assign o[38982] = i[38982];
  assign o[38981] = i[38981];
  assign o[38980] = i[38980];
  assign o[38979] = i[38979];
  assign o[38978] = i[38978];
  assign o[38977] = i[38977];
  assign o[38976] = i[38976];
  assign o[38975] = i[38975];
  assign o[38974] = i[38974];
  assign o[38973] = i[38973];
  assign o[38972] = i[38972];
  assign o[38971] = i[38971];
  assign o[38970] = i[38970];
  assign o[38969] = i[38969];
  assign o[38968] = i[38968];
  assign o[38967] = i[38967];
  assign o[38966] = i[38966];
  assign o[38965] = i[38965];
  assign o[38964] = i[38964];
  assign o[38963] = i[38963];
  assign o[38962] = i[38962];
  assign o[38961] = i[38961];
  assign o[38960] = i[38960];
  assign o[38959] = i[38959];
  assign o[38958] = i[38958];
  assign o[38957] = i[38957];
  assign o[38956] = i[38956];
  assign o[38955] = i[38955];
  assign o[38954] = i[38954];
  assign o[38953] = i[38953];
  assign o[38952] = i[38952];
  assign o[38951] = i[38951];
  assign o[38950] = i[38950];
  assign o[38949] = i[38949];
  assign o[38948] = i[38948];
  assign o[38947] = i[38947];
  assign o[38946] = i[38946];
  assign o[38945] = i[38945];
  assign o[38944] = i[38944];
  assign o[38943] = i[38943];
  assign o[38942] = i[38942];
  assign o[38941] = i[38941];
  assign o[38940] = i[38940];
  assign o[38939] = i[38939];
  assign o[38938] = i[38938];
  assign o[38937] = i[38937];
  assign o[38936] = i[38936];
  assign o[38935] = i[38935];
  assign o[38934] = i[38934];
  assign o[38933] = i[38933];
  assign o[38932] = i[38932];
  assign o[38931] = i[38931];
  assign o[38930] = i[38930];
  assign o[38929] = i[38929];
  assign o[38928] = i[38928];
  assign o[38927] = i[38927];
  assign o[38926] = i[38926];
  assign o[38925] = i[38925];
  assign o[38924] = i[38924];
  assign o[38923] = i[38923];
  assign o[38922] = i[38922];
  assign o[38921] = i[38921];
  assign o[38920] = i[38920];
  assign o[38919] = i[38919];
  assign o[38918] = i[38918];
  assign o[38917] = i[38917];
  assign o[38916] = i[38916];
  assign o[38915] = i[38915];
  assign o[38914] = i[38914];
  assign o[38913] = i[38913];
  assign o[38912] = i[38912];
  assign o[38911] = i[38911];
  assign o[38910] = i[38910];
  assign o[38909] = i[38909];
  assign o[38908] = i[38908];
  assign o[38907] = i[38907];
  assign o[38906] = i[38906];
  assign o[38905] = i[38905];
  assign o[38904] = i[38904];
  assign o[38903] = i[38903];
  assign o[38902] = i[38902];
  assign o[38901] = i[38901];
  assign o[38900] = i[38900];
  assign o[38899] = i[38899];
  assign o[38898] = i[38898];
  assign o[38897] = i[38897];
  assign o[38896] = i[38896];
  assign o[38895] = i[38895];
  assign o[38894] = i[38894];
  assign o[38893] = i[38893];
  assign o[38892] = i[38892];
  assign o[38891] = i[38891];
  assign o[38890] = i[38890];
  assign o[38889] = i[38889];
  assign o[38888] = i[38888];
  assign o[38887] = i[38887];
  assign o[38886] = i[38886];
  assign o[38885] = i[38885];
  assign o[38884] = i[38884];
  assign o[38883] = i[38883];
  assign o[38882] = i[38882];
  assign o[38881] = i[38881];
  assign o[38880] = i[38880];
  assign o[38879] = i[38879];
  assign o[38878] = i[38878];
  assign o[38877] = i[38877];
  assign o[38876] = i[38876];
  assign o[38875] = i[38875];
  assign o[38874] = i[38874];
  assign o[38873] = i[38873];
  assign o[38872] = i[38872];
  assign o[38871] = i[38871];
  assign o[38870] = i[38870];
  assign o[38869] = i[38869];
  assign o[38868] = i[38868];
  assign o[38867] = i[38867];
  assign o[38866] = i[38866];
  assign o[38865] = i[38865];
  assign o[38864] = i[38864];
  assign o[38863] = i[38863];
  assign o[38862] = i[38862];
  assign o[38861] = i[38861];
  assign o[38860] = i[38860];
  assign o[38859] = i[38859];
  assign o[38858] = i[38858];
  assign o[38857] = i[38857];
  assign o[38856] = i[38856];
  assign o[38855] = i[38855];
  assign o[38854] = i[38854];
  assign o[38853] = i[38853];
  assign o[38852] = i[38852];
  assign o[38851] = i[38851];
  assign o[38850] = i[38850];
  assign o[38849] = i[38849];
  assign o[38848] = i[38848];
  assign o[38847] = i[38847];
  assign o[38846] = i[38846];
  assign o[38845] = i[38845];
  assign o[38844] = i[38844];
  assign o[38843] = i[38843];
  assign o[38842] = i[38842];
  assign o[38841] = i[38841];
  assign o[38840] = i[38840];
  assign o[38839] = i[38839];
  assign o[38838] = i[38838];
  assign o[38837] = i[38837];
  assign o[38836] = i[38836];
  assign o[38835] = i[38835];
  assign o[38834] = i[38834];
  assign o[38833] = i[38833];
  assign o[38832] = i[38832];
  assign o[38831] = i[38831];
  assign o[38830] = i[38830];
  assign o[38829] = i[38829];
  assign o[38828] = i[38828];
  assign o[38827] = i[38827];
  assign o[38826] = i[38826];
  assign o[38825] = i[38825];
  assign o[38824] = i[38824];
  assign o[38823] = i[38823];
  assign o[38822] = i[38822];
  assign o[38821] = i[38821];
  assign o[38820] = i[38820];
  assign o[38819] = i[38819];
  assign o[38818] = i[38818];
  assign o[38817] = i[38817];
  assign o[38816] = i[38816];
  assign o[38815] = i[38815];
  assign o[38814] = i[38814];
  assign o[38813] = i[38813];
  assign o[38812] = i[38812];
  assign o[38811] = i[38811];
  assign o[38810] = i[38810];
  assign o[38809] = i[38809];
  assign o[38808] = i[38808];
  assign o[38807] = i[38807];
  assign o[38806] = i[38806];
  assign o[38805] = i[38805];
  assign o[38804] = i[38804];
  assign o[38803] = i[38803];
  assign o[38802] = i[38802];
  assign o[38801] = i[38801];
  assign o[38800] = i[38800];
  assign o[38799] = i[38799];
  assign o[38798] = i[38798];
  assign o[38797] = i[38797];
  assign o[38796] = i[38796];
  assign o[38795] = i[38795];
  assign o[38794] = i[38794];
  assign o[38793] = i[38793];
  assign o[38792] = i[38792];
  assign o[38791] = i[38791];
  assign o[38790] = i[38790];
  assign o[38789] = i[38789];
  assign o[38788] = i[38788];
  assign o[38787] = i[38787];
  assign o[38786] = i[38786];
  assign o[38785] = i[38785];
  assign o[38784] = i[38784];
  assign o[38783] = i[38783];
  assign o[38782] = i[38782];
  assign o[38781] = i[38781];
  assign o[38780] = i[38780];
  assign o[38779] = i[38779];
  assign o[38778] = i[38778];
  assign o[38777] = i[38777];
  assign o[38776] = i[38776];
  assign o[38775] = i[38775];
  assign o[38774] = i[38774];
  assign o[38773] = i[38773];
  assign o[38772] = i[38772];
  assign o[38771] = i[38771];
  assign o[38770] = i[38770];
  assign o[38769] = i[38769];
  assign o[38768] = i[38768];
  assign o[38767] = i[38767];
  assign o[38766] = i[38766];
  assign o[38765] = i[38765];
  assign o[38764] = i[38764];
  assign o[38763] = i[38763];
  assign o[38762] = i[38762];
  assign o[38761] = i[38761];
  assign o[38760] = i[38760];
  assign o[38759] = i[38759];
  assign o[38758] = i[38758];
  assign o[38757] = i[38757];
  assign o[38756] = i[38756];
  assign o[38755] = i[38755];
  assign o[38754] = i[38754];
  assign o[38753] = i[38753];
  assign o[38752] = i[38752];
  assign o[38751] = i[38751];
  assign o[38750] = i[38750];
  assign o[38749] = i[38749];
  assign o[38748] = i[38748];
  assign o[38747] = i[38747];
  assign o[38746] = i[38746];
  assign o[38745] = i[38745];
  assign o[38744] = i[38744];
  assign o[38743] = i[38743];
  assign o[38742] = i[38742];
  assign o[38741] = i[38741];
  assign o[38740] = i[38740];
  assign o[38739] = i[38739];
  assign o[38738] = i[38738];
  assign o[38737] = i[38737];
  assign o[38736] = i[38736];
  assign o[38735] = i[38735];
  assign o[38734] = i[38734];
  assign o[38733] = i[38733];
  assign o[38732] = i[38732];
  assign o[38731] = i[38731];
  assign o[38730] = i[38730];
  assign o[38729] = i[38729];
  assign o[38728] = i[38728];
  assign o[38727] = i[38727];
  assign o[38726] = i[38726];
  assign o[38725] = i[38725];
  assign o[38724] = i[38724];
  assign o[38723] = i[38723];
  assign o[38722] = i[38722];
  assign o[38721] = i[38721];
  assign o[38720] = i[38720];
  assign o[38719] = i[38719];
  assign o[38718] = i[38718];
  assign o[38717] = i[38717];
  assign o[38716] = i[38716];
  assign o[38715] = i[38715];
  assign o[38714] = i[38714];
  assign o[38713] = i[38713];
  assign o[38712] = i[38712];
  assign o[38711] = i[38711];
  assign o[38710] = i[38710];
  assign o[38709] = i[38709];
  assign o[38708] = i[38708];
  assign o[38707] = i[38707];
  assign o[38706] = i[38706];
  assign o[38705] = i[38705];
  assign o[38704] = i[38704];
  assign o[38703] = i[38703];
  assign o[38702] = i[38702];
  assign o[38701] = i[38701];
  assign o[38700] = i[38700];
  assign o[38699] = i[38699];
  assign o[38698] = i[38698];
  assign o[38697] = i[38697];
  assign o[38696] = i[38696];
  assign o[38695] = i[38695];
  assign o[38694] = i[38694];
  assign o[38693] = i[38693];
  assign o[38692] = i[38692];
  assign o[38691] = i[38691];
  assign o[38690] = i[38690];
  assign o[38689] = i[38689];
  assign o[38688] = i[38688];
  assign o[38687] = i[38687];
  assign o[38686] = i[38686];
  assign o[38685] = i[38685];
  assign o[38684] = i[38684];
  assign o[38683] = i[38683];
  assign o[38682] = i[38682];
  assign o[38681] = i[38681];
  assign o[38680] = i[38680];
  assign o[38679] = i[38679];
  assign o[38678] = i[38678];
  assign o[38677] = i[38677];
  assign o[38676] = i[38676];
  assign o[38675] = i[38675];
  assign o[38674] = i[38674];
  assign o[38673] = i[38673];
  assign o[38672] = i[38672];
  assign o[38671] = i[38671];
  assign o[38670] = i[38670];
  assign o[38669] = i[38669];
  assign o[38668] = i[38668];
  assign o[38667] = i[38667];
  assign o[38666] = i[38666];
  assign o[38665] = i[38665];
  assign o[38664] = i[38664];
  assign o[38663] = i[38663];
  assign o[38662] = i[38662];
  assign o[38661] = i[38661];
  assign o[38660] = i[38660];
  assign o[38659] = i[38659];
  assign o[38658] = i[38658];
  assign o[38657] = i[38657];
  assign o[38656] = i[38656];
  assign o[38655] = i[38655];
  assign o[38654] = i[38654];
  assign o[38653] = i[38653];
  assign o[38652] = i[38652];
  assign o[38651] = i[38651];
  assign o[38650] = i[38650];
  assign o[38649] = i[38649];
  assign o[38648] = i[38648];
  assign o[38647] = i[38647];
  assign o[38646] = i[38646];
  assign o[38645] = i[38645];
  assign o[38644] = i[38644];
  assign o[38643] = i[38643];
  assign o[38642] = i[38642];
  assign o[38641] = i[38641];
  assign o[38640] = i[38640];
  assign o[38639] = i[38639];
  assign o[38638] = i[38638];
  assign o[38637] = i[38637];
  assign o[38636] = i[38636];
  assign o[38635] = i[38635];
  assign o[38634] = i[38634];
  assign o[38633] = i[38633];
  assign o[38632] = i[38632];
  assign o[38631] = i[38631];
  assign o[38630] = i[38630];
  assign o[38629] = i[38629];
  assign o[38628] = i[38628];
  assign o[38627] = i[38627];
  assign o[38626] = i[38626];
  assign o[38625] = i[38625];
  assign o[38624] = i[38624];
  assign o[38623] = i[38623];
  assign o[38622] = i[38622];
  assign o[38621] = i[38621];
  assign o[38620] = i[38620];
  assign o[38619] = i[38619];
  assign o[38618] = i[38618];
  assign o[38617] = i[38617];
  assign o[38616] = i[38616];
  assign o[38615] = i[38615];
  assign o[38614] = i[38614];
  assign o[38613] = i[38613];
  assign o[38612] = i[38612];
  assign o[38611] = i[38611];
  assign o[38610] = i[38610];
  assign o[38609] = i[38609];
  assign o[38608] = i[38608];
  assign o[38607] = i[38607];
  assign o[38606] = i[38606];
  assign o[38605] = i[38605];
  assign o[38604] = i[38604];
  assign o[38603] = i[38603];
  assign o[38602] = i[38602];
  assign o[38601] = i[38601];
  assign o[38600] = i[38600];
  assign o[38599] = i[38599];
  assign o[38598] = i[38598];
  assign o[38597] = i[38597];
  assign o[38596] = i[38596];
  assign o[38595] = i[38595];
  assign o[38594] = i[38594];
  assign o[38593] = i[38593];
  assign o[38592] = i[38592];
  assign o[38591] = i[38591];
  assign o[38590] = i[38590];
  assign o[38589] = i[38589];
  assign o[38588] = i[38588];
  assign o[38587] = i[38587];
  assign o[38586] = i[38586];
  assign o[38585] = i[38585];
  assign o[38584] = i[38584];
  assign o[38583] = i[38583];
  assign o[38582] = i[38582];
  assign o[38581] = i[38581];
  assign o[38580] = i[38580];
  assign o[38579] = i[38579];
  assign o[38578] = i[38578];
  assign o[38577] = i[38577];
  assign o[38576] = i[38576];
  assign o[38575] = i[38575];
  assign o[38574] = i[38574];
  assign o[38573] = i[38573];
  assign o[38572] = i[38572];
  assign o[38571] = i[38571];
  assign o[38570] = i[38570];
  assign o[38569] = i[38569];
  assign o[38568] = i[38568];
  assign o[38567] = i[38567];
  assign o[38566] = i[38566];
  assign o[38565] = i[38565];
  assign o[38564] = i[38564];
  assign o[38563] = i[38563];
  assign o[38562] = i[38562];
  assign o[38561] = i[38561];
  assign o[38560] = i[38560];
  assign o[38559] = i[38559];
  assign o[38558] = i[38558];
  assign o[38557] = i[38557];
  assign o[38556] = i[38556];
  assign o[38555] = i[38555];
  assign o[38554] = i[38554];
  assign o[38553] = i[38553];
  assign o[38552] = i[38552];
  assign o[38551] = i[38551];
  assign o[38550] = i[38550];
  assign o[38549] = i[38549];
  assign o[38548] = i[38548];
  assign o[38547] = i[38547];
  assign o[38546] = i[38546];
  assign o[38545] = i[38545];
  assign o[38544] = i[38544];
  assign o[38543] = i[38543];
  assign o[38542] = i[38542];
  assign o[38541] = i[38541];
  assign o[38540] = i[38540];
  assign o[38539] = i[38539];
  assign o[38538] = i[38538];
  assign o[38537] = i[38537];
  assign o[38536] = i[38536];
  assign o[38535] = i[38535];
  assign o[38534] = i[38534];
  assign o[38533] = i[38533];
  assign o[38532] = i[38532];
  assign o[38531] = i[38531];
  assign o[38530] = i[38530];
  assign o[38529] = i[38529];
  assign o[38528] = i[38528];
  assign o[38527] = i[38527];
  assign o[38526] = i[38526];
  assign o[38525] = i[38525];
  assign o[38524] = i[38524];
  assign o[38523] = i[38523];
  assign o[38522] = i[38522];
  assign o[38521] = i[38521];
  assign o[38520] = i[38520];
  assign o[38519] = i[38519];
  assign o[38518] = i[38518];
  assign o[38517] = i[38517];
  assign o[38516] = i[38516];
  assign o[38515] = i[38515];
  assign o[38514] = i[38514];
  assign o[38513] = i[38513];
  assign o[38512] = i[38512];
  assign o[38511] = i[38511];
  assign o[38510] = i[38510];
  assign o[38509] = i[38509];
  assign o[38508] = i[38508];
  assign o[38507] = i[38507];
  assign o[38506] = i[38506];
  assign o[38505] = i[38505];
  assign o[38504] = i[38504];
  assign o[38503] = i[38503];
  assign o[38502] = i[38502];
  assign o[38501] = i[38501];
  assign o[38500] = i[38500];
  assign o[38499] = i[38499];
  assign o[38498] = i[38498];
  assign o[38497] = i[38497];
  assign o[38496] = i[38496];
  assign o[38495] = i[38495];
  assign o[38494] = i[38494];
  assign o[38493] = i[38493];
  assign o[38492] = i[38492];
  assign o[38491] = i[38491];
  assign o[38490] = i[38490];
  assign o[38489] = i[38489];
  assign o[38488] = i[38488];
  assign o[38487] = i[38487];
  assign o[38486] = i[38486];
  assign o[38485] = i[38485];
  assign o[38484] = i[38484];
  assign o[38483] = i[38483];
  assign o[38482] = i[38482];
  assign o[38481] = i[38481];
  assign o[38480] = i[38480];
  assign o[38479] = i[38479];
  assign o[38478] = i[38478];
  assign o[38477] = i[38477];
  assign o[38476] = i[38476];
  assign o[38475] = i[38475];
  assign o[38474] = i[38474];
  assign o[38473] = i[38473];
  assign o[38472] = i[38472];
  assign o[38471] = i[38471];
  assign o[38470] = i[38470];
  assign o[38469] = i[38469];
  assign o[38468] = i[38468];
  assign o[38467] = i[38467];
  assign o[38466] = i[38466];
  assign o[38465] = i[38465];
  assign o[38464] = i[38464];
  assign o[38463] = i[38463];
  assign o[38462] = i[38462];
  assign o[38461] = i[38461];
  assign o[38460] = i[38460];
  assign o[38459] = i[38459];
  assign o[38458] = i[38458];
  assign o[38457] = i[38457];
  assign o[38456] = i[38456];
  assign o[38455] = i[38455];
  assign o[38454] = i[38454];
  assign o[38453] = i[38453];
  assign o[38452] = i[38452];
  assign o[38451] = i[38451];
  assign o[38450] = i[38450];
  assign o[38449] = i[38449];
  assign o[38448] = i[38448];
  assign o[38447] = i[38447];
  assign o[38446] = i[38446];
  assign o[38445] = i[38445];
  assign o[38444] = i[38444];
  assign o[38443] = i[38443];
  assign o[38442] = i[38442];
  assign o[38441] = i[38441];
  assign o[38440] = i[38440];
  assign o[38439] = i[38439];
  assign o[38438] = i[38438];
  assign o[38437] = i[38437];
  assign o[38436] = i[38436];
  assign o[38435] = i[38435];
  assign o[38434] = i[38434];
  assign o[38433] = i[38433];
  assign o[38432] = i[38432];
  assign o[38431] = i[38431];
  assign o[38430] = i[38430];
  assign o[38429] = i[38429];
  assign o[38428] = i[38428];
  assign o[38427] = i[38427];
  assign o[38426] = i[38426];
  assign o[38425] = i[38425];
  assign o[38424] = i[38424];
  assign o[38423] = i[38423];
  assign o[38422] = i[38422];
  assign o[38421] = i[38421];
  assign o[38420] = i[38420];
  assign o[38419] = i[38419];
  assign o[38418] = i[38418];
  assign o[38417] = i[38417];
  assign o[38416] = i[38416];
  assign o[38415] = i[38415];
  assign o[38414] = i[38414];
  assign o[38413] = i[38413];
  assign o[38412] = i[38412];
  assign o[38411] = i[38411];
  assign o[38410] = i[38410];
  assign o[38409] = i[38409];
  assign o[38408] = i[38408];
  assign o[38407] = i[38407];
  assign o[38406] = i[38406];
  assign o[38405] = i[38405];
  assign o[38404] = i[38404];
  assign o[38403] = i[38403];
  assign o[38402] = i[38402];
  assign o[38401] = i[38401];
  assign o[38400] = i[38400];
  assign o[38399] = i[38399];
  assign o[38398] = i[38398];
  assign o[38397] = i[38397];
  assign o[38396] = i[38396];
  assign o[38395] = i[38395];
  assign o[38394] = i[38394];
  assign o[38393] = i[38393];
  assign o[38392] = i[38392];
  assign o[38391] = i[38391];
  assign o[38390] = i[38390];
  assign o[38389] = i[38389];
  assign o[38388] = i[38388];
  assign o[38387] = i[38387];
  assign o[38386] = i[38386];
  assign o[38385] = i[38385];
  assign o[38384] = i[38384];
  assign o[38383] = i[38383];
  assign o[38382] = i[38382];
  assign o[38381] = i[38381];
  assign o[38380] = i[38380];
  assign o[38379] = i[38379];
  assign o[38378] = i[38378];
  assign o[38377] = i[38377];
  assign o[38376] = i[38376];
  assign o[38375] = i[38375];
  assign o[38374] = i[38374];
  assign o[38373] = i[38373];
  assign o[38372] = i[38372];
  assign o[38371] = i[38371];
  assign o[38370] = i[38370];
  assign o[38369] = i[38369];
  assign o[38368] = i[38368];
  assign o[38367] = i[38367];
  assign o[38366] = i[38366];
  assign o[38365] = i[38365];
  assign o[38364] = i[38364];
  assign o[38363] = i[38363];
  assign o[38362] = i[38362];
  assign o[38361] = i[38361];
  assign o[38360] = i[38360];
  assign o[38359] = i[38359];
  assign o[38358] = i[38358];
  assign o[38357] = i[38357];
  assign o[38356] = i[38356];
  assign o[38355] = i[38355];
  assign o[38354] = i[38354];
  assign o[38353] = i[38353];
  assign o[38352] = i[38352];
  assign o[38351] = i[38351];
  assign o[38350] = i[38350];
  assign o[38349] = i[38349];
  assign o[38348] = i[38348];
  assign o[38347] = i[38347];
  assign o[38346] = i[38346];
  assign o[38345] = i[38345];
  assign o[38344] = i[38344];
  assign o[38343] = i[38343];
  assign o[38342] = i[38342];
  assign o[38341] = i[38341];
  assign o[38340] = i[38340];
  assign o[38339] = i[38339];
  assign o[38338] = i[38338];
  assign o[38337] = i[38337];
  assign o[38336] = i[38336];
  assign o[38335] = i[38335];
  assign o[38334] = i[38334];
  assign o[38333] = i[38333];
  assign o[38332] = i[38332];
  assign o[38331] = i[38331];
  assign o[38330] = i[38330];
  assign o[38329] = i[38329];
  assign o[38328] = i[38328];
  assign o[38327] = i[38327];
  assign o[38326] = i[38326];
  assign o[38325] = i[38325];
  assign o[38324] = i[38324];
  assign o[38323] = i[38323];
  assign o[38322] = i[38322];
  assign o[38321] = i[38321];
  assign o[38320] = i[38320];
  assign o[38319] = i[38319];
  assign o[38318] = i[38318];
  assign o[38317] = i[38317];
  assign o[38316] = i[38316];
  assign o[38315] = i[38315];
  assign o[38314] = i[38314];
  assign o[38313] = i[38313];
  assign o[38312] = i[38312];
  assign o[38311] = i[38311];
  assign o[38310] = i[38310];
  assign o[38309] = i[38309];
  assign o[38308] = i[38308];
  assign o[38307] = i[38307];
  assign o[38306] = i[38306];
  assign o[38305] = i[38305];
  assign o[38304] = i[38304];
  assign o[38303] = i[38303];
  assign o[38302] = i[38302];
  assign o[38301] = i[38301];
  assign o[38300] = i[38300];
  assign o[38299] = i[38299];
  assign o[38298] = i[38298];
  assign o[38297] = i[38297];
  assign o[38296] = i[38296];
  assign o[38295] = i[38295];
  assign o[38294] = i[38294];
  assign o[38293] = i[38293];
  assign o[38292] = i[38292];
  assign o[38291] = i[38291];
  assign o[38290] = i[38290];
  assign o[38289] = i[38289];
  assign o[38288] = i[38288];
  assign o[38287] = i[38287];
  assign o[38286] = i[38286];
  assign o[38285] = i[38285];
  assign o[38284] = i[38284];
  assign o[38283] = i[38283];
  assign o[38282] = i[38282];
  assign o[38281] = i[38281];
  assign o[38280] = i[38280];
  assign o[38279] = i[38279];
  assign o[38278] = i[38278];
  assign o[38277] = i[38277];
  assign o[38276] = i[38276];
  assign o[38275] = i[38275];
  assign o[38274] = i[38274];
  assign o[38273] = i[38273];
  assign o[38272] = i[38272];
  assign o[38271] = i[38271];
  assign o[38270] = i[38270];
  assign o[38269] = i[38269];
  assign o[38268] = i[38268];
  assign o[38267] = i[38267];
  assign o[38266] = i[38266];
  assign o[38265] = i[38265];
  assign o[38264] = i[38264];
  assign o[38263] = i[38263];
  assign o[38262] = i[38262];
  assign o[38261] = i[38261];
  assign o[38260] = i[38260];
  assign o[38259] = i[38259];
  assign o[38258] = i[38258];
  assign o[38257] = i[38257];
  assign o[38256] = i[38256];
  assign o[38255] = i[38255];
  assign o[38254] = i[38254];
  assign o[38253] = i[38253];
  assign o[38252] = i[38252];
  assign o[38251] = i[38251];
  assign o[38250] = i[38250];
  assign o[38249] = i[38249];
  assign o[38248] = i[38248];
  assign o[38247] = i[38247];
  assign o[38246] = i[38246];
  assign o[38245] = i[38245];
  assign o[38244] = i[38244];
  assign o[38243] = i[38243];
  assign o[38242] = i[38242];
  assign o[38241] = i[38241];
  assign o[38240] = i[38240];
  assign o[38239] = i[38239];
  assign o[38238] = i[38238];
  assign o[38237] = i[38237];
  assign o[38236] = i[38236];
  assign o[38235] = i[38235];
  assign o[38234] = i[38234];
  assign o[38233] = i[38233];
  assign o[38232] = i[38232];
  assign o[38231] = i[38231];
  assign o[38230] = i[38230];
  assign o[38229] = i[38229];
  assign o[38228] = i[38228];
  assign o[38227] = i[38227];
  assign o[38226] = i[38226];
  assign o[38225] = i[38225];
  assign o[38224] = i[38224];
  assign o[38223] = i[38223];
  assign o[38222] = i[38222];
  assign o[38221] = i[38221];
  assign o[38220] = i[38220];
  assign o[38219] = i[38219];
  assign o[38218] = i[38218];
  assign o[38217] = i[38217];
  assign o[38216] = i[38216];
  assign o[38215] = i[38215];
  assign o[38214] = i[38214];
  assign o[38213] = i[38213];
  assign o[38212] = i[38212];
  assign o[38211] = i[38211];
  assign o[38210] = i[38210];
  assign o[38209] = i[38209];
  assign o[38208] = i[38208];
  assign o[38207] = i[38207];
  assign o[38206] = i[38206];
  assign o[38205] = i[38205];
  assign o[38204] = i[38204];
  assign o[38203] = i[38203];
  assign o[38202] = i[38202];
  assign o[38201] = i[38201];
  assign o[38200] = i[38200];
  assign o[38199] = i[38199];
  assign o[38198] = i[38198];
  assign o[38197] = i[38197];
  assign o[38196] = i[38196];
  assign o[38195] = i[38195];
  assign o[38194] = i[38194];
  assign o[38193] = i[38193];
  assign o[38192] = i[38192];
  assign o[38191] = i[38191];
  assign o[38190] = i[38190];
  assign o[38189] = i[38189];
  assign o[38188] = i[38188];
  assign o[38187] = i[38187];
  assign o[38186] = i[38186];
  assign o[38185] = i[38185];
  assign o[38184] = i[38184];
  assign o[38183] = i[38183];
  assign o[38182] = i[38182];
  assign o[38181] = i[38181];
  assign o[38180] = i[38180];
  assign o[38179] = i[38179];
  assign o[38178] = i[38178];
  assign o[38177] = i[38177];
  assign o[38176] = i[38176];
  assign o[38175] = i[38175];
  assign o[38174] = i[38174];
  assign o[38173] = i[38173];
  assign o[38172] = i[38172];
  assign o[38171] = i[38171];
  assign o[38170] = i[38170];
  assign o[38169] = i[38169];
  assign o[38168] = i[38168];
  assign o[38167] = i[38167];
  assign o[38166] = i[38166];
  assign o[38165] = i[38165];
  assign o[38164] = i[38164];
  assign o[38163] = i[38163];
  assign o[38162] = i[38162];
  assign o[38161] = i[38161];
  assign o[38160] = i[38160];
  assign o[38159] = i[38159];
  assign o[38158] = i[38158];
  assign o[38157] = i[38157];
  assign o[38156] = i[38156];
  assign o[38155] = i[38155];
  assign o[38154] = i[38154];
  assign o[38153] = i[38153];
  assign o[38152] = i[38152];
  assign o[38151] = i[38151];
  assign o[38150] = i[38150];
  assign o[38149] = i[38149];
  assign o[38148] = i[38148];
  assign o[38147] = i[38147];
  assign o[38146] = i[38146];
  assign o[38145] = i[38145];
  assign o[38144] = i[38144];
  assign o[38143] = i[38143];
  assign o[38142] = i[38142];
  assign o[38141] = i[38141];
  assign o[38140] = i[38140];
  assign o[38139] = i[38139];
  assign o[38138] = i[38138];
  assign o[38137] = i[38137];
  assign o[38136] = i[38136];
  assign o[38135] = i[38135];
  assign o[38134] = i[38134];
  assign o[38133] = i[38133];
  assign o[38132] = i[38132];
  assign o[38131] = i[38131];
  assign o[38130] = i[38130];
  assign o[38129] = i[38129];
  assign o[38128] = i[38128];
  assign o[38127] = i[38127];
  assign o[38126] = i[38126];
  assign o[38125] = i[38125];
  assign o[38124] = i[38124];
  assign o[38123] = i[38123];
  assign o[38122] = i[38122];
  assign o[38121] = i[38121];
  assign o[38120] = i[38120];
  assign o[38119] = i[38119];
  assign o[38118] = i[38118];
  assign o[38117] = i[38117];
  assign o[38116] = i[38116];
  assign o[38115] = i[38115];
  assign o[38114] = i[38114];
  assign o[38113] = i[38113];
  assign o[38112] = i[38112];
  assign o[38111] = i[38111];
  assign o[38110] = i[38110];
  assign o[38109] = i[38109];
  assign o[38108] = i[38108];
  assign o[38107] = i[38107];
  assign o[38106] = i[38106];
  assign o[38105] = i[38105];
  assign o[38104] = i[38104];
  assign o[38103] = i[38103];
  assign o[38102] = i[38102];
  assign o[38101] = i[38101];
  assign o[38100] = i[38100];
  assign o[38099] = i[38099];
  assign o[38098] = i[38098];
  assign o[38097] = i[38097];
  assign o[38096] = i[38096];
  assign o[38095] = i[38095];
  assign o[38094] = i[38094];
  assign o[38093] = i[38093];
  assign o[38092] = i[38092];
  assign o[38091] = i[38091];
  assign o[38090] = i[38090];
  assign o[38089] = i[38089];
  assign o[38088] = i[38088];
  assign o[38087] = i[38087];
  assign o[38086] = i[38086];
  assign o[38085] = i[38085];
  assign o[38084] = i[38084];
  assign o[38083] = i[38083];
  assign o[38082] = i[38082];
  assign o[38081] = i[38081];
  assign o[38080] = i[38080];
  assign o[38079] = i[38079];
  assign o[38078] = i[38078];
  assign o[38077] = i[38077];
  assign o[38076] = i[38076];
  assign o[38075] = i[38075];
  assign o[38074] = i[38074];
  assign o[38073] = i[38073];
  assign o[38072] = i[38072];
  assign o[38071] = i[38071];
  assign o[38070] = i[38070];
  assign o[38069] = i[38069];
  assign o[38068] = i[38068];
  assign o[38067] = i[38067];
  assign o[38066] = i[38066];
  assign o[38065] = i[38065];
  assign o[38064] = i[38064];
  assign o[38063] = i[38063];
  assign o[38062] = i[38062];
  assign o[38061] = i[38061];
  assign o[38060] = i[38060];
  assign o[38059] = i[38059];
  assign o[38058] = i[38058];
  assign o[38057] = i[38057];
  assign o[38056] = i[38056];
  assign o[38055] = i[38055];
  assign o[38054] = i[38054];
  assign o[38053] = i[38053];
  assign o[38052] = i[38052];
  assign o[38051] = i[38051];
  assign o[38050] = i[38050];
  assign o[38049] = i[38049];
  assign o[38048] = i[38048];
  assign o[38047] = i[38047];
  assign o[38046] = i[38046];
  assign o[38045] = i[38045];
  assign o[38044] = i[38044];
  assign o[38043] = i[38043];
  assign o[38042] = i[38042];
  assign o[38041] = i[38041];
  assign o[38040] = i[38040];
  assign o[38039] = i[38039];
  assign o[38038] = i[38038];
  assign o[38037] = i[38037];
  assign o[38036] = i[38036];
  assign o[38035] = i[38035];
  assign o[38034] = i[38034];
  assign o[38033] = i[38033];
  assign o[38032] = i[38032];
  assign o[38031] = i[38031];
  assign o[38030] = i[38030];
  assign o[38029] = i[38029];
  assign o[38028] = i[38028];
  assign o[38027] = i[38027];
  assign o[38026] = i[38026];
  assign o[38025] = i[38025];
  assign o[38024] = i[38024];
  assign o[38023] = i[38023];
  assign o[38022] = i[38022];
  assign o[38021] = i[38021];
  assign o[38020] = i[38020];
  assign o[38019] = i[38019];
  assign o[38018] = i[38018];
  assign o[38017] = i[38017];
  assign o[38016] = i[38016];
  assign o[38015] = i[38015];
  assign o[38014] = i[38014];
  assign o[38013] = i[38013];
  assign o[38012] = i[38012];
  assign o[38011] = i[38011];
  assign o[38010] = i[38010];
  assign o[38009] = i[38009];
  assign o[38008] = i[38008];
  assign o[38007] = i[38007];
  assign o[38006] = i[38006];
  assign o[38005] = i[38005];
  assign o[38004] = i[38004];
  assign o[38003] = i[38003];
  assign o[38002] = i[38002];
  assign o[38001] = i[38001];
  assign o[38000] = i[38000];
  assign o[37999] = i[37999];
  assign o[37998] = i[37998];
  assign o[37997] = i[37997];
  assign o[37996] = i[37996];
  assign o[37995] = i[37995];
  assign o[37994] = i[37994];
  assign o[37993] = i[37993];
  assign o[37992] = i[37992];
  assign o[37991] = i[37991];
  assign o[37990] = i[37990];
  assign o[37989] = i[37989];
  assign o[37988] = i[37988];
  assign o[37987] = i[37987];
  assign o[37986] = i[37986];
  assign o[37985] = i[37985];
  assign o[37984] = i[37984];
  assign o[37983] = i[37983];
  assign o[37982] = i[37982];
  assign o[37981] = i[37981];
  assign o[37980] = i[37980];
  assign o[37979] = i[37979];
  assign o[37978] = i[37978];
  assign o[37977] = i[37977];
  assign o[37976] = i[37976];
  assign o[37975] = i[37975];
  assign o[37974] = i[37974];
  assign o[37973] = i[37973];
  assign o[37972] = i[37972];
  assign o[37971] = i[37971];
  assign o[37970] = i[37970];
  assign o[37969] = i[37969];
  assign o[37968] = i[37968];
  assign o[37967] = i[37967];
  assign o[37966] = i[37966];
  assign o[37965] = i[37965];
  assign o[37964] = i[37964];
  assign o[37963] = i[37963];
  assign o[37962] = i[37962];
  assign o[37961] = i[37961];
  assign o[37960] = i[37960];
  assign o[37959] = i[37959];
  assign o[37958] = i[37958];
  assign o[37957] = i[37957];
  assign o[37956] = i[37956];
  assign o[37955] = i[37955];
  assign o[37954] = i[37954];
  assign o[37953] = i[37953];
  assign o[37952] = i[37952];
  assign o[37951] = i[37951];
  assign o[37950] = i[37950];
  assign o[37949] = i[37949];
  assign o[37948] = i[37948];
  assign o[37947] = i[37947];
  assign o[37946] = i[37946];
  assign o[37945] = i[37945];
  assign o[37944] = i[37944];
  assign o[37943] = i[37943];
  assign o[37942] = i[37942];
  assign o[37941] = i[37941];
  assign o[37940] = i[37940];
  assign o[37939] = i[37939];
  assign o[37938] = i[37938];
  assign o[37937] = i[37937];
  assign o[37936] = i[37936];
  assign o[37935] = i[37935];
  assign o[37934] = i[37934];
  assign o[37933] = i[37933];
  assign o[37932] = i[37932];
  assign o[37931] = i[37931];
  assign o[37930] = i[37930];
  assign o[37929] = i[37929];
  assign o[37928] = i[37928];
  assign o[37927] = i[37927];
  assign o[37926] = i[37926];
  assign o[37925] = i[37925];
  assign o[37924] = i[37924];
  assign o[37923] = i[37923];
  assign o[37922] = i[37922];
  assign o[37921] = i[37921];
  assign o[37920] = i[37920];
  assign o[37919] = i[37919];
  assign o[37918] = i[37918];
  assign o[37917] = i[37917];
  assign o[37916] = i[37916];
  assign o[37915] = i[37915];
  assign o[37914] = i[37914];
  assign o[37913] = i[37913];
  assign o[37912] = i[37912];
  assign o[37911] = i[37911];
  assign o[37910] = i[37910];
  assign o[37909] = i[37909];
  assign o[37908] = i[37908];
  assign o[37907] = i[37907];
  assign o[37906] = i[37906];
  assign o[37905] = i[37905];
  assign o[37904] = i[37904];
  assign o[37903] = i[37903];
  assign o[37902] = i[37902];
  assign o[37901] = i[37901];
  assign o[37900] = i[37900];
  assign o[37899] = i[37899];
  assign o[37898] = i[37898];
  assign o[37897] = i[37897];
  assign o[37896] = i[37896];
  assign o[37895] = i[37895];
  assign o[37894] = i[37894];
  assign o[37893] = i[37893];
  assign o[37892] = i[37892];
  assign o[37891] = i[37891];
  assign o[37890] = i[37890];
  assign o[37889] = i[37889];
  assign o[37888] = i[37888];
  assign o[37887] = i[37887];
  assign o[37886] = i[37886];
  assign o[37885] = i[37885];
  assign o[37884] = i[37884];
  assign o[37883] = i[37883];
  assign o[37882] = i[37882];
  assign o[37881] = i[37881];
  assign o[37880] = i[37880];
  assign o[37879] = i[37879];
  assign o[37878] = i[37878];
  assign o[37877] = i[37877];
  assign o[37876] = i[37876];
  assign o[37875] = i[37875];
  assign o[37874] = i[37874];
  assign o[37873] = i[37873];
  assign o[37872] = i[37872];
  assign o[37871] = i[37871];
  assign o[37870] = i[37870];
  assign o[37869] = i[37869];
  assign o[37868] = i[37868];
  assign o[37867] = i[37867];
  assign o[37866] = i[37866];
  assign o[37865] = i[37865];
  assign o[37864] = i[37864];
  assign o[37863] = i[37863];
  assign o[37862] = i[37862];
  assign o[37861] = i[37861];
  assign o[37860] = i[37860];
  assign o[37859] = i[37859];
  assign o[37858] = i[37858];
  assign o[37857] = i[37857];
  assign o[37856] = i[37856];
  assign o[37855] = i[37855];
  assign o[37854] = i[37854];
  assign o[37853] = i[37853];
  assign o[37852] = i[37852];
  assign o[37851] = i[37851];
  assign o[37850] = i[37850];
  assign o[37849] = i[37849];
  assign o[37848] = i[37848];
  assign o[37847] = i[37847];
  assign o[37846] = i[37846];
  assign o[37845] = i[37845];
  assign o[37844] = i[37844];
  assign o[37843] = i[37843];
  assign o[37842] = i[37842];
  assign o[37841] = i[37841];
  assign o[37840] = i[37840];
  assign o[37839] = i[37839];
  assign o[37838] = i[37838];
  assign o[37837] = i[37837];
  assign o[37836] = i[37836];
  assign o[37835] = i[37835];
  assign o[37834] = i[37834];
  assign o[37833] = i[37833];
  assign o[37832] = i[37832];
  assign o[37831] = i[37831];
  assign o[37830] = i[37830];
  assign o[37829] = i[37829];
  assign o[37828] = i[37828];
  assign o[37827] = i[37827];
  assign o[37826] = i[37826];
  assign o[37825] = i[37825];
  assign o[37824] = i[37824];
  assign o[37823] = i[37823];
  assign o[37822] = i[37822];
  assign o[37821] = i[37821];
  assign o[37820] = i[37820];
  assign o[37819] = i[37819];
  assign o[37818] = i[37818];
  assign o[37817] = i[37817];
  assign o[37816] = i[37816];
  assign o[37815] = i[37815];
  assign o[37814] = i[37814];
  assign o[37813] = i[37813];
  assign o[37812] = i[37812];
  assign o[37811] = i[37811];
  assign o[37810] = i[37810];
  assign o[37809] = i[37809];
  assign o[37808] = i[37808];
  assign o[37807] = i[37807];
  assign o[37806] = i[37806];
  assign o[37805] = i[37805];
  assign o[37804] = i[37804];
  assign o[37803] = i[37803];
  assign o[37802] = i[37802];
  assign o[37801] = i[37801];
  assign o[37800] = i[37800];
  assign o[37799] = i[37799];
  assign o[37798] = i[37798];
  assign o[37797] = i[37797];
  assign o[37796] = i[37796];
  assign o[37795] = i[37795];
  assign o[37794] = i[37794];
  assign o[37793] = i[37793];
  assign o[37792] = i[37792];
  assign o[37791] = i[37791];
  assign o[37790] = i[37790];
  assign o[37789] = i[37789];
  assign o[37788] = i[37788];
  assign o[37787] = i[37787];
  assign o[37786] = i[37786];
  assign o[37785] = i[37785];
  assign o[37784] = i[37784];
  assign o[37783] = i[37783];
  assign o[37782] = i[37782];
  assign o[37781] = i[37781];
  assign o[37780] = i[37780];
  assign o[37779] = i[37779];
  assign o[37778] = i[37778];
  assign o[37777] = i[37777];
  assign o[37776] = i[37776];
  assign o[37775] = i[37775];
  assign o[37774] = i[37774];
  assign o[37773] = i[37773];
  assign o[37772] = i[37772];
  assign o[37771] = i[37771];
  assign o[37770] = i[37770];
  assign o[37769] = i[37769];
  assign o[37768] = i[37768];
  assign o[37767] = i[37767];
  assign o[37766] = i[37766];
  assign o[37765] = i[37765];
  assign o[37764] = i[37764];
  assign o[37763] = i[37763];
  assign o[37762] = i[37762];
  assign o[37761] = i[37761];
  assign o[37760] = i[37760];
  assign o[37759] = i[37759];
  assign o[37758] = i[37758];
  assign o[37757] = i[37757];
  assign o[37756] = i[37756];
  assign o[37755] = i[37755];
  assign o[37754] = i[37754];
  assign o[37753] = i[37753];
  assign o[37752] = i[37752];
  assign o[37751] = i[37751];
  assign o[37750] = i[37750];
  assign o[37749] = i[37749];
  assign o[37748] = i[37748];
  assign o[37747] = i[37747];
  assign o[37746] = i[37746];
  assign o[37745] = i[37745];
  assign o[37744] = i[37744];
  assign o[37743] = i[37743];
  assign o[37742] = i[37742];
  assign o[37741] = i[37741];
  assign o[37740] = i[37740];
  assign o[37739] = i[37739];
  assign o[37738] = i[37738];
  assign o[37737] = i[37737];
  assign o[37736] = i[37736];
  assign o[37735] = i[37735];
  assign o[37734] = i[37734];
  assign o[37733] = i[37733];
  assign o[37732] = i[37732];
  assign o[37731] = i[37731];
  assign o[37730] = i[37730];
  assign o[37729] = i[37729];
  assign o[37728] = i[37728];
  assign o[37727] = i[37727];
  assign o[37726] = i[37726];
  assign o[37725] = i[37725];
  assign o[37724] = i[37724];
  assign o[37723] = i[37723];
  assign o[37722] = i[37722];
  assign o[37721] = i[37721];
  assign o[37720] = i[37720];
  assign o[37719] = i[37719];
  assign o[37718] = i[37718];
  assign o[37717] = i[37717];
  assign o[37716] = i[37716];
  assign o[37715] = i[37715];
  assign o[37714] = i[37714];
  assign o[37713] = i[37713];
  assign o[37712] = i[37712];
  assign o[37711] = i[37711];
  assign o[37710] = i[37710];
  assign o[37709] = i[37709];
  assign o[37708] = i[37708];
  assign o[37707] = i[37707];
  assign o[37706] = i[37706];
  assign o[37705] = i[37705];
  assign o[37704] = i[37704];
  assign o[37703] = i[37703];
  assign o[37702] = i[37702];
  assign o[37701] = i[37701];
  assign o[37700] = i[37700];
  assign o[37699] = i[37699];
  assign o[37698] = i[37698];
  assign o[37697] = i[37697];
  assign o[37696] = i[37696];
  assign o[37695] = i[37695];
  assign o[37694] = i[37694];
  assign o[37693] = i[37693];
  assign o[37692] = i[37692];
  assign o[37691] = i[37691];
  assign o[37690] = i[37690];
  assign o[37689] = i[37689];
  assign o[37688] = i[37688];
  assign o[37687] = i[37687];
  assign o[37686] = i[37686];
  assign o[37685] = i[37685];
  assign o[37684] = i[37684];
  assign o[37683] = i[37683];
  assign o[37682] = i[37682];
  assign o[37681] = i[37681];
  assign o[37680] = i[37680];
  assign o[37679] = i[37679];
  assign o[37678] = i[37678];
  assign o[37677] = i[37677];
  assign o[37676] = i[37676];
  assign o[37675] = i[37675];
  assign o[37674] = i[37674];
  assign o[37673] = i[37673];
  assign o[37672] = i[37672];
  assign o[37671] = i[37671];
  assign o[37670] = i[37670];
  assign o[37669] = i[37669];
  assign o[37668] = i[37668];
  assign o[37667] = i[37667];
  assign o[37666] = i[37666];
  assign o[37665] = i[37665];
  assign o[37664] = i[37664];
  assign o[37663] = i[37663];
  assign o[37662] = i[37662];
  assign o[37661] = i[37661];
  assign o[37660] = i[37660];
  assign o[37659] = i[37659];
  assign o[37658] = i[37658];
  assign o[37657] = i[37657];
  assign o[37656] = i[37656];
  assign o[37655] = i[37655];
  assign o[37654] = i[37654];
  assign o[37653] = i[37653];
  assign o[37652] = i[37652];
  assign o[37651] = i[37651];
  assign o[37650] = i[37650];
  assign o[37649] = i[37649];
  assign o[37648] = i[37648];
  assign o[37647] = i[37647];
  assign o[37646] = i[37646];
  assign o[37645] = i[37645];
  assign o[37644] = i[37644];
  assign o[37643] = i[37643];
  assign o[37642] = i[37642];
  assign o[37641] = i[37641];
  assign o[37640] = i[37640];
  assign o[37639] = i[37639];
  assign o[37638] = i[37638];
  assign o[37637] = i[37637];
  assign o[37636] = i[37636];
  assign o[37635] = i[37635];
  assign o[37634] = i[37634];
  assign o[37633] = i[37633];
  assign o[37632] = i[37632];
  assign o[37631] = i[37631];
  assign o[37630] = i[37630];
  assign o[37629] = i[37629];
  assign o[37628] = i[37628];
  assign o[37627] = i[37627];
  assign o[37626] = i[37626];
  assign o[37625] = i[37625];
  assign o[37624] = i[37624];
  assign o[37623] = i[37623];
  assign o[37622] = i[37622];
  assign o[37621] = i[37621];
  assign o[37620] = i[37620];
  assign o[37619] = i[37619];
  assign o[37618] = i[37618];
  assign o[37617] = i[37617];
  assign o[37616] = i[37616];
  assign o[37615] = i[37615];
  assign o[37614] = i[37614];
  assign o[37613] = i[37613];
  assign o[37612] = i[37612];
  assign o[37611] = i[37611];
  assign o[37610] = i[37610];
  assign o[37609] = i[37609];
  assign o[37608] = i[37608];
  assign o[37607] = i[37607];
  assign o[37606] = i[37606];
  assign o[37605] = i[37605];
  assign o[37604] = i[37604];
  assign o[37603] = i[37603];
  assign o[37602] = i[37602];
  assign o[37601] = i[37601];
  assign o[37600] = i[37600];
  assign o[37599] = i[37599];
  assign o[37598] = i[37598];
  assign o[37597] = i[37597];
  assign o[37596] = i[37596];
  assign o[37595] = i[37595];
  assign o[37594] = i[37594];
  assign o[37593] = i[37593];
  assign o[37592] = i[37592];
  assign o[37591] = i[37591];
  assign o[37590] = i[37590];
  assign o[37589] = i[37589];
  assign o[37588] = i[37588];
  assign o[37587] = i[37587];
  assign o[37586] = i[37586];
  assign o[37585] = i[37585];
  assign o[37584] = i[37584];
  assign o[37583] = i[37583];
  assign o[37582] = i[37582];
  assign o[37581] = i[37581];
  assign o[37580] = i[37580];
  assign o[37579] = i[37579];
  assign o[37578] = i[37578];
  assign o[37577] = i[37577];
  assign o[37576] = i[37576];
  assign o[37575] = i[37575];
  assign o[37574] = i[37574];
  assign o[37573] = i[37573];
  assign o[37572] = i[37572];
  assign o[37571] = i[37571];
  assign o[37570] = i[37570];
  assign o[37569] = i[37569];
  assign o[37568] = i[37568];
  assign o[37567] = i[37567];
  assign o[37566] = i[37566];
  assign o[37565] = i[37565];
  assign o[37564] = i[37564];
  assign o[37563] = i[37563];
  assign o[37562] = i[37562];
  assign o[37561] = i[37561];
  assign o[37560] = i[37560];
  assign o[37559] = i[37559];
  assign o[37558] = i[37558];
  assign o[37557] = i[37557];
  assign o[37556] = i[37556];
  assign o[37555] = i[37555];
  assign o[37554] = i[37554];
  assign o[37553] = i[37553];
  assign o[37552] = i[37552];
  assign o[37551] = i[37551];
  assign o[37550] = i[37550];
  assign o[37549] = i[37549];
  assign o[37548] = i[37548];
  assign o[37547] = i[37547];
  assign o[37546] = i[37546];
  assign o[37545] = i[37545];
  assign o[37544] = i[37544];
  assign o[37543] = i[37543];
  assign o[37542] = i[37542];
  assign o[37541] = i[37541];
  assign o[37540] = i[37540];
  assign o[37539] = i[37539];
  assign o[37538] = i[37538];
  assign o[37537] = i[37537];
  assign o[37536] = i[37536];
  assign o[37535] = i[37535];
  assign o[37534] = i[37534];
  assign o[37533] = i[37533];
  assign o[37532] = i[37532];
  assign o[37531] = i[37531];
  assign o[37530] = i[37530];
  assign o[37529] = i[37529];
  assign o[37528] = i[37528];
  assign o[37527] = i[37527];
  assign o[37526] = i[37526];
  assign o[37525] = i[37525];
  assign o[37524] = i[37524];
  assign o[37523] = i[37523];
  assign o[37522] = i[37522];
  assign o[37521] = i[37521];
  assign o[37520] = i[37520];
  assign o[37519] = i[37519];
  assign o[37518] = i[37518];
  assign o[37517] = i[37517];
  assign o[37516] = i[37516];
  assign o[37515] = i[37515];
  assign o[37514] = i[37514];
  assign o[37513] = i[37513];
  assign o[37512] = i[37512];
  assign o[37511] = i[37511];
  assign o[37510] = i[37510];
  assign o[37509] = i[37509];
  assign o[37508] = i[37508];
  assign o[37507] = i[37507];
  assign o[37506] = i[37506];
  assign o[37505] = i[37505];
  assign o[37504] = i[37504];
  assign o[37503] = i[37503];
  assign o[37502] = i[37502];
  assign o[37501] = i[37501];
  assign o[37500] = i[37500];
  assign o[37499] = i[37499];
  assign o[37498] = i[37498];
  assign o[37497] = i[37497];
  assign o[37496] = i[37496];
  assign o[37495] = i[37495];
  assign o[37494] = i[37494];
  assign o[37493] = i[37493];
  assign o[37492] = i[37492];
  assign o[37491] = i[37491];
  assign o[37490] = i[37490];
  assign o[37489] = i[37489];
  assign o[37488] = i[37488];
  assign o[37487] = i[37487];
  assign o[37486] = i[37486];
  assign o[37485] = i[37485];
  assign o[37484] = i[37484];
  assign o[37483] = i[37483];
  assign o[37482] = i[37482];
  assign o[37481] = i[37481];
  assign o[37480] = i[37480];
  assign o[37479] = i[37479];
  assign o[37478] = i[37478];
  assign o[37477] = i[37477];
  assign o[37476] = i[37476];
  assign o[37475] = i[37475];
  assign o[37474] = i[37474];
  assign o[37473] = i[37473];
  assign o[37472] = i[37472];
  assign o[37471] = i[37471];
  assign o[37470] = i[37470];
  assign o[37469] = i[37469];
  assign o[37468] = i[37468];
  assign o[37467] = i[37467];
  assign o[37466] = i[37466];
  assign o[37465] = i[37465];
  assign o[37464] = i[37464];
  assign o[37463] = i[37463];
  assign o[37462] = i[37462];
  assign o[37461] = i[37461];
  assign o[37460] = i[37460];
  assign o[37459] = i[37459];
  assign o[37458] = i[37458];
  assign o[37457] = i[37457];
  assign o[37456] = i[37456];
  assign o[37455] = i[37455];
  assign o[37454] = i[37454];
  assign o[37453] = i[37453];
  assign o[37452] = i[37452];
  assign o[37451] = i[37451];
  assign o[37450] = i[37450];
  assign o[37449] = i[37449];
  assign o[37448] = i[37448];
  assign o[37447] = i[37447];
  assign o[37446] = i[37446];
  assign o[37445] = i[37445];
  assign o[37444] = i[37444];
  assign o[37443] = i[37443];
  assign o[37442] = i[37442];
  assign o[37441] = i[37441];
  assign o[37440] = i[37440];
  assign o[37439] = i[37439];
  assign o[37438] = i[37438];
  assign o[37437] = i[37437];
  assign o[37436] = i[37436];
  assign o[37435] = i[37435];
  assign o[37434] = i[37434];
  assign o[37433] = i[37433];
  assign o[37432] = i[37432];
  assign o[37431] = i[37431];
  assign o[37430] = i[37430];
  assign o[37429] = i[37429];
  assign o[37428] = i[37428];
  assign o[37427] = i[37427];
  assign o[37426] = i[37426];
  assign o[37425] = i[37425];
  assign o[37424] = i[37424];
  assign o[37423] = i[37423];
  assign o[37422] = i[37422];
  assign o[37421] = i[37421];
  assign o[37420] = i[37420];
  assign o[37419] = i[37419];
  assign o[37418] = i[37418];
  assign o[37417] = i[37417];
  assign o[37416] = i[37416];
  assign o[37415] = i[37415];
  assign o[37414] = i[37414];
  assign o[37413] = i[37413];
  assign o[37412] = i[37412];
  assign o[37411] = i[37411];
  assign o[37410] = i[37410];
  assign o[37409] = i[37409];
  assign o[37408] = i[37408];
  assign o[37407] = i[37407];
  assign o[37406] = i[37406];
  assign o[37405] = i[37405];
  assign o[37404] = i[37404];
  assign o[37403] = i[37403];
  assign o[37402] = i[37402];
  assign o[37401] = i[37401];
  assign o[37400] = i[37400];
  assign o[37399] = i[37399];
  assign o[37398] = i[37398];
  assign o[37397] = i[37397];
  assign o[37396] = i[37396];
  assign o[37395] = i[37395];
  assign o[37394] = i[37394];
  assign o[37393] = i[37393];
  assign o[37392] = i[37392];
  assign o[37391] = i[37391];
  assign o[37390] = i[37390];
  assign o[37389] = i[37389];
  assign o[37388] = i[37388];
  assign o[37387] = i[37387];
  assign o[37386] = i[37386];
  assign o[37385] = i[37385];
  assign o[37384] = i[37384];
  assign o[37383] = i[37383];
  assign o[37382] = i[37382];
  assign o[37381] = i[37381];
  assign o[37380] = i[37380];
  assign o[37379] = i[37379];
  assign o[37378] = i[37378];
  assign o[37377] = i[37377];
  assign o[37376] = i[37376];
  assign o[37375] = i[37375];
  assign o[37374] = i[37374];
  assign o[37373] = i[37373];
  assign o[37372] = i[37372];
  assign o[37371] = i[37371];
  assign o[37370] = i[37370];
  assign o[37369] = i[37369];
  assign o[37368] = i[37368];
  assign o[37367] = i[37367];
  assign o[37366] = i[37366];
  assign o[37365] = i[37365];
  assign o[37364] = i[37364];
  assign o[37363] = i[37363];
  assign o[37362] = i[37362];
  assign o[37361] = i[37361];
  assign o[37360] = i[37360];
  assign o[37359] = i[37359];
  assign o[37358] = i[37358];
  assign o[37357] = i[37357];
  assign o[37356] = i[37356];
  assign o[37355] = i[37355];
  assign o[37354] = i[37354];
  assign o[37353] = i[37353];
  assign o[37352] = i[37352];
  assign o[37351] = i[37351];
  assign o[37350] = i[37350];
  assign o[37349] = i[37349];
  assign o[37348] = i[37348];
  assign o[37347] = i[37347];
  assign o[37346] = i[37346];
  assign o[37345] = i[37345];
  assign o[37344] = i[37344];
  assign o[37343] = i[37343];
  assign o[37342] = i[37342];
  assign o[37341] = i[37341];
  assign o[37340] = i[37340];
  assign o[37339] = i[37339];
  assign o[37338] = i[37338];
  assign o[37337] = i[37337];
  assign o[37336] = i[37336];
  assign o[37335] = i[37335];
  assign o[37334] = i[37334];
  assign o[37333] = i[37333];
  assign o[37332] = i[37332];
  assign o[37331] = i[37331];
  assign o[37330] = i[37330];
  assign o[37329] = i[37329];
  assign o[37328] = i[37328];
  assign o[37327] = i[37327];
  assign o[37326] = i[37326];
  assign o[37325] = i[37325];
  assign o[37324] = i[37324];
  assign o[37323] = i[37323];
  assign o[37322] = i[37322];
  assign o[37321] = i[37321];
  assign o[37320] = i[37320];
  assign o[37319] = i[37319];
  assign o[37318] = i[37318];
  assign o[37317] = i[37317];
  assign o[37316] = i[37316];
  assign o[37315] = i[37315];
  assign o[37314] = i[37314];
  assign o[37313] = i[37313];
  assign o[37312] = i[37312];
  assign o[37311] = i[37311];
  assign o[37310] = i[37310];
  assign o[37309] = i[37309];
  assign o[37308] = i[37308];
  assign o[37307] = i[37307];
  assign o[37306] = i[37306];
  assign o[37305] = i[37305];
  assign o[37304] = i[37304];
  assign o[37303] = i[37303];
  assign o[37302] = i[37302];
  assign o[37301] = i[37301];
  assign o[37300] = i[37300];
  assign o[37299] = i[37299];
  assign o[37298] = i[37298];
  assign o[37297] = i[37297];
  assign o[37296] = i[37296];
  assign o[37295] = i[37295];
  assign o[37294] = i[37294];
  assign o[37293] = i[37293];
  assign o[37292] = i[37292];
  assign o[37291] = i[37291];
  assign o[37290] = i[37290];
  assign o[37289] = i[37289];
  assign o[37288] = i[37288];
  assign o[37287] = i[37287];
  assign o[37286] = i[37286];
  assign o[37285] = i[37285];
  assign o[37284] = i[37284];
  assign o[37283] = i[37283];
  assign o[37282] = i[37282];
  assign o[37281] = i[37281];
  assign o[37280] = i[37280];
  assign o[37279] = i[37279];
  assign o[37278] = i[37278];
  assign o[37277] = i[37277];
  assign o[37276] = i[37276];
  assign o[37275] = i[37275];
  assign o[37274] = i[37274];
  assign o[37273] = i[37273];
  assign o[37272] = i[37272];
  assign o[37271] = i[37271];
  assign o[37270] = i[37270];
  assign o[37269] = i[37269];
  assign o[37268] = i[37268];
  assign o[37267] = i[37267];
  assign o[37266] = i[37266];
  assign o[37265] = i[37265];
  assign o[37264] = i[37264];
  assign o[37263] = i[37263];
  assign o[37262] = i[37262];
  assign o[37261] = i[37261];
  assign o[37260] = i[37260];
  assign o[37259] = i[37259];
  assign o[37258] = i[37258];
  assign o[37257] = i[37257];
  assign o[37256] = i[37256];
  assign o[37255] = i[37255];
  assign o[37254] = i[37254];
  assign o[37253] = i[37253];
  assign o[37252] = i[37252];
  assign o[37251] = i[37251];
  assign o[37250] = i[37250];
  assign o[37249] = i[37249];
  assign o[37248] = i[37248];
  assign o[37247] = i[37247];
  assign o[37246] = i[37246];
  assign o[37245] = i[37245];
  assign o[37244] = i[37244];
  assign o[37243] = i[37243];
  assign o[37242] = i[37242];
  assign o[37241] = i[37241];
  assign o[37240] = i[37240];
  assign o[37239] = i[37239];
  assign o[37238] = i[37238];
  assign o[37237] = i[37237];
  assign o[37236] = i[37236];
  assign o[37235] = i[37235];
  assign o[37234] = i[37234];
  assign o[37233] = i[37233];
  assign o[37232] = i[37232];
  assign o[37231] = i[37231];
  assign o[37230] = i[37230];
  assign o[37229] = i[37229];
  assign o[37228] = i[37228];
  assign o[37227] = i[37227];
  assign o[37226] = i[37226];
  assign o[37225] = i[37225];
  assign o[37224] = i[37224];
  assign o[37223] = i[37223];
  assign o[37222] = i[37222];
  assign o[37221] = i[37221];
  assign o[37220] = i[37220];
  assign o[37219] = i[37219];
  assign o[37218] = i[37218];
  assign o[37217] = i[37217];
  assign o[37216] = i[37216];
  assign o[37215] = i[37215];
  assign o[37214] = i[37214];
  assign o[37213] = i[37213];
  assign o[37212] = i[37212];
  assign o[37211] = i[37211];
  assign o[37210] = i[37210];
  assign o[37209] = i[37209];
  assign o[37208] = i[37208];
  assign o[37207] = i[37207];
  assign o[37206] = i[37206];
  assign o[37205] = i[37205];
  assign o[37204] = i[37204];
  assign o[37203] = i[37203];
  assign o[37202] = i[37202];
  assign o[37201] = i[37201];
  assign o[37200] = i[37200];
  assign o[37199] = i[37199];
  assign o[37198] = i[37198];
  assign o[37197] = i[37197];
  assign o[37196] = i[37196];
  assign o[37195] = i[37195];
  assign o[37194] = i[37194];
  assign o[37193] = i[37193];
  assign o[37192] = i[37192];
  assign o[37191] = i[37191];
  assign o[37190] = i[37190];
  assign o[37189] = i[37189];
  assign o[37188] = i[37188];
  assign o[37187] = i[37187];
  assign o[37186] = i[37186];
  assign o[37185] = i[37185];
  assign o[37184] = i[37184];
  assign o[37183] = i[37183];
  assign o[37182] = i[37182];
  assign o[37181] = i[37181];
  assign o[37180] = i[37180];
  assign o[37179] = i[37179];
  assign o[37178] = i[37178];
  assign o[37177] = i[37177];
  assign o[37176] = i[37176];
  assign o[37175] = i[37175];
  assign o[37174] = i[37174];
  assign o[37173] = i[37173];
  assign o[37172] = i[37172];
  assign o[37171] = i[37171];
  assign o[37170] = i[37170];
  assign o[37169] = i[37169];
  assign o[37168] = i[37168];
  assign o[37167] = i[37167];
  assign o[37166] = i[37166];
  assign o[37165] = i[37165];
  assign o[37164] = i[37164];
  assign o[37163] = i[37163];
  assign o[37162] = i[37162];
  assign o[37161] = i[37161];
  assign o[37160] = i[37160];
  assign o[37159] = i[37159];
  assign o[37158] = i[37158];
  assign o[37157] = i[37157];
  assign o[37156] = i[37156];
  assign o[37155] = i[37155];
  assign o[37154] = i[37154];
  assign o[37153] = i[37153];
  assign o[37152] = i[37152];
  assign o[37151] = i[37151];
  assign o[37150] = i[37150];
  assign o[37149] = i[37149];
  assign o[37148] = i[37148];
  assign o[37147] = i[37147];
  assign o[37146] = i[37146];
  assign o[37145] = i[37145];
  assign o[37144] = i[37144];
  assign o[37143] = i[37143];
  assign o[37142] = i[37142];
  assign o[37141] = i[37141];
  assign o[37140] = i[37140];
  assign o[37139] = i[37139];
  assign o[37138] = i[37138];
  assign o[37137] = i[37137];
  assign o[37136] = i[37136];
  assign o[37135] = i[37135];
  assign o[37134] = i[37134];
  assign o[37133] = i[37133];
  assign o[37132] = i[37132];
  assign o[37131] = i[37131];
  assign o[37130] = i[37130];
  assign o[37129] = i[37129];
  assign o[37128] = i[37128];
  assign o[37127] = i[37127];
  assign o[37126] = i[37126];
  assign o[37125] = i[37125];
  assign o[37124] = i[37124];
  assign o[37123] = i[37123];
  assign o[37122] = i[37122];
  assign o[37121] = i[37121];
  assign o[37120] = i[37120];
  assign o[37119] = i[37119];
  assign o[37118] = i[37118];
  assign o[37117] = i[37117];
  assign o[37116] = i[37116];
  assign o[37115] = i[37115];
  assign o[37114] = i[37114];
  assign o[37113] = i[37113];
  assign o[37112] = i[37112];
  assign o[37111] = i[37111];
  assign o[37110] = i[37110];
  assign o[37109] = i[37109];
  assign o[37108] = i[37108];
  assign o[37107] = i[37107];
  assign o[37106] = i[37106];
  assign o[37105] = i[37105];
  assign o[37104] = i[37104];
  assign o[37103] = i[37103];
  assign o[37102] = i[37102];
  assign o[37101] = i[37101];
  assign o[37100] = i[37100];
  assign o[37099] = i[37099];
  assign o[37098] = i[37098];
  assign o[37097] = i[37097];
  assign o[37096] = i[37096];
  assign o[37095] = i[37095];
  assign o[37094] = i[37094];
  assign o[37093] = i[37093];
  assign o[37092] = i[37092];
  assign o[37091] = i[37091];
  assign o[37090] = i[37090];
  assign o[37089] = i[37089];
  assign o[37088] = i[37088];
  assign o[37087] = i[37087];
  assign o[37086] = i[37086];
  assign o[37085] = i[37085];
  assign o[37084] = i[37084];
  assign o[37083] = i[37083];
  assign o[37082] = i[37082];
  assign o[37081] = i[37081];
  assign o[37080] = i[37080];
  assign o[37079] = i[37079];
  assign o[37078] = i[37078];
  assign o[37077] = i[37077];
  assign o[37076] = i[37076];
  assign o[37075] = i[37075];
  assign o[37074] = i[37074];
  assign o[37073] = i[37073];
  assign o[37072] = i[37072];
  assign o[37071] = i[37071];
  assign o[37070] = i[37070];
  assign o[37069] = i[37069];
  assign o[37068] = i[37068];
  assign o[37067] = i[37067];
  assign o[37066] = i[37066];
  assign o[37065] = i[37065];
  assign o[37064] = i[37064];
  assign o[37063] = i[37063];
  assign o[37062] = i[37062];
  assign o[37061] = i[37061];
  assign o[37060] = i[37060];
  assign o[37059] = i[37059];
  assign o[37058] = i[37058];
  assign o[37057] = i[37057];
  assign o[37056] = i[37056];
  assign o[37055] = i[37055];
  assign o[37054] = i[37054];
  assign o[37053] = i[37053];
  assign o[37052] = i[37052];
  assign o[37051] = i[37051];
  assign o[37050] = i[37050];
  assign o[37049] = i[37049];
  assign o[37048] = i[37048];
  assign o[37047] = i[37047];
  assign o[37046] = i[37046];
  assign o[37045] = i[37045];
  assign o[37044] = i[37044];
  assign o[37043] = i[37043];
  assign o[37042] = i[37042];
  assign o[37041] = i[37041];
  assign o[37040] = i[37040];
  assign o[37039] = i[37039];
  assign o[37038] = i[37038];
  assign o[37037] = i[37037];
  assign o[37036] = i[37036];
  assign o[37035] = i[37035];
  assign o[37034] = i[37034];
  assign o[37033] = i[37033];
  assign o[37032] = i[37032];
  assign o[37031] = i[37031];
  assign o[37030] = i[37030];
  assign o[37029] = i[37029];
  assign o[37028] = i[37028];
  assign o[37027] = i[37027];
  assign o[37026] = i[37026];
  assign o[37025] = i[37025];
  assign o[37024] = i[37024];
  assign o[37023] = i[37023];
  assign o[37022] = i[37022];
  assign o[37021] = i[37021];
  assign o[37020] = i[37020];
  assign o[37019] = i[37019];
  assign o[37018] = i[37018];
  assign o[37017] = i[37017];
  assign o[37016] = i[37016];
  assign o[37015] = i[37015];
  assign o[37014] = i[37014];
  assign o[37013] = i[37013];
  assign o[37012] = i[37012];
  assign o[37011] = i[37011];
  assign o[37010] = i[37010];
  assign o[37009] = i[37009];
  assign o[37008] = i[37008];
  assign o[37007] = i[37007];
  assign o[37006] = i[37006];
  assign o[37005] = i[37005];
  assign o[37004] = i[37004];
  assign o[37003] = i[37003];
  assign o[37002] = i[37002];
  assign o[37001] = i[37001];
  assign o[37000] = i[37000];
  assign o[36999] = i[36999];
  assign o[36998] = i[36998];
  assign o[36997] = i[36997];
  assign o[36996] = i[36996];
  assign o[36995] = i[36995];
  assign o[36994] = i[36994];
  assign o[36993] = i[36993];
  assign o[36992] = i[36992];
  assign o[36991] = i[36991];
  assign o[36990] = i[36990];
  assign o[36989] = i[36989];
  assign o[36988] = i[36988];
  assign o[36987] = i[36987];
  assign o[36986] = i[36986];
  assign o[36985] = i[36985];
  assign o[36984] = i[36984];
  assign o[36983] = i[36983];
  assign o[36982] = i[36982];
  assign o[36981] = i[36981];
  assign o[36980] = i[36980];
  assign o[36979] = i[36979];
  assign o[36978] = i[36978];
  assign o[36977] = i[36977];
  assign o[36976] = i[36976];
  assign o[36975] = i[36975];
  assign o[36974] = i[36974];
  assign o[36973] = i[36973];
  assign o[36972] = i[36972];
  assign o[36971] = i[36971];
  assign o[36970] = i[36970];
  assign o[36969] = i[36969];
  assign o[36968] = i[36968];
  assign o[36967] = i[36967];
  assign o[36966] = i[36966];
  assign o[36965] = i[36965];
  assign o[36964] = i[36964];
  assign o[36963] = i[36963];
  assign o[36962] = i[36962];
  assign o[36961] = i[36961];
  assign o[36960] = i[36960];
  assign o[36959] = i[36959];
  assign o[36958] = i[36958];
  assign o[36957] = i[36957];
  assign o[36956] = i[36956];
  assign o[36955] = i[36955];
  assign o[36954] = i[36954];
  assign o[36953] = i[36953];
  assign o[36952] = i[36952];
  assign o[36951] = i[36951];
  assign o[36950] = i[36950];
  assign o[36949] = i[36949];
  assign o[36948] = i[36948];
  assign o[36947] = i[36947];
  assign o[36946] = i[36946];
  assign o[36945] = i[36945];
  assign o[36944] = i[36944];
  assign o[36943] = i[36943];
  assign o[36942] = i[36942];
  assign o[36941] = i[36941];
  assign o[36940] = i[36940];
  assign o[36939] = i[36939];
  assign o[36938] = i[36938];
  assign o[36937] = i[36937];
  assign o[36936] = i[36936];
  assign o[36935] = i[36935];
  assign o[36934] = i[36934];
  assign o[36933] = i[36933];
  assign o[36932] = i[36932];
  assign o[36931] = i[36931];
  assign o[36930] = i[36930];
  assign o[36929] = i[36929];
  assign o[36928] = i[36928];
  assign o[36927] = i[36927];
  assign o[36926] = i[36926];
  assign o[36925] = i[36925];
  assign o[36924] = i[36924];
  assign o[36923] = i[36923];
  assign o[36922] = i[36922];
  assign o[36921] = i[36921];
  assign o[36920] = i[36920];
  assign o[36919] = i[36919];
  assign o[36918] = i[36918];
  assign o[36917] = i[36917];
  assign o[36916] = i[36916];
  assign o[36915] = i[36915];
  assign o[36914] = i[36914];
  assign o[36913] = i[36913];
  assign o[36912] = i[36912];
  assign o[36911] = i[36911];
  assign o[36910] = i[36910];
  assign o[36909] = i[36909];
  assign o[36908] = i[36908];
  assign o[36907] = i[36907];
  assign o[36906] = i[36906];
  assign o[36905] = i[36905];
  assign o[36904] = i[36904];
  assign o[36903] = i[36903];
  assign o[36902] = i[36902];
  assign o[36901] = i[36901];
  assign o[36900] = i[36900];
  assign o[36899] = i[36899];
  assign o[36898] = i[36898];
  assign o[36897] = i[36897];
  assign o[36896] = i[36896];
  assign o[36895] = i[36895];
  assign o[36894] = i[36894];
  assign o[36893] = i[36893];
  assign o[36892] = i[36892];
  assign o[36891] = i[36891];
  assign o[36890] = i[36890];
  assign o[36889] = i[36889];
  assign o[36888] = i[36888];
  assign o[36887] = i[36887];
  assign o[36886] = i[36886];
  assign o[36885] = i[36885];
  assign o[36884] = i[36884];
  assign o[36883] = i[36883];
  assign o[36882] = i[36882];
  assign o[36881] = i[36881];
  assign o[36880] = i[36880];
  assign o[36879] = i[36879];
  assign o[36878] = i[36878];
  assign o[36877] = i[36877];
  assign o[36876] = i[36876];
  assign o[36875] = i[36875];
  assign o[36874] = i[36874];
  assign o[36873] = i[36873];
  assign o[36872] = i[36872];
  assign o[36871] = i[36871];
  assign o[36870] = i[36870];
  assign o[36869] = i[36869];
  assign o[36868] = i[36868];
  assign o[36867] = i[36867];
  assign o[36866] = i[36866];
  assign o[36865] = i[36865];
  assign o[36864] = i[36864];
  assign o[36863] = i[36863];
  assign o[36862] = i[36862];
  assign o[36861] = i[36861];
  assign o[36860] = i[36860];
  assign o[36859] = i[36859];
  assign o[36858] = i[36858];
  assign o[36857] = i[36857];
  assign o[36856] = i[36856];
  assign o[36855] = i[36855];
  assign o[36854] = i[36854];
  assign o[36853] = i[36853];
  assign o[36852] = i[36852];
  assign o[36851] = i[36851];
  assign o[36850] = i[36850];
  assign o[36849] = i[36849];
  assign o[36848] = i[36848];
  assign o[36847] = i[36847];
  assign o[36846] = i[36846];
  assign o[36845] = i[36845];
  assign o[36844] = i[36844];
  assign o[36843] = i[36843];
  assign o[36842] = i[36842];
  assign o[36841] = i[36841];
  assign o[36840] = i[36840];
  assign o[36839] = i[36839];
  assign o[36838] = i[36838];
  assign o[36837] = i[36837];
  assign o[36836] = i[36836];
  assign o[36835] = i[36835];
  assign o[36834] = i[36834];
  assign o[36833] = i[36833];
  assign o[36832] = i[36832];
  assign o[36831] = i[36831];
  assign o[36830] = i[36830];
  assign o[36829] = i[36829];
  assign o[36828] = i[36828];
  assign o[36827] = i[36827];
  assign o[36826] = i[36826];
  assign o[36825] = i[36825];
  assign o[36824] = i[36824];
  assign o[36823] = i[36823];
  assign o[36822] = i[36822];
  assign o[36821] = i[36821];
  assign o[36820] = i[36820];
  assign o[36819] = i[36819];
  assign o[36818] = i[36818];
  assign o[36817] = i[36817];
  assign o[36816] = i[36816];
  assign o[36815] = i[36815];
  assign o[36814] = i[36814];
  assign o[36813] = i[36813];
  assign o[36812] = i[36812];
  assign o[36811] = i[36811];
  assign o[36810] = i[36810];
  assign o[36809] = i[36809];
  assign o[36808] = i[36808];
  assign o[36807] = i[36807];
  assign o[36806] = i[36806];
  assign o[36805] = i[36805];
  assign o[36804] = i[36804];
  assign o[36803] = i[36803];
  assign o[36802] = i[36802];
  assign o[36801] = i[36801];
  assign o[36800] = i[36800];
  assign o[36799] = i[36799];
  assign o[36798] = i[36798];
  assign o[36797] = i[36797];
  assign o[36796] = i[36796];
  assign o[36795] = i[36795];
  assign o[36794] = i[36794];
  assign o[36793] = i[36793];
  assign o[36792] = i[36792];
  assign o[36791] = i[36791];
  assign o[36790] = i[36790];
  assign o[36789] = i[36789];
  assign o[36788] = i[36788];
  assign o[36787] = i[36787];
  assign o[36786] = i[36786];
  assign o[36785] = i[36785];
  assign o[36784] = i[36784];
  assign o[36783] = i[36783];
  assign o[36782] = i[36782];
  assign o[36781] = i[36781];
  assign o[36780] = i[36780];
  assign o[36779] = i[36779];
  assign o[36778] = i[36778];
  assign o[36777] = i[36777];
  assign o[36776] = i[36776];
  assign o[36775] = i[36775];
  assign o[36774] = i[36774];
  assign o[36773] = i[36773];
  assign o[36772] = i[36772];
  assign o[36771] = i[36771];
  assign o[36770] = i[36770];
  assign o[36769] = i[36769];
  assign o[36768] = i[36768];
  assign o[36767] = i[36767];
  assign o[36766] = i[36766];
  assign o[36765] = i[36765];
  assign o[36764] = i[36764];
  assign o[36763] = i[36763];
  assign o[36762] = i[36762];
  assign o[36761] = i[36761];
  assign o[36760] = i[36760];
  assign o[36759] = i[36759];
  assign o[36758] = i[36758];
  assign o[36757] = i[36757];
  assign o[36756] = i[36756];
  assign o[36755] = i[36755];
  assign o[36754] = i[36754];
  assign o[36753] = i[36753];
  assign o[36752] = i[36752];
  assign o[36751] = i[36751];
  assign o[36750] = i[36750];
  assign o[36749] = i[36749];
  assign o[36748] = i[36748];
  assign o[36747] = i[36747];
  assign o[36746] = i[36746];
  assign o[36745] = i[36745];
  assign o[36744] = i[36744];
  assign o[36743] = i[36743];
  assign o[36742] = i[36742];
  assign o[36741] = i[36741];
  assign o[36740] = i[36740];
  assign o[36739] = i[36739];
  assign o[36738] = i[36738];
  assign o[36737] = i[36737];
  assign o[36736] = i[36736];
  assign o[36735] = i[36735];
  assign o[36734] = i[36734];
  assign o[36733] = i[36733];
  assign o[36732] = i[36732];
  assign o[36731] = i[36731];
  assign o[36730] = i[36730];
  assign o[36729] = i[36729];
  assign o[36728] = i[36728];
  assign o[36727] = i[36727];
  assign o[36726] = i[36726];
  assign o[36725] = i[36725];
  assign o[36724] = i[36724];
  assign o[36723] = i[36723];
  assign o[36722] = i[36722];
  assign o[36721] = i[36721];
  assign o[36720] = i[36720];
  assign o[36719] = i[36719];
  assign o[36718] = i[36718];
  assign o[36717] = i[36717];
  assign o[36716] = i[36716];
  assign o[36715] = i[36715];
  assign o[36714] = i[36714];
  assign o[36713] = i[36713];
  assign o[36712] = i[36712];
  assign o[36711] = i[36711];
  assign o[36710] = i[36710];
  assign o[36709] = i[36709];
  assign o[36708] = i[36708];
  assign o[36707] = i[36707];
  assign o[36706] = i[36706];
  assign o[36705] = i[36705];
  assign o[36704] = i[36704];
  assign o[36703] = i[36703];
  assign o[36702] = i[36702];
  assign o[36701] = i[36701];
  assign o[36700] = i[36700];
  assign o[36699] = i[36699];
  assign o[36698] = i[36698];
  assign o[36697] = i[36697];
  assign o[36696] = i[36696];
  assign o[36695] = i[36695];
  assign o[36694] = i[36694];
  assign o[36693] = i[36693];
  assign o[36692] = i[36692];
  assign o[36691] = i[36691];
  assign o[36690] = i[36690];
  assign o[36689] = i[36689];
  assign o[36688] = i[36688];
  assign o[36687] = i[36687];
  assign o[36686] = i[36686];
  assign o[36685] = i[36685];
  assign o[36684] = i[36684];
  assign o[36683] = i[36683];
  assign o[36682] = i[36682];
  assign o[36681] = i[36681];
  assign o[36680] = i[36680];
  assign o[36679] = i[36679];
  assign o[36678] = i[36678];
  assign o[36677] = i[36677];
  assign o[36676] = i[36676];
  assign o[36675] = i[36675];
  assign o[36674] = i[36674];
  assign o[36673] = i[36673];
  assign o[36672] = i[36672];
  assign o[36671] = i[36671];
  assign o[36670] = i[36670];
  assign o[36669] = i[36669];
  assign o[36668] = i[36668];
  assign o[36667] = i[36667];
  assign o[36666] = i[36666];
  assign o[36665] = i[36665];
  assign o[36664] = i[36664];
  assign o[36663] = i[36663];
  assign o[36662] = i[36662];
  assign o[36661] = i[36661];
  assign o[36660] = i[36660];
  assign o[36659] = i[36659];
  assign o[36658] = i[36658];
  assign o[36657] = i[36657];
  assign o[36656] = i[36656];
  assign o[36655] = i[36655];
  assign o[36654] = i[36654];
  assign o[36653] = i[36653];
  assign o[36652] = i[36652];
  assign o[36651] = i[36651];
  assign o[36650] = i[36650];
  assign o[36649] = i[36649];
  assign o[36648] = i[36648];
  assign o[36647] = i[36647];
  assign o[36646] = i[36646];
  assign o[36645] = i[36645];
  assign o[36644] = i[36644];
  assign o[36643] = i[36643];
  assign o[36642] = i[36642];
  assign o[36641] = i[36641];
  assign o[36640] = i[36640];
  assign o[36639] = i[36639];
  assign o[36638] = i[36638];
  assign o[36637] = i[36637];
  assign o[36636] = i[36636];
  assign o[36635] = i[36635];
  assign o[36634] = i[36634];
  assign o[36633] = i[36633];
  assign o[36632] = i[36632];
  assign o[36631] = i[36631];
  assign o[36630] = i[36630];
  assign o[36629] = i[36629];
  assign o[36628] = i[36628];
  assign o[36627] = i[36627];
  assign o[36626] = i[36626];
  assign o[36625] = i[36625];
  assign o[36624] = i[36624];
  assign o[36623] = i[36623];
  assign o[36622] = i[36622];
  assign o[36621] = i[36621];
  assign o[36620] = i[36620];
  assign o[36619] = i[36619];
  assign o[36618] = i[36618];
  assign o[36617] = i[36617];
  assign o[36616] = i[36616];
  assign o[36615] = i[36615];
  assign o[36614] = i[36614];
  assign o[36613] = i[36613];
  assign o[36612] = i[36612];
  assign o[36611] = i[36611];
  assign o[36610] = i[36610];
  assign o[36609] = i[36609];
  assign o[36608] = i[36608];
  assign o[36607] = i[36607];
  assign o[36606] = i[36606];
  assign o[36605] = i[36605];
  assign o[36604] = i[36604];
  assign o[36603] = i[36603];
  assign o[36602] = i[36602];
  assign o[36601] = i[36601];
  assign o[36600] = i[36600];
  assign o[36599] = i[36599];
  assign o[36598] = i[36598];
  assign o[36597] = i[36597];
  assign o[36596] = i[36596];
  assign o[36595] = i[36595];
  assign o[36594] = i[36594];
  assign o[36593] = i[36593];
  assign o[36592] = i[36592];
  assign o[36591] = i[36591];
  assign o[36590] = i[36590];
  assign o[36589] = i[36589];
  assign o[36588] = i[36588];
  assign o[36587] = i[36587];
  assign o[36586] = i[36586];
  assign o[36585] = i[36585];
  assign o[36584] = i[36584];
  assign o[36583] = i[36583];
  assign o[36582] = i[36582];
  assign o[36581] = i[36581];
  assign o[36580] = i[36580];
  assign o[36579] = i[36579];
  assign o[36578] = i[36578];
  assign o[36577] = i[36577];
  assign o[36576] = i[36576];
  assign o[36575] = i[36575];
  assign o[36574] = i[36574];
  assign o[36573] = i[36573];
  assign o[36572] = i[36572];
  assign o[36571] = i[36571];
  assign o[36570] = i[36570];
  assign o[36569] = i[36569];
  assign o[36568] = i[36568];
  assign o[36567] = i[36567];
  assign o[36566] = i[36566];
  assign o[36565] = i[36565];
  assign o[36564] = i[36564];
  assign o[36563] = i[36563];
  assign o[36562] = i[36562];
  assign o[36561] = i[36561];
  assign o[36560] = i[36560];
  assign o[36559] = i[36559];
  assign o[36558] = i[36558];
  assign o[36557] = i[36557];
  assign o[36556] = i[36556];
  assign o[36555] = i[36555];
  assign o[36554] = i[36554];
  assign o[36553] = i[36553];
  assign o[36552] = i[36552];
  assign o[36551] = i[36551];
  assign o[36550] = i[36550];
  assign o[36549] = i[36549];
  assign o[36548] = i[36548];
  assign o[36547] = i[36547];
  assign o[36546] = i[36546];
  assign o[36545] = i[36545];
  assign o[36544] = i[36544];
  assign o[36543] = i[36543];
  assign o[36542] = i[36542];
  assign o[36541] = i[36541];
  assign o[36540] = i[36540];
  assign o[36539] = i[36539];
  assign o[36538] = i[36538];
  assign o[36537] = i[36537];
  assign o[36536] = i[36536];
  assign o[36535] = i[36535];
  assign o[36534] = i[36534];
  assign o[36533] = i[36533];
  assign o[36532] = i[36532];
  assign o[36531] = i[36531];
  assign o[36530] = i[36530];
  assign o[36529] = i[36529];
  assign o[36528] = i[36528];
  assign o[36527] = i[36527];
  assign o[36526] = i[36526];
  assign o[36525] = i[36525];
  assign o[36524] = i[36524];
  assign o[36523] = i[36523];
  assign o[36522] = i[36522];
  assign o[36521] = i[36521];
  assign o[36520] = i[36520];
  assign o[36519] = i[36519];
  assign o[36518] = i[36518];
  assign o[36517] = i[36517];
  assign o[36516] = i[36516];
  assign o[36515] = i[36515];
  assign o[36514] = i[36514];
  assign o[36513] = i[36513];
  assign o[36512] = i[36512];
  assign o[36511] = i[36511];
  assign o[36510] = i[36510];
  assign o[36509] = i[36509];
  assign o[36508] = i[36508];
  assign o[36507] = i[36507];
  assign o[36506] = i[36506];
  assign o[36505] = i[36505];
  assign o[36504] = i[36504];
  assign o[36503] = i[36503];
  assign o[36502] = i[36502];
  assign o[36501] = i[36501];
  assign o[36500] = i[36500];
  assign o[36499] = i[36499];
  assign o[36498] = i[36498];
  assign o[36497] = i[36497];
  assign o[36496] = i[36496];
  assign o[36495] = i[36495];
  assign o[36494] = i[36494];
  assign o[36493] = i[36493];
  assign o[36492] = i[36492];
  assign o[36491] = i[36491];
  assign o[36490] = i[36490];
  assign o[36489] = i[36489];
  assign o[36488] = i[36488];
  assign o[36487] = i[36487];
  assign o[36486] = i[36486];
  assign o[36485] = i[36485];
  assign o[36484] = i[36484];
  assign o[36483] = i[36483];
  assign o[36482] = i[36482];
  assign o[36481] = i[36481];
  assign o[36480] = i[36480];
  assign o[36479] = i[36479];
  assign o[36478] = i[36478];
  assign o[36477] = i[36477];
  assign o[36476] = i[36476];
  assign o[36475] = i[36475];
  assign o[36474] = i[36474];
  assign o[36473] = i[36473];
  assign o[36472] = i[36472];
  assign o[36471] = i[36471];
  assign o[36470] = i[36470];
  assign o[36469] = i[36469];
  assign o[36468] = i[36468];
  assign o[36467] = i[36467];
  assign o[36466] = i[36466];
  assign o[36465] = i[36465];
  assign o[36464] = i[36464];
  assign o[36463] = i[36463];
  assign o[36462] = i[36462];
  assign o[36461] = i[36461];
  assign o[36460] = i[36460];
  assign o[36459] = i[36459];
  assign o[36458] = i[36458];
  assign o[36457] = i[36457];
  assign o[36456] = i[36456];
  assign o[36455] = i[36455];
  assign o[36454] = i[36454];
  assign o[36453] = i[36453];
  assign o[36452] = i[36452];
  assign o[36451] = i[36451];
  assign o[36450] = i[36450];
  assign o[36449] = i[36449];
  assign o[36448] = i[36448];
  assign o[36447] = i[36447];
  assign o[36446] = i[36446];
  assign o[36445] = i[36445];
  assign o[36444] = i[36444];
  assign o[36443] = i[36443];
  assign o[36442] = i[36442];
  assign o[36441] = i[36441];
  assign o[36440] = i[36440];
  assign o[36439] = i[36439];
  assign o[36438] = i[36438];
  assign o[36437] = i[36437];
  assign o[36436] = i[36436];
  assign o[36435] = i[36435];
  assign o[36434] = i[36434];
  assign o[36433] = i[36433];
  assign o[36432] = i[36432];
  assign o[36431] = i[36431];
  assign o[36430] = i[36430];
  assign o[36429] = i[36429];
  assign o[36428] = i[36428];
  assign o[36427] = i[36427];
  assign o[36426] = i[36426];
  assign o[36425] = i[36425];
  assign o[36424] = i[36424];
  assign o[36423] = i[36423];
  assign o[36422] = i[36422];
  assign o[36421] = i[36421];
  assign o[36420] = i[36420];
  assign o[36419] = i[36419];
  assign o[36418] = i[36418];
  assign o[36417] = i[36417];
  assign o[36416] = i[36416];
  assign o[36415] = i[36415];
  assign o[36414] = i[36414];
  assign o[36413] = i[36413];
  assign o[36412] = i[36412];
  assign o[36411] = i[36411];
  assign o[36410] = i[36410];
  assign o[36409] = i[36409];
  assign o[36408] = i[36408];
  assign o[36407] = i[36407];
  assign o[36406] = i[36406];
  assign o[36405] = i[36405];
  assign o[36404] = i[36404];
  assign o[36403] = i[36403];
  assign o[36402] = i[36402];
  assign o[36401] = i[36401];
  assign o[36400] = i[36400];
  assign o[36399] = i[36399];
  assign o[36398] = i[36398];
  assign o[36397] = i[36397];
  assign o[36396] = i[36396];
  assign o[36395] = i[36395];
  assign o[36394] = i[36394];
  assign o[36393] = i[36393];
  assign o[36392] = i[36392];
  assign o[36391] = i[36391];
  assign o[36390] = i[36390];
  assign o[36389] = i[36389];
  assign o[36388] = i[36388];
  assign o[36387] = i[36387];
  assign o[36386] = i[36386];
  assign o[36385] = i[36385];
  assign o[36384] = i[36384];
  assign o[36383] = i[36383];
  assign o[36382] = i[36382];
  assign o[36381] = i[36381];
  assign o[36380] = i[36380];
  assign o[36379] = i[36379];
  assign o[36378] = i[36378];
  assign o[36377] = i[36377];
  assign o[36376] = i[36376];
  assign o[36375] = i[36375];
  assign o[36374] = i[36374];
  assign o[36373] = i[36373];
  assign o[36372] = i[36372];
  assign o[36371] = i[36371];
  assign o[36370] = i[36370];
  assign o[36369] = i[36369];
  assign o[36368] = i[36368];
  assign o[36367] = i[36367];
  assign o[36366] = i[36366];
  assign o[36365] = i[36365];
  assign o[36364] = i[36364];
  assign o[36363] = i[36363];
  assign o[36362] = i[36362];
  assign o[36361] = i[36361];
  assign o[36360] = i[36360];
  assign o[36359] = i[36359];
  assign o[36358] = i[36358];
  assign o[36357] = i[36357];
  assign o[36356] = i[36356];
  assign o[36355] = i[36355];
  assign o[36354] = i[36354];
  assign o[36353] = i[36353];
  assign o[36352] = i[36352];
  assign o[36351] = i[36351];
  assign o[36350] = i[36350];
  assign o[36349] = i[36349];
  assign o[36348] = i[36348];
  assign o[36347] = i[36347];
  assign o[36346] = i[36346];
  assign o[36345] = i[36345];
  assign o[36344] = i[36344];
  assign o[36343] = i[36343];
  assign o[36342] = i[36342];
  assign o[36341] = i[36341];
  assign o[36340] = i[36340];
  assign o[36339] = i[36339];
  assign o[36338] = i[36338];
  assign o[36337] = i[36337];
  assign o[36336] = i[36336];
  assign o[36335] = i[36335];
  assign o[36334] = i[36334];
  assign o[36333] = i[36333];
  assign o[36332] = i[36332];
  assign o[36331] = i[36331];
  assign o[36330] = i[36330];
  assign o[36329] = i[36329];
  assign o[36328] = i[36328];
  assign o[36327] = i[36327];
  assign o[36326] = i[36326];
  assign o[36325] = i[36325];
  assign o[36324] = i[36324];
  assign o[36323] = i[36323];
  assign o[36322] = i[36322];
  assign o[36321] = i[36321];
  assign o[36320] = i[36320];
  assign o[36319] = i[36319];
  assign o[36318] = i[36318];
  assign o[36317] = i[36317];
  assign o[36316] = i[36316];
  assign o[36315] = i[36315];
  assign o[36314] = i[36314];
  assign o[36313] = i[36313];
  assign o[36312] = i[36312];
  assign o[36311] = i[36311];
  assign o[36310] = i[36310];
  assign o[36309] = i[36309];
  assign o[36308] = i[36308];
  assign o[36307] = i[36307];
  assign o[36306] = i[36306];
  assign o[36305] = i[36305];
  assign o[36304] = i[36304];
  assign o[36303] = i[36303];
  assign o[36302] = i[36302];
  assign o[36301] = i[36301];
  assign o[36300] = i[36300];
  assign o[36299] = i[36299];
  assign o[36298] = i[36298];
  assign o[36297] = i[36297];
  assign o[36296] = i[36296];
  assign o[36295] = i[36295];
  assign o[36294] = i[36294];
  assign o[36293] = i[36293];
  assign o[36292] = i[36292];
  assign o[36291] = i[36291];
  assign o[36290] = i[36290];
  assign o[36289] = i[36289];
  assign o[36288] = i[36288];
  assign o[36287] = i[36287];
  assign o[36286] = i[36286];
  assign o[36285] = i[36285];
  assign o[36284] = i[36284];
  assign o[36283] = i[36283];
  assign o[36282] = i[36282];
  assign o[36281] = i[36281];
  assign o[36280] = i[36280];
  assign o[36279] = i[36279];
  assign o[36278] = i[36278];
  assign o[36277] = i[36277];
  assign o[36276] = i[36276];
  assign o[36275] = i[36275];
  assign o[36274] = i[36274];
  assign o[36273] = i[36273];
  assign o[36272] = i[36272];
  assign o[36271] = i[36271];
  assign o[36270] = i[36270];
  assign o[36269] = i[36269];
  assign o[36268] = i[36268];
  assign o[36267] = i[36267];
  assign o[36266] = i[36266];
  assign o[36265] = i[36265];
  assign o[36264] = i[36264];
  assign o[36263] = i[36263];
  assign o[36262] = i[36262];
  assign o[36261] = i[36261];
  assign o[36260] = i[36260];
  assign o[36259] = i[36259];
  assign o[36258] = i[36258];
  assign o[36257] = i[36257];
  assign o[36256] = i[36256];
  assign o[36255] = i[36255];
  assign o[36254] = i[36254];
  assign o[36253] = i[36253];
  assign o[36252] = i[36252];
  assign o[36251] = i[36251];
  assign o[36250] = i[36250];
  assign o[36249] = i[36249];
  assign o[36248] = i[36248];
  assign o[36247] = i[36247];
  assign o[36246] = i[36246];
  assign o[36245] = i[36245];
  assign o[36244] = i[36244];
  assign o[36243] = i[36243];
  assign o[36242] = i[36242];
  assign o[36241] = i[36241];
  assign o[36240] = i[36240];
  assign o[36239] = i[36239];
  assign o[36238] = i[36238];
  assign o[36237] = i[36237];
  assign o[36236] = i[36236];
  assign o[36235] = i[36235];
  assign o[36234] = i[36234];
  assign o[36233] = i[36233];
  assign o[36232] = i[36232];
  assign o[36231] = i[36231];
  assign o[36230] = i[36230];
  assign o[36229] = i[36229];
  assign o[36228] = i[36228];
  assign o[36227] = i[36227];
  assign o[36226] = i[36226];
  assign o[36225] = i[36225];
  assign o[36224] = i[36224];
  assign o[36223] = i[36223];
  assign o[36222] = i[36222];
  assign o[36221] = i[36221];
  assign o[36220] = i[36220];
  assign o[36219] = i[36219];
  assign o[36218] = i[36218];
  assign o[36217] = i[36217];
  assign o[36216] = i[36216];
  assign o[36215] = i[36215];
  assign o[36214] = i[36214];
  assign o[36213] = i[36213];
  assign o[36212] = i[36212];
  assign o[36211] = i[36211];
  assign o[36210] = i[36210];
  assign o[36209] = i[36209];
  assign o[36208] = i[36208];
  assign o[36207] = i[36207];
  assign o[36206] = i[36206];
  assign o[36205] = i[36205];
  assign o[36204] = i[36204];
  assign o[36203] = i[36203];
  assign o[36202] = i[36202];
  assign o[36201] = i[36201];
  assign o[36200] = i[36200];
  assign o[36199] = i[36199];
  assign o[36198] = i[36198];
  assign o[36197] = i[36197];
  assign o[36196] = i[36196];
  assign o[36195] = i[36195];
  assign o[36194] = i[36194];
  assign o[36193] = i[36193];
  assign o[36192] = i[36192];
  assign o[36191] = i[36191];
  assign o[36190] = i[36190];
  assign o[36189] = i[36189];
  assign o[36188] = i[36188];
  assign o[36187] = i[36187];
  assign o[36186] = i[36186];
  assign o[36185] = i[36185];
  assign o[36184] = i[36184];
  assign o[36183] = i[36183];
  assign o[36182] = i[36182];
  assign o[36181] = i[36181];
  assign o[36180] = i[36180];
  assign o[36179] = i[36179];
  assign o[36178] = i[36178];
  assign o[36177] = i[36177];
  assign o[36176] = i[36176];
  assign o[36175] = i[36175];
  assign o[36174] = i[36174];
  assign o[36173] = i[36173];
  assign o[36172] = i[36172];
  assign o[36171] = i[36171];
  assign o[36170] = i[36170];
  assign o[36169] = i[36169];
  assign o[36168] = i[36168];
  assign o[36167] = i[36167];
  assign o[36166] = i[36166];
  assign o[36165] = i[36165];
  assign o[36164] = i[36164];
  assign o[36163] = i[36163];
  assign o[36162] = i[36162];
  assign o[36161] = i[36161];
  assign o[36160] = i[36160];
  assign o[36159] = i[36159];
  assign o[36158] = i[36158];
  assign o[36157] = i[36157];
  assign o[36156] = i[36156];
  assign o[36155] = i[36155];
  assign o[36154] = i[36154];
  assign o[36153] = i[36153];
  assign o[36152] = i[36152];
  assign o[36151] = i[36151];
  assign o[36150] = i[36150];
  assign o[36149] = i[36149];
  assign o[36148] = i[36148];
  assign o[36147] = i[36147];
  assign o[36146] = i[36146];
  assign o[36145] = i[36145];
  assign o[36144] = i[36144];
  assign o[36143] = i[36143];
  assign o[36142] = i[36142];
  assign o[36141] = i[36141];
  assign o[36140] = i[36140];
  assign o[36139] = i[36139];
  assign o[36138] = i[36138];
  assign o[36137] = i[36137];
  assign o[36136] = i[36136];
  assign o[36135] = i[36135];
  assign o[36134] = i[36134];
  assign o[36133] = i[36133];
  assign o[36132] = i[36132];
  assign o[36131] = i[36131];
  assign o[36130] = i[36130];
  assign o[36129] = i[36129];
  assign o[36128] = i[36128];
  assign o[36127] = i[36127];
  assign o[36126] = i[36126];
  assign o[36125] = i[36125];
  assign o[36124] = i[36124];
  assign o[36123] = i[36123];
  assign o[36122] = i[36122];
  assign o[36121] = i[36121];
  assign o[36120] = i[36120];
  assign o[36119] = i[36119];
  assign o[36118] = i[36118];
  assign o[36117] = i[36117];
  assign o[36116] = i[36116];
  assign o[36115] = i[36115];
  assign o[36114] = i[36114];
  assign o[36113] = i[36113];
  assign o[36112] = i[36112];
  assign o[36111] = i[36111];
  assign o[36110] = i[36110];
  assign o[36109] = i[36109];
  assign o[36108] = i[36108];
  assign o[36107] = i[36107];
  assign o[36106] = i[36106];
  assign o[36105] = i[36105];
  assign o[36104] = i[36104];
  assign o[36103] = i[36103];
  assign o[36102] = i[36102];
  assign o[36101] = i[36101];
  assign o[36100] = i[36100];
  assign o[36099] = i[36099];
  assign o[36098] = i[36098];
  assign o[36097] = i[36097];
  assign o[36096] = i[36096];
  assign o[36095] = i[36095];
  assign o[36094] = i[36094];
  assign o[36093] = i[36093];
  assign o[36092] = i[36092];
  assign o[36091] = i[36091];
  assign o[36090] = i[36090];
  assign o[36089] = i[36089];
  assign o[36088] = i[36088];
  assign o[36087] = i[36087];
  assign o[36086] = i[36086];
  assign o[36085] = i[36085];
  assign o[36084] = i[36084];
  assign o[36083] = i[36083];
  assign o[36082] = i[36082];
  assign o[36081] = i[36081];
  assign o[36080] = i[36080];
  assign o[36079] = i[36079];
  assign o[36078] = i[36078];
  assign o[36077] = i[36077];
  assign o[36076] = i[36076];
  assign o[36075] = i[36075];
  assign o[36074] = i[36074];
  assign o[36073] = i[36073];
  assign o[36072] = i[36072];
  assign o[36071] = i[36071];
  assign o[36070] = i[36070];
  assign o[36069] = i[36069];
  assign o[36068] = i[36068];
  assign o[36067] = i[36067];
  assign o[36066] = i[36066];
  assign o[36065] = i[36065];
  assign o[36064] = i[36064];
  assign o[36063] = i[36063];
  assign o[36062] = i[36062];
  assign o[36061] = i[36061];
  assign o[36060] = i[36060];
  assign o[36059] = i[36059];
  assign o[36058] = i[36058];
  assign o[36057] = i[36057];
  assign o[36056] = i[36056];
  assign o[36055] = i[36055];
  assign o[36054] = i[36054];
  assign o[36053] = i[36053];
  assign o[36052] = i[36052];
  assign o[36051] = i[36051];
  assign o[36050] = i[36050];
  assign o[36049] = i[36049];
  assign o[36048] = i[36048];
  assign o[36047] = i[36047];
  assign o[36046] = i[36046];
  assign o[36045] = i[36045];
  assign o[36044] = i[36044];
  assign o[36043] = i[36043];
  assign o[36042] = i[36042];
  assign o[36041] = i[36041];
  assign o[36040] = i[36040];
  assign o[36039] = i[36039];
  assign o[36038] = i[36038];
  assign o[36037] = i[36037];
  assign o[36036] = i[36036];
  assign o[36035] = i[36035];
  assign o[36034] = i[36034];
  assign o[36033] = i[36033];
  assign o[36032] = i[36032];
  assign o[36031] = i[36031];
  assign o[36030] = i[36030];
  assign o[36029] = i[36029];
  assign o[36028] = i[36028];
  assign o[36027] = i[36027];
  assign o[36026] = i[36026];
  assign o[36025] = i[36025];
  assign o[36024] = i[36024];
  assign o[36023] = i[36023];
  assign o[36022] = i[36022];
  assign o[36021] = i[36021];
  assign o[36020] = i[36020];
  assign o[36019] = i[36019];
  assign o[36018] = i[36018];
  assign o[36017] = i[36017];
  assign o[36016] = i[36016];
  assign o[36015] = i[36015];
  assign o[36014] = i[36014];
  assign o[36013] = i[36013];
  assign o[36012] = i[36012];
  assign o[36011] = i[36011];
  assign o[36010] = i[36010];
  assign o[36009] = i[36009];
  assign o[36008] = i[36008];
  assign o[36007] = i[36007];
  assign o[36006] = i[36006];
  assign o[36005] = i[36005];
  assign o[36004] = i[36004];
  assign o[36003] = i[36003];
  assign o[36002] = i[36002];
  assign o[36001] = i[36001];
  assign o[36000] = i[36000];
  assign o[35999] = i[35999];
  assign o[35998] = i[35998];
  assign o[35997] = i[35997];
  assign o[35996] = i[35996];
  assign o[35995] = i[35995];
  assign o[35994] = i[35994];
  assign o[35993] = i[35993];
  assign o[35992] = i[35992];
  assign o[35991] = i[35991];
  assign o[35990] = i[35990];
  assign o[35989] = i[35989];
  assign o[35988] = i[35988];
  assign o[35987] = i[35987];
  assign o[35986] = i[35986];
  assign o[35985] = i[35985];
  assign o[35984] = i[35984];
  assign o[35983] = i[35983];
  assign o[35982] = i[35982];
  assign o[35981] = i[35981];
  assign o[35980] = i[35980];
  assign o[35979] = i[35979];
  assign o[35978] = i[35978];
  assign o[35977] = i[35977];
  assign o[35976] = i[35976];
  assign o[35975] = i[35975];
  assign o[35974] = i[35974];
  assign o[35973] = i[35973];
  assign o[35972] = i[35972];
  assign o[35971] = i[35971];
  assign o[35970] = i[35970];
  assign o[35969] = i[35969];
  assign o[35968] = i[35968];
  assign o[35967] = i[35967];
  assign o[35966] = i[35966];
  assign o[35965] = i[35965];
  assign o[35964] = i[35964];
  assign o[35963] = i[35963];
  assign o[35962] = i[35962];
  assign o[35961] = i[35961];
  assign o[35960] = i[35960];
  assign o[35959] = i[35959];
  assign o[35958] = i[35958];
  assign o[35957] = i[35957];
  assign o[35956] = i[35956];
  assign o[35955] = i[35955];
  assign o[35954] = i[35954];
  assign o[35953] = i[35953];
  assign o[35952] = i[35952];
  assign o[35951] = i[35951];
  assign o[35950] = i[35950];
  assign o[35949] = i[35949];
  assign o[35948] = i[35948];
  assign o[35947] = i[35947];
  assign o[35946] = i[35946];
  assign o[35945] = i[35945];
  assign o[35944] = i[35944];
  assign o[35943] = i[35943];
  assign o[35942] = i[35942];
  assign o[35941] = i[35941];
  assign o[35940] = i[35940];
  assign o[35939] = i[35939];
  assign o[35938] = i[35938];
  assign o[35937] = i[35937];
  assign o[35936] = i[35936];
  assign o[35935] = i[35935];
  assign o[35934] = i[35934];
  assign o[35933] = i[35933];
  assign o[35932] = i[35932];
  assign o[35931] = i[35931];
  assign o[35930] = i[35930];
  assign o[35929] = i[35929];
  assign o[35928] = i[35928];
  assign o[35927] = i[35927];
  assign o[35926] = i[35926];
  assign o[35925] = i[35925];
  assign o[35924] = i[35924];
  assign o[35923] = i[35923];
  assign o[35922] = i[35922];
  assign o[35921] = i[35921];
  assign o[35920] = i[35920];
  assign o[35919] = i[35919];
  assign o[35918] = i[35918];
  assign o[35917] = i[35917];
  assign o[35916] = i[35916];
  assign o[35915] = i[35915];
  assign o[35914] = i[35914];
  assign o[35913] = i[35913];
  assign o[35912] = i[35912];
  assign o[35911] = i[35911];
  assign o[35910] = i[35910];
  assign o[35909] = i[35909];
  assign o[35908] = i[35908];
  assign o[35907] = i[35907];
  assign o[35906] = i[35906];
  assign o[35905] = i[35905];
  assign o[35904] = i[35904];
  assign o[35903] = i[35903];
  assign o[35902] = i[35902];
  assign o[35901] = i[35901];
  assign o[35900] = i[35900];
  assign o[35899] = i[35899];
  assign o[35898] = i[35898];
  assign o[35897] = i[35897];
  assign o[35896] = i[35896];
  assign o[35895] = i[35895];
  assign o[35894] = i[35894];
  assign o[35893] = i[35893];
  assign o[35892] = i[35892];
  assign o[35891] = i[35891];
  assign o[35890] = i[35890];
  assign o[35889] = i[35889];
  assign o[35888] = i[35888];
  assign o[35887] = i[35887];
  assign o[35886] = i[35886];
  assign o[35885] = i[35885];
  assign o[35884] = i[35884];
  assign o[35883] = i[35883];
  assign o[35882] = i[35882];
  assign o[35881] = i[35881];
  assign o[35880] = i[35880];
  assign o[35879] = i[35879];
  assign o[35878] = i[35878];
  assign o[35877] = i[35877];
  assign o[35876] = i[35876];
  assign o[35875] = i[35875];
  assign o[35874] = i[35874];
  assign o[35873] = i[35873];
  assign o[35872] = i[35872];
  assign o[35871] = i[35871];
  assign o[35870] = i[35870];
  assign o[35869] = i[35869];
  assign o[35868] = i[35868];
  assign o[35867] = i[35867];
  assign o[35866] = i[35866];
  assign o[35865] = i[35865];
  assign o[35864] = i[35864];
  assign o[35863] = i[35863];
  assign o[35862] = i[35862];
  assign o[35861] = i[35861];
  assign o[35860] = i[35860];
  assign o[35859] = i[35859];
  assign o[35858] = i[35858];
  assign o[35857] = i[35857];
  assign o[35856] = i[35856];
  assign o[35855] = i[35855];
  assign o[35854] = i[35854];
  assign o[35853] = i[35853];
  assign o[35852] = i[35852];
  assign o[35851] = i[35851];
  assign o[35850] = i[35850];
  assign o[35849] = i[35849];
  assign o[35848] = i[35848];
  assign o[35847] = i[35847];
  assign o[35846] = i[35846];
  assign o[35845] = i[35845];
  assign o[35844] = i[35844];
  assign o[35843] = i[35843];
  assign o[35842] = i[35842];
  assign o[35841] = i[35841];
  assign o[35840] = i[35840];
  assign o[35839] = i[35839];
  assign o[35838] = i[35838];
  assign o[35837] = i[35837];
  assign o[35836] = i[35836];
  assign o[35835] = i[35835];
  assign o[35834] = i[35834];
  assign o[35833] = i[35833];
  assign o[35832] = i[35832];
  assign o[35831] = i[35831];
  assign o[35830] = i[35830];
  assign o[35829] = i[35829];
  assign o[35828] = i[35828];
  assign o[35827] = i[35827];
  assign o[35826] = i[35826];
  assign o[35825] = i[35825];
  assign o[35824] = i[35824];
  assign o[35823] = i[35823];
  assign o[35822] = i[35822];
  assign o[35821] = i[35821];
  assign o[35820] = i[35820];
  assign o[35819] = i[35819];
  assign o[35818] = i[35818];
  assign o[35817] = i[35817];
  assign o[35816] = i[35816];
  assign o[35815] = i[35815];
  assign o[35814] = i[35814];
  assign o[35813] = i[35813];
  assign o[35812] = i[35812];
  assign o[35811] = i[35811];
  assign o[35810] = i[35810];
  assign o[35809] = i[35809];
  assign o[35808] = i[35808];
  assign o[35807] = i[35807];
  assign o[35806] = i[35806];
  assign o[35805] = i[35805];
  assign o[35804] = i[35804];
  assign o[35803] = i[35803];
  assign o[35802] = i[35802];
  assign o[35801] = i[35801];
  assign o[35800] = i[35800];
  assign o[35799] = i[35799];
  assign o[35798] = i[35798];
  assign o[35797] = i[35797];
  assign o[35796] = i[35796];
  assign o[35795] = i[35795];
  assign o[35794] = i[35794];
  assign o[35793] = i[35793];
  assign o[35792] = i[35792];
  assign o[35791] = i[35791];
  assign o[35790] = i[35790];
  assign o[35789] = i[35789];
  assign o[35788] = i[35788];
  assign o[35787] = i[35787];
  assign o[35786] = i[35786];
  assign o[35785] = i[35785];
  assign o[35784] = i[35784];
  assign o[35783] = i[35783];
  assign o[35782] = i[35782];
  assign o[35781] = i[35781];
  assign o[35780] = i[35780];
  assign o[35779] = i[35779];
  assign o[35778] = i[35778];
  assign o[35777] = i[35777];
  assign o[35776] = i[35776];
  assign o[35775] = i[35775];
  assign o[35774] = i[35774];
  assign o[35773] = i[35773];
  assign o[35772] = i[35772];
  assign o[35771] = i[35771];
  assign o[35770] = i[35770];
  assign o[35769] = i[35769];
  assign o[35768] = i[35768];
  assign o[35767] = i[35767];
  assign o[35766] = i[35766];
  assign o[35765] = i[35765];
  assign o[35764] = i[35764];
  assign o[35763] = i[35763];
  assign o[35762] = i[35762];
  assign o[35761] = i[35761];
  assign o[35760] = i[35760];
  assign o[35759] = i[35759];
  assign o[35758] = i[35758];
  assign o[35757] = i[35757];
  assign o[35756] = i[35756];
  assign o[35755] = i[35755];
  assign o[35754] = i[35754];
  assign o[35753] = i[35753];
  assign o[35752] = i[35752];
  assign o[35751] = i[35751];
  assign o[35750] = i[35750];
  assign o[35749] = i[35749];
  assign o[35748] = i[35748];
  assign o[35747] = i[35747];
  assign o[35746] = i[35746];
  assign o[35745] = i[35745];
  assign o[35744] = i[35744];
  assign o[35743] = i[35743];
  assign o[35742] = i[35742];
  assign o[35741] = i[35741];
  assign o[35740] = i[35740];
  assign o[35739] = i[35739];
  assign o[35738] = i[35738];
  assign o[35737] = i[35737];
  assign o[35736] = i[35736];
  assign o[35735] = i[35735];
  assign o[35734] = i[35734];
  assign o[35733] = i[35733];
  assign o[35732] = i[35732];
  assign o[35731] = i[35731];
  assign o[35730] = i[35730];
  assign o[35729] = i[35729];
  assign o[35728] = i[35728];
  assign o[35727] = i[35727];
  assign o[35726] = i[35726];
  assign o[35725] = i[35725];
  assign o[35724] = i[35724];
  assign o[35723] = i[35723];
  assign o[35722] = i[35722];
  assign o[35721] = i[35721];
  assign o[35720] = i[35720];
  assign o[35719] = i[35719];
  assign o[35718] = i[35718];
  assign o[35717] = i[35717];
  assign o[35716] = i[35716];
  assign o[35715] = i[35715];
  assign o[35714] = i[35714];
  assign o[35713] = i[35713];
  assign o[35712] = i[35712];
  assign o[35711] = i[35711];
  assign o[35710] = i[35710];
  assign o[35709] = i[35709];
  assign o[35708] = i[35708];
  assign o[35707] = i[35707];
  assign o[35706] = i[35706];
  assign o[35705] = i[35705];
  assign o[35704] = i[35704];
  assign o[35703] = i[35703];
  assign o[35702] = i[35702];
  assign o[35701] = i[35701];
  assign o[35700] = i[35700];
  assign o[35699] = i[35699];
  assign o[35698] = i[35698];
  assign o[35697] = i[35697];
  assign o[35696] = i[35696];
  assign o[35695] = i[35695];
  assign o[35694] = i[35694];
  assign o[35693] = i[35693];
  assign o[35692] = i[35692];
  assign o[35691] = i[35691];
  assign o[35690] = i[35690];
  assign o[35689] = i[35689];
  assign o[35688] = i[35688];
  assign o[35687] = i[35687];
  assign o[35686] = i[35686];
  assign o[35685] = i[35685];
  assign o[35684] = i[35684];
  assign o[35683] = i[35683];
  assign o[35682] = i[35682];
  assign o[35681] = i[35681];
  assign o[35680] = i[35680];
  assign o[35679] = i[35679];
  assign o[35678] = i[35678];
  assign o[35677] = i[35677];
  assign o[35676] = i[35676];
  assign o[35675] = i[35675];
  assign o[35674] = i[35674];
  assign o[35673] = i[35673];
  assign o[35672] = i[35672];
  assign o[35671] = i[35671];
  assign o[35670] = i[35670];
  assign o[35669] = i[35669];
  assign o[35668] = i[35668];
  assign o[35667] = i[35667];
  assign o[35666] = i[35666];
  assign o[35665] = i[35665];
  assign o[35664] = i[35664];
  assign o[35663] = i[35663];
  assign o[35662] = i[35662];
  assign o[35661] = i[35661];
  assign o[35660] = i[35660];
  assign o[35659] = i[35659];
  assign o[35658] = i[35658];
  assign o[35657] = i[35657];
  assign o[35656] = i[35656];
  assign o[35655] = i[35655];
  assign o[35654] = i[35654];
  assign o[35653] = i[35653];
  assign o[35652] = i[35652];
  assign o[35651] = i[35651];
  assign o[35650] = i[35650];
  assign o[35649] = i[35649];
  assign o[35648] = i[35648];
  assign o[35647] = i[35647];
  assign o[35646] = i[35646];
  assign o[35645] = i[35645];
  assign o[35644] = i[35644];
  assign o[35643] = i[35643];
  assign o[35642] = i[35642];
  assign o[35641] = i[35641];
  assign o[35640] = i[35640];
  assign o[35639] = i[35639];
  assign o[35638] = i[35638];
  assign o[35637] = i[35637];
  assign o[35636] = i[35636];
  assign o[35635] = i[35635];
  assign o[35634] = i[35634];
  assign o[35633] = i[35633];
  assign o[35632] = i[35632];
  assign o[35631] = i[35631];
  assign o[35630] = i[35630];
  assign o[35629] = i[35629];
  assign o[35628] = i[35628];
  assign o[35627] = i[35627];
  assign o[35626] = i[35626];
  assign o[35625] = i[35625];
  assign o[35624] = i[35624];
  assign o[35623] = i[35623];
  assign o[35622] = i[35622];
  assign o[35621] = i[35621];
  assign o[35620] = i[35620];
  assign o[35619] = i[35619];
  assign o[35618] = i[35618];
  assign o[35617] = i[35617];
  assign o[35616] = i[35616];
  assign o[35615] = i[35615];
  assign o[35614] = i[35614];
  assign o[35613] = i[35613];
  assign o[35612] = i[35612];
  assign o[35611] = i[35611];
  assign o[35610] = i[35610];
  assign o[35609] = i[35609];
  assign o[35608] = i[35608];
  assign o[35607] = i[35607];
  assign o[35606] = i[35606];
  assign o[35605] = i[35605];
  assign o[35604] = i[35604];
  assign o[35603] = i[35603];
  assign o[35602] = i[35602];
  assign o[35601] = i[35601];
  assign o[35600] = i[35600];
  assign o[35599] = i[35599];
  assign o[35598] = i[35598];
  assign o[35597] = i[35597];
  assign o[35596] = i[35596];
  assign o[35595] = i[35595];
  assign o[35594] = i[35594];
  assign o[35593] = i[35593];
  assign o[35592] = i[35592];
  assign o[35591] = i[35591];
  assign o[35590] = i[35590];
  assign o[35589] = i[35589];
  assign o[35588] = i[35588];
  assign o[35587] = i[35587];
  assign o[35586] = i[35586];
  assign o[35585] = i[35585];
  assign o[35584] = i[35584];
  assign o[35583] = i[35583];
  assign o[35582] = i[35582];
  assign o[35581] = i[35581];
  assign o[35580] = i[35580];
  assign o[35579] = i[35579];
  assign o[35578] = i[35578];
  assign o[35577] = i[35577];
  assign o[35576] = i[35576];
  assign o[35575] = i[35575];
  assign o[35574] = i[35574];
  assign o[35573] = i[35573];
  assign o[35572] = i[35572];
  assign o[35571] = i[35571];
  assign o[35570] = i[35570];
  assign o[35569] = i[35569];
  assign o[35568] = i[35568];
  assign o[35567] = i[35567];
  assign o[35566] = i[35566];
  assign o[35565] = i[35565];
  assign o[35564] = i[35564];
  assign o[35563] = i[35563];
  assign o[35562] = i[35562];
  assign o[35561] = i[35561];
  assign o[35560] = i[35560];
  assign o[35559] = i[35559];
  assign o[35558] = i[35558];
  assign o[35557] = i[35557];
  assign o[35556] = i[35556];
  assign o[35555] = i[35555];
  assign o[35554] = i[35554];
  assign o[35553] = i[35553];
  assign o[35552] = i[35552];
  assign o[35551] = i[35551];
  assign o[35550] = i[35550];
  assign o[35549] = i[35549];
  assign o[35548] = i[35548];
  assign o[35547] = i[35547];
  assign o[35546] = i[35546];
  assign o[35545] = i[35545];
  assign o[35544] = i[35544];
  assign o[35543] = i[35543];
  assign o[35542] = i[35542];
  assign o[35541] = i[35541];
  assign o[35540] = i[35540];
  assign o[35539] = i[35539];
  assign o[35538] = i[35538];
  assign o[35537] = i[35537];
  assign o[35536] = i[35536];
  assign o[35535] = i[35535];
  assign o[35534] = i[35534];
  assign o[35533] = i[35533];
  assign o[35532] = i[35532];
  assign o[35531] = i[35531];
  assign o[35530] = i[35530];
  assign o[35529] = i[35529];
  assign o[35528] = i[35528];
  assign o[35527] = i[35527];
  assign o[35526] = i[35526];
  assign o[35525] = i[35525];
  assign o[35524] = i[35524];
  assign o[35523] = i[35523];
  assign o[35522] = i[35522];
  assign o[35521] = i[35521];
  assign o[35520] = i[35520];
  assign o[35519] = i[35519];
  assign o[35518] = i[35518];
  assign o[35517] = i[35517];
  assign o[35516] = i[35516];
  assign o[35515] = i[35515];
  assign o[35514] = i[35514];
  assign o[35513] = i[35513];
  assign o[35512] = i[35512];
  assign o[35511] = i[35511];
  assign o[35510] = i[35510];
  assign o[35509] = i[35509];
  assign o[35508] = i[35508];
  assign o[35507] = i[35507];
  assign o[35506] = i[35506];
  assign o[35505] = i[35505];
  assign o[35504] = i[35504];
  assign o[35503] = i[35503];
  assign o[35502] = i[35502];
  assign o[35501] = i[35501];
  assign o[35500] = i[35500];
  assign o[35499] = i[35499];
  assign o[35498] = i[35498];
  assign o[35497] = i[35497];
  assign o[35496] = i[35496];
  assign o[35495] = i[35495];
  assign o[35494] = i[35494];
  assign o[35493] = i[35493];
  assign o[35492] = i[35492];
  assign o[35491] = i[35491];
  assign o[35490] = i[35490];
  assign o[35489] = i[35489];
  assign o[35488] = i[35488];
  assign o[35487] = i[35487];
  assign o[35486] = i[35486];
  assign o[35485] = i[35485];
  assign o[35484] = i[35484];
  assign o[35483] = i[35483];
  assign o[35482] = i[35482];
  assign o[35481] = i[35481];
  assign o[35480] = i[35480];
  assign o[35479] = i[35479];
  assign o[35478] = i[35478];
  assign o[35477] = i[35477];
  assign o[35476] = i[35476];
  assign o[35475] = i[35475];
  assign o[35474] = i[35474];
  assign o[35473] = i[35473];
  assign o[35472] = i[35472];
  assign o[35471] = i[35471];
  assign o[35470] = i[35470];
  assign o[35469] = i[35469];
  assign o[35468] = i[35468];
  assign o[35467] = i[35467];
  assign o[35466] = i[35466];
  assign o[35465] = i[35465];
  assign o[35464] = i[35464];
  assign o[35463] = i[35463];
  assign o[35462] = i[35462];
  assign o[35461] = i[35461];
  assign o[35460] = i[35460];
  assign o[35459] = i[35459];
  assign o[35458] = i[35458];
  assign o[35457] = i[35457];
  assign o[35456] = i[35456];
  assign o[35455] = i[35455];
  assign o[35454] = i[35454];
  assign o[35453] = i[35453];
  assign o[35452] = i[35452];
  assign o[35451] = i[35451];
  assign o[35450] = i[35450];
  assign o[35449] = i[35449];
  assign o[35448] = i[35448];
  assign o[35447] = i[35447];
  assign o[35446] = i[35446];
  assign o[35445] = i[35445];
  assign o[35444] = i[35444];
  assign o[35443] = i[35443];
  assign o[35442] = i[35442];
  assign o[35441] = i[35441];
  assign o[35440] = i[35440];
  assign o[35439] = i[35439];
  assign o[35438] = i[35438];
  assign o[35437] = i[35437];
  assign o[35436] = i[35436];
  assign o[35435] = i[35435];
  assign o[35434] = i[35434];
  assign o[35433] = i[35433];
  assign o[35432] = i[35432];
  assign o[35431] = i[35431];
  assign o[35430] = i[35430];
  assign o[35429] = i[35429];
  assign o[35428] = i[35428];
  assign o[35427] = i[35427];
  assign o[35426] = i[35426];
  assign o[35425] = i[35425];
  assign o[35424] = i[35424];
  assign o[35423] = i[35423];
  assign o[35422] = i[35422];
  assign o[35421] = i[35421];
  assign o[35420] = i[35420];
  assign o[35419] = i[35419];
  assign o[35418] = i[35418];
  assign o[35417] = i[35417];
  assign o[35416] = i[35416];
  assign o[35415] = i[35415];
  assign o[35414] = i[35414];
  assign o[35413] = i[35413];
  assign o[35412] = i[35412];
  assign o[35411] = i[35411];
  assign o[35410] = i[35410];
  assign o[35409] = i[35409];
  assign o[35408] = i[35408];
  assign o[35407] = i[35407];
  assign o[35406] = i[35406];
  assign o[35405] = i[35405];
  assign o[35404] = i[35404];
  assign o[35403] = i[35403];
  assign o[35402] = i[35402];
  assign o[35401] = i[35401];
  assign o[35400] = i[35400];
  assign o[35399] = i[35399];
  assign o[35398] = i[35398];
  assign o[35397] = i[35397];
  assign o[35396] = i[35396];
  assign o[35395] = i[35395];
  assign o[35394] = i[35394];
  assign o[35393] = i[35393];
  assign o[35392] = i[35392];
  assign o[35391] = i[35391];
  assign o[35390] = i[35390];
  assign o[35389] = i[35389];
  assign o[35388] = i[35388];
  assign o[35387] = i[35387];
  assign o[35386] = i[35386];
  assign o[35385] = i[35385];
  assign o[35384] = i[35384];
  assign o[35383] = i[35383];
  assign o[35382] = i[35382];
  assign o[35381] = i[35381];
  assign o[35380] = i[35380];
  assign o[35379] = i[35379];
  assign o[35378] = i[35378];
  assign o[35377] = i[35377];
  assign o[35376] = i[35376];
  assign o[35375] = i[35375];
  assign o[35374] = i[35374];
  assign o[35373] = i[35373];
  assign o[35372] = i[35372];
  assign o[35371] = i[35371];
  assign o[35370] = i[35370];
  assign o[35369] = i[35369];
  assign o[35368] = i[35368];
  assign o[35367] = i[35367];
  assign o[35366] = i[35366];
  assign o[35365] = i[35365];
  assign o[35364] = i[35364];
  assign o[35363] = i[35363];
  assign o[35362] = i[35362];
  assign o[35361] = i[35361];
  assign o[35360] = i[35360];
  assign o[35359] = i[35359];
  assign o[35358] = i[35358];
  assign o[35357] = i[35357];
  assign o[35356] = i[35356];
  assign o[35355] = i[35355];
  assign o[35354] = i[35354];
  assign o[35353] = i[35353];
  assign o[35352] = i[35352];
  assign o[35351] = i[35351];
  assign o[35350] = i[35350];
  assign o[35349] = i[35349];
  assign o[35348] = i[35348];
  assign o[35347] = i[35347];
  assign o[35346] = i[35346];
  assign o[35345] = i[35345];
  assign o[35344] = i[35344];
  assign o[35343] = i[35343];
  assign o[35342] = i[35342];
  assign o[35341] = i[35341];
  assign o[35340] = i[35340];
  assign o[35339] = i[35339];
  assign o[35338] = i[35338];
  assign o[35337] = i[35337];
  assign o[35336] = i[35336];
  assign o[35335] = i[35335];
  assign o[35334] = i[35334];
  assign o[35333] = i[35333];
  assign o[35332] = i[35332];
  assign o[35331] = i[35331];
  assign o[35330] = i[35330];
  assign o[35329] = i[35329];
  assign o[35328] = i[35328];
  assign o[35327] = i[35327];
  assign o[35326] = i[35326];
  assign o[35325] = i[35325];
  assign o[35324] = i[35324];
  assign o[35323] = i[35323];
  assign o[35322] = i[35322];
  assign o[35321] = i[35321];
  assign o[35320] = i[35320];
  assign o[35319] = i[35319];
  assign o[35318] = i[35318];
  assign o[35317] = i[35317];
  assign o[35316] = i[35316];
  assign o[35315] = i[35315];
  assign o[35314] = i[35314];
  assign o[35313] = i[35313];
  assign o[35312] = i[35312];
  assign o[35311] = i[35311];
  assign o[35310] = i[35310];
  assign o[35309] = i[35309];
  assign o[35308] = i[35308];
  assign o[35307] = i[35307];
  assign o[35306] = i[35306];
  assign o[35305] = i[35305];
  assign o[35304] = i[35304];
  assign o[35303] = i[35303];
  assign o[35302] = i[35302];
  assign o[35301] = i[35301];
  assign o[35300] = i[35300];
  assign o[35299] = i[35299];
  assign o[35298] = i[35298];
  assign o[35297] = i[35297];
  assign o[35296] = i[35296];
  assign o[35295] = i[35295];
  assign o[35294] = i[35294];
  assign o[35293] = i[35293];
  assign o[35292] = i[35292];
  assign o[35291] = i[35291];
  assign o[35290] = i[35290];
  assign o[35289] = i[35289];
  assign o[35288] = i[35288];
  assign o[35287] = i[35287];
  assign o[35286] = i[35286];
  assign o[35285] = i[35285];
  assign o[35284] = i[35284];
  assign o[35283] = i[35283];
  assign o[35282] = i[35282];
  assign o[35281] = i[35281];
  assign o[35280] = i[35280];
  assign o[35279] = i[35279];
  assign o[35278] = i[35278];
  assign o[35277] = i[35277];
  assign o[35276] = i[35276];
  assign o[35275] = i[35275];
  assign o[35274] = i[35274];
  assign o[35273] = i[35273];
  assign o[35272] = i[35272];
  assign o[35271] = i[35271];
  assign o[35270] = i[35270];
  assign o[35269] = i[35269];
  assign o[35268] = i[35268];
  assign o[35267] = i[35267];
  assign o[35266] = i[35266];
  assign o[35265] = i[35265];
  assign o[35264] = i[35264];
  assign o[35263] = i[35263];
  assign o[35262] = i[35262];
  assign o[35261] = i[35261];
  assign o[35260] = i[35260];
  assign o[35259] = i[35259];
  assign o[35258] = i[35258];
  assign o[35257] = i[35257];
  assign o[35256] = i[35256];
  assign o[35255] = i[35255];
  assign o[35254] = i[35254];
  assign o[35253] = i[35253];
  assign o[35252] = i[35252];
  assign o[35251] = i[35251];
  assign o[35250] = i[35250];
  assign o[35249] = i[35249];
  assign o[35248] = i[35248];
  assign o[35247] = i[35247];
  assign o[35246] = i[35246];
  assign o[35245] = i[35245];
  assign o[35244] = i[35244];
  assign o[35243] = i[35243];
  assign o[35242] = i[35242];
  assign o[35241] = i[35241];
  assign o[35240] = i[35240];
  assign o[35239] = i[35239];
  assign o[35238] = i[35238];
  assign o[35237] = i[35237];
  assign o[35236] = i[35236];
  assign o[35235] = i[35235];
  assign o[35234] = i[35234];
  assign o[35233] = i[35233];
  assign o[35232] = i[35232];
  assign o[35231] = i[35231];
  assign o[35230] = i[35230];
  assign o[35229] = i[35229];
  assign o[35228] = i[35228];
  assign o[35227] = i[35227];
  assign o[35226] = i[35226];
  assign o[35225] = i[35225];
  assign o[35224] = i[35224];
  assign o[35223] = i[35223];
  assign o[35222] = i[35222];
  assign o[35221] = i[35221];
  assign o[35220] = i[35220];
  assign o[35219] = i[35219];
  assign o[35218] = i[35218];
  assign o[35217] = i[35217];
  assign o[35216] = i[35216];
  assign o[35215] = i[35215];
  assign o[35214] = i[35214];
  assign o[35213] = i[35213];
  assign o[35212] = i[35212];
  assign o[35211] = i[35211];
  assign o[35210] = i[35210];
  assign o[35209] = i[35209];
  assign o[35208] = i[35208];
  assign o[35207] = i[35207];
  assign o[35206] = i[35206];
  assign o[35205] = i[35205];
  assign o[35204] = i[35204];
  assign o[35203] = i[35203];
  assign o[35202] = i[35202];
  assign o[35201] = i[35201];
  assign o[35200] = i[35200];
  assign o[35199] = i[35199];
  assign o[35198] = i[35198];
  assign o[35197] = i[35197];
  assign o[35196] = i[35196];
  assign o[35195] = i[35195];
  assign o[35194] = i[35194];
  assign o[35193] = i[35193];
  assign o[35192] = i[35192];
  assign o[35191] = i[35191];
  assign o[35190] = i[35190];
  assign o[35189] = i[35189];
  assign o[35188] = i[35188];
  assign o[35187] = i[35187];
  assign o[35186] = i[35186];
  assign o[35185] = i[35185];
  assign o[35184] = i[35184];
  assign o[35183] = i[35183];
  assign o[35182] = i[35182];
  assign o[35181] = i[35181];
  assign o[35180] = i[35180];
  assign o[35179] = i[35179];
  assign o[35178] = i[35178];
  assign o[35177] = i[35177];
  assign o[35176] = i[35176];
  assign o[35175] = i[35175];
  assign o[35174] = i[35174];
  assign o[35173] = i[35173];
  assign o[35172] = i[35172];
  assign o[35171] = i[35171];
  assign o[35170] = i[35170];
  assign o[35169] = i[35169];
  assign o[35168] = i[35168];
  assign o[35167] = i[35167];
  assign o[35166] = i[35166];
  assign o[35165] = i[35165];
  assign o[35164] = i[35164];
  assign o[35163] = i[35163];
  assign o[35162] = i[35162];
  assign o[35161] = i[35161];
  assign o[35160] = i[35160];
  assign o[35159] = i[35159];
  assign o[35158] = i[35158];
  assign o[35157] = i[35157];
  assign o[35156] = i[35156];
  assign o[35155] = i[35155];
  assign o[35154] = i[35154];
  assign o[35153] = i[35153];
  assign o[35152] = i[35152];
  assign o[35151] = i[35151];
  assign o[35150] = i[35150];
  assign o[35149] = i[35149];
  assign o[35148] = i[35148];
  assign o[35147] = i[35147];
  assign o[35146] = i[35146];
  assign o[35145] = i[35145];
  assign o[35144] = i[35144];
  assign o[35143] = i[35143];
  assign o[35142] = i[35142];
  assign o[35141] = i[35141];
  assign o[35140] = i[35140];
  assign o[35139] = i[35139];
  assign o[35138] = i[35138];
  assign o[35137] = i[35137];
  assign o[35136] = i[35136];
  assign o[35135] = i[35135];
  assign o[35134] = i[35134];
  assign o[35133] = i[35133];
  assign o[35132] = i[35132];
  assign o[35131] = i[35131];
  assign o[35130] = i[35130];
  assign o[35129] = i[35129];
  assign o[35128] = i[35128];
  assign o[35127] = i[35127];
  assign o[35126] = i[35126];
  assign o[35125] = i[35125];
  assign o[35124] = i[35124];
  assign o[35123] = i[35123];
  assign o[35122] = i[35122];
  assign o[35121] = i[35121];
  assign o[35120] = i[35120];
  assign o[35119] = i[35119];
  assign o[35118] = i[35118];
  assign o[35117] = i[35117];
  assign o[35116] = i[35116];
  assign o[35115] = i[35115];
  assign o[35114] = i[35114];
  assign o[35113] = i[35113];
  assign o[35112] = i[35112];
  assign o[35111] = i[35111];
  assign o[35110] = i[35110];
  assign o[35109] = i[35109];
  assign o[35108] = i[35108];
  assign o[35107] = i[35107];
  assign o[35106] = i[35106];
  assign o[35105] = i[35105];
  assign o[35104] = i[35104];
  assign o[35103] = i[35103];
  assign o[35102] = i[35102];
  assign o[35101] = i[35101];
  assign o[35100] = i[35100];
  assign o[35099] = i[35099];
  assign o[35098] = i[35098];
  assign o[35097] = i[35097];
  assign o[35096] = i[35096];
  assign o[35095] = i[35095];
  assign o[35094] = i[35094];
  assign o[35093] = i[35093];
  assign o[35092] = i[35092];
  assign o[35091] = i[35091];
  assign o[35090] = i[35090];
  assign o[35089] = i[35089];
  assign o[35088] = i[35088];
  assign o[35087] = i[35087];
  assign o[35086] = i[35086];
  assign o[35085] = i[35085];
  assign o[35084] = i[35084];
  assign o[35083] = i[35083];
  assign o[35082] = i[35082];
  assign o[35081] = i[35081];
  assign o[35080] = i[35080];
  assign o[35079] = i[35079];
  assign o[35078] = i[35078];
  assign o[35077] = i[35077];
  assign o[35076] = i[35076];
  assign o[35075] = i[35075];
  assign o[35074] = i[35074];
  assign o[35073] = i[35073];
  assign o[35072] = i[35072];
  assign o[35071] = i[35071];
  assign o[35070] = i[35070];
  assign o[35069] = i[35069];
  assign o[35068] = i[35068];
  assign o[35067] = i[35067];
  assign o[35066] = i[35066];
  assign o[35065] = i[35065];
  assign o[35064] = i[35064];
  assign o[35063] = i[35063];
  assign o[35062] = i[35062];
  assign o[35061] = i[35061];
  assign o[35060] = i[35060];
  assign o[35059] = i[35059];
  assign o[35058] = i[35058];
  assign o[35057] = i[35057];
  assign o[35056] = i[35056];
  assign o[35055] = i[35055];
  assign o[35054] = i[35054];
  assign o[35053] = i[35053];
  assign o[35052] = i[35052];
  assign o[35051] = i[35051];
  assign o[35050] = i[35050];
  assign o[35049] = i[35049];
  assign o[35048] = i[35048];
  assign o[35047] = i[35047];
  assign o[35046] = i[35046];
  assign o[35045] = i[35045];
  assign o[35044] = i[35044];
  assign o[35043] = i[35043];
  assign o[35042] = i[35042];
  assign o[35041] = i[35041];
  assign o[35040] = i[35040];
  assign o[35039] = i[35039];
  assign o[35038] = i[35038];
  assign o[35037] = i[35037];
  assign o[35036] = i[35036];
  assign o[35035] = i[35035];
  assign o[35034] = i[35034];
  assign o[35033] = i[35033];
  assign o[35032] = i[35032];
  assign o[35031] = i[35031];
  assign o[35030] = i[35030];
  assign o[35029] = i[35029];
  assign o[35028] = i[35028];
  assign o[35027] = i[35027];
  assign o[35026] = i[35026];
  assign o[35025] = i[35025];
  assign o[35024] = i[35024];
  assign o[35023] = i[35023];
  assign o[35022] = i[35022];
  assign o[35021] = i[35021];
  assign o[35020] = i[35020];
  assign o[35019] = i[35019];
  assign o[35018] = i[35018];
  assign o[35017] = i[35017];
  assign o[35016] = i[35016];
  assign o[35015] = i[35015];
  assign o[35014] = i[35014];
  assign o[35013] = i[35013];
  assign o[35012] = i[35012];
  assign o[35011] = i[35011];
  assign o[35010] = i[35010];
  assign o[35009] = i[35009];
  assign o[35008] = i[35008];
  assign o[35007] = i[35007];
  assign o[35006] = i[35006];
  assign o[35005] = i[35005];
  assign o[35004] = i[35004];
  assign o[35003] = i[35003];
  assign o[35002] = i[35002];
  assign o[35001] = i[35001];
  assign o[35000] = i[35000];
  assign o[34999] = i[34999];
  assign o[34998] = i[34998];
  assign o[34997] = i[34997];
  assign o[34996] = i[34996];
  assign o[34995] = i[34995];
  assign o[34994] = i[34994];
  assign o[34993] = i[34993];
  assign o[34992] = i[34992];
  assign o[34991] = i[34991];
  assign o[34990] = i[34990];
  assign o[34989] = i[34989];
  assign o[34988] = i[34988];
  assign o[34987] = i[34987];
  assign o[34986] = i[34986];
  assign o[34985] = i[34985];
  assign o[34984] = i[34984];
  assign o[34983] = i[34983];
  assign o[34982] = i[34982];
  assign o[34981] = i[34981];
  assign o[34980] = i[34980];
  assign o[34979] = i[34979];
  assign o[34978] = i[34978];
  assign o[34977] = i[34977];
  assign o[34976] = i[34976];
  assign o[34975] = i[34975];
  assign o[34974] = i[34974];
  assign o[34973] = i[34973];
  assign o[34972] = i[34972];
  assign o[34971] = i[34971];
  assign o[34970] = i[34970];
  assign o[34969] = i[34969];
  assign o[34968] = i[34968];
  assign o[34967] = i[34967];
  assign o[34966] = i[34966];
  assign o[34965] = i[34965];
  assign o[34964] = i[34964];
  assign o[34963] = i[34963];
  assign o[34962] = i[34962];
  assign o[34961] = i[34961];
  assign o[34960] = i[34960];
  assign o[34959] = i[34959];
  assign o[34958] = i[34958];
  assign o[34957] = i[34957];
  assign o[34956] = i[34956];
  assign o[34955] = i[34955];
  assign o[34954] = i[34954];
  assign o[34953] = i[34953];
  assign o[34952] = i[34952];
  assign o[34951] = i[34951];
  assign o[34950] = i[34950];
  assign o[34949] = i[34949];
  assign o[34948] = i[34948];
  assign o[34947] = i[34947];
  assign o[34946] = i[34946];
  assign o[34945] = i[34945];
  assign o[34944] = i[34944];
  assign o[34943] = i[34943];
  assign o[34942] = i[34942];
  assign o[34941] = i[34941];
  assign o[34940] = i[34940];
  assign o[34939] = i[34939];
  assign o[34938] = i[34938];
  assign o[34937] = i[34937];
  assign o[34936] = i[34936];
  assign o[34935] = i[34935];
  assign o[34934] = i[34934];
  assign o[34933] = i[34933];
  assign o[34932] = i[34932];
  assign o[34931] = i[34931];
  assign o[34930] = i[34930];
  assign o[34929] = i[34929];
  assign o[34928] = i[34928];
  assign o[34927] = i[34927];
  assign o[34926] = i[34926];
  assign o[34925] = i[34925];
  assign o[34924] = i[34924];
  assign o[34923] = i[34923];
  assign o[34922] = i[34922];
  assign o[34921] = i[34921];
  assign o[34920] = i[34920];
  assign o[34919] = i[34919];
  assign o[34918] = i[34918];
  assign o[34917] = i[34917];
  assign o[34916] = i[34916];
  assign o[34915] = i[34915];
  assign o[34914] = i[34914];
  assign o[34913] = i[34913];
  assign o[34912] = i[34912];
  assign o[34911] = i[34911];
  assign o[34910] = i[34910];
  assign o[34909] = i[34909];
  assign o[34908] = i[34908];
  assign o[34907] = i[34907];
  assign o[34906] = i[34906];
  assign o[34905] = i[34905];
  assign o[34904] = i[34904];
  assign o[34903] = i[34903];
  assign o[34902] = i[34902];
  assign o[34901] = i[34901];
  assign o[34900] = i[34900];
  assign o[34899] = i[34899];
  assign o[34898] = i[34898];
  assign o[34897] = i[34897];
  assign o[34896] = i[34896];
  assign o[34895] = i[34895];
  assign o[34894] = i[34894];
  assign o[34893] = i[34893];
  assign o[34892] = i[34892];
  assign o[34891] = i[34891];
  assign o[34890] = i[34890];
  assign o[34889] = i[34889];
  assign o[34888] = i[34888];
  assign o[34887] = i[34887];
  assign o[34886] = i[34886];
  assign o[34885] = i[34885];
  assign o[34884] = i[34884];
  assign o[34883] = i[34883];
  assign o[34882] = i[34882];
  assign o[34881] = i[34881];
  assign o[34880] = i[34880];
  assign o[34879] = i[34879];
  assign o[34878] = i[34878];
  assign o[34877] = i[34877];
  assign o[34876] = i[34876];
  assign o[34875] = i[34875];
  assign o[34874] = i[34874];
  assign o[34873] = i[34873];
  assign o[34872] = i[34872];
  assign o[34871] = i[34871];
  assign o[34870] = i[34870];
  assign o[34869] = i[34869];
  assign o[34868] = i[34868];
  assign o[34867] = i[34867];
  assign o[34866] = i[34866];
  assign o[34865] = i[34865];
  assign o[34864] = i[34864];
  assign o[34863] = i[34863];
  assign o[34862] = i[34862];
  assign o[34861] = i[34861];
  assign o[34860] = i[34860];
  assign o[34859] = i[34859];
  assign o[34858] = i[34858];
  assign o[34857] = i[34857];
  assign o[34856] = i[34856];
  assign o[34855] = i[34855];
  assign o[34854] = i[34854];
  assign o[34853] = i[34853];
  assign o[34852] = i[34852];
  assign o[34851] = i[34851];
  assign o[34850] = i[34850];
  assign o[34849] = i[34849];
  assign o[34848] = i[34848];
  assign o[34847] = i[34847];
  assign o[34846] = i[34846];
  assign o[34845] = i[34845];
  assign o[34844] = i[34844];
  assign o[34843] = i[34843];
  assign o[34842] = i[34842];
  assign o[34841] = i[34841];
  assign o[34840] = i[34840];
  assign o[34839] = i[34839];
  assign o[34838] = i[34838];
  assign o[34837] = i[34837];
  assign o[34836] = i[34836];
  assign o[34835] = i[34835];
  assign o[34834] = i[34834];
  assign o[34833] = i[34833];
  assign o[34832] = i[34832];
  assign o[34831] = i[34831];
  assign o[34830] = i[34830];
  assign o[34829] = i[34829];
  assign o[34828] = i[34828];
  assign o[34827] = i[34827];
  assign o[34826] = i[34826];
  assign o[34825] = i[34825];
  assign o[34824] = i[34824];
  assign o[34823] = i[34823];
  assign o[34822] = i[34822];
  assign o[34821] = i[34821];
  assign o[34820] = i[34820];
  assign o[34819] = i[34819];
  assign o[34818] = i[34818];
  assign o[34817] = i[34817];
  assign o[34816] = i[34816];
  assign o[34815] = i[34815];
  assign o[34814] = i[34814];
  assign o[34813] = i[34813];
  assign o[34812] = i[34812];
  assign o[34811] = i[34811];
  assign o[34810] = i[34810];
  assign o[34809] = i[34809];
  assign o[34808] = i[34808];
  assign o[34807] = i[34807];
  assign o[34806] = i[34806];
  assign o[34805] = i[34805];
  assign o[34804] = i[34804];
  assign o[34803] = i[34803];
  assign o[34802] = i[34802];
  assign o[34801] = i[34801];
  assign o[34800] = i[34800];
  assign o[34799] = i[34799];
  assign o[34798] = i[34798];
  assign o[34797] = i[34797];
  assign o[34796] = i[34796];
  assign o[34795] = i[34795];
  assign o[34794] = i[34794];
  assign o[34793] = i[34793];
  assign o[34792] = i[34792];
  assign o[34791] = i[34791];
  assign o[34790] = i[34790];
  assign o[34789] = i[34789];
  assign o[34788] = i[34788];
  assign o[34787] = i[34787];
  assign o[34786] = i[34786];
  assign o[34785] = i[34785];
  assign o[34784] = i[34784];
  assign o[34783] = i[34783];
  assign o[34782] = i[34782];
  assign o[34781] = i[34781];
  assign o[34780] = i[34780];
  assign o[34779] = i[34779];
  assign o[34778] = i[34778];
  assign o[34777] = i[34777];
  assign o[34776] = i[34776];
  assign o[34775] = i[34775];
  assign o[34774] = i[34774];
  assign o[34773] = i[34773];
  assign o[34772] = i[34772];
  assign o[34771] = i[34771];
  assign o[34770] = i[34770];
  assign o[34769] = i[34769];
  assign o[34768] = i[34768];
  assign o[34767] = i[34767];
  assign o[34766] = i[34766];
  assign o[34765] = i[34765];
  assign o[34764] = i[34764];
  assign o[34763] = i[34763];
  assign o[34762] = i[34762];
  assign o[34761] = i[34761];
  assign o[34760] = i[34760];
  assign o[34759] = i[34759];
  assign o[34758] = i[34758];
  assign o[34757] = i[34757];
  assign o[34756] = i[34756];
  assign o[34755] = i[34755];
  assign o[34754] = i[34754];
  assign o[34753] = i[34753];
  assign o[34752] = i[34752];
  assign o[34751] = i[34751];
  assign o[34750] = i[34750];
  assign o[34749] = i[34749];
  assign o[34748] = i[34748];
  assign o[34747] = i[34747];
  assign o[34746] = i[34746];
  assign o[34745] = i[34745];
  assign o[34744] = i[34744];
  assign o[34743] = i[34743];
  assign o[34742] = i[34742];
  assign o[34741] = i[34741];
  assign o[34740] = i[34740];
  assign o[34739] = i[34739];
  assign o[34738] = i[34738];
  assign o[34737] = i[34737];
  assign o[34736] = i[34736];
  assign o[34735] = i[34735];
  assign o[34734] = i[34734];
  assign o[34733] = i[34733];
  assign o[34732] = i[34732];
  assign o[34731] = i[34731];
  assign o[34730] = i[34730];
  assign o[34729] = i[34729];
  assign o[34728] = i[34728];
  assign o[34727] = i[34727];
  assign o[34726] = i[34726];
  assign o[34725] = i[34725];
  assign o[34724] = i[34724];
  assign o[34723] = i[34723];
  assign o[34722] = i[34722];
  assign o[34721] = i[34721];
  assign o[34720] = i[34720];
  assign o[34719] = i[34719];
  assign o[34718] = i[34718];
  assign o[34717] = i[34717];
  assign o[34716] = i[34716];
  assign o[34715] = i[34715];
  assign o[34714] = i[34714];
  assign o[34713] = i[34713];
  assign o[34712] = i[34712];
  assign o[34711] = i[34711];
  assign o[34710] = i[34710];
  assign o[34709] = i[34709];
  assign o[34708] = i[34708];
  assign o[34707] = i[34707];
  assign o[34706] = i[34706];
  assign o[34705] = i[34705];
  assign o[34704] = i[34704];
  assign o[34703] = i[34703];
  assign o[34702] = i[34702];
  assign o[34701] = i[34701];
  assign o[34700] = i[34700];
  assign o[34699] = i[34699];
  assign o[34698] = i[34698];
  assign o[34697] = i[34697];
  assign o[34696] = i[34696];
  assign o[34695] = i[34695];
  assign o[34694] = i[34694];
  assign o[34693] = i[34693];
  assign o[34692] = i[34692];
  assign o[34691] = i[34691];
  assign o[34690] = i[34690];
  assign o[34689] = i[34689];
  assign o[34688] = i[34688];
  assign o[34687] = i[34687];
  assign o[34686] = i[34686];
  assign o[34685] = i[34685];
  assign o[34684] = i[34684];
  assign o[34683] = i[34683];
  assign o[34682] = i[34682];
  assign o[34681] = i[34681];
  assign o[34680] = i[34680];
  assign o[34679] = i[34679];
  assign o[34678] = i[34678];
  assign o[34677] = i[34677];
  assign o[34676] = i[34676];
  assign o[34675] = i[34675];
  assign o[34674] = i[34674];
  assign o[34673] = i[34673];
  assign o[34672] = i[34672];
  assign o[34671] = i[34671];
  assign o[34670] = i[34670];
  assign o[34669] = i[34669];
  assign o[34668] = i[34668];
  assign o[34667] = i[34667];
  assign o[34666] = i[34666];
  assign o[34665] = i[34665];
  assign o[34664] = i[34664];
  assign o[34663] = i[34663];
  assign o[34662] = i[34662];
  assign o[34661] = i[34661];
  assign o[34660] = i[34660];
  assign o[34659] = i[34659];
  assign o[34658] = i[34658];
  assign o[34657] = i[34657];
  assign o[34656] = i[34656];
  assign o[34655] = i[34655];
  assign o[34654] = i[34654];
  assign o[34653] = i[34653];
  assign o[34652] = i[34652];
  assign o[34651] = i[34651];
  assign o[34650] = i[34650];
  assign o[34649] = i[34649];
  assign o[34648] = i[34648];
  assign o[34647] = i[34647];
  assign o[34646] = i[34646];
  assign o[34645] = i[34645];
  assign o[34644] = i[34644];
  assign o[34643] = i[34643];
  assign o[34642] = i[34642];
  assign o[34641] = i[34641];
  assign o[34640] = i[34640];
  assign o[34639] = i[34639];
  assign o[34638] = i[34638];
  assign o[34637] = i[34637];
  assign o[34636] = i[34636];
  assign o[34635] = i[34635];
  assign o[34634] = i[34634];
  assign o[34633] = i[34633];
  assign o[34632] = i[34632];
  assign o[34631] = i[34631];
  assign o[34630] = i[34630];
  assign o[34629] = i[34629];
  assign o[34628] = i[34628];
  assign o[34627] = i[34627];
  assign o[34626] = i[34626];
  assign o[34625] = i[34625];
  assign o[34624] = i[34624];
  assign o[34623] = i[34623];
  assign o[34622] = i[34622];
  assign o[34621] = i[34621];
  assign o[34620] = i[34620];
  assign o[34619] = i[34619];
  assign o[34618] = i[34618];
  assign o[34617] = i[34617];
  assign o[34616] = i[34616];
  assign o[34615] = i[34615];
  assign o[34614] = i[34614];
  assign o[34613] = i[34613];
  assign o[34612] = i[34612];
  assign o[34611] = i[34611];
  assign o[34610] = i[34610];
  assign o[34609] = i[34609];
  assign o[34608] = i[34608];
  assign o[34607] = i[34607];
  assign o[34606] = i[34606];
  assign o[34605] = i[34605];
  assign o[34604] = i[34604];
  assign o[34603] = i[34603];
  assign o[34602] = i[34602];
  assign o[34601] = i[34601];
  assign o[34600] = i[34600];
  assign o[34599] = i[34599];
  assign o[34598] = i[34598];
  assign o[34597] = i[34597];
  assign o[34596] = i[34596];
  assign o[34595] = i[34595];
  assign o[34594] = i[34594];
  assign o[34593] = i[34593];
  assign o[34592] = i[34592];
  assign o[34591] = i[34591];
  assign o[34590] = i[34590];
  assign o[34589] = i[34589];
  assign o[34588] = i[34588];
  assign o[34587] = i[34587];
  assign o[34586] = i[34586];
  assign o[34585] = i[34585];
  assign o[34584] = i[34584];
  assign o[34583] = i[34583];
  assign o[34582] = i[34582];
  assign o[34581] = i[34581];
  assign o[34580] = i[34580];
  assign o[34579] = i[34579];
  assign o[34578] = i[34578];
  assign o[34577] = i[34577];
  assign o[34576] = i[34576];
  assign o[34575] = i[34575];
  assign o[34574] = i[34574];
  assign o[34573] = i[34573];
  assign o[34572] = i[34572];
  assign o[34571] = i[34571];
  assign o[34570] = i[34570];
  assign o[34569] = i[34569];
  assign o[34568] = i[34568];
  assign o[34567] = i[34567];
  assign o[34566] = i[34566];
  assign o[34565] = i[34565];
  assign o[34564] = i[34564];
  assign o[34563] = i[34563];
  assign o[34562] = i[34562];
  assign o[34561] = i[34561];
  assign o[34560] = i[34560];
  assign o[34559] = i[34559];
  assign o[34558] = i[34558];
  assign o[34557] = i[34557];
  assign o[34556] = i[34556];
  assign o[34555] = i[34555];
  assign o[34554] = i[34554];
  assign o[34553] = i[34553];
  assign o[34552] = i[34552];
  assign o[34551] = i[34551];
  assign o[34550] = i[34550];
  assign o[34549] = i[34549];
  assign o[34548] = i[34548];
  assign o[34547] = i[34547];
  assign o[34546] = i[34546];
  assign o[34545] = i[34545];
  assign o[34544] = i[34544];
  assign o[34543] = i[34543];
  assign o[34542] = i[34542];
  assign o[34541] = i[34541];
  assign o[34540] = i[34540];
  assign o[34539] = i[34539];
  assign o[34538] = i[34538];
  assign o[34537] = i[34537];
  assign o[34536] = i[34536];
  assign o[34535] = i[34535];
  assign o[34534] = i[34534];
  assign o[34533] = i[34533];
  assign o[34532] = i[34532];
  assign o[34531] = i[34531];
  assign o[34530] = i[34530];
  assign o[34529] = i[34529];
  assign o[34528] = i[34528];
  assign o[34527] = i[34527];
  assign o[34526] = i[34526];
  assign o[34525] = i[34525];
  assign o[34524] = i[34524];
  assign o[34523] = i[34523];
  assign o[34522] = i[34522];
  assign o[34521] = i[34521];
  assign o[34520] = i[34520];
  assign o[34519] = i[34519];
  assign o[34518] = i[34518];
  assign o[34517] = i[34517];
  assign o[34516] = i[34516];
  assign o[34515] = i[34515];
  assign o[34514] = i[34514];
  assign o[34513] = i[34513];
  assign o[34512] = i[34512];
  assign o[34511] = i[34511];
  assign o[34510] = i[34510];
  assign o[34509] = i[34509];
  assign o[34508] = i[34508];
  assign o[34507] = i[34507];
  assign o[34506] = i[34506];
  assign o[34505] = i[34505];
  assign o[34504] = i[34504];
  assign o[34503] = i[34503];
  assign o[34502] = i[34502];
  assign o[34501] = i[34501];
  assign o[34500] = i[34500];
  assign o[34499] = i[34499];
  assign o[34498] = i[34498];
  assign o[34497] = i[34497];
  assign o[34496] = i[34496];
  assign o[34495] = i[34495];
  assign o[34494] = i[34494];
  assign o[34493] = i[34493];
  assign o[34492] = i[34492];
  assign o[34491] = i[34491];
  assign o[34490] = i[34490];
  assign o[34489] = i[34489];
  assign o[34488] = i[34488];
  assign o[34487] = i[34487];
  assign o[34486] = i[34486];
  assign o[34485] = i[34485];
  assign o[34484] = i[34484];
  assign o[34483] = i[34483];
  assign o[34482] = i[34482];
  assign o[34481] = i[34481];
  assign o[34480] = i[34480];
  assign o[34479] = i[34479];
  assign o[34478] = i[34478];
  assign o[34477] = i[34477];
  assign o[34476] = i[34476];
  assign o[34475] = i[34475];
  assign o[34474] = i[34474];
  assign o[34473] = i[34473];
  assign o[34472] = i[34472];
  assign o[34471] = i[34471];
  assign o[34470] = i[34470];
  assign o[34469] = i[34469];
  assign o[34468] = i[34468];
  assign o[34467] = i[34467];
  assign o[34466] = i[34466];
  assign o[34465] = i[34465];
  assign o[34464] = i[34464];
  assign o[34463] = i[34463];
  assign o[34462] = i[34462];
  assign o[34461] = i[34461];
  assign o[34460] = i[34460];
  assign o[34459] = i[34459];
  assign o[34458] = i[34458];
  assign o[34457] = i[34457];
  assign o[34456] = i[34456];
  assign o[34455] = i[34455];
  assign o[34454] = i[34454];
  assign o[34453] = i[34453];
  assign o[34452] = i[34452];
  assign o[34451] = i[34451];
  assign o[34450] = i[34450];
  assign o[34449] = i[34449];
  assign o[34448] = i[34448];
  assign o[34447] = i[34447];
  assign o[34446] = i[34446];
  assign o[34445] = i[34445];
  assign o[34444] = i[34444];
  assign o[34443] = i[34443];
  assign o[34442] = i[34442];
  assign o[34441] = i[34441];
  assign o[34440] = i[34440];
  assign o[34439] = i[34439];
  assign o[34438] = i[34438];
  assign o[34437] = i[34437];
  assign o[34436] = i[34436];
  assign o[34435] = i[34435];
  assign o[34434] = i[34434];
  assign o[34433] = i[34433];
  assign o[34432] = i[34432];
  assign o[34431] = i[34431];
  assign o[34430] = i[34430];
  assign o[34429] = i[34429];
  assign o[34428] = i[34428];
  assign o[34427] = i[34427];
  assign o[34426] = i[34426];
  assign o[34425] = i[34425];
  assign o[34424] = i[34424];
  assign o[34423] = i[34423];
  assign o[34422] = i[34422];
  assign o[34421] = i[34421];
  assign o[34420] = i[34420];
  assign o[34419] = i[34419];
  assign o[34418] = i[34418];
  assign o[34417] = i[34417];
  assign o[34416] = i[34416];
  assign o[34415] = i[34415];
  assign o[34414] = i[34414];
  assign o[34413] = i[34413];
  assign o[34412] = i[34412];
  assign o[34411] = i[34411];
  assign o[34410] = i[34410];
  assign o[34409] = i[34409];
  assign o[34408] = i[34408];
  assign o[34407] = i[34407];
  assign o[34406] = i[34406];
  assign o[34405] = i[34405];
  assign o[34404] = i[34404];
  assign o[34403] = i[34403];
  assign o[34402] = i[34402];
  assign o[34401] = i[34401];
  assign o[34400] = i[34400];
  assign o[34399] = i[34399];
  assign o[34398] = i[34398];
  assign o[34397] = i[34397];
  assign o[34396] = i[34396];
  assign o[34395] = i[34395];
  assign o[34394] = i[34394];
  assign o[34393] = i[34393];
  assign o[34392] = i[34392];
  assign o[34391] = i[34391];
  assign o[34390] = i[34390];
  assign o[34389] = i[34389];
  assign o[34388] = i[34388];
  assign o[34387] = i[34387];
  assign o[34386] = i[34386];
  assign o[34385] = i[34385];
  assign o[34384] = i[34384];
  assign o[34383] = i[34383];
  assign o[34382] = i[34382];
  assign o[34381] = i[34381];
  assign o[34380] = i[34380];
  assign o[34379] = i[34379];
  assign o[34378] = i[34378];
  assign o[34377] = i[34377];
  assign o[34376] = i[34376];
  assign o[34375] = i[34375];
  assign o[34374] = i[34374];
  assign o[34373] = i[34373];
  assign o[34372] = i[34372];
  assign o[34371] = i[34371];
  assign o[34370] = i[34370];
  assign o[34369] = i[34369];
  assign o[34368] = i[34368];
  assign o[34367] = i[34367];
  assign o[34366] = i[34366];
  assign o[34365] = i[34365];
  assign o[34364] = i[34364];
  assign o[34363] = i[34363];
  assign o[34362] = i[34362];
  assign o[34361] = i[34361];
  assign o[34360] = i[34360];
  assign o[34359] = i[34359];
  assign o[34358] = i[34358];
  assign o[34357] = i[34357];
  assign o[34356] = i[34356];
  assign o[34355] = i[34355];
  assign o[34354] = i[34354];
  assign o[34353] = i[34353];
  assign o[34352] = i[34352];
  assign o[34351] = i[34351];
  assign o[34350] = i[34350];
  assign o[34349] = i[34349];
  assign o[34348] = i[34348];
  assign o[34347] = i[34347];
  assign o[34346] = i[34346];
  assign o[34345] = i[34345];
  assign o[34344] = i[34344];
  assign o[34343] = i[34343];
  assign o[34342] = i[34342];
  assign o[34341] = i[34341];
  assign o[34340] = i[34340];
  assign o[34339] = i[34339];
  assign o[34338] = i[34338];
  assign o[34337] = i[34337];
  assign o[34336] = i[34336];
  assign o[34335] = i[34335];
  assign o[34334] = i[34334];
  assign o[34333] = i[34333];
  assign o[34332] = i[34332];
  assign o[34331] = i[34331];
  assign o[34330] = i[34330];
  assign o[34329] = i[34329];
  assign o[34328] = i[34328];
  assign o[34327] = i[34327];
  assign o[34326] = i[34326];
  assign o[34325] = i[34325];
  assign o[34324] = i[34324];
  assign o[34323] = i[34323];
  assign o[34322] = i[34322];
  assign o[34321] = i[34321];
  assign o[34320] = i[34320];
  assign o[34319] = i[34319];
  assign o[34318] = i[34318];
  assign o[34317] = i[34317];
  assign o[34316] = i[34316];
  assign o[34315] = i[34315];
  assign o[34314] = i[34314];
  assign o[34313] = i[34313];
  assign o[34312] = i[34312];
  assign o[34311] = i[34311];
  assign o[34310] = i[34310];
  assign o[34309] = i[34309];
  assign o[34308] = i[34308];
  assign o[34307] = i[34307];
  assign o[34306] = i[34306];
  assign o[34305] = i[34305];
  assign o[34304] = i[34304];
  assign o[34303] = i[34303];
  assign o[34302] = i[34302];
  assign o[34301] = i[34301];
  assign o[34300] = i[34300];
  assign o[34299] = i[34299];
  assign o[34298] = i[34298];
  assign o[34297] = i[34297];
  assign o[34296] = i[34296];
  assign o[34295] = i[34295];
  assign o[34294] = i[34294];
  assign o[34293] = i[34293];
  assign o[34292] = i[34292];
  assign o[34291] = i[34291];
  assign o[34290] = i[34290];
  assign o[34289] = i[34289];
  assign o[34288] = i[34288];
  assign o[34287] = i[34287];
  assign o[34286] = i[34286];
  assign o[34285] = i[34285];
  assign o[34284] = i[34284];
  assign o[34283] = i[34283];
  assign o[34282] = i[34282];
  assign o[34281] = i[34281];
  assign o[34280] = i[34280];
  assign o[34279] = i[34279];
  assign o[34278] = i[34278];
  assign o[34277] = i[34277];
  assign o[34276] = i[34276];
  assign o[34275] = i[34275];
  assign o[34274] = i[34274];
  assign o[34273] = i[34273];
  assign o[34272] = i[34272];
  assign o[34271] = i[34271];
  assign o[34270] = i[34270];
  assign o[34269] = i[34269];
  assign o[34268] = i[34268];
  assign o[34267] = i[34267];
  assign o[34266] = i[34266];
  assign o[34265] = i[34265];
  assign o[34264] = i[34264];
  assign o[34263] = i[34263];
  assign o[34262] = i[34262];
  assign o[34261] = i[34261];
  assign o[34260] = i[34260];
  assign o[34259] = i[34259];
  assign o[34258] = i[34258];
  assign o[34257] = i[34257];
  assign o[34256] = i[34256];
  assign o[34255] = i[34255];
  assign o[34254] = i[34254];
  assign o[34253] = i[34253];
  assign o[34252] = i[34252];
  assign o[34251] = i[34251];
  assign o[34250] = i[34250];
  assign o[34249] = i[34249];
  assign o[34248] = i[34248];
  assign o[34247] = i[34247];
  assign o[34246] = i[34246];
  assign o[34245] = i[34245];
  assign o[34244] = i[34244];
  assign o[34243] = i[34243];
  assign o[34242] = i[34242];
  assign o[34241] = i[34241];
  assign o[34240] = i[34240];
  assign o[34239] = i[34239];
  assign o[34238] = i[34238];
  assign o[34237] = i[34237];
  assign o[34236] = i[34236];
  assign o[34235] = i[34235];
  assign o[34234] = i[34234];
  assign o[34233] = i[34233];
  assign o[34232] = i[34232];
  assign o[34231] = i[34231];
  assign o[34230] = i[34230];
  assign o[34229] = i[34229];
  assign o[34228] = i[34228];
  assign o[34227] = i[34227];
  assign o[34226] = i[34226];
  assign o[34225] = i[34225];
  assign o[34224] = i[34224];
  assign o[34223] = i[34223];
  assign o[34222] = i[34222];
  assign o[34221] = i[34221];
  assign o[34220] = i[34220];
  assign o[34219] = i[34219];
  assign o[34218] = i[34218];
  assign o[34217] = i[34217];
  assign o[34216] = i[34216];
  assign o[34215] = i[34215];
  assign o[34214] = i[34214];
  assign o[34213] = i[34213];
  assign o[34212] = i[34212];
  assign o[34211] = i[34211];
  assign o[34210] = i[34210];
  assign o[34209] = i[34209];
  assign o[34208] = i[34208];
  assign o[34207] = i[34207];
  assign o[34206] = i[34206];
  assign o[34205] = i[34205];
  assign o[34204] = i[34204];
  assign o[34203] = i[34203];
  assign o[34202] = i[34202];
  assign o[34201] = i[34201];
  assign o[34200] = i[34200];
  assign o[34199] = i[34199];
  assign o[34198] = i[34198];
  assign o[34197] = i[34197];
  assign o[34196] = i[34196];
  assign o[34195] = i[34195];
  assign o[34194] = i[34194];
  assign o[34193] = i[34193];
  assign o[34192] = i[34192];
  assign o[34191] = i[34191];
  assign o[34190] = i[34190];
  assign o[34189] = i[34189];
  assign o[34188] = i[34188];
  assign o[34187] = i[34187];
  assign o[34186] = i[34186];
  assign o[34185] = i[34185];
  assign o[34184] = i[34184];
  assign o[34183] = i[34183];
  assign o[34182] = i[34182];
  assign o[34181] = i[34181];
  assign o[34180] = i[34180];
  assign o[34179] = i[34179];
  assign o[34178] = i[34178];
  assign o[34177] = i[34177];
  assign o[34176] = i[34176];
  assign o[34175] = i[34175];
  assign o[34174] = i[34174];
  assign o[34173] = i[34173];
  assign o[34172] = i[34172];
  assign o[34171] = i[34171];
  assign o[34170] = i[34170];
  assign o[34169] = i[34169];
  assign o[34168] = i[34168];
  assign o[34167] = i[34167];
  assign o[34166] = i[34166];
  assign o[34165] = i[34165];
  assign o[34164] = i[34164];
  assign o[34163] = i[34163];
  assign o[34162] = i[34162];
  assign o[34161] = i[34161];
  assign o[34160] = i[34160];
  assign o[34159] = i[34159];
  assign o[34158] = i[34158];
  assign o[34157] = i[34157];
  assign o[34156] = i[34156];
  assign o[34155] = i[34155];
  assign o[34154] = i[34154];
  assign o[34153] = i[34153];
  assign o[34152] = i[34152];
  assign o[34151] = i[34151];
  assign o[34150] = i[34150];
  assign o[34149] = i[34149];
  assign o[34148] = i[34148];
  assign o[34147] = i[34147];
  assign o[34146] = i[34146];
  assign o[34145] = i[34145];
  assign o[34144] = i[34144];
  assign o[34143] = i[34143];
  assign o[34142] = i[34142];
  assign o[34141] = i[34141];
  assign o[34140] = i[34140];
  assign o[34139] = i[34139];
  assign o[34138] = i[34138];
  assign o[34137] = i[34137];
  assign o[34136] = i[34136];
  assign o[34135] = i[34135];
  assign o[34134] = i[34134];
  assign o[34133] = i[34133];
  assign o[34132] = i[34132];
  assign o[34131] = i[34131];
  assign o[34130] = i[34130];
  assign o[34129] = i[34129];
  assign o[34128] = i[34128];
  assign o[34127] = i[34127];
  assign o[34126] = i[34126];
  assign o[34125] = i[34125];
  assign o[34124] = i[34124];
  assign o[34123] = i[34123];
  assign o[34122] = i[34122];
  assign o[34121] = i[34121];
  assign o[34120] = i[34120];
  assign o[34119] = i[34119];
  assign o[34118] = i[34118];
  assign o[34117] = i[34117];
  assign o[34116] = i[34116];
  assign o[34115] = i[34115];
  assign o[34114] = i[34114];
  assign o[34113] = i[34113];
  assign o[34112] = i[34112];
  assign o[34111] = i[34111];
  assign o[34110] = i[34110];
  assign o[34109] = i[34109];
  assign o[34108] = i[34108];
  assign o[34107] = i[34107];
  assign o[34106] = i[34106];
  assign o[34105] = i[34105];
  assign o[34104] = i[34104];
  assign o[34103] = i[34103];
  assign o[34102] = i[34102];
  assign o[34101] = i[34101];
  assign o[34100] = i[34100];
  assign o[34099] = i[34099];
  assign o[34098] = i[34098];
  assign o[34097] = i[34097];
  assign o[34096] = i[34096];
  assign o[34095] = i[34095];
  assign o[34094] = i[34094];
  assign o[34093] = i[34093];
  assign o[34092] = i[34092];
  assign o[34091] = i[34091];
  assign o[34090] = i[34090];
  assign o[34089] = i[34089];
  assign o[34088] = i[34088];
  assign o[34087] = i[34087];
  assign o[34086] = i[34086];
  assign o[34085] = i[34085];
  assign o[34084] = i[34084];
  assign o[34083] = i[34083];
  assign o[34082] = i[34082];
  assign o[34081] = i[34081];
  assign o[34080] = i[34080];
  assign o[34079] = i[34079];
  assign o[34078] = i[34078];
  assign o[34077] = i[34077];
  assign o[34076] = i[34076];
  assign o[34075] = i[34075];
  assign o[34074] = i[34074];
  assign o[34073] = i[34073];
  assign o[34072] = i[34072];
  assign o[34071] = i[34071];
  assign o[34070] = i[34070];
  assign o[34069] = i[34069];
  assign o[34068] = i[34068];
  assign o[34067] = i[34067];
  assign o[34066] = i[34066];
  assign o[34065] = i[34065];
  assign o[34064] = i[34064];
  assign o[34063] = i[34063];
  assign o[34062] = i[34062];
  assign o[34061] = i[34061];
  assign o[34060] = i[34060];
  assign o[34059] = i[34059];
  assign o[34058] = i[34058];
  assign o[34057] = i[34057];
  assign o[34056] = i[34056];
  assign o[34055] = i[34055];
  assign o[34054] = i[34054];
  assign o[34053] = i[34053];
  assign o[34052] = i[34052];
  assign o[34051] = i[34051];
  assign o[34050] = i[34050];
  assign o[34049] = i[34049];
  assign o[34048] = i[34048];
  assign o[34047] = i[34047];
  assign o[34046] = i[34046];
  assign o[34045] = i[34045];
  assign o[34044] = i[34044];
  assign o[34043] = i[34043];
  assign o[34042] = i[34042];
  assign o[34041] = i[34041];
  assign o[34040] = i[34040];
  assign o[34039] = i[34039];
  assign o[34038] = i[34038];
  assign o[34037] = i[34037];
  assign o[34036] = i[34036];
  assign o[34035] = i[34035];
  assign o[34034] = i[34034];
  assign o[34033] = i[34033];
  assign o[34032] = i[34032];
  assign o[34031] = i[34031];
  assign o[34030] = i[34030];
  assign o[34029] = i[34029];
  assign o[34028] = i[34028];
  assign o[34027] = i[34027];
  assign o[34026] = i[34026];
  assign o[34025] = i[34025];
  assign o[34024] = i[34024];
  assign o[34023] = i[34023];
  assign o[34022] = i[34022];
  assign o[34021] = i[34021];
  assign o[34020] = i[34020];
  assign o[34019] = i[34019];
  assign o[34018] = i[34018];
  assign o[34017] = i[34017];
  assign o[34016] = i[34016];
  assign o[34015] = i[34015];
  assign o[34014] = i[34014];
  assign o[34013] = i[34013];
  assign o[34012] = i[34012];
  assign o[34011] = i[34011];
  assign o[34010] = i[34010];
  assign o[34009] = i[34009];
  assign o[34008] = i[34008];
  assign o[34007] = i[34007];
  assign o[34006] = i[34006];
  assign o[34005] = i[34005];
  assign o[34004] = i[34004];
  assign o[34003] = i[34003];
  assign o[34002] = i[34002];
  assign o[34001] = i[34001];
  assign o[34000] = i[34000];
  assign o[33999] = i[33999];
  assign o[33998] = i[33998];
  assign o[33997] = i[33997];
  assign o[33996] = i[33996];
  assign o[33995] = i[33995];
  assign o[33994] = i[33994];
  assign o[33993] = i[33993];
  assign o[33992] = i[33992];
  assign o[33991] = i[33991];
  assign o[33990] = i[33990];
  assign o[33989] = i[33989];
  assign o[33988] = i[33988];
  assign o[33987] = i[33987];
  assign o[33986] = i[33986];
  assign o[33985] = i[33985];
  assign o[33984] = i[33984];
  assign o[33983] = i[33983];
  assign o[33982] = i[33982];
  assign o[33981] = i[33981];
  assign o[33980] = i[33980];
  assign o[33979] = i[33979];
  assign o[33978] = i[33978];
  assign o[33977] = i[33977];
  assign o[33976] = i[33976];
  assign o[33975] = i[33975];
  assign o[33974] = i[33974];
  assign o[33973] = i[33973];
  assign o[33972] = i[33972];
  assign o[33971] = i[33971];
  assign o[33970] = i[33970];
  assign o[33969] = i[33969];
  assign o[33968] = i[33968];
  assign o[33967] = i[33967];
  assign o[33966] = i[33966];
  assign o[33965] = i[33965];
  assign o[33964] = i[33964];
  assign o[33963] = i[33963];
  assign o[33962] = i[33962];
  assign o[33961] = i[33961];
  assign o[33960] = i[33960];
  assign o[33959] = i[33959];
  assign o[33958] = i[33958];
  assign o[33957] = i[33957];
  assign o[33956] = i[33956];
  assign o[33955] = i[33955];
  assign o[33954] = i[33954];
  assign o[33953] = i[33953];
  assign o[33952] = i[33952];
  assign o[33951] = i[33951];
  assign o[33950] = i[33950];
  assign o[33949] = i[33949];
  assign o[33948] = i[33948];
  assign o[33947] = i[33947];
  assign o[33946] = i[33946];
  assign o[33945] = i[33945];
  assign o[33944] = i[33944];
  assign o[33943] = i[33943];
  assign o[33942] = i[33942];
  assign o[33941] = i[33941];
  assign o[33940] = i[33940];
  assign o[33939] = i[33939];
  assign o[33938] = i[33938];
  assign o[33937] = i[33937];
  assign o[33936] = i[33936];
  assign o[33935] = i[33935];
  assign o[33934] = i[33934];
  assign o[33933] = i[33933];
  assign o[33932] = i[33932];
  assign o[33931] = i[33931];
  assign o[33930] = i[33930];
  assign o[33929] = i[33929];
  assign o[33928] = i[33928];
  assign o[33927] = i[33927];
  assign o[33926] = i[33926];
  assign o[33925] = i[33925];
  assign o[33924] = i[33924];
  assign o[33923] = i[33923];
  assign o[33922] = i[33922];
  assign o[33921] = i[33921];
  assign o[33920] = i[33920];
  assign o[33919] = i[33919];
  assign o[33918] = i[33918];
  assign o[33917] = i[33917];
  assign o[33916] = i[33916];
  assign o[33915] = i[33915];
  assign o[33914] = i[33914];
  assign o[33913] = i[33913];
  assign o[33912] = i[33912];
  assign o[33911] = i[33911];
  assign o[33910] = i[33910];
  assign o[33909] = i[33909];
  assign o[33908] = i[33908];
  assign o[33907] = i[33907];
  assign o[33906] = i[33906];
  assign o[33905] = i[33905];
  assign o[33904] = i[33904];
  assign o[33903] = i[33903];
  assign o[33902] = i[33902];
  assign o[33901] = i[33901];
  assign o[33900] = i[33900];
  assign o[33899] = i[33899];
  assign o[33898] = i[33898];
  assign o[33897] = i[33897];
  assign o[33896] = i[33896];
  assign o[33895] = i[33895];
  assign o[33894] = i[33894];
  assign o[33893] = i[33893];
  assign o[33892] = i[33892];
  assign o[33891] = i[33891];
  assign o[33890] = i[33890];
  assign o[33889] = i[33889];
  assign o[33888] = i[33888];
  assign o[33887] = i[33887];
  assign o[33886] = i[33886];
  assign o[33885] = i[33885];
  assign o[33884] = i[33884];
  assign o[33883] = i[33883];
  assign o[33882] = i[33882];
  assign o[33881] = i[33881];
  assign o[33880] = i[33880];
  assign o[33879] = i[33879];
  assign o[33878] = i[33878];
  assign o[33877] = i[33877];
  assign o[33876] = i[33876];
  assign o[33875] = i[33875];
  assign o[33874] = i[33874];
  assign o[33873] = i[33873];
  assign o[33872] = i[33872];
  assign o[33871] = i[33871];
  assign o[33870] = i[33870];
  assign o[33869] = i[33869];
  assign o[33868] = i[33868];
  assign o[33867] = i[33867];
  assign o[33866] = i[33866];
  assign o[33865] = i[33865];
  assign o[33864] = i[33864];
  assign o[33863] = i[33863];
  assign o[33862] = i[33862];
  assign o[33861] = i[33861];
  assign o[33860] = i[33860];
  assign o[33859] = i[33859];
  assign o[33858] = i[33858];
  assign o[33857] = i[33857];
  assign o[33856] = i[33856];
  assign o[33855] = i[33855];
  assign o[33854] = i[33854];
  assign o[33853] = i[33853];
  assign o[33852] = i[33852];
  assign o[33851] = i[33851];
  assign o[33850] = i[33850];
  assign o[33849] = i[33849];
  assign o[33848] = i[33848];
  assign o[33847] = i[33847];
  assign o[33846] = i[33846];
  assign o[33845] = i[33845];
  assign o[33844] = i[33844];
  assign o[33843] = i[33843];
  assign o[33842] = i[33842];
  assign o[33841] = i[33841];
  assign o[33840] = i[33840];
  assign o[33839] = i[33839];
  assign o[33838] = i[33838];
  assign o[33837] = i[33837];
  assign o[33836] = i[33836];
  assign o[33835] = i[33835];
  assign o[33834] = i[33834];
  assign o[33833] = i[33833];
  assign o[33832] = i[33832];
  assign o[33831] = i[33831];
  assign o[33830] = i[33830];
  assign o[33829] = i[33829];
  assign o[33828] = i[33828];
  assign o[33827] = i[33827];
  assign o[33826] = i[33826];
  assign o[33825] = i[33825];
  assign o[33824] = i[33824];
  assign o[33823] = i[33823];
  assign o[33822] = i[33822];
  assign o[33821] = i[33821];
  assign o[33820] = i[33820];
  assign o[33819] = i[33819];
  assign o[33818] = i[33818];
  assign o[33817] = i[33817];
  assign o[33816] = i[33816];
  assign o[33815] = i[33815];
  assign o[33814] = i[33814];
  assign o[33813] = i[33813];
  assign o[33812] = i[33812];
  assign o[33811] = i[33811];
  assign o[33810] = i[33810];
  assign o[33809] = i[33809];
  assign o[33808] = i[33808];
  assign o[33807] = i[33807];
  assign o[33806] = i[33806];
  assign o[33805] = i[33805];
  assign o[33804] = i[33804];
  assign o[33803] = i[33803];
  assign o[33802] = i[33802];
  assign o[33801] = i[33801];
  assign o[33800] = i[33800];
  assign o[33799] = i[33799];
  assign o[33798] = i[33798];
  assign o[33797] = i[33797];
  assign o[33796] = i[33796];
  assign o[33795] = i[33795];
  assign o[33794] = i[33794];
  assign o[33793] = i[33793];
  assign o[33792] = i[33792];
  assign o[33791] = i[33791];
  assign o[33790] = i[33790];
  assign o[33789] = i[33789];
  assign o[33788] = i[33788];
  assign o[33787] = i[33787];
  assign o[33786] = i[33786];
  assign o[33785] = i[33785];
  assign o[33784] = i[33784];
  assign o[33783] = i[33783];
  assign o[33782] = i[33782];
  assign o[33781] = i[33781];
  assign o[33780] = i[33780];
  assign o[33779] = i[33779];
  assign o[33778] = i[33778];
  assign o[33777] = i[33777];
  assign o[33776] = i[33776];
  assign o[33775] = i[33775];
  assign o[33774] = i[33774];
  assign o[33773] = i[33773];
  assign o[33772] = i[33772];
  assign o[33771] = i[33771];
  assign o[33770] = i[33770];
  assign o[33769] = i[33769];
  assign o[33768] = i[33768];
  assign o[33767] = i[33767];
  assign o[33766] = i[33766];
  assign o[33765] = i[33765];
  assign o[33764] = i[33764];
  assign o[33763] = i[33763];
  assign o[33762] = i[33762];
  assign o[33761] = i[33761];
  assign o[33760] = i[33760];
  assign o[33759] = i[33759];
  assign o[33758] = i[33758];
  assign o[33757] = i[33757];
  assign o[33756] = i[33756];
  assign o[33755] = i[33755];
  assign o[33754] = i[33754];
  assign o[33753] = i[33753];
  assign o[33752] = i[33752];
  assign o[33751] = i[33751];
  assign o[33750] = i[33750];
  assign o[33749] = i[33749];
  assign o[33748] = i[33748];
  assign o[33747] = i[33747];
  assign o[33746] = i[33746];
  assign o[33745] = i[33745];
  assign o[33744] = i[33744];
  assign o[33743] = i[33743];
  assign o[33742] = i[33742];
  assign o[33741] = i[33741];
  assign o[33740] = i[33740];
  assign o[33739] = i[33739];
  assign o[33738] = i[33738];
  assign o[33737] = i[33737];
  assign o[33736] = i[33736];
  assign o[33735] = i[33735];
  assign o[33734] = i[33734];
  assign o[33733] = i[33733];
  assign o[33732] = i[33732];
  assign o[33731] = i[33731];
  assign o[33730] = i[33730];
  assign o[33729] = i[33729];
  assign o[33728] = i[33728];
  assign o[33727] = i[33727];
  assign o[33726] = i[33726];
  assign o[33725] = i[33725];
  assign o[33724] = i[33724];
  assign o[33723] = i[33723];
  assign o[33722] = i[33722];
  assign o[33721] = i[33721];
  assign o[33720] = i[33720];
  assign o[33719] = i[33719];
  assign o[33718] = i[33718];
  assign o[33717] = i[33717];
  assign o[33716] = i[33716];
  assign o[33715] = i[33715];
  assign o[33714] = i[33714];
  assign o[33713] = i[33713];
  assign o[33712] = i[33712];
  assign o[33711] = i[33711];
  assign o[33710] = i[33710];
  assign o[33709] = i[33709];
  assign o[33708] = i[33708];
  assign o[33707] = i[33707];
  assign o[33706] = i[33706];
  assign o[33705] = i[33705];
  assign o[33704] = i[33704];
  assign o[33703] = i[33703];
  assign o[33702] = i[33702];
  assign o[33701] = i[33701];
  assign o[33700] = i[33700];
  assign o[33699] = i[33699];
  assign o[33698] = i[33698];
  assign o[33697] = i[33697];
  assign o[33696] = i[33696];
  assign o[33695] = i[33695];
  assign o[33694] = i[33694];
  assign o[33693] = i[33693];
  assign o[33692] = i[33692];
  assign o[33691] = i[33691];
  assign o[33690] = i[33690];
  assign o[33689] = i[33689];
  assign o[33688] = i[33688];
  assign o[33687] = i[33687];
  assign o[33686] = i[33686];
  assign o[33685] = i[33685];
  assign o[33684] = i[33684];
  assign o[33683] = i[33683];
  assign o[33682] = i[33682];
  assign o[33681] = i[33681];
  assign o[33680] = i[33680];
  assign o[33679] = i[33679];
  assign o[33678] = i[33678];
  assign o[33677] = i[33677];
  assign o[33676] = i[33676];
  assign o[33675] = i[33675];
  assign o[33674] = i[33674];
  assign o[33673] = i[33673];
  assign o[33672] = i[33672];
  assign o[33671] = i[33671];
  assign o[33670] = i[33670];
  assign o[33669] = i[33669];
  assign o[33668] = i[33668];
  assign o[33667] = i[33667];
  assign o[33666] = i[33666];
  assign o[33665] = i[33665];
  assign o[33664] = i[33664];
  assign o[33663] = i[33663];
  assign o[33662] = i[33662];
  assign o[33661] = i[33661];
  assign o[33660] = i[33660];
  assign o[33659] = i[33659];
  assign o[33658] = i[33658];
  assign o[33657] = i[33657];
  assign o[33656] = i[33656];
  assign o[33655] = i[33655];
  assign o[33654] = i[33654];
  assign o[33653] = i[33653];
  assign o[33652] = i[33652];
  assign o[33651] = i[33651];
  assign o[33650] = i[33650];
  assign o[33649] = i[33649];
  assign o[33648] = i[33648];
  assign o[33647] = i[33647];
  assign o[33646] = i[33646];
  assign o[33645] = i[33645];
  assign o[33644] = i[33644];
  assign o[33643] = i[33643];
  assign o[33642] = i[33642];
  assign o[33641] = i[33641];
  assign o[33640] = i[33640];
  assign o[33639] = i[33639];
  assign o[33638] = i[33638];
  assign o[33637] = i[33637];
  assign o[33636] = i[33636];
  assign o[33635] = i[33635];
  assign o[33634] = i[33634];
  assign o[33633] = i[33633];
  assign o[33632] = i[33632];
  assign o[33631] = i[33631];
  assign o[33630] = i[33630];
  assign o[33629] = i[33629];
  assign o[33628] = i[33628];
  assign o[33627] = i[33627];
  assign o[33626] = i[33626];
  assign o[33625] = i[33625];
  assign o[33624] = i[33624];
  assign o[33623] = i[33623];
  assign o[33622] = i[33622];
  assign o[33621] = i[33621];
  assign o[33620] = i[33620];
  assign o[33619] = i[33619];
  assign o[33618] = i[33618];
  assign o[33617] = i[33617];
  assign o[33616] = i[33616];
  assign o[33615] = i[33615];
  assign o[33614] = i[33614];
  assign o[33613] = i[33613];
  assign o[33612] = i[33612];
  assign o[33611] = i[33611];
  assign o[33610] = i[33610];
  assign o[33609] = i[33609];
  assign o[33608] = i[33608];
  assign o[33607] = i[33607];
  assign o[33606] = i[33606];
  assign o[33605] = i[33605];
  assign o[33604] = i[33604];
  assign o[33603] = i[33603];
  assign o[33602] = i[33602];
  assign o[33601] = i[33601];
  assign o[33600] = i[33600];
  assign o[33599] = i[33599];
  assign o[33598] = i[33598];
  assign o[33597] = i[33597];
  assign o[33596] = i[33596];
  assign o[33595] = i[33595];
  assign o[33594] = i[33594];
  assign o[33593] = i[33593];
  assign o[33592] = i[33592];
  assign o[33591] = i[33591];
  assign o[33590] = i[33590];
  assign o[33589] = i[33589];
  assign o[33588] = i[33588];
  assign o[33587] = i[33587];
  assign o[33586] = i[33586];
  assign o[33585] = i[33585];
  assign o[33584] = i[33584];
  assign o[33583] = i[33583];
  assign o[33582] = i[33582];
  assign o[33581] = i[33581];
  assign o[33580] = i[33580];
  assign o[33579] = i[33579];
  assign o[33578] = i[33578];
  assign o[33577] = i[33577];
  assign o[33576] = i[33576];
  assign o[33575] = i[33575];
  assign o[33574] = i[33574];
  assign o[33573] = i[33573];
  assign o[33572] = i[33572];
  assign o[33571] = i[33571];
  assign o[33570] = i[33570];
  assign o[33569] = i[33569];
  assign o[33568] = i[33568];
  assign o[33567] = i[33567];
  assign o[33566] = i[33566];
  assign o[33565] = i[33565];
  assign o[33564] = i[33564];
  assign o[33563] = i[33563];
  assign o[33562] = i[33562];
  assign o[33561] = i[33561];
  assign o[33560] = i[33560];
  assign o[33559] = i[33559];
  assign o[33558] = i[33558];
  assign o[33557] = i[33557];
  assign o[33556] = i[33556];
  assign o[33555] = i[33555];
  assign o[33554] = i[33554];
  assign o[33553] = i[33553];
  assign o[33552] = i[33552];
  assign o[33551] = i[33551];
  assign o[33550] = i[33550];
  assign o[33549] = i[33549];
  assign o[33548] = i[33548];
  assign o[33547] = i[33547];
  assign o[33546] = i[33546];
  assign o[33545] = i[33545];
  assign o[33544] = i[33544];
  assign o[33543] = i[33543];
  assign o[33542] = i[33542];
  assign o[33541] = i[33541];
  assign o[33540] = i[33540];
  assign o[33539] = i[33539];
  assign o[33538] = i[33538];
  assign o[33537] = i[33537];
  assign o[33536] = i[33536];
  assign o[33535] = i[33535];
  assign o[33534] = i[33534];
  assign o[33533] = i[33533];
  assign o[33532] = i[33532];
  assign o[33531] = i[33531];
  assign o[33530] = i[33530];
  assign o[33529] = i[33529];
  assign o[33528] = i[33528];
  assign o[33527] = i[33527];
  assign o[33526] = i[33526];
  assign o[33525] = i[33525];
  assign o[33524] = i[33524];
  assign o[33523] = i[33523];
  assign o[33522] = i[33522];
  assign o[33521] = i[33521];
  assign o[33520] = i[33520];
  assign o[33519] = i[33519];
  assign o[33518] = i[33518];
  assign o[33517] = i[33517];
  assign o[33516] = i[33516];
  assign o[33515] = i[33515];
  assign o[33514] = i[33514];
  assign o[33513] = i[33513];
  assign o[33512] = i[33512];
  assign o[33511] = i[33511];
  assign o[33510] = i[33510];
  assign o[33509] = i[33509];
  assign o[33508] = i[33508];
  assign o[33507] = i[33507];
  assign o[33506] = i[33506];
  assign o[33505] = i[33505];
  assign o[33504] = i[33504];
  assign o[33503] = i[33503];
  assign o[33502] = i[33502];
  assign o[33501] = i[33501];
  assign o[33500] = i[33500];
  assign o[33499] = i[33499];
  assign o[33498] = i[33498];
  assign o[33497] = i[33497];
  assign o[33496] = i[33496];
  assign o[33495] = i[33495];
  assign o[33494] = i[33494];
  assign o[33493] = i[33493];
  assign o[33492] = i[33492];
  assign o[33491] = i[33491];
  assign o[33490] = i[33490];
  assign o[33489] = i[33489];
  assign o[33488] = i[33488];
  assign o[33487] = i[33487];
  assign o[33486] = i[33486];
  assign o[33485] = i[33485];
  assign o[33484] = i[33484];
  assign o[33483] = i[33483];
  assign o[33482] = i[33482];
  assign o[33481] = i[33481];
  assign o[33480] = i[33480];
  assign o[33479] = i[33479];
  assign o[33478] = i[33478];
  assign o[33477] = i[33477];
  assign o[33476] = i[33476];
  assign o[33475] = i[33475];
  assign o[33474] = i[33474];
  assign o[33473] = i[33473];
  assign o[33472] = i[33472];
  assign o[33471] = i[33471];
  assign o[33470] = i[33470];
  assign o[33469] = i[33469];
  assign o[33468] = i[33468];
  assign o[33467] = i[33467];
  assign o[33466] = i[33466];
  assign o[33465] = i[33465];
  assign o[33464] = i[33464];
  assign o[33463] = i[33463];
  assign o[33462] = i[33462];
  assign o[33461] = i[33461];
  assign o[33460] = i[33460];
  assign o[33459] = i[33459];
  assign o[33458] = i[33458];
  assign o[33457] = i[33457];
  assign o[33456] = i[33456];
  assign o[33455] = i[33455];
  assign o[33454] = i[33454];
  assign o[33453] = i[33453];
  assign o[33452] = i[33452];
  assign o[33451] = i[33451];
  assign o[33450] = i[33450];
  assign o[33449] = i[33449];
  assign o[33448] = i[33448];
  assign o[33447] = i[33447];
  assign o[33446] = i[33446];
  assign o[33445] = i[33445];
  assign o[33444] = i[33444];
  assign o[33443] = i[33443];
  assign o[33442] = i[33442];
  assign o[33441] = i[33441];
  assign o[33440] = i[33440];
  assign o[33439] = i[33439];
  assign o[33438] = i[33438];
  assign o[33437] = i[33437];
  assign o[33436] = i[33436];
  assign o[33435] = i[33435];
  assign o[33434] = i[33434];
  assign o[33433] = i[33433];
  assign o[33432] = i[33432];
  assign o[33431] = i[33431];
  assign o[33430] = i[33430];
  assign o[33429] = i[33429];
  assign o[33428] = i[33428];
  assign o[33427] = i[33427];
  assign o[33426] = i[33426];
  assign o[33425] = i[33425];
  assign o[33424] = i[33424];
  assign o[33423] = i[33423];
  assign o[33422] = i[33422];
  assign o[33421] = i[33421];
  assign o[33420] = i[33420];
  assign o[33419] = i[33419];
  assign o[33418] = i[33418];
  assign o[33417] = i[33417];
  assign o[33416] = i[33416];
  assign o[33415] = i[33415];
  assign o[33414] = i[33414];
  assign o[33413] = i[33413];
  assign o[33412] = i[33412];
  assign o[33411] = i[33411];
  assign o[33410] = i[33410];
  assign o[33409] = i[33409];
  assign o[33408] = i[33408];
  assign o[33407] = i[33407];
  assign o[33406] = i[33406];
  assign o[33405] = i[33405];
  assign o[33404] = i[33404];
  assign o[33403] = i[33403];
  assign o[33402] = i[33402];
  assign o[33401] = i[33401];
  assign o[33400] = i[33400];
  assign o[33399] = i[33399];
  assign o[33398] = i[33398];
  assign o[33397] = i[33397];
  assign o[33396] = i[33396];
  assign o[33395] = i[33395];
  assign o[33394] = i[33394];
  assign o[33393] = i[33393];
  assign o[33392] = i[33392];
  assign o[33391] = i[33391];
  assign o[33390] = i[33390];
  assign o[33389] = i[33389];
  assign o[33388] = i[33388];
  assign o[33387] = i[33387];
  assign o[33386] = i[33386];
  assign o[33385] = i[33385];
  assign o[33384] = i[33384];
  assign o[33383] = i[33383];
  assign o[33382] = i[33382];
  assign o[33381] = i[33381];
  assign o[33380] = i[33380];
  assign o[33379] = i[33379];
  assign o[33378] = i[33378];
  assign o[33377] = i[33377];
  assign o[33376] = i[33376];
  assign o[33375] = i[33375];
  assign o[33374] = i[33374];
  assign o[33373] = i[33373];
  assign o[33372] = i[33372];
  assign o[33371] = i[33371];
  assign o[33370] = i[33370];
  assign o[33369] = i[33369];
  assign o[33368] = i[33368];
  assign o[33367] = i[33367];
  assign o[33366] = i[33366];
  assign o[33365] = i[33365];
  assign o[33364] = i[33364];
  assign o[33363] = i[33363];
  assign o[33362] = i[33362];
  assign o[33361] = i[33361];
  assign o[33360] = i[33360];
  assign o[33359] = i[33359];
  assign o[33358] = i[33358];
  assign o[33357] = i[33357];
  assign o[33356] = i[33356];
  assign o[33355] = i[33355];
  assign o[33354] = i[33354];
  assign o[33353] = i[33353];
  assign o[33352] = i[33352];
  assign o[33351] = i[33351];
  assign o[33350] = i[33350];
  assign o[33349] = i[33349];
  assign o[33348] = i[33348];
  assign o[33347] = i[33347];
  assign o[33346] = i[33346];
  assign o[33345] = i[33345];
  assign o[33344] = i[33344];
  assign o[33343] = i[33343];
  assign o[33342] = i[33342];
  assign o[33341] = i[33341];
  assign o[33340] = i[33340];
  assign o[33339] = i[33339];
  assign o[33338] = i[33338];
  assign o[33337] = i[33337];
  assign o[33336] = i[33336];
  assign o[33335] = i[33335];
  assign o[33334] = i[33334];
  assign o[33333] = i[33333];
  assign o[33332] = i[33332];
  assign o[33331] = i[33331];
  assign o[33330] = i[33330];
  assign o[33329] = i[33329];
  assign o[33328] = i[33328];
  assign o[33327] = i[33327];
  assign o[33326] = i[33326];
  assign o[33325] = i[33325];
  assign o[33324] = i[33324];
  assign o[33323] = i[33323];
  assign o[33322] = i[33322];
  assign o[33321] = i[33321];
  assign o[33320] = i[33320];
  assign o[33319] = i[33319];
  assign o[33318] = i[33318];
  assign o[33317] = i[33317];
  assign o[33316] = i[33316];
  assign o[33315] = i[33315];
  assign o[33314] = i[33314];
  assign o[33313] = i[33313];
  assign o[33312] = i[33312];
  assign o[33311] = i[33311];
  assign o[33310] = i[33310];
  assign o[33309] = i[33309];
  assign o[33308] = i[33308];
  assign o[33307] = i[33307];
  assign o[33306] = i[33306];
  assign o[33305] = i[33305];
  assign o[33304] = i[33304];
  assign o[33303] = i[33303];
  assign o[33302] = i[33302];
  assign o[33301] = i[33301];
  assign o[33300] = i[33300];
  assign o[33299] = i[33299];
  assign o[33298] = i[33298];
  assign o[33297] = i[33297];
  assign o[33296] = i[33296];
  assign o[33295] = i[33295];
  assign o[33294] = i[33294];
  assign o[33293] = i[33293];
  assign o[33292] = i[33292];
  assign o[33291] = i[33291];
  assign o[33290] = i[33290];
  assign o[33289] = i[33289];
  assign o[33288] = i[33288];
  assign o[33287] = i[33287];
  assign o[33286] = i[33286];
  assign o[33285] = i[33285];
  assign o[33284] = i[33284];
  assign o[33283] = i[33283];
  assign o[33282] = i[33282];
  assign o[33281] = i[33281];
  assign o[33280] = i[33280];
  assign o[33279] = i[33279];
  assign o[33278] = i[33278];
  assign o[33277] = i[33277];
  assign o[33276] = i[33276];
  assign o[33275] = i[33275];
  assign o[33274] = i[33274];
  assign o[33273] = i[33273];
  assign o[33272] = i[33272];
  assign o[33271] = i[33271];
  assign o[33270] = i[33270];
  assign o[33269] = i[33269];
  assign o[33268] = i[33268];
  assign o[33267] = i[33267];
  assign o[33266] = i[33266];
  assign o[33265] = i[33265];
  assign o[33264] = i[33264];
  assign o[33263] = i[33263];
  assign o[33262] = i[33262];
  assign o[33261] = i[33261];
  assign o[33260] = i[33260];
  assign o[33259] = i[33259];
  assign o[33258] = i[33258];
  assign o[33257] = i[33257];
  assign o[33256] = i[33256];
  assign o[33255] = i[33255];
  assign o[33254] = i[33254];
  assign o[33253] = i[33253];
  assign o[33252] = i[33252];
  assign o[33251] = i[33251];
  assign o[33250] = i[33250];
  assign o[33249] = i[33249];
  assign o[33248] = i[33248];
  assign o[33247] = i[33247];
  assign o[33246] = i[33246];
  assign o[33245] = i[33245];
  assign o[33244] = i[33244];
  assign o[33243] = i[33243];
  assign o[33242] = i[33242];
  assign o[33241] = i[33241];
  assign o[33240] = i[33240];
  assign o[33239] = i[33239];
  assign o[33238] = i[33238];
  assign o[33237] = i[33237];
  assign o[33236] = i[33236];
  assign o[33235] = i[33235];
  assign o[33234] = i[33234];
  assign o[33233] = i[33233];
  assign o[33232] = i[33232];
  assign o[33231] = i[33231];
  assign o[33230] = i[33230];
  assign o[33229] = i[33229];
  assign o[33228] = i[33228];
  assign o[33227] = i[33227];
  assign o[33226] = i[33226];
  assign o[33225] = i[33225];
  assign o[33224] = i[33224];
  assign o[33223] = i[33223];
  assign o[33222] = i[33222];
  assign o[33221] = i[33221];
  assign o[33220] = i[33220];
  assign o[33219] = i[33219];
  assign o[33218] = i[33218];
  assign o[33217] = i[33217];
  assign o[33216] = i[33216];
  assign o[33215] = i[33215];
  assign o[33214] = i[33214];
  assign o[33213] = i[33213];
  assign o[33212] = i[33212];
  assign o[33211] = i[33211];
  assign o[33210] = i[33210];
  assign o[33209] = i[33209];
  assign o[33208] = i[33208];
  assign o[33207] = i[33207];
  assign o[33206] = i[33206];
  assign o[33205] = i[33205];
  assign o[33204] = i[33204];
  assign o[33203] = i[33203];
  assign o[33202] = i[33202];
  assign o[33201] = i[33201];
  assign o[33200] = i[33200];
  assign o[33199] = i[33199];
  assign o[33198] = i[33198];
  assign o[33197] = i[33197];
  assign o[33196] = i[33196];
  assign o[33195] = i[33195];
  assign o[33194] = i[33194];
  assign o[33193] = i[33193];
  assign o[33192] = i[33192];
  assign o[33191] = i[33191];
  assign o[33190] = i[33190];
  assign o[33189] = i[33189];
  assign o[33188] = i[33188];
  assign o[33187] = i[33187];
  assign o[33186] = i[33186];
  assign o[33185] = i[33185];
  assign o[33184] = i[33184];
  assign o[33183] = i[33183];
  assign o[33182] = i[33182];
  assign o[33181] = i[33181];
  assign o[33180] = i[33180];
  assign o[33179] = i[33179];
  assign o[33178] = i[33178];
  assign o[33177] = i[33177];
  assign o[33176] = i[33176];
  assign o[33175] = i[33175];
  assign o[33174] = i[33174];
  assign o[33173] = i[33173];
  assign o[33172] = i[33172];
  assign o[33171] = i[33171];
  assign o[33170] = i[33170];
  assign o[33169] = i[33169];
  assign o[33168] = i[33168];
  assign o[33167] = i[33167];
  assign o[33166] = i[33166];
  assign o[33165] = i[33165];
  assign o[33164] = i[33164];
  assign o[33163] = i[33163];
  assign o[33162] = i[33162];
  assign o[33161] = i[33161];
  assign o[33160] = i[33160];
  assign o[33159] = i[33159];
  assign o[33158] = i[33158];
  assign o[33157] = i[33157];
  assign o[33156] = i[33156];
  assign o[33155] = i[33155];
  assign o[33154] = i[33154];
  assign o[33153] = i[33153];
  assign o[33152] = i[33152];
  assign o[33151] = i[33151];
  assign o[33150] = i[33150];
  assign o[33149] = i[33149];
  assign o[33148] = i[33148];
  assign o[33147] = i[33147];
  assign o[33146] = i[33146];
  assign o[33145] = i[33145];
  assign o[33144] = i[33144];
  assign o[33143] = i[33143];
  assign o[33142] = i[33142];
  assign o[33141] = i[33141];
  assign o[33140] = i[33140];
  assign o[33139] = i[33139];
  assign o[33138] = i[33138];
  assign o[33137] = i[33137];
  assign o[33136] = i[33136];
  assign o[33135] = i[33135];
  assign o[33134] = i[33134];
  assign o[33133] = i[33133];
  assign o[33132] = i[33132];
  assign o[33131] = i[33131];
  assign o[33130] = i[33130];
  assign o[33129] = i[33129];
  assign o[33128] = i[33128];
  assign o[33127] = i[33127];
  assign o[33126] = i[33126];
  assign o[33125] = i[33125];
  assign o[33124] = i[33124];
  assign o[33123] = i[33123];
  assign o[33122] = i[33122];
  assign o[33121] = i[33121];
  assign o[33120] = i[33120];
  assign o[33119] = i[33119];
  assign o[33118] = i[33118];
  assign o[33117] = i[33117];
  assign o[33116] = i[33116];
  assign o[33115] = i[33115];
  assign o[33114] = i[33114];
  assign o[33113] = i[33113];
  assign o[33112] = i[33112];
  assign o[33111] = i[33111];
  assign o[33110] = i[33110];
  assign o[33109] = i[33109];
  assign o[33108] = i[33108];
  assign o[33107] = i[33107];
  assign o[33106] = i[33106];
  assign o[33105] = i[33105];
  assign o[33104] = i[33104];
  assign o[33103] = i[33103];
  assign o[33102] = i[33102];
  assign o[33101] = i[33101];
  assign o[33100] = i[33100];
  assign o[33099] = i[33099];
  assign o[33098] = i[33098];
  assign o[33097] = i[33097];
  assign o[33096] = i[33096];
  assign o[33095] = i[33095];
  assign o[33094] = i[33094];
  assign o[33093] = i[33093];
  assign o[33092] = i[33092];
  assign o[33091] = i[33091];
  assign o[33090] = i[33090];
  assign o[33089] = i[33089];
  assign o[33088] = i[33088];
  assign o[33087] = i[33087];
  assign o[33086] = i[33086];
  assign o[33085] = i[33085];
  assign o[33084] = i[33084];
  assign o[33083] = i[33083];
  assign o[33082] = i[33082];
  assign o[33081] = i[33081];
  assign o[33080] = i[33080];
  assign o[33079] = i[33079];
  assign o[33078] = i[33078];
  assign o[33077] = i[33077];
  assign o[33076] = i[33076];
  assign o[33075] = i[33075];
  assign o[33074] = i[33074];
  assign o[33073] = i[33073];
  assign o[33072] = i[33072];
  assign o[33071] = i[33071];
  assign o[33070] = i[33070];
  assign o[33069] = i[33069];
  assign o[33068] = i[33068];
  assign o[33067] = i[33067];
  assign o[33066] = i[33066];
  assign o[33065] = i[33065];
  assign o[33064] = i[33064];
  assign o[33063] = i[33063];
  assign o[33062] = i[33062];
  assign o[33061] = i[33061];
  assign o[33060] = i[33060];
  assign o[33059] = i[33059];
  assign o[33058] = i[33058];
  assign o[33057] = i[33057];
  assign o[33056] = i[33056];
  assign o[33055] = i[33055];
  assign o[33054] = i[33054];
  assign o[33053] = i[33053];
  assign o[33052] = i[33052];
  assign o[33051] = i[33051];
  assign o[33050] = i[33050];
  assign o[33049] = i[33049];
  assign o[33048] = i[33048];
  assign o[33047] = i[33047];
  assign o[33046] = i[33046];
  assign o[33045] = i[33045];
  assign o[33044] = i[33044];
  assign o[33043] = i[33043];
  assign o[33042] = i[33042];
  assign o[33041] = i[33041];
  assign o[33040] = i[33040];
  assign o[33039] = i[33039];
  assign o[33038] = i[33038];
  assign o[33037] = i[33037];
  assign o[33036] = i[33036];
  assign o[33035] = i[33035];
  assign o[33034] = i[33034];
  assign o[33033] = i[33033];
  assign o[33032] = i[33032];
  assign o[33031] = i[33031];
  assign o[33030] = i[33030];
  assign o[33029] = i[33029];
  assign o[33028] = i[33028];
  assign o[33027] = i[33027];
  assign o[33026] = i[33026];
  assign o[33025] = i[33025];
  assign o[33024] = i[33024];
  assign o[33023] = i[33023];
  assign o[33022] = i[33022];
  assign o[33021] = i[33021];
  assign o[33020] = i[33020];
  assign o[33019] = i[33019];
  assign o[33018] = i[33018];
  assign o[33017] = i[33017];
  assign o[33016] = i[33016];
  assign o[33015] = i[33015];
  assign o[33014] = i[33014];
  assign o[33013] = i[33013];
  assign o[33012] = i[33012];
  assign o[33011] = i[33011];
  assign o[33010] = i[33010];
  assign o[33009] = i[33009];
  assign o[33008] = i[33008];
  assign o[33007] = i[33007];
  assign o[33006] = i[33006];
  assign o[33005] = i[33005];
  assign o[33004] = i[33004];
  assign o[33003] = i[33003];
  assign o[33002] = i[33002];
  assign o[33001] = i[33001];
  assign o[33000] = i[33000];
  assign o[32999] = i[32999];
  assign o[32998] = i[32998];
  assign o[32997] = i[32997];
  assign o[32996] = i[32996];
  assign o[32995] = i[32995];
  assign o[32994] = i[32994];
  assign o[32993] = i[32993];
  assign o[32992] = i[32992];
  assign o[32991] = i[32991];
  assign o[32990] = i[32990];
  assign o[32989] = i[32989];
  assign o[32988] = i[32988];
  assign o[32987] = i[32987];
  assign o[32986] = i[32986];
  assign o[32985] = i[32985];
  assign o[32984] = i[32984];
  assign o[32983] = i[32983];
  assign o[32982] = i[32982];
  assign o[32981] = i[32981];
  assign o[32980] = i[32980];
  assign o[32979] = i[32979];
  assign o[32978] = i[32978];
  assign o[32977] = i[32977];
  assign o[32976] = i[32976];
  assign o[32975] = i[32975];
  assign o[32974] = i[32974];
  assign o[32973] = i[32973];
  assign o[32972] = i[32972];
  assign o[32971] = i[32971];
  assign o[32970] = i[32970];
  assign o[32969] = i[32969];
  assign o[32968] = i[32968];
  assign o[32967] = i[32967];
  assign o[32966] = i[32966];
  assign o[32965] = i[32965];
  assign o[32964] = i[32964];
  assign o[32963] = i[32963];
  assign o[32962] = i[32962];
  assign o[32961] = i[32961];
  assign o[32960] = i[32960];
  assign o[32959] = i[32959];
  assign o[32958] = i[32958];
  assign o[32957] = i[32957];
  assign o[32956] = i[32956];
  assign o[32955] = i[32955];
  assign o[32954] = i[32954];
  assign o[32953] = i[32953];
  assign o[32952] = i[32952];
  assign o[32951] = i[32951];
  assign o[32950] = i[32950];
  assign o[32949] = i[32949];
  assign o[32948] = i[32948];
  assign o[32947] = i[32947];
  assign o[32946] = i[32946];
  assign o[32945] = i[32945];
  assign o[32944] = i[32944];
  assign o[32943] = i[32943];
  assign o[32942] = i[32942];
  assign o[32941] = i[32941];
  assign o[32940] = i[32940];
  assign o[32939] = i[32939];
  assign o[32938] = i[32938];
  assign o[32937] = i[32937];
  assign o[32936] = i[32936];
  assign o[32935] = i[32935];
  assign o[32934] = i[32934];
  assign o[32933] = i[32933];
  assign o[32932] = i[32932];
  assign o[32931] = i[32931];
  assign o[32930] = i[32930];
  assign o[32929] = i[32929];
  assign o[32928] = i[32928];
  assign o[32927] = i[32927];
  assign o[32926] = i[32926];
  assign o[32925] = i[32925];
  assign o[32924] = i[32924];
  assign o[32923] = i[32923];
  assign o[32922] = i[32922];
  assign o[32921] = i[32921];
  assign o[32920] = i[32920];
  assign o[32919] = i[32919];
  assign o[32918] = i[32918];
  assign o[32917] = i[32917];
  assign o[32916] = i[32916];
  assign o[32915] = i[32915];
  assign o[32914] = i[32914];
  assign o[32913] = i[32913];
  assign o[32912] = i[32912];
  assign o[32911] = i[32911];
  assign o[32910] = i[32910];
  assign o[32909] = i[32909];
  assign o[32908] = i[32908];
  assign o[32907] = i[32907];
  assign o[32906] = i[32906];
  assign o[32905] = i[32905];
  assign o[32904] = i[32904];
  assign o[32903] = i[32903];
  assign o[32902] = i[32902];
  assign o[32901] = i[32901];
  assign o[32900] = i[32900];
  assign o[32899] = i[32899];
  assign o[32898] = i[32898];
  assign o[32897] = i[32897];
  assign o[32896] = i[32896];
  assign o[32895] = i[32895];
  assign o[32894] = i[32894];
  assign o[32893] = i[32893];
  assign o[32892] = i[32892];
  assign o[32891] = i[32891];
  assign o[32890] = i[32890];
  assign o[32889] = i[32889];
  assign o[32888] = i[32888];
  assign o[32887] = i[32887];
  assign o[32886] = i[32886];
  assign o[32885] = i[32885];
  assign o[32884] = i[32884];
  assign o[32883] = i[32883];
  assign o[32882] = i[32882];
  assign o[32881] = i[32881];
  assign o[32880] = i[32880];
  assign o[32879] = i[32879];
  assign o[32878] = i[32878];
  assign o[32877] = i[32877];
  assign o[32876] = i[32876];
  assign o[32875] = i[32875];
  assign o[32874] = i[32874];
  assign o[32873] = i[32873];
  assign o[32872] = i[32872];
  assign o[32871] = i[32871];
  assign o[32870] = i[32870];
  assign o[32869] = i[32869];
  assign o[32868] = i[32868];
  assign o[32867] = i[32867];
  assign o[32866] = i[32866];
  assign o[32865] = i[32865];
  assign o[32864] = i[32864];
  assign o[32863] = i[32863];
  assign o[32862] = i[32862];
  assign o[32861] = i[32861];
  assign o[32860] = i[32860];
  assign o[32859] = i[32859];
  assign o[32858] = i[32858];
  assign o[32857] = i[32857];
  assign o[32856] = i[32856];
  assign o[32855] = i[32855];
  assign o[32854] = i[32854];
  assign o[32853] = i[32853];
  assign o[32852] = i[32852];
  assign o[32851] = i[32851];
  assign o[32850] = i[32850];
  assign o[32849] = i[32849];
  assign o[32848] = i[32848];
  assign o[32847] = i[32847];
  assign o[32846] = i[32846];
  assign o[32845] = i[32845];
  assign o[32844] = i[32844];
  assign o[32843] = i[32843];
  assign o[32842] = i[32842];
  assign o[32841] = i[32841];
  assign o[32840] = i[32840];
  assign o[32839] = i[32839];
  assign o[32838] = i[32838];
  assign o[32837] = i[32837];
  assign o[32836] = i[32836];
  assign o[32835] = i[32835];
  assign o[32834] = i[32834];
  assign o[32833] = i[32833];
  assign o[32832] = i[32832];
  assign o[32831] = i[32831];
  assign o[32830] = i[32830];
  assign o[32829] = i[32829];
  assign o[32828] = i[32828];
  assign o[32827] = i[32827];
  assign o[32826] = i[32826];
  assign o[32825] = i[32825];
  assign o[32824] = i[32824];
  assign o[32823] = i[32823];
  assign o[32822] = i[32822];
  assign o[32821] = i[32821];
  assign o[32820] = i[32820];
  assign o[32819] = i[32819];
  assign o[32818] = i[32818];
  assign o[32817] = i[32817];
  assign o[32816] = i[32816];
  assign o[32815] = i[32815];
  assign o[32814] = i[32814];
  assign o[32813] = i[32813];
  assign o[32812] = i[32812];
  assign o[32811] = i[32811];
  assign o[32810] = i[32810];
  assign o[32809] = i[32809];
  assign o[32808] = i[32808];
  assign o[32807] = i[32807];
  assign o[32806] = i[32806];
  assign o[32805] = i[32805];
  assign o[32804] = i[32804];
  assign o[32803] = i[32803];
  assign o[32802] = i[32802];
  assign o[32801] = i[32801];
  assign o[32800] = i[32800];
  assign o[32799] = i[32799];
  assign o[32798] = i[32798];
  assign o[32797] = i[32797];
  assign o[32796] = i[32796];
  assign o[32795] = i[32795];
  assign o[32794] = i[32794];
  assign o[32793] = i[32793];
  assign o[32792] = i[32792];
  assign o[32791] = i[32791];
  assign o[32790] = i[32790];
  assign o[32789] = i[32789];
  assign o[32788] = i[32788];
  assign o[32787] = i[32787];
  assign o[32786] = i[32786];
  assign o[32785] = i[32785];
  assign o[32784] = i[32784];
  assign o[32783] = i[32783];
  assign o[32782] = i[32782];
  assign o[32781] = i[32781];
  assign o[32780] = i[32780];
  assign o[32779] = i[32779];
  assign o[32778] = i[32778];
  assign o[32777] = i[32777];
  assign o[32776] = i[32776];
  assign o[32775] = i[32775];
  assign o[32774] = i[32774];
  assign o[32773] = i[32773];
  assign o[32772] = i[32772];
  assign o[32771] = i[32771];
  assign o[32770] = i[32770];
  assign o[32769] = i[32769];
  assign o[32768] = i[32768];
  assign o[32767] = i[32767];
  assign o[32766] = i[32766];
  assign o[32765] = i[32765];
  assign o[32764] = i[32764];
  assign o[32763] = i[32763];
  assign o[32762] = i[32762];
  assign o[32761] = i[32761];
  assign o[32760] = i[32760];
  assign o[32759] = i[32759];
  assign o[32758] = i[32758];
  assign o[32757] = i[32757];
  assign o[32756] = i[32756];
  assign o[32755] = i[32755];
  assign o[32754] = i[32754];
  assign o[32753] = i[32753];
  assign o[32752] = i[32752];
  assign o[32751] = i[32751];
  assign o[32750] = i[32750];
  assign o[32749] = i[32749];
  assign o[32748] = i[32748];
  assign o[32747] = i[32747];
  assign o[32746] = i[32746];
  assign o[32745] = i[32745];
  assign o[32744] = i[32744];
  assign o[32743] = i[32743];
  assign o[32742] = i[32742];
  assign o[32741] = i[32741];
  assign o[32740] = i[32740];
  assign o[32739] = i[32739];
  assign o[32738] = i[32738];
  assign o[32737] = i[32737];
  assign o[32736] = i[32736];
  assign o[32735] = i[32735];
  assign o[32734] = i[32734];
  assign o[32733] = i[32733];
  assign o[32732] = i[32732];
  assign o[32731] = i[32731];
  assign o[32730] = i[32730];
  assign o[32729] = i[32729];
  assign o[32728] = i[32728];
  assign o[32727] = i[32727];
  assign o[32726] = i[32726];
  assign o[32725] = i[32725];
  assign o[32724] = i[32724];
  assign o[32723] = i[32723];
  assign o[32722] = i[32722];
  assign o[32721] = i[32721];
  assign o[32720] = i[32720];
  assign o[32719] = i[32719];
  assign o[32718] = i[32718];
  assign o[32717] = i[32717];
  assign o[32716] = i[32716];
  assign o[32715] = i[32715];
  assign o[32714] = i[32714];
  assign o[32713] = i[32713];
  assign o[32712] = i[32712];
  assign o[32711] = i[32711];
  assign o[32710] = i[32710];
  assign o[32709] = i[32709];
  assign o[32708] = i[32708];
  assign o[32707] = i[32707];
  assign o[32706] = i[32706];
  assign o[32705] = i[32705];
  assign o[32704] = i[32704];
  assign o[32703] = i[32703];
  assign o[32702] = i[32702];
  assign o[32701] = i[32701];
  assign o[32700] = i[32700];
  assign o[32699] = i[32699];
  assign o[32698] = i[32698];
  assign o[32697] = i[32697];
  assign o[32696] = i[32696];
  assign o[32695] = i[32695];
  assign o[32694] = i[32694];
  assign o[32693] = i[32693];
  assign o[32692] = i[32692];
  assign o[32691] = i[32691];
  assign o[32690] = i[32690];
  assign o[32689] = i[32689];
  assign o[32688] = i[32688];
  assign o[32687] = i[32687];
  assign o[32686] = i[32686];
  assign o[32685] = i[32685];
  assign o[32684] = i[32684];
  assign o[32683] = i[32683];
  assign o[32682] = i[32682];
  assign o[32681] = i[32681];
  assign o[32680] = i[32680];
  assign o[32679] = i[32679];
  assign o[32678] = i[32678];
  assign o[32677] = i[32677];
  assign o[32676] = i[32676];
  assign o[32675] = i[32675];
  assign o[32674] = i[32674];
  assign o[32673] = i[32673];
  assign o[32672] = i[32672];
  assign o[32671] = i[32671];
  assign o[32670] = i[32670];
  assign o[32669] = i[32669];
  assign o[32668] = i[32668];
  assign o[32667] = i[32667];
  assign o[32666] = i[32666];
  assign o[32665] = i[32665];
  assign o[32664] = i[32664];
  assign o[32663] = i[32663];
  assign o[32662] = i[32662];
  assign o[32661] = i[32661];
  assign o[32660] = i[32660];
  assign o[32659] = i[32659];
  assign o[32658] = i[32658];
  assign o[32657] = i[32657];
  assign o[32656] = i[32656];
  assign o[32655] = i[32655];
  assign o[32654] = i[32654];
  assign o[32653] = i[32653];
  assign o[32652] = i[32652];
  assign o[32651] = i[32651];
  assign o[32650] = i[32650];
  assign o[32649] = i[32649];
  assign o[32648] = i[32648];
  assign o[32647] = i[32647];
  assign o[32646] = i[32646];
  assign o[32645] = i[32645];
  assign o[32644] = i[32644];
  assign o[32643] = i[32643];
  assign o[32642] = i[32642];
  assign o[32641] = i[32641];
  assign o[32640] = i[32640];
  assign o[32639] = i[32639];
  assign o[32638] = i[32638];
  assign o[32637] = i[32637];
  assign o[32636] = i[32636];
  assign o[32635] = i[32635];
  assign o[32634] = i[32634];
  assign o[32633] = i[32633];
  assign o[32632] = i[32632];
  assign o[32631] = i[32631];
  assign o[32630] = i[32630];
  assign o[32629] = i[32629];
  assign o[32628] = i[32628];
  assign o[32627] = i[32627];
  assign o[32626] = i[32626];
  assign o[32625] = i[32625];
  assign o[32624] = i[32624];
  assign o[32623] = i[32623];
  assign o[32622] = i[32622];
  assign o[32621] = i[32621];
  assign o[32620] = i[32620];
  assign o[32619] = i[32619];
  assign o[32618] = i[32618];
  assign o[32617] = i[32617];
  assign o[32616] = i[32616];
  assign o[32615] = i[32615];
  assign o[32614] = i[32614];
  assign o[32613] = i[32613];
  assign o[32612] = i[32612];
  assign o[32611] = i[32611];
  assign o[32610] = i[32610];
  assign o[32609] = i[32609];
  assign o[32608] = i[32608];
  assign o[32607] = i[32607];
  assign o[32606] = i[32606];
  assign o[32605] = i[32605];
  assign o[32604] = i[32604];
  assign o[32603] = i[32603];
  assign o[32602] = i[32602];
  assign o[32601] = i[32601];
  assign o[32600] = i[32600];
  assign o[32599] = i[32599];
  assign o[32598] = i[32598];
  assign o[32597] = i[32597];
  assign o[32596] = i[32596];
  assign o[32595] = i[32595];
  assign o[32594] = i[32594];
  assign o[32593] = i[32593];
  assign o[32592] = i[32592];
  assign o[32591] = i[32591];
  assign o[32590] = i[32590];
  assign o[32589] = i[32589];
  assign o[32588] = i[32588];
  assign o[32587] = i[32587];
  assign o[32586] = i[32586];
  assign o[32585] = i[32585];
  assign o[32584] = i[32584];
  assign o[32583] = i[32583];
  assign o[32582] = i[32582];
  assign o[32581] = i[32581];
  assign o[32580] = i[32580];
  assign o[32579] = i[32579];
  assign o[32578] = i[32578];
  assign o[32577] = i[32577];
  assign o[32576] = i[32576];
  assign o[32575] = i[32575];
  assign o[32574] = i[32574];
  assign o[32573] = i[32573];
  assign o[32572] = i[32572];
  assign o[32571] = i[32571];
  assign o[32570] = i[32570];
  assign o[32569] = i[32569];
  assign o[32568] = i[32568];
  assign o[32567] = i[32567];
  assign o[32566] = i[32566];
  assign o[32565] = i[32565];
  assign o[32564] = i[32564];
  assign o[32563] = i[32563];
  assign o[32562] = i[32562];
  assign o[32561] = i[32561];
  assign o[32560] = i[32560];
  assign o[32559] = i[32559];
  assign o[32558] = i[32558];
  assign o[32557] = i[32557];
  assign o[32556] = i[32556];
  assign o[32555] = i[32555];
  assign o[32554] = i[32554];
  assign o[32553] = i[32553];
  assign o[32552] = i[32552];
  assign o[32551] = i[32551];
  assign o[32550] = i[32550];
  assign o[32549] = i[32549];
  assign o[32548] = i[32548];
  assign o[32547] = i[32547];
  assign o[32546] = i[32546];
  assign o[32545] = i[32545];
  assign o[32544] = i[32544];
  assign o[32543] = i[32543];
  assign o[32542] = i[32542];
  assign o[32541] = i[32541];
  assign o[32540] = i[32540];
  assign o[32539] = i[32539];
  assign o[32538] = i[32538];
  assign o[32537] = i[32537];
  assign o[32536] = i[32536];
  assign o[32535] = i[32535];
  assign o[32534] = i[32534];
  assign o[32533] = i[32533];
  assign o[32532] = i[32532];
  assign o[32531] = i[32531];
  assign o[32530] = i[32530];
  assign o[32529] = i[32529];
  assign o[32528] = i[32528];
  assign o[32527] = i[32527];
  assign o[32526] = i[32526];
  assign o[32525] = i[32525];
  assign o[32524] = i[32524];
  assign o[32523] = i[32523];
  assign o[32522] = i[32522];
  assign o[32521] = i[32521];
  assign o[32520] = i[32520];
  assign o[32519] = i[32519];
  assign o[32518] = i[32518];
  assign o[32517] = i[32517];
  assign o[32516] = i[32516];
  assign o[32515] = i[32515];
  assign o[32514] = i[32514];
  assign o[32513] = i[32513];
  assign o[32512] = i[32512];
  assign o[32511] = i[32511];
  assign o[32510] = i[32510];
  assign o[32509] = i[32509];
  assign o[32508] = i[32508];
  assign o[32507] = i[32507];
  assign o[32506] = i[32506];
  assign o[32505] = i[32505];
  assign o[32504] = i[32504];
  assign o[32503] = i[32503];
  assign o[32502] = i[32502];
  assign o[32501] = i[32501];
  assign o[32500] = i[32500];
  assign o[32499] = i[32499];
  assign o[32498] = i[32498];
  assign o[32497] = i[32497];
  assign o[32496] = i[32496];
  assign o[32495] = i[32495];
  assign o[32494] = i[32494];
  assign o[32493] = i[32493];
  assign o[32492] = i[32492];
  assign o[32491] = i[32491];
  assign o[32490] = i[32490];
  assign o[32489] = i[32489];
  assign o[32488] = i[32488];
  assign o[32487] = i[32487];
  assign o[32486] = i[32486];
  assign o[32485] = i[32485];
  assign o[32484] = i[32484];
  assign o[32483] = i[32483];
  assign o[32482] = i[32482];
  assign o[32481] = i[32481];
  assign o[32480] = i[32480];
  assign o[32479] = i[32479];
  assign o[32478] = i[32478];
  assign o[32477] = i[32477];
  assign o[32476] = i[32476];
  assign o[32475] = i[32475];
  assign o[32474] = i[32474];
  assign o[32473] = i[32473];
  assign o[32472] = i[32472];
  assign o[32471] = i[32471];
  assign o[32470] = i[32470];
  assign o[32469] = i[32469];
  assign o[32468] = i[32468];
  assign o[32467] = i[32467];
  assign o[32466] = i[32466];
  assign o[32465] = i[32465];
  assign o[32464] = i[32464];
  assign o[32463] = i[32463];
  assign o[32462] = i[32462];
  assign o[32461] = i[32461];
  assign o[32460] = i[32460];
  assign o[32459] = i[32459];
  assign o[32458] = i[32458];
  assign o[32457] = i[32457];
  assign o[32456] = i[32456];
  assign o[32455] = i[32455];
  assign o[32454] = i[32454];
  assign o[32453] = i[32453];
  assign o[32452] = i[32452];
  assign o[32451] = i[32451];
  assign o[32450] = i[32450];
  assign o[32449] = i[32449];
  assign o[32448] = i[32448];
  assign o[32447] = i[32447];
  assign o[32446] = i[32446];
  assign o[32445] = i[32445];
  assign o[32444] = i[32444];
  assign o[32443] = i[32443];
  assign o[32442] = i[32442];
  assign o[32441] = i[32441];
  assign o[32440] = i[32440];
  assign o[32439] = i[32439];
  assign o[32438] = i[32438];
  assign o[32437] = i[32437];
  assign o[32436] = i[32436];
  assign o[32435] = i[32435];
  assign o[32434] = i[32434];
  assign o[32433] = i[32433];
  assign o[32432] = i[32432];
  assign o[32431] = i[32431];
  assign o[32430] = i[32430];
  assign o[32429] = i[32429];
  assign o[32428] = i[32428];
  assign o[32427] = i[32427];
  assign o[32426] = i[32426];
  assign o[32425] = i[32425];
  assign o[32424] = i[32424];
  assign o[32423] = i[32423];
  assign o[32422] = i[32422];
  assign o[32421] = i[32421];
  assign o[32420] = i[32420];
  assign o[32419] = i[32419];
  assign o[32418] = i[32418];
  assign o[32417] = i[32417];
  assign o[32416] = i[32416];
  assign o[32415] = i[32415];
  assign o[32414] = i[32414];
  assign o[32413] = i[32413];
  assign o[32412] = i[32412];
  assign o[32411] = i[32411];
  assign o[32410] = i[32410];
  assign o[32409] = i[32409];
  assign o[32408] = i[32408];
  assign o[32407] = i[32407];
  assign o[32406] = i[32406];
  assign o[32405] = i[32405];
  assign o[32404] = i[32404];
  assign o[32403] = i[32403];
  assign o[32402] = i[32402];
  assign o[32401] = i[32401];
  assign o[32400] = i[32400];
  assign o[32399] = i[32399];
  assign o[32398] = i[32398];
  assign o[32397] = i[32397];
  assign o[32396] = i[32396];
  assign o[32395] = i[32395];
  assign o[32394] = i[32394];
  assign o[32393] = i[32393];
  assign o[32392] = i[32392];
  assign o[32391] = i[32391];
  assign o[32390] = i[32390];
  assign o[32389] = i[32389];
  assign o[32388] = i[32388];
  assign o[32387] = i[32387];
  assign o[32386] = i[32386];
  assign o[32385] = i[32385];
  assign o[32384] = i[32384];
  assign o[32383] = i[32383];
  assign o[32382] = i[32382];
  assign o[32381] = i[32381];
  assign o[32380] = i[32380];
  assign o[32379] = i[32379];
  assign o[32378] = i[32378];
  assign o[32377] = i[32377];
  assign o[32376] = i[32376];
  assign o[32375] = i[32375];
  assign o[32374] = i[32374];
  assign o[32373] = i[32373];
  assign o[32372] = i[32372];
  assign o[32371] = i[32371];
  assign o[32370] = i[32370];
  assign o[32369] = i[32369];
  assign o[32368] = i[32368];
  assign o[32367] = i[32367];
  assign o[32366] = i[32366];
  assign o[32365] = i[32365];
  assign o[32364] = i[32364];
  assign o[32363] = i[32363];
  assign o[32362] = i[32362];
  assign o[32361] = i[32361];
  assign o[32360] = i[32360];
  assign o[32359] = i[32359];
  assign o[32358] = i[32358];
  assign o[32357] = i[32357];
  assign o[32356] = i[32356];
  assign o[32355] = i[32355];
  assign o[32354] = i[32354];
  assign o[32353] = i[32353];
  assign o[32352] = i[32352];
  assign o[32351] = i[32351];
  assign o[32350] = i[32350];
  assign o[32349] = i[32349];
  assign o[32348] = i[32348];
  assign o[32347] = i[32347];
  assign o[32346] = i[32346];
  assign o[32345] = i[32345];
  assign o[32344] = i[32344];
  assign o[32343] = i[32343];
  assign o[32342] = i[32342];
  assign o[32341] = i[32341];
  assign o[32340] = i[32340];
  assign o[32339] = i[32339];
  assign o[32338] = i[32338];
  assign o[32337] = i[32337];
  assign o[32336] = i[32336];
  assign o[32335] = i[32335];
  assign o[32334] = i[32334];
  assign o[32333] = i[32333];
  assign o[32332] = i[32332];
  assign o[32331] = i[32331];
  assign o[32330] = i[32330];
  assign o[32329] = i[32329];
  assign o[32328] = i[32328];
  assign o[32327] = i[32327];
  assign o[32326] = i[32326];
  assign o[32325] = i[32325];
  assign o[32324] = i[32324];
  assign o[32323] = i[32323];
  assign o[32322] = i[32322];
  assign o[32321] = i[32321];
  assign o[32320] = i[32320];
  assign o[32319] = i[32319];
  assign o[32318] = i[32318];
  assign o[32317] = i[32317];
  assign o[32316] = i[32316];
  assign o[32315] = i[32315];
  assign o[32314] = i[32314];
  assign o[32313] = i[32313];
  assign o[32312] = i[32312];
  assign o[32311] = i[32311];
  assign o[32310] = i[32310];
  assign o[32309] = i[32309];
  assign o[32308] = i[32308];
  assign o[32307] = i[32307];
  assign o[32306] = i[32306];
  assign o[32305] = i[32305];
  assign o[32304] = i[32304];
  assign o[32303] = i[32303];
  assign o[32302] = i[32302];
  assign o[32301] = i[32301];
  assign o[32300] = i[32300];
  assign o[32299] = i[32299];
  assign o[32298] = i[32298];
  assign o[32297] = i[32297];
  assign o[32296] = i[32296];
  assign o[32295] = i[32295];
  assign o[32294] = i[32294];
  assign o[32293] = i[32293];
  assign o[32292] = i[32292];
  assign o[32291] = i[32291];
  assign o[32290] = i[32290];
  assign o[32289] = i[32289];
  assign o[32288] = i[32288];
  assign o[32287] = i[32287];
  assign o[32286] = i[32286];
  assign o[32285] = i[32285];
  assign o[32284] = i[32284];
  assign o[32283] = i[32283];
  assign o[32282] = i[32282];
  assign o[32281] = i[32281];
  assign o[32280] = i[32280];
  assign o[32279] = i[32279];
  assign o[32278] = i[32278];
  assign o[32277] = i[32277];
  assign o[32276] = i[32276];
  assign o[32275] = i[32275];
  assign o[32274] = i[32274];
  assign o[32273] = i[32273];
  assign o[32272] = i[32272];
  assign o[32271] = i[32271];
  assign o[32270] = i[32270];
  assign o[32269] = i[32269];
  assign o[32268] = i[32268];
  assign o[32267] = i[32267];
  assign o[32266] = i[32266];
  assign o[32265] = i[32265];
  assign o[32264] = i[32264];
  assign o[32263] = i[32263];
  assign o[32262] = i[32262];
  assign o[32261] = i[32261];
  assign o[32260] = i[32260];
  assign o[32259] = i[32259];
  assign o[32258] = i[32258];
  assign o[32257] = i[32257];
  assign o[32256] = i[32256];
  assign o[32255] = i[32255];
  assign o[32254] = i[32254];
  assign o[32253] = i[32253];
  assign o[32252] = i[32252];
  assign o[32251] = i[32251];
  assign o[32250] = i[32250];
  assign o[32249] = i[32249];
  assign o[32248] = i[32248];
  assign o[32247] = i[32247];
  assign o[32246] = i[32246];
  assign o[32245] = i[32245];
  assign o[32244] = i[32244];
  assign o[32243] = i[32243];
  assign o[32242] = i[32242];
  assign o[32241] = i[32241];
  assign o[32240] = i[32240];
  assign o[32239] = i[32239];
  assign o[32238] = i[32238];
  assign o[32237] = i[32237];
  assign o[32236] = i[32236];
  assign o[32235] = i[32235];
  assign o[32234] = i[32234];
  assign o[32233] = i[32233];
  assign o[32232] = i[32232];
  assign o[32231] = i[32231];
  assign o[32230] = i[32230];
  assign o[32229] = i[32229];
  assign o[32228] = i[32228];
  assign o[32227] = i[32227];
  assign o[32226] = i[32226];
  assign o[32225] = i[32225];
  assign o[32224] = i[32224];
  assign o[32223] = i[32223];
  assign o[32222] = i[32222];
  assign o[32221] = i[32221];
  assign o[32220] = i[32220];
  assign o[32219] = i[32219];
  assign o[32218] = i[32218];
  assign o[32217] = i[32217];
  assign o[32216] = i[32216];
  assign o[32215] = i[32215];
  assign o[32214] = i[32214];
  assign o[32213] = i[32213];
  assign o[32212] = i[32212];
  assign o[32211] = i[32211];
  assign o[32210] = i[32210];
  assign o[32209] = i[32209];
  assign o[32208] = i[32208];
  assign o[32207] = i[32207];
  assign o[32206] = i[32206];
  assign o[32205] = i[32205];
  assign o[32204] = i[32204];
  assign o[32203] = i[32203];
  assign o[32202] = i[32202];
  assign o[32201] = i[32201];
  assign o[32200] = i[32200];
  assign o[32199] = i[32199];
  assign o[32198] = i[32198];
  assign o[32197] = i[32197];
  assign o[32196] = i[32196];
  assign o[32195] = i[32195];
  assign o[32194] = i[32194];
  assign o[32193] = i[32193];
  assign o[32192] = i[32192];
  assign o[32191] = i[32191];
  assign o[32190] = i[32190];
  assign o[32189] = i[32189];
  assign o[32188] = i[32188];
  assign o[32187] = i[32187];
  assign o[32186] = i[32186];
  assign o[32185] = i[32185];
  assign o[32184] = i[32184];
  assign o[32183] = i[32183];
  assign o[32182] = i[32182];
  assign o[32181] = i[32181];
  assign o[32180] = i[32180];
  assign o[32179] = i[32179];
  assign o[32178] = i[32178];
  assign o[32177] = i[32177];
  assign o[32176] = i[32176];
  assign o[32175] = i[32175];
  assign o[32174] = i[32174];
  assign o[32173] = i[32173];
  assign o[32172] = i[32172];
  assign o[32171] = i[32171];
  assign o[32170] = i[32170];
  assign o[32169] = i[32169];
  assign o[32168] = i[32168];
  assign o[32167] = i[32167];
  assign o[32166] = i[32166];
  assign o[32165] = i[32165];
  assign o[32164] = i[32164];
  assign o[32163] = i[32163];
  assign o[32162] = i[32162];
  assign o[32161] = i[32161];
  assign o[32160] = i[32160];
  assign o[32159] = i[32159];
  assign o[32158] = i[32158];
  assign o[32157] = i[32157];
  assign o[32156] = i[32156];
  assign o[32155] = i[32155];
  assign o[32154] = i[32154];
  assign o[32153] = i[32153];
  assign o[32152] = i[32152];
  assign o[32151] = i[32151];
  assign o[32150] = i[32150];
  assign o[32149] = i[32149];
  assign o[32148] = i[32148];
  assign o[32147] = i[32147];
  assign o[32146] = i[32146];
  assign o[32145] = i[32145];
  assign o[32144] = i[32144];
  assign o[32143] = i[32143];
  assign o[32142] = i[32142];
  assign o[32141] = i[32141];
  assign o[32140] = i[32140];
  assign o[32139] = i[32139];
  assign o[32138] = i[32138];
  assign o[32137] = i[32137];
  assign o[32136] = i[32136];
  assign o[32135] = i[32135];
  assign o[32134] = i[32134];
  assign o[32133] = i[32133];
  assign o[32132] = i[32132];
  assign o[32131] = i[32131];
  assign o[32130] = i[32130];
  assign o[32129] = i[32129];
  assign o[32128] = i[32128];
  assign o[32127] = i[32127];
  assign o[32126] = i[32126];
  assign o[32125] = i[32125];
  assign o[32124] = i[32124];
  assign o[32123] = i[32123];
  assign o[32122] = i[32122];
  assign o[32121] = i[32121];
  assign o[32120] = i[32120];
  assign o[32119] = i[32119];
  assign o[32118] = i[32118];
  assign o[32117] = i[32117];
  assign o[32116] = i[32116];
  assign o[32115] = i[32115];
  assign o[32114] = i[32114];
  assign o[32113] = i[32113];
  assign o[32112] = i[32112];
  assign o[32111] = i[32111];
  assign o[32110] = i[32110];
  assign o[32109] = i[32109];
  assign o[32108] = i[32108];
  assign o[32107] = i[32107];
  assign o[32106] = i[32106];
  assign o[32105] = i[32105];
  assign o[32104] = i[32104];
  assign o[32103] = i[32103];
  assign o[32102] = i[32102];
  assign o[32101] = i[32101];
  assign o[32100] = i[32100];
  assign o[32099] = i[32099];
  assign o[32098] = i[32098];
  assign o[32097] = i[32097];
  assign o[32096] = i[32096];
  assign o[32095] = i[32095];
  assign o[32094] = i[32094];
  assign o[32093] = i[32093];
  assign o[32092] = i[32092];
  assign o[32091] = i[32091];
  assign o[32090] = i[32090];
  assign o[32089] = i[32089];
  assign o[32088] = i[32088];
  assign o[32087] = i[32087];
  assign o[32086] = i[32086];
  assign o[32085] = i[32085];
  assign o[32084] = i[32084];
  assign o[32083] = i[32083];
  assign o[32082] = i[32082];
  assign o[32081] = i[32081];
  assign o[32080] = i[32080];
  assign o[32079] = i[32079];
  assign o[32078] = i[32078];
  assign o[32077] = i[32077];
  assign o[32076] = i[32076];
  assign o[32075] = i[32075];
  assign o[32074] = i[32074];
  assign o[32073] = i[32073];
  assign o[32072] = i[32072];
  assign o[32071] = i[32071];
  assign o[32070] = i[32070];
  assign o[32069] = i[32069];
  assign o[32068] = i[32068];
  assign o[32067] = i[32067];
  assign o[32066] = i[32066];
  assign o[32065] = i[32065];
  assign o[32064] = i[32064];
  assign o[32063] = i[32063];
  assign o[32062] = i[32062];
  assign o[32061] = i[32061];
  assign o[32060] = i[32060];
  assign o[32059] = i[32059];
  assign o[32058] = i[32058];
  assign o[32057] = i[32057];
  assign o[32056] = i[32056];
  assign o[32055] = i[32055];
  assign o[32054] = i[32054];
  assign o[32053] = i[32053];
  assign o[32052] = i[32052];
  assign o[32051] = i[32051];
  assign o[32050] = i[32050];
  assign o[32049] = i[32049];
  assign o[32048] = i[32048];
  assign o[32047] = i[32047];
  assign o[32046] = i[32046];
  assign o[32045] = i[32045];
  assign o[32044] = i[32044];
  assign o[32043] = i[32043];
  assign o[32042] = i[32042];
  assign o[32041] = i[32041];
  assign o[32040] = i[32040];
  assign o[32039] = i[32039];
  assign o[32038] = i[32038];
  assign o[32037] = i[32037];
  assign o[32036] = i[32036];
  assign o[32035] = i[32035];
  assign o[32034] = i[32034];
  assign o[32033] = i[32033];
  assign o[32032] = i[32032];
  assign o[32031] = i[32031];
  assign o[32030] = i[32030];
  assign o[32029] = i[32029];
  assign o[32028] = i[32028];
  assign o[32027] = i[32027];
  assign o[32026] = i[32026];
  assign o[32025] = i[32025];
  assign o[32024] = i[32024];
  assign o[32023] = i[32023];
  assign o[32022] = i[32022];
  assign o[32021] = i[32021];
  assign o[32020] = i[32020];
  assign o[32019] = i[32019];
  assign o[32018] = i[32018];
  assign o[32017] = i[32017];
  assign o[32016] = i[32016];
  assign o[32015] = i[32015];
  assign o[32014] = i[32014];
  assign o[32013] = i[32013];
  assign o[32012] = i[32012];
  assign o[32011] = i[32011];
  assign o[32010] = i[32010];
  assign o[32009] = i[32009];
  assign o[32008] = i[32008];
  assign o[32007] = i[32007];
  assign o[32006] = i[32006];
  assign o[32005] = i[32005];
  assign o[32004] = i[32004];
  assign o[32003] = i[32003];
  assign o[32002] = i[32002];
  assign o[32001] = i[32001];
  assign o[32000] = i[32000];
  assign o[31999] = i[31999];
  assign o[31998] = i[31998];
  assign o[31997] = i[31997];
  assign o[31996] = i[31996];
  assign o[31995] = i[31995];
  assign o[31994] = i[31994];
  assign o[31993] = i[31993];
  assign o[31992] = i[31992];
  assign o[31991] = i[31991];
  assign o[31990] = i[31990];
  assign o[31989] = i[31989];
  assign o[31988] = i[31988];
  assign o[31987] = i[31987];
  assign o[31986] = i[31986];
  assign o[31985] = i[31985];
  assign o[31984] = i[31984];
  assign o[31983] = i[31983];
  assign o[31982] = i[31982];
  assign o[31981] = i[31981];
  assign o[31980] = i[31980];
  assign o[31979] = i[31979];
  assign o[31978] = i[31978];
  assign o[31977] = i[31977];
  assign o[31976] = i[31976];
  assign o[31975] = i[31975];
  assign o[31974] = i[31974];
  assign o[31973] = i[31973];
  assign o[31972] = i[31972];
  assign o[31971] = i[31971];
  assign o[31970] = i[31970];
  assign o[31969] = i[31969];
  assign o[31968] = i[31968];
  assign o[31967] = i[31967];
  assign o[31966] = i[31966];
  assign o[31965] = i[31965];
  assign o[31964] = i[31964];
  assign o[31963] = i[31963];
  assign o[31962] = i[31962];
  assign o[31961] = i[31961];
  assign o[31960] = i[31960];
  assign o[31959] = i[31959];
  assign o[31958] = i[31958];
  assign o[31957] = i[31957];
  assign o[31956] = i[31956];
  assign o[31955] = i[31955];
  assign o[31954] = i[31954];
  assign o[31953] = i[31953];
  assign o[31952] = i[31952];
  assign o[31951] = i[31951];
  assign o[31950] = i[31950];
  assign o[31949] = i[31949];
  assign o[31948] = i[31948];
  assign o[31947] = i[31947];
  assign o[31946] = i[31946];
  assign o[31945] = i[31945];
  assign o[31944] = i[31944];
  assign o[31943] = i[31943];
  assign o[31942] = i[31942];
  assign o[31941] = i[31941];
  assign o[31940] = i[31940];
  assign o[31939] = i[31939];
  assign o[31938] = i[31938];
  assign o[31937] = i[31937];
  assign o[31936] = i[31936];
  assign o[31935] = i[31935];
  assign o[31934] = i[31934];
  assign o[31933] = i[31933];
  assign o[31932] = i[31932];
  assign o[31931] = i[31931];
  assign o[31930] = i[31930];
  assign o[31929] = i[31929];
  assign o[31928] = i[31928];
  assign o[31927] = i[31927];
  assign o[31926] = i[31926];
  assign o[31925] = i[31925];
  assign o[31924] = i[31924];
  assign o[31923] = i[31923];
  assign o[31922] = i[31922];
  assign o[31921] = i[31921];
  assign o[31920] = i[31920];
  assign o[31919] = i[31919];
  assign o[31918] = i[31918];
  assign o[31917] = i[31917];
  assign o[31916] = i[31916];
  assign o[31915] = i[31915];
  assign o[31914] = i[31914];
  assign o[31913] = i[31913];
  assign o[31912] = i[31912];
  assign o[31911] = i[31911];
  assign o[31910] = i[31910];
  assign o[31909] = i[31909];
  assign o[31908] = i[31908];
  assign o[31907] = i[31907];
  assign o[31906] = i[31906];
  assign o[31905] = i[31905];
  assign o[31904] = i[31904];
  assign o[31903] = i[31903];
  assign o[31902] = i[31902];
  assign o[31901] = i[31901];
  assign o[31900] = i[31900];
  assign o[31899] = i[31899];
  assign o[31898] = i[31898];
  assign o[31897] = i[31897];
  assign o[31896] = i[31896];
  assign o[31895] = i[31895];
  assign o[31894] = i[31894];
  assign o[31893] = i[31893];
  assign o[31892] = i[31892];
  assign o[31891] = i[31891];
  assign o[31890] = i[31890];
  assign o[31889] = i[31889];
  assign o[31888] = i[31888];
  assign o[31887] = i[31887];
  assign o[31886] = i[31886];
  assign o[31885] = i[31885];
  assign o[31884] = i[31884];
  assign o[31883] = i[31883];
  assign o[31882] = i[31882];
  assign o[31881] = i[31881];
  assign o[31880] = i[31880];
  assign o[31879] = i[31879];
  assign o[31878] = i[31878];
  assign o[31877] = i[31877];
  assign o[31876] = i[31876];
  assign o[31875] = i[31875];
  assign o[31874] = i[31874];
  assign o[31873] = i[31873];
  assign o[31872] = i[31872];
  assign o[31871] = i[31871];
  assign o[31870] = i[31870];
  assign o[31869] = i[31869];
  assign o[31868] = i[31868];
  assign o[31867] = i[31867];
  assign o[31866] = i[31866];
  assign o[31865] = i[31865];
  assign o[31864] = i[31864];
  assign o[31863] = i[31863];
  assign o[31862] = i[31862];
  assign o[31861] = i[31861];
  assign o[31860] = i[31860];
  assign o[31859] = i[31859];
  assign o[31858] = i[31858];
  assign o[31857] = i[31857];
  assign o[31856] = i[31856];
  assign o[31855] = i[31855];
  assign o[31854] = i[31854];
  assign o[31853] = i[31853];
  assign o[31852] = i[31852];
  assign o[31851] = i[31851];
  assign o[31850] = i[31850];
  assign o[31849] = i[31849];
  assign o[31848] = i[31848];
  assign o[31847] = i[31847];
  assign o[31846] = i[31846];
  assign o[31845] = i[31845];
  assign o[31844] = i[31844];
  assign o[31843] = i[31843];
  assign o[31842] = i[31842];
  assign o[31841] = i[31841];
  assign o[31840] = i[31840];
  assign o[31839] = i[31839];
  assign o[31838] = i[31838];
  assign o[31837] = i[31837];
  assign o[31836] = i[31836];
  assign o[31835] = i[31835];
  assign o[31834] = i[31834];
  assign o[31833] = i[31833];
  assign o[31832] = i[31832];
  assign o[31831] = i[31831];
  assign o[31830] = i[31830];
  assign o[31829] = i[31829];
  assign o[31828] = i[31828];
  assign o[31827] = i[31827];
  assign o[31826] = i[31826];
  assign o[31825] = i[31825];
  assign o[31824] = i[31824];
  assign o[31823] = i[31823];
  assign o[31822] = i[31822];
  assign o[31821] = i[31821];
  assign o[31820] = i[31820];
  assign o[31819] = i[31819];
  assign o[31818] = i[31818];
  assign o[31817] = i[31817];
  assign o[31816] = i[31816];
  assign o[31815] = i[31815];
  assign o[31814] = i[31814];
  assign o[31813] = i[31813];
  assign o[31812] = i[31812];
  assign o[31811] = i[31811];
  assign o[31810] = i[31810];
  assign o[31809] = i[31809];
  assign o[31808] = i[31808];
  assign o[31807] = i[31807];
  assign o[31806] = i[31806];
  assign o[31805] = i[31805];
  assign o[31804] = i[31804];
  assign o[31803] = i[31803];
  assign o[31802] = i[31802];
  assign o[31801] = i[31801];
  assign o[31800] = i[31800];
  assign o[31799] = i[31799];
  assign o[31798] = i[31798];
  assign o[31797] = i[31797];
  assign o[31796] = i[31796];
  assign o[31795] = i[31795];
  assign o[31794] = i[31794];
  assign o[31793] = i[31793];
  assign o[31792] = i[31792];
  assign o[31791] = i[31791];
  assign o[31790] = i[31790];
  assign o[31789] = i[31789];
  assign o[31788] = i[31788];
  assign o[31787] = i[31787];
  assign o[31786] = i[31786];
  assign o[31785] = i[31785];
  assign o[31784] = i[31784];
  assign o[31783] = i[31783];
  assign o[31782] = i[31782];
  assign o[31781] = i[31781];
  assign o[31780] = i[31780];
  assign o[31779] = i[31779];
  assign o[31778] = i[31778];
  assign o[31777] = i[31777];
  assign o[31776] = i[31776];
  assign o[31775] = i[31775];
  assign o[31774] = i[31774];
  assign o[31773] = i[31773];
  assign o[31772] = i[31772];
  assign o[31771] = i[31771];
  assign o[31770] = i[31770];
  assign o[31769] = i[31769];
  assign o[31768] = i[31768];
  assign o[31767] = i[31767];
  assign o[31766] = i[31766];
  assign o[31765] = i[31765];
  assign o[31764] = i[31764];
  assign o[31763] = i[31763];
  assign o[31762] = i[31762];
  assign o[31761] = i[31761];
  assign o[31760] = i[31760];
  assign o[31759] = i[31759];
  assign o[31758] = i[31758];
  assign o[31757] = i[31757];
  assign o[31756] = i[31756];
  assign o[31755] = i[31755];
  assign o[31754] = i[31754];
  assign o[31753] = i[31753];
  assign o[31752] = i[31752];
  assign o[31751] = i[31751];
  assign o[31750] = i[31750];
  assign o[31749] = i[31749];
  assign o[31748] = i[31748];
  assign o[31747] = i[31747];
  assign o[31746] = i[31746];
  assign o[31745] = i[31745];
  assign o[31744] = i[31744];
  assign o[31743] = i[31743];
  assign o[31742] = i[31742];
  assign o[31741] = i[31741];
  assign o[31740] = i[31740];
  assign o[31739] = i[31739];
  assign o[31738] = i[31738];
  assign o[31737] = i[31737];
  assign o[31736] = i[31736];
  assign o[31735] = i[31735];
  assign o[31734] = i[31734];
  assign o[31733] = i[31733];
  assign o[31732] = i[31732];
  assign o[31731] = i[31731];
  assign o[31730] = i[31730];
  assign o[31729] = i[31729];
  assign o[31728] = i[31728];
  assign o[31727] = i[31727];
  assign o[31726] = i[31726];
  assign o[31725] = i[31725];
  assign o[31724] = i[31724];
  assign o[31723] = i[31723];
  assign o[31722] = i[31722];
  assign o[31721] = i[31721];
  assign o[31720] = i[31720];
  assign o[31719] = i[31719];
  assign o[31718] = i[31718];
  assign o[31717] = i[31717];
  assign o[31716] = i[31716];
  assign o[31715] = i[31715];
  assign o[31714] = i[31714];
  assign o[31713] = i[31713];
  assign o[31712] = i[31712];
  assign o[31711] = i[31711];
  assign o[31710] = i[31710];
  assign o[31709] = i[31709];
  assign o[31708] = i[31708];
  assign o[31707] = i[31707];
  assign o[31706] = i[31706];
  assign o[31705] = i[31705];
  assign o[31704] = i[31704];
  assign o[31703] = i[31703];
  assign o[31702] = i[31702];
  assign o[31701] = i[31701];
  assign o[31700] = i[31700];
  assign o[31699] = i[31699];
  assign o[31698] = i[31698];
  assign o[31697] = i[31697];
  assign o[31696] = i[31696];
  assign o[31695] = i[31695];
  assign o[31694] = i[31694];
  assign o[31693] = i[31693];
  assign o[31692] = i[31692];
  assign o[31691] = i[31691];
  assign o[31690] = i[31690];
  assign o[31689] = i[31689];
  assign o[31688] = i[31688];
  assign o[31687] = i[31687];
  assign o[31686] = i[31686];
  assign o[31685] = i[31685];
  assign o[31684] = i[31684];
  assign o[31683] = i[31683];
  assign o[31682] = i[31682];
  assign o[31681] = i[31681];
  assign o[31680] = i[31680];
  assign o[31679] = i[31679];
  assign o[31678] = i[31678];
  assign o[31677] = i[31677];
  assign o[31676] = i[31676];
  assign o[31675] = i[31675];
  assign o[31674] = i[31674];
  assign o[31673] = i[31673];
  assign o[31672] = i[31672];
  assign o[31671] = i[31671];
  assign o[31670] = i[31670];
  assign o[31669] = i[31669];
  assign o[31668] = i[31668];
  assign o[31667] = i[31667];
  assign o[31666] = i[31666];
  assign o[31665] = i[31665];
  assign o[31664] = i[31664];
  assign o[31663] = i[31663];
  assign o[31662] = i[31662];
  assign o[31661] = i[31661];
  assign o[31660] = i[31660];
  assign o[31659] = i[31659];
  assign o[31658] = i[31658];
  assign o[31657] = i[31657];
  assign o[31656] = i[31656];
  assign o[31655] = i[31655];
  assign o[31654] = i[31654];
  assign o[31653] = i[31653];
  assign o[31652] = i[31652];
  assign o[31651] = i[31651];
  assign o[31650] = i[31650];
  assign o[31649] = i[31649];
  assign o[31648] = i[31648];
  assign o[31647] = i[31647];
  assign o[31646] = i[31646];
  assign o[31645] = i[31645];
  assign o[31644] = i[31644];
  assign o[31643] = i[31643];
  assign o[31642] = i[31642];
  assign o[31641] = i[31641];
  assign o[31640] = i[31640];
  assign o[31639] = i[31639];
  assign o[31638] = i[31638];
  assign o[31637] = i[31637];
  assign o[31636] = i[31636];
  assign o[31635] = i[31635];
  assign o[31634] = i[31634];
  assign o[31633] = i[31633];
  assign o[31632] = i[31632];
  assign o[31631] = i[31631];
  assign o[31630] = i[31630];
  assign o[31629] = i[31629];
  assign o[31628] = i[31628];
  assign o[31627] = i[31627];
  assign o[31626] = i[31626];
  assign o[31625] = i[31625];
  assign o[31624] = i[31624];
  assign o[31623] = i[31623];
  assign o[31622] = i[31622];
  assign o[31621] = i[31621];
  assign o[31620] = i[31620];
  assign o[31619] = i[31619];
  assign o[31618] = i[31618];
  assign o[31617] = i[31617];
  assign o[31616] = i[31616];
  assign o[31615] = i[31615];
  assign o[31614] = i[31614];
  assign o[31613] = i[31613];
  assign o[31612] = i[31612];
  assign o[31611] = i[31611];
  assign o[31610] = i[31610];
  assign o[31609] = i[31609];
  assign o[31608] = i[31608];
  assign o[31607] = i[31607];
  assign o[31606] = i[31606];
  assign o[31605] = i[31605];
  assign o[31604] = i[31604];
  assign o[31603] = i[31603];
  assign o[31602] = i[31602];
  assign o[31601] = i[31601];
  assign o[31600] = i[31600];
  assign o[31599] = i[31599];
  assign o[31598] = i[31598];
  assign o[31597] = i[31597];
  assign o[31596] = i[31596];
  assign o[31595] = i[31595];
  assign o[31594] = i[31594];
  assign o[31593] = i[31593];
  assign o[31592] = i[31592];
  assign o[31591] = i[31591];
  assign o[31590] = i[31590];
  assign o[31589] = i[31589];
  assign o[31588] = i[31588];
  assign o[31587] = i[31587];
  assign o[31586] = i[31586];
  assign o[31585] = i[31585];
  assign o[31584] = i[31584];
  assign o[31583] = i[31583];
  assign o[31582] = i[31582];
  assign o[31581] = i[31581];
  assign o[31580] = i[31580];
  assign o[31579] = i[31579];
  assign o[31578] = i[31578];
  assign o[31577] = i[31577];
  assign o[31576] = i[31576];
  assign o[31575] = i[31575];
  assign o[31574] = i[31574];
  assign o[31573] = i[31573];
  assign o[31572] = i[31572];
  assign o[31571] = i[31571];
  assign o[31570] = i[31570];
  assign o[31569] = i[31569];
  assign o[31568] = i[31568];
  assign o[31567] = i[31567];
  assign o[31566] = i[31566];
  assign o[31565] = i[31565];
  assign o[31564] = i[31564];
  assign o[31563] = i[31563];
  assign o[31562] = i[31562];
  assign o[31561] = i[31561];
  assign o[31560] = i[31560];
  assign o[31559] = i[31559];
  assign o[31558] = i[31558];
  assign o[31557] = i[31557];
  assign o[31556] = i[31556];
  assign o[31555] = i[31555];
  assign o[31554] = i[31554];
  assign o[31553] = i[31553];
  assign o[31552] = i[31552];
  assign o[31551] = i[31551];
  assign o[31550] = i[31550];
  assign o[31549] = i[31549];
  assign o[31548] = i[31548];
  assign o[31547] = i[31547];
  assign o[31546] = i[31546];
  assign o[31545] = i[31545];
  assign o[31544] = i[31544];
  assign o[31543] = i[31543];
  assign o[31542] = i[31542];
  assign o[31541] = i[31541];
  assign o[31540] = i[31540];
  assign o[31539] = i[31539];
  assign o[31538] = i[31538];
  assign o[31537] = i[31537];
  assign o[31536] = i[31536];
  assign o[31535] = i[31535];
  assign o[31534] = i[31534];
  assign o[31533] = i[31533];
  assign o[31532] = i[31532];
  assign o[31531] = i[31531];
  assign o[31530] = i[31530];
  assign o[31529] = i[31529];
  assign o[31528] = i[31528];
  assign o[31527] = i[31527];
  assign o[31526] = i[31526];
  assign o[31525] = i[31525];
  assign o[31524] = i[31524];
  assign o[31523] = i[31523];
  assign o[31522] = i[31522];
  assign o[31521] = i[31521];
  assign o[31520] = i[31520];
  assign o[31519] = i[31519];
  assign o[31518] = i[31518];
  assign o[31517] = i[31517];
  assign o[31516] = i[31516];
  assign o[31515] = i[31515];
  assign o[31514] = i[31514];
  assign o[31513] = i[31513];
  assign o[31512] = i[31512];
  assign o[31511] = i[31511];
  assign o[31510] = i[31510];
  assign o[31509] = i[31509];
  assign o[31508] = i[31508];
  assign o[31507] = i[31507];
  assign o[31506] = i[31506];
  assign o[31505] = i[31505];
  assign o[31504] = i[31504];
  assign o[31503] = i[31503];
  assign o[31502] = i[31502];
  assign o[31501] = i[31501];
  assign o[31500] = i[31500];
  assign o[31499] = i[31499];
  assign o[31498] = i[31498];
  assign o[31497] = i[31497];
  assign o[31496] = i[31496];
  assign o[31495] = i[31495];
  assign o[31494] = i[31494];
  assign o[31493] = i[31493];
  assign o[31492] = i[31492];
  assign o[31491] = i[31491];
  assign o[31490] = i[31490];
  assign o[31489] = i[31489];
  assign o[31488] = i[31488];
  assign o[31487] = i[31487];
  assign o[31486] = i[31486];
  assign o[31485] = i[31485];
  assign o[31484] = i[31484];
  assign o[31483] = i[31483];
  assign o[31482] = i[31482];
  assign o[31481] = i[31481];
  assign o[31480] = i[31480];
  assign o[31479] = i[31479];
  assign o[31478] = i[31478];
  assign o[31477] = i[31477];
  assign o[31476] = i[31476];
  assign o[31475] = i[31475];
  assign o[31474] = i[31474];
  assign o[31473] = i[31473];
  assign o[31472] = i[31472];
  assign o[31471] = i[31471];
  assign o[31470] = i[31470];
  assign o[31469] = i[31469];
  assign o[31468] = i[31468];
  assign o[31467] = i[31467];
  assign o[31466] = i[31466];
  assign o[31465] = i[31465];
  assign o[31464] = i[31464];
  assign o[31463] = i[31463];
  assign o[31462] = i[31462];
  assign o[31461] = i[31461];
  assign o[31460] = i[31460];
  assign o[31459] = i[31459];
  assign o[31458] = i[31458];
  assign o[31457] = i[31457];
  assign o[31456] = i[31456];
  assign o[31455] = i[31455];
  assign o[31454] = i[31454];
  assign o[31453] = i[31453];
  assign o[31452] = i[31452];
  assign o[31451] = i[31451];
  assign o[31450] = i[31450];
  assign o[31449] = i[31449];
  assign o[31448] = i[31448];
  assign o[31447] = i[31447];
  assign o[31446] = i[31446];
  assign o[31445] = i[31445];
  assign o[31444] = i[31444];
  assign o[31443] = i[31443];
  assign o[31442] = i[31442];
  assign o[31441] = i[31441];
  assign o[31440] = i[31440];
  assign o[31439] = i[31439];
  assign o[31438] = i[31438];
  assign o[31437] = i[31437];
  assign o[31436] = i[31436];
  assign o[31435] = i[31435];
  assign o[31434] = i[31434];
  assign o[31433] = i[31433];
  assign o[31432] = i[31432];
  assign o[31431] = i[31431];
  assign o[31430] = i[31430];
  assign o[31429] = i[31429];
  assign o[31428] = i[31428];
  assign o[31427] = i[31427];
  assign o[31426] = i[31426];
  assign o[31425] = i[31425];
  assign o[31424] = i[31424];
  assign o[31423] = i[31423];
  assign o[31422] = i[31422];
  assign o[31421] = i[31421];
  assign o[31420] = i[31420];
  assign o[31419] = i[31419];
  assign o[31418] = i[31418];
  assign o[31417] = i[31417];
  assign o[31416] = i[31416];
  assign o[31415] = i[31415];
  assign o[31414] = i[31414];
  assign o[31413] = i[31413];
  assign o[31412] = i[31412];
  assign o[31411] = i[31411];
  assign o[31410] = i[31410];
  assign o[31409] = i[31409];
  assign o[31408] = i[31408];
  assign o[31407] = i[31407];
  assign o[31406] = i[31406];
  assign o[31405] = i[31405];
  assign o[31404] = i[31404];
  assign o[31403] = i[31403];
  assign o[31402] = i[31402];
  assign o[31401] = i[31401];
  assign o[31400] = i[31400];
  assign o[31399] = i[31399];
  assign o[31398] = i[31398];
  assign o[31397] = i[31397];
  assign o[31396] = i[31396];
  assign o[31395] = i[31395];
  assign o[31394] = i[31394];
  assign o[31393] = i[31393];
  assign o[31392] = i[31392];
  assign o[31391] = i[31391];
  assign o[31390] = i[31390];
  assign o[31389] = i[31389];
  assign o[31388] = i[31388];
  assign o[31387] = i[31387];
  assign o[31386] = i[31386];
  assign o[31385] = i[31385];
  assign o[31384] = i[31384];
  assign o[31383] = i[31383];
  assign o[31382] = i[31382];
  assign o[31381] = i[31381];
  assign o[31380] = i[31380];
  assign o[31379] = i[31379];
  assign o[31378] = i[31378];
  assign o[31377] = i[31377];
  assign o[31376] = i[31376];
  assign o[31375] = i[31375];
  assign o[31374] = i[31374];
  assign o[31373] = i[31373];
  assign o[31372] = i[31372];
  assign o[31371] = i[31371];
  assign o[31370] = i[31370];
  assign o[31369] = i[31369];
  assign o[31368] = i[31368];
  assign o[31367] = i[31367];
  assign o[31366] = i[31366];
  assign o[31365] = i[31365];
  assign o[31364] = i[31364];
  assign o[31363] = i[31363];
  assign o[31362] = i[31362];
  assign o[31361] = i[31361];
  assign o[31360] = i[31360];
  assign o[31359] = i[31359];
  assign o[31358] = i[31358];
  assign o[31357] = i[31357];
  assign o[31356] = i[31356];
  assign o[31355] = i[31355];
  assign o[31354] = i[31354];
  assign o[31353] = i[31353];
  assign o[31352] = i[31352];
  assign o[31351] = i[31351];
  assign o[31350] = i[31350];
  assign o[31349] = i[31349];
  assign o[31348] = i[31348];
  assign o[31347] = i[31347];
  assign o[31346] = i[31346];
  assign o[31345] = i[31345];
  assign o[31344] = i[31344];
  assign o[31343] = i[31343];
  assign o[31342] = i[31342];
  assign o[31341] = i[31341];
  assign o[31340] = i[31340];
  assign o[31339] = i[31339];
  assign o[31338] = i[31338];
  assign o[31337] = i[31337];
  assign o[31336] = i[31336];
  assign o[31335] = i[31335];
  assign o[31334] = i[31334];
  assign o[31333] = i[31333];
  assign o[31332] = i[31332];
  assign o[31331] = i[31331];
  assign o[31330] = i[31330];
  assign o[31329] = i[31329];
  assign o[31328] = i[31328];
  assign o[31327] = i[31327];
  assign o[31326] = i[31326];
  assign o[31325] = i[31325];
  assign o[31324] = i[31324];
  assign o[31323] = i[31323];
  assign o[31322] = i[31322];
  assign o[31321] = i[31321];
  assign o[31320] = i[31320];
  assign o[31319] = i[31319];
  assign o[31318] = i[31318];
  assign o[31317] = i[31317];
  assign o[31316] = i[31316];
  assign o[31315] = i[31315];
  assign o[31314] = i[31314];
  assign o[31313] = i[31313];
  assign o[31312] = i[31312];
  assign o[31311] = i[31311];
  assign o[31310] = i[31310];
  assign o[31309] = i[31309];
  assign o[31308] = i[31308];
  assign o[31307] = i[31307];
  assign o[31306] = i[31306];
  assign o[31305] = i[31305];
  assign o[31304] = i[31304];
  assign o[31303] = i[31303];
  assign o[31302] = i[31302];
  assign o[31301] = i[31301];
  assign o[31300] = i[31300];
  assign o[31299] = i[31299];
  assign o[31298] = i[31298];
  assign o[31297] = i[31297];
  assign o[31296] = i[31296];
  assign o[31295] = i[31295];
  assign o[31294] = i[31294];
  assign o[31293] = i[31293];
  assign o[31292] = i[31292];
  assign o[31291] = i[31291];
  assign o[31290] = i[31290];
  assign o[31289] = i[31289];
  assign o[31288] = i[31288];
  assign o[31287] = i[31287];
  assign o[31286] = i[31286];
  assign o[31285] = i[31285];
  assign o[31284] = i[31284];
  assign o[31283] = i[31283];
  assign o[31282] = i[31282];
  assign o[31281] = i[31281];
  assign o[31280] = i[31280];
  assign o[31279] = i[31279];
  assign o[31278] = i[31278];
  assign o[31277] = i[31277];
  assign o[31276] = i[31276];
  assign o[31275] = i[31275];
  assign o[31274] = i[31274];
  assign o[31273] = i[31273];
  assign o[31272] = i[31272];
  assign o[31271] = i[31271];
  assign o[31270] = i[31270];
  assign o[31269] = i[31269];
  assign o[31268] = i[31268];
  assign o[31267] = i[31267];
  assign o[31266] = i[31266];
  assign o[31265] = i[31265];
  assign o[31264] = i[31264];
  assign o[31263] = i[31263];
  assign o[31262] = i[31262];
  assign o[31261] = i[31261];
  assign o[31260] = i[31260];
  assign o[31259] = i[31259];
  assign o[31258] = i[31258];
  assign o[31257] = i[31257];
  assign o[31256] = i[31256];
  assign o[31255] = i[31255];
  assign o[31254] = i[31254];
  assign o[31253] = i[31253];
  assign o[31252] = i[31252];
  assign o[31251] = i[31251];
  assign o[31250] = i[31250];
  assign o[31249] = i[31249];
  assign o[31248] = i[31248];
  assign o[31247] = i[31247];
  assign o[31246] = i[31246];
  assign o[31245] = i[31245];
  assign o[31244] = i[31244];
  assign o[31243] = i[31243];
  assign o[31242] = i[31242];
  assign o[31241] = i[31241];
  assign o[31240] = i[31240];
  assign o[31239] = i[31239];
  assign o[31238] = i[31238];
  assign o[31237] = i[31237];
  assign o[31236] = i[31236];
  assign o[31235] = i[31235];
  assign o[31234] = i[31234];
  assign o[31233] = i[31233];
  assign o[31232] = i[31232];
  assign o[31231] = i[31231];
  assign o[31230] = i[31230];
  assign o[31229] = i[31229];
  assign o[31228] = i[31228];
  assign o[31227] = i[31227];
  assign o[31226] = i[31226];
  assign o[31225] = i[31225];
  assign o[31224] = i[31224];
  assign o[31223] = i[31223];
  assign o[31222] = i[31222];
  assign o[31221] = i[31221];
  assign o[31220] = i[31220];
  assign o[31219] = i[31219];
  assign o[31218] = i[31218];
  assign o[31217] = i[31217];
  assign o[31216] = i[31216];
  assign o[31215] = i[31215];
  assign o[31214] = i[31214];
  assign o[31213] = i[31213];
  assign o[31212] = i[31212];
  assign o[31211] = i[31211];
  assign o[31210] = i[31210];
  assign o[31209] = i[31209];
  assign o[31208] = i[31208];
  assign o[31207] = i[31207];
  assign o[31206] = i[31206];
  assign o[31205] = i[31205];
  assign o[31204] = i[31204];
  assign o[31203] = i[31203];
  assign o[31202] = i[31202];
  assign o[31201] = i[31201];
  assign o[31200] = i[31200];
  assign o[31199] = i[31199];
  assign o[31198] = i[31198];
  assign o[31197] = i[31197];
  assign o[31196] = i[31196];
  assign o[31195] = i[31195];
  assign o[31194] = i[31194];
  assign o[31193] = i[31193];
  assign o[31192] = i[31192];
  assign o[31191] = i[31191];
  assign o[31190] = i[31190];
  assign o[31189] = i[31189];
  assign o[31188] = i[31188];
  assign o[31187] = i[31187];
  assign o[31186] = i[31186];
  assign o[31185] = i[31185];
  assign o[31184] = i[31184];
  assign o[31183] = i[31183];
  assign o[31182] = i[31182];
  assign o[31181] = i[31181];
  assign o[31180] = i[31180];
  assign o[31179] = i[31179];
  assign o[31178] = i[31178];
  assign o[31177] = i[31177];
  assign o[31176] = i[31176];
  assign o[31175] = i[31175];
  assign o[31174] = i[31174];
  assign o[31173] = i[31173];
  assign o[31172] = i[31172];
  assign o[31171] = i[31171];
  assign o[31170] = i[31170];
  assign o[31169] = i[31169];
  assign o[31168] = i[31168];
  assign o[31167] = i[31167];
  assign o[31166] = i[31166];
  assign o[31165] = i[31165];
  assign o[31164] = i[31164];
  assign o[31163] = i[31163];
  assign o[31162] = i[31162];
  assign o[31161] = i[31161];
  assign o[31160] = i[31160];
  assign o[31159] = i[31159];
  assign o[31158] = i[31158];
  assign o[31157] = i[31157];
  assign o[31156] = i[31156];
  assign o[31155] = i[31155];
  assign o[31154] = i[31154];
  assign o[31153] = i[31153];
  assign o[31152] = i[31152];
  assign o[31151] = i[31151];
  assign o[31150] = i[31150];
  assign o[31149] = i[31149];
  assign o[31148] = i[31148];
  assign o[31147] = i[31147];
  assign o[31146] = i[31146];
  assign o[31145] = i[31145];
  assign o[31144] = i[31144];
  assign o[31143] = i[31143];
  assign o[31142] = i[31142];
  assign o[31141] = i[31141];
  assign o[31140] = i[31140];
  assign o[31139] = i[31139];
  assign o[31138] = i[31138];
  assign o[31137] = i[31137];
  assign o[31136] = i[31136];
  assign o[31135] = i[31135];
  assign o[31134] = i[31134];
  assign o[31133] = i[31133];
  assign o[31132] = i[31132];
  assign o[31131] = i[31131];
  assign o[31130] = i[31130];
  assign o[31129] = i[31129];
  assign o[31128] = i[31128];
  assign o[31127] = i[31127];
  assign o[31126] = i[31126];
  assign o[31125] = i[31125];
  assign o[31124] = i[31124];
  assign o[31123] = i[31123];
  assign o[31122] = i[31122];
  assign o[31121] = i[31121];
  assign o[31120] = i[31120];
  assign o[31119] = i[31119];
  assign o[31118] = i[31118];
  assign o[31117] = i[31117];
  assign o[31116] = i[31116];
  assign o[31115] = i[31115];
  assign o[31114] = i[31114];
  assign o[31113] = i[31113];
  assign o[31112] = i[31112];
  assign o[31111] = i[31111];
  assign o[31110] = i[31110];
  assign o[31109] = i[31109];
  assign o[31108] = i[31108];
  assign o[31107] = i[31107];
  assign o[31106] = i[31106];
  assign o[31105] = i[31105];
  assign o[31104] = i[31104];
  assign o[31103] = i[31103];
  assign o[31102] = i[31102];
  assign o[31101] = i[31101];
  assign o[31100] = i[31100];
  assign o[31099] = i[31099];
  assign o[31098] = i[31098];
  assign o[31097] = i[31097];
  assign o[31096] = i[31096];
  assign o[31095] = i[31095];
  assign o[31094] = i[31094];
  assign o[31093] = i[31093];
  assign o[31092] = i[31092];
  assign o[31091] = i[31091];
  assign o[31090] = i[31090];
  assign o[31089] = i[31089];
  assign o[31088] = i[31088];
  assign o[31087] = i[31087];
  assign o[31086] = i[31086];
  assign o[31085] = i[31085];
  assign o[31084] = i[31084];
  assign o[31083] = i[31083];
  assign o[31082] = i[31082];
  assign o[31081] = i[31081];
  assign o[31080] = i[31080];
  assign o[31079] = i[31079];
  assign o[31078] = i[31078];
  assign o[31077] = i[31077];
  assign o[31076] = i[31076];
  assign o[31075] = i[31075];
  assign o[31074] = i[31074];
  assign o[31073] = i[31073];
  assign o[31072] = i[31072];
  assign o[31071] = i[31071];
  assign o[31070] = i[31070];
  assign o[31069] = i[31069];
  assign o[31068] = i[31068];
  assign o[31067] = i[31067];
  assign o[31066] = i[31066];
  assign o[31065] = i[31065];
  assign o[31064] = i[31064];
  assign o[31063] = i[31063];
  assign o[31062] = i[31062];
  assign o[31061] = i[31061];
  assign o[31060] = i[31060];
  assign o[31059] = i[31059];
  assign o[31058] = i[31058];
  assign o[31057] = i[31057];
  assign o[31056] = i[31056];
  assign o[31055] = i[31055];
  assign o[31054] = i[31054];
  assign o[31053] = i[31053];
  assign o[31052] = i[31052];
  assign o[31051] = i[31051];
  assign o[31050] = i[31050];
  assign o[31049] = i[31049];
  assign o[31048] = i[31048];
  assign o[31047] = i[31047];
  assign o[31046] = i[31046];
  assign o[31045] = i[31045];
  assign o[31044] = i[31044];
  assign o[31043] = i[31043];
  assign o[31042] = i[31042];
  assign o[31041] = i[31041];
  assign o[31040] = i[31040];
  assign o[31039] = i[31039];
  assign o[31038] = i[31038];
  assign o[31037] = i[31037];
  assign o[31036] = i[31036];
  assign o[31035] = i[31035];
  assign o[31034] = i[31034];
  assign o[31033] = i[31033];
  assign o[31032] = i[31032];
  assign o[31031] = i[31031];
  assign o[31030] = i[31030];
  assign o[31029] = i[31029];
  assign o[31028] = i[31028];
  assign o[31027] = i[31027];
  assign o[31026] = i[31026];
  assign o[31025] = i[31025];
  assign o[31024] = i[31024];
  assign o[31023] = i[31023];
  assign o[31022] = i[31022];
  assign o[31021] = i[31021];
  assign o[31020] = i[31020];
  assign o[31019] = i[31019];
  assign o[31018] = i[31018];
  assign o[31017] = i[31017];
  assign o[31016] = i[31016];
  assign o[31015] = i[31015];
  assign o[31014] = i[31014];
  assign o[31013] = i[31013];
  assign o[31012] = i[31012];
  assign o[31011] = i[31011];
  assign o[31010] = i[31010];
  assign o[31009] = i[31009];
  assign o[31008] = i[31008];
  assign o[31007] = i[31007];
  assign o[31006] = i[31006];
  assign o[31005] = i[31005];
  assign o[31004] = i[31004];
  assign o[31003] = i[31003];
  assign o[31002] = i[31002];
  assign o[31001] = i[31001];
  assign o[31000] = i[31000];
  assign o[30999] = i[30999];
  assign o[30998] = i[30998];
  assign o[30997] = i[30997];
  assign o[30996] = i[30996];
  assign o[30995] = i[30995];
  assign o[30994] = i[30994];
  assign o[30993] = i[30993];
  assign o[30992] = i[30992];
  assign o[30991] = i[30991];
  assign o[30990] = i[30990];
  assign o[30989] = i[30989];
  assign o[30988] = i[30988];
  assign o[30987] = i[30987];
  assign o[30986] = i[30986];
  assign o[30985] = i[30985];
  assign o[30984] = i[30984];
  assign o[30983] = i[30983];
  assign o[30982] = i[30982];
  assign o[30981] = i[30981];
  assign o[30980] = i[30980];
  assign o[30979] = i[30979];
  assign o[30978] = i[30978];
  assign o[30977] = i[30977];
  assign o[30976] = i[30976];
  assign o[30975] = i[30975];
  assign o[30974] = i[30974];
  assign o[30973] = i[30973];
  assign o[30972] = i[30972];
  assign o[30971] = i[30971];
  assign o[30970] = i[30970];
  assign o[30969] = i[30969];
  assign o[30968] = i[30968];
  assign o[30967] = i[30967];
  assign o[30966] = i[30966];
  assign o[30965] = i[30965];
  assign o[30964] = i[30964];
  assign o[30963] = i[30963];
  assign o[30962] = i[30962];
  assign o[30961] = i[30961];
  assign o[30960] = i[30960];
  assign o[30959] = i[30959];
  assign o[30958] = i[30958];
  assign o[30957] = i[30957];
  assign o[30956] = i[30956];
  assign o[30955] = i[30955];
  assign o[30954] = i[30954];
  assign o[30953] = i[30953];
  assign o[30952] = i[30952];
  assign o[30951] = i[30951];
  assign o[30950] = i[30950];
  assign o[30949] = i[30949];
  assign o[30948] = i[30948];
  assign o[30947] = i[30947];
  assign o[30946] = i[30946];
  assign o[30945] = i[30945];
  assign o[30944] = i[30944];
  assign o[30943] = i[30943];
  assign o[30942] = i[30942];
  assign o[30941] = i[30941];
  assign o[30940] = i[30940];
  assign o[30939] = i[30939];
  assign o[30938] = i[30938];
  assign o[30937] = i[30937];
  assign o[30936] = i[30936];
  assign o[30935] = i[30935];
  assign o[30934] = i[30934];
  assign o[30933] = i[30933];
  assign o[30932] = i[30932];
  assign o[30931] = i[30931];
  assign o[30930] = i[30930];
  assign o[30929] = i[30929];
  assign o[30928] = i[30928];
  assign o[30927] = i[30927];
  assign o[30926] = i[30926];
  assign o[30925] = i[30925];
  assign o[30924] = i[30924];
  assign o[30923] = i[30923];
  assign o[30922] = i[30922];
  assign o[30921] = i[30921];
  assign o[30920] = i[30920];
  assign o[30919] = i[30919];
  assign o[30918] = i[30918];
  assign o[30917] = i[30917];
  assign o[30916] = i[30916];
  assign o[30915] = i[30915];
  assign o[30914] = i[30914];
  assign o[30913] = i[30913];
  assign o[30912] = i[30912];
  assign o[30911] = i[30911];
  assign o[30910] = i[30910];
  assign o[30909] = i[30909];
  assign o[30908] = i[30908];
  assign o[30907] = i[30907];
  assign o[30906] = i[30906];
  assign o[30905] = i[30905];
  assign o[30904] = i[30904];
  assign o[30903] = i[30903];
  assign o[30902] = i[30902];
  assign o[30901] = i[30901];
  assign o[30900] = i[30900];
  assign o[30899] = i[30899];
  assign o[30898] = i[30898];
  assign o[30897] = i[30897];
  assign o[30896] = i[30896];
  assign o[30895] = i[30895];
  assign o[30894] = i[30894];
  assign o[30893] = i[30893];
  assign o[30892] = i[30892];
  assign o[30891] = i[30891];
  assign o[30890] = i[30890];
  assign o[30889] = i[30889];
  assign o[30888] = i[30888];
  assign o[30887] = i[30887];
  assign o[30886] = i[30886];
  assign o[30885] = i[30885];
  assign o[30884] = i[30884];
  assign o[30883] = i[30883];
  assign o[30882] = i[30882];
  assign o[30881] = i[30881];
  assign o[30880] = i[30880];
  assign o[30879] = i[30879];
  assign o[30878] = i[30878];
  assign o[30877] = i[30877];
  assign o[30876] = i[30876];
  assign o[30875] = i[30875];
  assign o[30874] = i[30874];
  assign o[30873] = i[30873];
  assign o[30872] = i[30872];
  assign o[30871] = i[30871];
  assign o[30870] = i[30870];
  assign o[30869] = i[30869];
  assign o[30868] = i[30868];
  assign o[30867] = i[30867];
  assign o[30866] = i[30866];
  assign o[30865] = i[30865];
  assign o[30864] = i[30864];
  assign o[30863] = i[30863];
  assign o[30862] = i[30862];
  assign o[30861] = i[30861];
  assign o[30860] = i[30860];
  assign o[30859] = i[30859];
  assign o[30858] = i[30858];
  assign o[30857] = i[30857];
  assign o[30856] = i[30856];
  assign o[30855] = i[30855];
  assign o[30854] = i[30854];
  assign o[30853] = i[30853];
  assign o[30852] = i[30852];
  assign o[30851] = i[30851];
  assign o[30850] = i[30850];
  assign o[30849] = i[30849];
  assign o[30848] = i[30848];
  assign o[30847] = i[30847];
  assign o[30846] = i[30846];
  assign o[30845] = i[30845];
  assign o[30844] = i[30844];
  assign o[30843] = i[30843];
  assign o[30842] = i[30842];
  assign o[30841] = i[30841];
  assign o[30840] = i[30840];
  assign o[30839] = i[30839];
  assign o[30838] = i[30838];
  assign o[30837] = i[30837];
  assign o[30836] = i[30836];
  assign o[30835] = i[30835];
  assign o[30834] = i[30834];
  assign o[30833] = i[30833];
  assign o[30832] = i[30832];
  assign o[30831] = i[30831];
  assign o[30830] = i[30830];
  assign o[30829] = i[30829];
  assign o[30828] = i[30828];
  assign o[30827] = i[30827];
  assign o[30826] = i[30826];
  assign o[30825] = i[30825];
  assign o[30824] = i[30824];
  assign o[30823] = i[30823];
  assign o[30822] = i[30822];
  assign o[30821] = i[30821];
  assign o[30820] = i[30820];
  assign o[30819] = i[30819];
  assign o[30818] = i[30818];
  assign o[30817] = i[30817];
  assign o[30816] = i[30816];
  assign o[30815] = i[30815];
  assign o[30814] = i[30814];
  assign o[30813] = i[30813];
  assign o[30812] = i[30812];
  assign o[30811] = i[30811];
  assign o[30810] = i[30810];
  assign o[30809] = i[30809];
  assign o[30808] = i[30808];
  assign o[30807] = i[30807];
  assign o[30806] = i[30806];
  assign o[30805] = i[30805];
  assign o[30804] = i[30804];
  assign o[30803] = i[30803];
  assign o[30802] = i[30802];
  assign o[30801] = i[30801];
  assign o[30800] = i[30800];
  assign o[30799] = i[30799];
  assign o[30798] = i[30798];
  assign o[30797] = i[30797];
  assign o[30796] = i[30796];
  assign o[30795] = i[30795];
  assign o[30794] = i[30794];
  assign o[30793] = i[30793];
  assign o[30792] = i[30792];
  assign o[30791] = i[30791];
  assign o[30790] = i[30790];
  assign o[30789] = i[30789];
  assign o[30788] = i[30788];
  assign o[30787] = i[30787];
  assign o[30786] = i[30786];
  assign o[30785] = i[30785];
  assign o[30784] = i[30784];
  assign o[30783] = i[30783];
  assign o[30782] = i[30782];
  assign o[30781] = i[30781];
  assign o[30780] = i[30780];
  assign o[30779] = i[30779];
  assign o[30778] = i[30778];
  assign o[30777] = i[30777];
  assign o[30776] = i[30776];
  assign o[30775] = i[30775];
  assign o[30774] = i[30774];
  assign o[30773] = i[30773];
  assign o[30772] = i[30772];
  assign o[30771] = i[30771];
  assign o[30770] = i[30770];
  assign o[30769] = i[30769];
  assign o[30768] = i[30768];
  assign o[30767] = i[30767];
  assign o[30766] = i[30766];
  assign o[30765] = i[30765];
  assign o[30764] = i[30764];
  assign o[30763] = i[30763];
  assign o[30762] = i[30762];
  assign o[30761] = i[30761];
  assign o[30760] = i[30760];
  assign o[30759] = i[30759];
  assign o[30758] = i[30758];
  assign o[30757] = i[30757];
  assign o[30756] = i[30756];
  assign o[30755] = i[30755];
  assign o[30754] = i[30754];
  assign o[30753] = i[30753];
  assign o[30752] = i[30752];
  assign o[30751] = i[30751];
  assign o[30750] = i[30750];
  assign o[30749] = i[30749];
  assign o[30748] = i[30748];
  assign o[30747] = i[30747];
  assign o[30746] = i[30746];
  assign o[30745] = i[30745];
  assign o[30744] = i[30744];
  assign o[30743] = i[30743];
  assign o[30742] = i[30742];
  assign o[30741] = i[30741];
  assign o[30740] = i[30740];
  assign o[30739] = i[30739];
  assign o[30738] = i[30738];
  assign o[30737] = i[30737];
  assign o[30736] = i[30736];
  assign o[30735] = i[30735];
  assign o[30734] = i[30734];
  assign o[30733] = i[30733];
  assign o[30732] = i[30732];
  assign o[30731] = i[30731];
  assign o[30730] = i[30730];
  assign o[30729] = i[30729];
  assign o[30728] = i[30728];
  assign o[30727] = i[30727];
  assign o[30726] = i[30726];
  assign o[30725] = i[30725];
  assign o[30724] = i[30724];
  assign o[30723] = i[30723];
  assign o[30722] = i[30722];
  assign o[30721] = i[30721];
  assign o[30720] = i[30720];
  assign o[30719] = i[30719];
  assign o[30718] = i[30718];
  assign o[30717] = i[30717];
  assign o[30716] = i[30716];
  assign o[30715] = i[30715];
  assign o[30714] = i[30714];
  assign o[30713] = i[30713];
  assign o[30712] = i[30712];
  assign o[30711] = i[30711];
  assign o[30710] = i[30710];
  assign o[30709] = i[30709];
  assign o[30708] = i[30708];
  assign o[30707] = i[30707];
  assign o[30706] = i[30706];
  assign o[30705] = i[30705];
  assign o[30704] = i[30704];
  assign o[30703] = i[30703];
  assign o[30702] = i[30702];
  assign o[30701] = i[30701];
  assign o[30700] = i[30700];
  assign o[30699] = i[30699];
  assign o[30698] = i[30698];
  assign o[30697] = i[30697];
  assign o[30696] = i[30696];
  assign o[30695] = i[30695];
  assign o[30694] = i[30694];
  assign o[30693] = i[30693];
  assign o[30692] = i[30692];
  assign o[30691] = i[30691];
  assign o[30690] = i[30690];
  assign o[30689] = i[30689];
  assign o[30688] = i[30688];
  assign o[30687] = i[30687];
  assign o[30686] = i[30686];
  assign o[30685] = i[30685];
  assign o[30684] = i[30684];
  assign o[30683] = i[30683];
  assign o[30682] = i[30682];
  assign o[30681] = i[30681];
  assign o[30680] = i[30680];
  assign o[30679] = i[30679];
  assign o[30678] = i[30678];
  assign o[30677] = i[30677];
  assign o[30676] = i[30676];
  assign o[30675] = i[30675];
  assign o[30674] = i[30674];
  assign o[30673] = i[30673];
  assign o[30672] = i[30672];
  assign o[30671] = i[30671];
  assign o[30670] = i[30670];
  assign o[30669] = i[30669];
  assign o[30668] = i[30668];
  assign o[30667] = i[30667];
  assign o[30666] = i[30666];
  assign o[30665] = i[30665];
  assign o[30664] = i[30664];
  assign o[30663] = i[30663];
  assign o[30662] = i[30662];
  assign o[30661] = i[30661];
  assign o[30660] = i[30660];
  assign o[30659] = i[30659];
  assign o[30658] = i[30658];
  assign o[30657] = i[30657];
  assign o[30656] = i[30656];
  assign o[30655] = i[30655];
  assign o[30654] = i[30654];
  assign o[30653] = i[30653];
  assign o[30652] = i[30652];
  assign o[30651] = i[30651];
  assign o[30650] = i[30650];
  assign o[30649] = i[30649];
  assign o[30648] = i[30648];
  assign o[30647] = i[30647];
  assign o[30646] = i[30646];
  assign o[30645] = i[30645];
  assign o[30644] = i[30644];
  assign o[30643] = i[30643];
  assign o[30642] = i[30642];
  assign o[30641] = i[30641];
  assign o[30640] = i[30640];
  assign o[30639] = i[30639];
  assign o[30638] = i[30638];
  assign o[30637] = i[30637];
  assign o[30636] = i[30636];
  assign o[30635] = i[30635];
  assign o[30634] = i[30634];
  assign o[30633] = i[30633];
  assign o[30632] = i[30632];
  assign o[30631] = i[30631];
  assign o[30630] = i[30630];
  assign o[30629] = i[30629];
  assign o[30628] = i[30628];
  assign o[30627] = i[30627];
  assign o[30626] = i[30626];
  assign o[30625] = i[30625];
  assign o[30624] = i[30624];
  assign o[30623] = i[30623];
  assign o[30622] = i[30622];
  assign o[30621] = i[30621];
  assign o[30620] = i[30620];
  assign o[30619] = i[30619];
  assign o[30618] = i[30618];
  assign o[30617] = i[30617];
  assign o[30616] = i[30616];
  assign o[30615] = i[30615];
  assign o[30614] = i[30614];
  assign o[30613] = i[30613];
  assign o[30612] = i[30612];
  assign o[30611] = i[30611];
  assign o[30610] = i[30610];
  assign o[30609] = i[30609];
  assign o[30608] = i[30608];
  assign o[30607] = i[30607];
  assign o[30606] = i[30606];
  assign o[30605] = i[30605];
  assign o[30604] = i[30604];
  assign o[30603] = i[30603];
  assign o[30602] = i[30602];
  assign o[30601] = i[30601];
  assign o[30600] = i[30600];
  assign o[30599] = i[30599];
  assign o[30598] = i[30598];
  assign o[30597] = i[30597];
  assign o[30596] = i[30596];
  assign o[30595] = i[30595];
  assign o[30594] = i[30594];
  assign o[30593] = i[30593];
  assign o[30592] = i[30592];
  assign o[30591] = i[30591];
  assign o[30590] = i[30590];
  assign o[30589] = i[30589];
  assign o[30588] = i[30588];
  assign o[30587] = i[30587];
  assign o[30586] = i[30586];
  assign o[30585] = i[30585];
  assign o[30584] = i[30584];
  assign o[30583] = i[30583];
  assign o[30582] = i[30582];
  assign o[30581] = i[30581];
  assign o[30580] = i[30580];
  assign o[30579] = i[30579];
  assign o[30578] = i[30578];
  assign o[30577] = i[30577];
  assign o[30576] = i[30576];
  assign o[30575] = i[30575];
  assign o[30574] = i[30574];
  assign o[30573] = i[30573];
  assign o[30572] = i[30572];
  assign o[30571] = i[30571];
  assign o[30570] = i[30570];
  assign o[30569] = i[30569];
  assign o[30568] = i[30568];
  assign o[30567] = i[30567];
  assign o[30566] = i[30566];
  assign o[30565] = i[30565];
  assign o[30564] = i[30564];
  assign o[30563] = i[30563];
  assign o[30562] = i[30562];
  assign o[30561] = i[30561];
  assign o[30560] = i[30560];
  assign o[30559] = i[30559];
  assign o[30558] = i[30558];
  assign o[30557] = i[30557];
  assign o[30556] = i[30556];
  assign o[30555] = i[30555];
  assign o[30554] = i[30554];
  assign o[30553] = i[30553];
  assign o[30552] = i[30552];
  assign o[30551] = i[30551];
  assign o[30550] = i[30550];
  assign o[30549] = i[30549];
  assign o[30548] = i[30548];
  assign o[30547] = i[30547];
  assign o[30546] = i[30546];
  assign o[30545] = i[30545];
  assign o[30544] = i[30544];
  assign o[30543] = i[30543];
  assign o[30542] = i[30542];
  assign o[30541] = i[30541];
  assign o[30540] = i[30540];
  assign o[30539] = i[30539];
  assign o[30538] = i[30538];
  assign o[30537] = i[30537];
  assign o[30536] = i[30536];
  assign o[30535] = i[30535];
  assign o[30534] = i[30534];
  assign o[30533] = i[30533];
  assign o[30532] = i[30532];
  assign o[30531] = i[30531];
  assign o[30530] = i[30530];
  assign o[30529] = i[30529];
  assign o[30528] = i[30528];
  assign o[30527] = i[30527];
  assign o[30526] = i[30526];
  assign o[30525] = i[30525];
  assign o[30524] = i[30524];
  assign o[30523] = i[30523];
  assign o[30522] = i[30522];
  assign o[30521] = i[30521];
  assign o[30520] = i[30520];
  assign o[30519] = i[30519];
  assign o[30518] = i[30518];
  assign o[30517] = i[30517];
  assign o[30516] = i[30516];
  assign o[30515] = i[30515];
  assign o[30514] = i[30514];
  assign o[30513] = i[30513];
  assign o[30512] = i[30512];
  assign o[30511] = i[30511];
  assign o[30510] = i[30510];
  assign o[30509] = i[30509];
  assign o[30508] = i[30508];
  assign o[30507] = i[30507];
  assign o[30506] = i[30506];
  assign o[30505] = i[30505];
  assign o[30504] = i[30504];
  assign o[30503] = i[30503];
  assign o[30502] = i[30502];
  assign o[30501] = i[30501];
  assign o[30500] = i[30500];
  assign o[30499] = i[30499];
  assign o[30498] = i[30498];
  assign o[30497] = i[30497];
  assign o[30496] = i[30496];
  assign o[30495] = i[30495];
  assign o[30494] = i[30494];
  assign o[30493] = i[30493];
  assign o[30492] = i[30492];
  assign o[30491] = i[30491];
  assign o[30490] = i[30490];
  assign o[30489] = i[30489];
  assign o[30488] = i[30488];
  assign o[30487] = i[30487];
  assign o[30486] = i[30486];
  assign o[30485] = i[30485];
  assign o[30484] = i[30484];
  assign o[30483] = i[30483];
  assign o[30482] = i[30482];
  assign o[30481] = i[30481];
  assign o[30480] = i[30480];
  assign o[30479] = i[30479];
  assign o[30478] = i[30478];
  assign o[30477] = i[30477];
  assign o[30476] = i[30476];
  assign o[30475] = i[30475];
  assign o[30474] = i[30474];
  assign o[30473] = i[30473];
  assign o[30472] = i[30472];
  assign o[30471] = i[30471];
  assign o[30470] = i[30470];
  assign o[30469] = i[30469];
  assign o[30468] = i[30468];
  assign o[30467] = i[30467];
  assign o[30466] = i[30466];
  assign o[30465] = i[30465];
  assign o[30464] = i[30464];
  assign o[30463] = i[30463];
  assign o[30462] = i[30462];
  assign o[30461] = i[30461];
  assign o[30460] = i[30460];
  assign o[30459] = i[30459];
  assign o[30458] = i[30458];
  assign o[30457] = i[30457];
  assign o[30456] = i[30456];
  assign o[30455] = i[30455];
  assign o[30454] = i[30454];
  assign o[30453] = i[30453];
  assign o[30452] = i[30452];
  assign o[30451] = i[30451];
  assign o[30450] = i[30450];
  assign o[30449] = i[30449];
  assign o[30448] = i[30448];
  assign o[30447] = i[30447];
  assign o[30446] = i[30446];
  assign o[30445] = i[30445];
  assign o[30444] = i[30444];
  assign o[30443] = i[30443];
  assign o[30442] = i[30442];
  assign o[30441] = i[30441];
  assign o[30440] = i[30440];
  assign o[30439] = i[30439];
  assign o[30438] = i[30438];
  assign o[30437] = i[30437];
  assign o[30436] = i[30436];
  assign o[30435] = i[30435];
  assign o[30434] = i[30434];
  assign o[30433] = i[30433];
  assign o[30432] = i[30432];
  assign o[30431] = i[30431];
  assign o[30430] = i[30430];
  assign o[30429] = i[30429];
  assign o[30428] = i[30428];
  assign o[30427] = i[30427];
  assign o[30426] = i[30426];
  assign o[30425] = i[30425];
  assign o[30424] = i[30424];
  assign o[30423] = i[30423];
  assign o[30422] = i[30422];
  assign o[30421] = i[30421];
  assign o[30420] = i[30420];
  assign o[30419] = i[30419];
  assign o[30418] = i[30418];
  assign o[30417] = i[30417];
  assign o[30416] = i[30416];
  assign o[30415] = i[30415];
  assign o[30414] = i[30414];
  assign o[30413] = i[30413];
  assign o[30412] = i[30412];
  assign o[30411] = i[30411];
  assign o[30410] = i[30410];
  assign o[30409] = i[30409];
  assign o[30408] = i[30408];
  assign o[30407] = i[30407];
  assign o[30406] = i[30406];
  assign o[30405] = i[30405];
  assign o[30404] = i[30404];
  assign o[30403] = i[30403];
  assign o[30402] = i[30402];
  assign o[30401] = i[30401];
  assign o[30400] = i[30400];
  assign o[30399] = i[30399];
  assign o[30398] = i[30398];
  assign o[30397] = i[30397];
  assign o[30396] = i[30396];
  assign o[30395] = i[30395];
  assign o[30394] = i[30394];
  assign o[30393] = i[30393];
  assign o[30392] = i[30392];
  assign o[30391] = i[30391];
  assign o[30390] = i[30390];
  assign o[30389] = i[30389];
  assign o[30388] = i[30388];
  assign o[30387] = i[30387];
  assign o[30386] = i[30386];
  assign o[30385] = i[30385];
  assign o[30384] = i[30384];
  assign o[30383] = i[30383];
  assign o[30382] = i[30382];
  assign o[30381] = i[30381];
  assign o[30380] = i[30380];
  assign o[30379] = i[30379];
  assign o[30378] = i[30378];
  assign o[30377] = i[30377];
  assign o[30376] = i[30376];
  assign o[30375] = i[30375];
  assign o[30374] = i[30374];
  assign o[30373] = i[30373];
  assign o[30372] = i[30372];
  assign o[30371] = i[30371];
  assign o[30370] = i[30370];
  assign o[30369] = i[30369];
  assign o[30368] = i[30368];
  assign o[30367] = i[30367];
  assign o[30366] = i[30366];
  assign o[30365] = i[30365];
  assign o[30364] = i[30364];
  assign o[30363] = i[30363];
  assign o[30362] = i[30362];
  assign o[30361] = i[30361];
  assign o[30360] = i[30360];
  assign o[30359] = i[30359];
  assign o[30358] = i[30358];
  assign o[30357] = i[30357];
  assign o[30356] = i[30356];
  assign o[30355] = i[30355];
  assign o[30354] = i[30354];
  assign o[30353] = i[30353];
  assign o[30352] = i[30352];
  assign o[30351] = i[30351];
  assign o[30350] = i[30350];
  assign o[30349] = i[30349];
  assign o[30348] = i[30348];
  assign o[30347] = i[30347];
  assign o[30346] = i[30346];
  assign o[30345] = i[30345];
  assign o[30344] = i[30344];
  assign o[30343] = i[30343];
  assign o[30342] = i[30342];
  assign o[30341] = i[30341];
  assign o[30340] = i[30340];
  assign o[30339] = i[30339];
  assign o[30338] = i[30338];
  assign o[30337] = i[30337];
  assign o[30336] = i[30336];
  assign o[30335] = i[30335];
  assign o[30334] = i[30334];
  assign o[30333] = i[30333];
  assign o[30332] = i[30332];
  assign o[30331] = i[30331];
  assign o[30330] = i[30330];
  assign o[30329] = i[30329];
  assign o[30328] = i[30328];
  assign o[30327] = i[30327];
  assign o[30326] = i[30326];
  assign o[30325] = i[30325];
  assign o[30324] = i[30324];
  assign o[30323] = i[30323];
  assign o[30322] = i[30322];
  assign o[30321] = i[30321];
  assign o[30320] = i[30320];
  assign o[30319] = i[30319];
  assign o[30318] = i[30318];
  assign o[30317] = i[30317];
  assign o[30316] = i[30316];
  assign o[30315] = i[30315];
  assign o[30314] = i[30314];
  assign o[30313] = i[30313];
  assign o[30312] = i[30312];
  assign o[30311] = i[30311];
  assign o[30310] = i[30310];
  assign o[30309] = i[30309];
  assign o[30308] = i[30308];
  assign o[30307] = i[30307];
  assign o[30306] = i[30306];
  assign o[30305] = i[30305];
  assign o[30304] = i[30304];
  assign o[30303] = i[30303];
  assign o[30302] = i[30302];
  assign o[30301] = i[30301];
  assign o[30300] = i[30300];
  assign o[30299] = i[30299];
  assign o[30298] = i[30298];
  assign o[30297] = i[30297];
  assign o[30296] = i[30296];
  assign o[30295] = i[30295];
  assign o[30294] = i[30294];
  assign o[30293] = i[30293];
  assign o[30292] = i[30292];
  assign o[30291] = i[30291];
  assign o[30290] = i[30290];
  assign o[30289] = i[30289];
  assign o[30288] = i[30288];
  assign o[30287] = i[30287];
  assign o[30286] = i[30286];
  assign o[30285] = i[30285];
  assign o[30284] = i[30284];
  assign o[30283] = i[30283];
  assign o[30282] = i[30282];
  assign o[30281] = i[30281];
  assign o[30280] = i[30280];
  assign o[30279] = i[30279];
  assign o[30278] = i[30278];
  assign o[30277] = i[30277];
  assign o[30276] = i[30276];
  assign o[30275] = i[30275];
  assign o[30274] = i[30274];
  assign o[30273] = i[30273];
  assign o[30272] = i[30272];
  assign o[30271] = i[30271];
  assign o[30270] = i[30270];
  assign o[30269] = i[30269];
  assign o[30268] = i[30268];
  assign o[30267] = i[30267];
  assign o[30266] = i[30266];
  assign o[30265] = i[30265];
  assign o[30264] = i[30264];
  assign o[30263] = i[30263];
  assign o[30262] = i[30262];
  assign o[30261] = i[30261];
  assign o[30260] = i[30260];
  assign o[30259] = i[30259];
  assign o[30258] = i[30258];
  assign o[30257] = i[30257];
  assign o[30256] = i[30256];
  assign o[30255] = i[30255];
  assign o[30254] = i[30254];
  assign o[30253] = i[30253];
  assign o[30252] = i[30252];
  assign o[30251] = i[30251];
  assign o[30250] = i[30250];
  assign o[30249] = i[30249];
  assign o[30248] = i[30248];
  assign o[30247] = i[30247];
  assign o[30246] = i[30246];
  assign o[30245] = i[30245];
  assign o[30244] = i[30244];
  assign o[30243] = i[30243];
  assign o[30242] = i[30242];
  assign o[30241] = i[30241];
  assign o[30240] = i[30240];
  assign o[30239] = i[30239];
  assign o[30238] = i[30238];
  assign o[30237] = i[30237];
  assign o[30236] = i[30236];
  assign o[30235] = i[30235];
  assign o[30234] = i[30234];
  assign o[30233] = i[30233];
  assign o[30232] = i[30232];
  assign o[30231] = i[30231];
  assign o[30230] = i[30230];
  assign o[30229] = i[30229];
  assign o[30228] = i[30228];
  assign o[30227] = i[30227];
  assign o[30226] = i[30226];
  assign o[30225] = i[30225];
  assign o[30224] = i[30224];
  assign o[30223] = i[30223];
  assign o[30222] = i[30222];
  assign o[30221] = i[30221];
  assign o[30220] = i[30220];
  assign o[30219] = i[30219];
  assign o[30218] = i[30218];
  assign o[30217] = i[30217];
  assign o[30216] = i[30216];
  assign o[30215] = i[30215];
  assign o[30214] = i[30214];
  assign o[30213] = i[30213];
  assign o[30212] = i[30212];
  assign o[30211] = i[30211];
  assign o[30210] = i[30210];
  assign o[30209] = i[30209];
  assign o[30208] = i[30208];
  assign o[30207] = i[30207];
  assign o[30206] = i[30206];
  assign o[30205] = i[30205];
  assign o[30204] = i[30204];
  assign o[30203] = i[30203];
  assign o[30202] = i[30202];
  assign o[30201] = i[30201];
  assign o[30200] = i[30200];
  assign o[30199] = i[30199];
  assign o[30198] = i[30198];
  assign o[30197] = i[30197];
  assign o[30196] = i[30196];
  assign o[30195] = i[30195];
  assign o[30194] = i[30194];
  assign o[30193] = i[30193];
  assign o[30192] = i[30192];
  assign o[30191] = i[30191];
  assign o[30190] = i[30190];
  assign o[30189] = i[30189];
  assign o[30188] = i[30188];
  assign o[30187] = i[30187];
  assign o[30186] = i[30186];
  assign o[30185] = i[30185];
  assign o[30184] = i[30184];
  assign o[30183] = i[30183];
  assign o[30182] = i[30182];
  assign o[30181] = i[30181];
  assign o[30180] = i[30180];
  assign o[30179] = i[30179];
  assign o[30178] = i[30178];
  assign o[30177] = i[30177];
  assign o[30176] = i[30176];
  assign o[30175] = i[30175];
  assign o[30174] = i[30174];
  assign o[30173] = i[30173];
  assign o[30172] = i[30172];
  assign o[30171] = i[30171];
  assign o[30170] = i[30170];
  assign o[30169] = i[30169];
  assign o[30168] = i[30168];
  assign o[30167] = i[30167];
  assign o[30166] = i[30166];
  assign o[30165] = i[30165];
  assign o[30164] = i[30164];
  assign o[30163] = i[30163];
  assign o[30162] = i[30162];
  assign o[30161] = i[30161];
  assign o[30160] = i[30160];
  assign o[30159] = i[30159];
  assign o[30158] = i[30158];
  assign o[30157] = i[30157];
  assign o[30156] = i[30156];
  assign o[30155] = i[30155];
  assign o[30154] = i[30154];
  assign o[30153] = i[30153];
  assign o[30152] = i[30152];
  assign o[30151] = i[30151];
  assign o[30150] = i[30150];
  assign o[30149] = i[30149];
  assign o[30148] = i[30148];
  assign o[30147] = i[30147];
  assign o[30146] = i[30146];
  assign o[30145] = i[30145];
  assign o[30144] = i[30144];
  assign o[30143] = i[30143];
  assign o[30142] = i[30142];
  assign o[30141] = i[30141];
  assign o[30140] = i[30140];
  assign o[30139] = i[30139];
  assign o[30138] = i[30138];
  assign o[30137] = i[30137];
  assign o[30136] = i[30136];
  assign o[30135] = i[30135];
  assign o[30134] = i[30134];
  assign o[30133] = i[30133];
  assign o[30132] = i[30132];
  assign o[30131] = i[30131];
  assign o[30130] = i[30130];
  assign o[30129] = i[30129];
  assign o[30128] = i[30128];
  assign o[30127] = i[30127];
  assign o[30126] = i[30126];
  assign o[30125] = i[30125];
  assign o[30124] = i[30124];
  assign o[30123] = i[30123];
  assign o[30122] = i[30122];
  assign o[30121] = i[30121];
  assign o[30120] = i[30120];
  assign o[30119] = i[30119];
  assign o[30118] = i[30118];
  assign o[30117] = i[30117];
  assign o[30116] = i[30116];
  assign o[30115] = i[30115];
  assign o[30114] = i[30114];
  assign o[30113] = i[30113];
  assign o[30112] = i[30112];
  assign o[30111] = i[30111];
  assign o[30110] = i[30110];
  assign o[30109] = i[30109];
  assign o[30108] = i[30108];
  assign o[30107] = i[30107];
  assign o[30106] = i[30106];
  assign o[30105] = i[30105];
  assign o[30104] = i[30104];
  assign o[30103] = i[30103];
  assign o[30102] = i[30102];
  assign o[30101] = i[30101];
  assign o[30100] = i[30100];
  assign o[30099] = i[30099];
  assign o[30098] = i[30098];
  assign o[30097] = i[30097];
  assign o[30096] = i[30096];
  assign o[30095] = i[30095];
  assign o[30094] = i[30094];
  assign o[30093] = i[30093];
  assign o[30092] = i[30092];
  assign o[30091] = i[30091];
  assign o[30090] = i[30090];
  assign o[30089] = i[30089];
  assign o[30088] = i[30088];
  assign o[30087] = i[30087];
  assign o[30086] = i[30086];
  assign o[30085] = i[30085];
  assign o[30084] = i[30084];
  assign o[30083] = i[30083];
  assign o[30082] = i[30082];
  assign o[30081] = i[30081];
  assign o[30080] = i[30080];
  assign o[30079] = i[30079];
  assign o[30078] = i[30078];
  assign o[30077] = i[30077];
  assign o[30076] = i[30076];
  assign o[30075] = i[30075];
  assign o[30074] = i[30074];
  assign o[30073] = i[30073];
  assign o[30072] = i[30072];
  assign o[30071] = i[30071];
  assign o[30070] = i[30070];
  assign o[30069] = i[30069];
  assign o[30068] = i[30068];
  assign o[30067] = i[30067];
  assign o[30066] = i[30066];
  assign o[30065] = i[30065];
  assign o[30064] = i[30064];
  assign o[30063] = i[30063];
  assign o[30062] = i[30062];
  assign o[30061] = i[30061];
  assign o[30060] = i[30060];
  assign o[30059] = i[30059];
  assign o[30058] = i[30058];
  assign o[30057] = i[30057];
  assign o[30056] = i[30056];
  assign o[30055] = i[30055];
  assign o[30054] = i[30054];
  assign o[30053] = i[30053];
  assign o[30052] = i[30052];
  assign o[30051] = i[30051];
  assign o[30050] = i[30050];
  assign o[30049] = i[30049];
  assign o[30048] = i[30048];
  assign o[30047] = i[30047];
  assign o[30046] = i[30046];
  assign o[30045] = i[30045];
  assign o[30044] = i[30044];
  assign o[30043] = i[30043];
  assign o[30042] = i[30042];
  assign o[30041] = i[30041];
  assign o[30040] = i[30040];
  assign o[30039] = i[30039];
  assign o[30038] = i[30038];
  assign o[30037] = i[30037];
  assign o[30036] = i[30036];
  assign o[30035] = i[30035];
  assign o[30034] = i[30034];
  assign o[30033] = i[30033];
  assign o[30032] = i[30032];
  assign o[30031] = i[30031];
  assign o[30030] = i[30030];
  assign o[30029] = i[30029];
  assign o[30028] = i[30028];
  assign o[30027] = i[30027];
  assign o[30026] = i[30026];
  assign o[30025] = i[30025];
  assign o[30024] = i[30024];
  assign o[30023] = i[30023];
  assign o[30022] = i[30022];
  assign o[30021] = i[30021];
  assign o[30020] = i[30020];
  assign o[30019] = i[30019];
  assign o[30018] = i[30018];
  assign o[30017] = i[30017];
  assign o[30016] = i[30016];
  assign o[30015] = i[30015];
  assign o[30014] = i[30014];
  assign o[30013] = i[30013];
  assign o[30012] = i[30012];
  assign o[30011] = i[30011];
  assign o[30010] = i[30010];
  assign o[30009] = i[30009];
  assign o[30008] = i[30008];
  assign o[30007] = i[30007];
  assign o[30006] = i[30006];
  assign o[30005] = i[30005];
  assign o[30004] = i[30004];
  assign o[30003] = i[30003];
  assign o[30002] = i[30002];
  assign o[30001] = i[30001];
  assign o[30000] = i[30000];
  assign o[29999] = i[29999];
  assign o[29998] = i[29998];
  assign o[29997] = i[29997];
  assign o[29996] = i[29996];
  assign o[29995] = i[29995];
  assign o[29994] = i[29994];
  assign o[29993] = i[29993];
  assign o[29992] = i[29992];
  assign o[29991] = i[29991];
  assign o[29990] = i[29990];
  assign o[29989] = i[29989];
  assign o[29988] = i[29988];
  assign o[29987] = i[29987];
  assign o[29986] = i[29986];
  assign o[29985] = i[29985];
  assign o[29984] = i[29984];
  assign o[29983] = i[29983];
  assign o[29982] = i[29982];
  assign o[29981] = i[29981];
  assign o[29980] = i[29980];
  assign o[29979] = i[29979];
  assign o[29978] = i[29978];
  assign o[29977] = i[29977];
  assign o[29976] = i[29976];
  assign o[29975] = i[29975];
  assign o[29974] = i[29974];
  assign o[29973] = i[29973];
  assign o[29972] = i[29972];
  assign o[29971] = i[29971];
  assign o[29970] = i[29970];
  assign o[29969] = i[29969];
  assign o[29968] = i[29968];
  assign o[29967] = i[29967];
  assign o[29966] = i[29966];
  assign o[29965] = i[29965];
  assign o[29964] = i[29964];
  assign o[29963] = i[29963];
  assign o[29962] = i[29962];
  assign o[29961] = i[29961];
  assign o[29960] = i[29960];
  assign o[29959] = i[29959];
  assign o[29958] = i[29958];
  assign o[29957] = i[29957];
  assign o[29956] = i[29956];
  assign o[29955] = i[29955];
  assign o[29954] = i[29954];
  assign o[29953] = i[29953];
  assign o[29952] = i[29952];
  assign o[29951] = i[29951];
  assign o[29950] = i[29950];
  assign o[29949] = i[29949];
  assign o[29948] = i[29948];
  assign o[29947] = i[29947];
  assign o[29946] = i[29946];
  assign o[29945] = i[29945];
  assign o[29944] = i[29944];
  assign o[29943] = i[29943];
  assign o[29942] = i[29942];
  assign o[29941] = i[29941];
  assign o[29940] = i[29940];
  assign o[29939] = i[29939];
  assign o[29938] = i[29938];
  assign o[29937] = i[29937];
  assign o[29936] = i[29936];
  assign o[29935] = i[29935];
  assign o[29934] = i[29934];
  assign o[29933] = i[29933];
  assign o[29932] = i[29932];
  assign o[29931] = i[29931];
  assign o[29930] = i[29930];
  assign o[29929] = i[29929];
  assign o[29928] = i[29928];
  assign o[29927] = i[29927];
  assign o[29926] = i[29926];
  assign o[29925] = i[29925];
  assign o[29924] = i[29924];
  assign o[29923] = i[29923];
  assign o[29922] = i[29922];
  assign o[29921] = i[29921];
  assign o[29920] = i[29920];
  assign o[29919] = i[29919];
  assign o[29918] = i[29918];
  assign o[29917] = i[29917];
  assign o[29916] = i[29916];
  assign o[29915] = i[29915];
  assign o[29914] = i[29914];
  assign o[29913] = i[29913];
  assign o[29912] = i[29912];
  assign o[29911] = i[29911];
  assign o[29910] = i[29910];
  assign o[29909] = i[29909];
  assign o[29908] = i[29908];
  assign o[29907] = i[29907];
  assign o[29906] = i[29906];
  assign o[29905] = i[29905];
  assign o[29904] = i[29904];
  assign o[29903] = i[29903];
  assign o[29902] = i[29902];
  assign o[29901] = i[29901];
  assign o[29900] = i[29900];
  assign o[29899] = i[29899];
  assign o[29898] = i[29898];
  assign o[29897] = i[29897];
  assign o[29896] = i[29896];
  assign o[29895] = i[29895];
  assign o[29894] = i[29894];
  assign o[29893] = i[29893];
  assign o[29892] = i[29892];
  assign o[29891] = i[29891];
  assign o[29890] = i[29890];
  assign o[29889] = i[29889];
  assign o[29888] = i[29888];
  assign o[29887] = i[29887];
  assign o[29886] = i[29886];
  assign o[29885] = i[29885];
  assign o[29884] = i[29884];
  assign o[29883] = i[29883];
  assign o[29882] = i[29882];
  assign o[29881] = i[29881];
  assign o[29880] = i[29880];
  assign o[29879] = i[29879];
  assign o[29878] = i[29878];
  assign o[29877] = i[29877];
  assign o[29876] = i[29876];
  assign o[29875] = i[29875];
  assign o[29874] = i[29874];
  assign o[29873] = i[29873];
  assign o[29872] = i[29872];
  assign o[29871] = i[29871];
  assign o[29870] = i[29870];
  assign o[29869] = i[29869];
  assign o[29868] = i[29868];
  assign o[29867] = i[29867];
  assign o[29866] = i[29866];
  assign o[29865] = i[29865];
  assign o[29864] = i[29864];
  assign o[29863] = i[29863];
  assign o[29862] = i[29862];
  assign o[29861] = i[29861];
  assign o[29860] = i[29860];
  assign o[29859] = i[29859];
  assign o[29858] = i[29858];
  assign o[29857] = i[29857];
  assign o[29856] = i[29856];
  assign o[29855] = i[29855];
  assign o[29854] = i[29854];
  assign o[29853] = i[29853];
  assign o[29852] = i[29852];
  assign o[29851] = i[29851];
  assign o[29850] = i[29850];
  assign o[29849] = i[29849];
  assign o[29848] = i[29848];
  assign o[29847] = i[29847];
  assign o[29846] = i[29846];
  assign o[29845] = i[29845];
  assign o[29844] = i[29844];
  assign o[29843] = i[29843];
  assign o[29842] = i[29842];
  assign o[29841] = i[29841];
  assign o[29840] = i[29840];
  assign o[29839] = i[29839];
  assign o[29838] = i[29838];
  assign o[29837] = i[29837];
  assign o[29836] = i[29836];
  assign o[29835] = i[29835];
  assign o[29834] = i[29834];
  assign o[29833] = i[29833];
  assign o[29832] = i[29832];
  assign o[29831] = i[29831];
  assign o[29830] = i[29830];
  assign o[29829] = i[29829];
  assign o[29828] = i[29828];
  assign o[29827] = i[29827];
  assign o[29826] = i[29826];
  assign o[29825] = i[29825];
  assign o[29824] = i[29824];
  assign o[29823] = i[29823];
  assign o[29822] = i[29822];
  assign o[29821] = i[29821];
  assign o[29820] = i[29820];
  assign o[29819] = i[29819];
  assign o[29818] = i[29818];
  assign o[29817] = i[29817];
  assign o[29816] = i[29816];
  assign o[29815] = i[29815];
  assign o[29814] = i[29814];
  assign o[29813] = i[29813];
  assign o[29812] = i[29812];
  assign o[29811] = i[29811];
  assign o[29810] = i[29810];
  assign o[29809] = i[29809];
  assign o[29808] = i[29808];
  assign o[29807] = i[29807];
  assign o[29806] = i[29806];
  assign o[29805] = i[29805];
  assign o[29804] = i[29804];
  assign o[29803] = i[29803];
  assign o[29802] = i[29802];
  assign o[29801] = i[29801];
  assign o[29800] = i[29800];
  assign o[29799] = i[29799];
  assign o[29798] = i[29798];
  assign o[29797] = i[29797];
  assign o[29796] = i[29796];
  assign o[29795] = i[29795];
  assign o[29794] = i[29794];
  assign o[29793] = i[29793];
  assign o[29792] = i[29792];
  assign o[29791] = i[29791];
  assign o[29790] = i[29790];
  assign o[29789] = i[29789];
  assign o[29788] = i[29788];
  assign o[29787] = i[29787];
  assign o[29786] = i[29786];
  assign o[29785] = i[29785];
  assign o[29784] = i[29784];
  assign o[29783] = i[29783];
  assign o[29782] = i[29782];
  assign o[29781] = i[29781];
  assign o[29780] = i[29780];
  assign o[29779] = i[29779];
  assign o[29778] = i[29778];
  assign o[29777] = i[29777];
  assign o[29776] = i[29776];
  assign o[29775] = i[29775];
  assign o[29774] = i[29774];
  assign o[29773] = i[29773];
  assign o[29772] = i[29772];
  assign o[29771] = i[29771];
  assign o[29770] = i[29770];
  assign o[29769] = i[29769];
  assign o[29768] = i[29768];
  assign o[29767] = i[29767];
  assign o[29766] = i[29766];
  assign o[29765] = i[29765];
  assign o[29764] = i[29764];
  assign o[29763] = i[29763];
  assign o[29762] = i[29762];
  assign o[29761] = i[29761];
  assign o[29760] = i[29760];
  assign o[29759] = i[29759];
  assign o[29758] = i[29758];
  assign o[29757] = i[29757];
  assign o[29756] = i[29756];
  assign o[29755] = i[29755];
  assign o[29754] = i[29754];
  assign o[29753] = i[29753];
  assign o[29752] = i[29752];
  assign o[29751] = i[29751];
  assign o[29750] = i[29750];
  assign o[29749] = i[29749];
  assign o[29748] = i[29748];
  assign o[29747] = i[29747];
  assign o[29746] = i[29746];
  assign o[29745] = i[29745];
  assign o[29744] = i[29744];
  assign o[29743] = i[29743];
  assign o[29742] = i[29742];
  assign o[29741] = i[29741];
  assign o[29740] = i[29740];
  assign o[29739] = i[29739];
  assign o[29738] = i[29738];
  assign o[29737] = i[29737];
  assign o[29736] = i[29736];
  assign o[29735] = i[29735];
  assign o[29734] = i[29734];
  assign o[29733] = i[29733];
  assign o[29732] = i[29732];
  assign o[29731] = i[29731];
  assign o[29730] = i[29730];
  assign o[29729] = i[29729];
  assign o[29728] = i[29728];
  assign o[29727] = i[29727];
  assign o[29726] = i[29726];
  assign o[29725] = i[29725];
  assign o[29724] = i[29724];
  assign o[29723] = i[29723];
  assign o[29722] = i[29722];
  assign o[29721] = i[29721];
  assign o[29720] = i[29720];
  assign o[29719] = i[29719];
  assign o[29718] = i[29718];
  assign o[29717] = i[29717];
  assign o[29716] = i[29716];
  assign o[29715] = i[29715];
  assign o[29714] = i[29714];
  assign o[29713] = i[29713];
  assign o[29712] = i[29712];
  assign o[29711] = i[29711];
  assign o[29710] = i[29710];
  assign o[29709] = i[29709];
  assign o[29708] = i[29708];
  assign o[29707] = i[29707];
  assign o[29706] = i[29706];
  assign o[29705] = i[29705];
  assign o[29704] = i[29704];
  assign o[29703] = i[29703];
  assign o[29702] = i[29702];
  assign o[29701] = i[29701];
  assign o[29700] = i[29700];
  assign o[29699] = i[29699];
  assign o[29698] = i[29698];
  assign o[29697] = i[29697];
  assign o[29696] = i[29696];
  assign o[29695] = i[29695];
  assign o[29694] = i[29694];
  assign o[29693] = i[29693];
  assign o[29692] = i[29692];
  assign o[29691] = i[29691];
  assign o[29690] = i[29690];
  assign o[29689] = i[29689];
  assign o[29688] = i[29688];
  assign o[29687] = i[29687];
  assign o[29686] = i[29686];
  assign o[29685] = i[29685];
  assign o[29684] = i[29684];
  assign o[29683] = i[29683];
  assign o[29682] = i[29682];
  assign o[29681] = i[29681];
  assign o[29680] = i[29680];
  assign o[29679] = i[29679];
  assign o[29678] = i[29678];
  assign o[29677] = i[29677];
  assign o[29676] = i[29676];
  assign o[29675] = i[29675];
  assign o[29674] = i[29674];
  assign o[29673] = i[29673];
  assign o[29672] = i[29672];
  assign o[29671] = i[29671];
  assign o[29670] = i[29670];
  assign o[29669] = i[29669];
  assign o[29668] = i[29668];
  assign o[29667] = i[29667];
  assign o[29666] = i[29666];
  assign o[29665] = i[29665];
  assign o[29664] = i[29664];
  assign o[29663] = i[29663];
  assign o[29662] = i[29662];
  assign o[29661] = i[29661];
  assign o[29660] = i[29660];
  assign o[29659] = i[29659];
  assign o[29658] = i[29658];
  assign o[29657] = i[29657];
  assign o[29656] = i[29656];
  assign o[29655] = i[29655];
  assign o[29654] = i[29654];
  assign o[29653] = i[29653];
  assign o[29652] = i[29652];
  assign o[29651] = i[29651];
  assign o[29650] = i[29650];
  assign o[29649] = i[29649];
  assign o[29648] = i[29648];
  assign o[29647] = i[29647];
  assign o[29646] = i[29646];
  assign o[29645] = i[29645];
  assign o[29644] = i[29644];
  assign o[29643] = i[29643];
  assign o[29642] = i[29642];
  assign o[29641] = i[29641];
  assign o[29640] = i[29640];
  assign o[29639] = i[29639];
  assign o[29638] = i[29638];
  assign o[29637] = i[29637];
  assign o[29636] = i[29636];
  assign o[29635] = i[29635];
  assign o[29634] = i[29634];
  assign o[29633] = i[29633];
  assign o[29632] = i[29632];
  assign o[29631] = i[29631];
  assign o[29630] = i[29630];
  assign o[29629] = i[29629];
  assign o[29628] = i[29628];
  assign o[29627] = i[29627];
  assign o[29626] = i[29626];
  assign o[29625] = i[29625];
  assign o[29624] = i[29624];
  assign o[29623] = i[29623];
  assign o[29622] = i[29622];
  assign o[29621] = i[29621];
  assign o[29620] = i[29620];
  assign o[29619] = i[29619];
  assign o[29618] = i[29618];
  assign o[29617] = i[29617];
  assign o[29616] = i[29616];
  assign o[29615] = i[29615];
  assign o[29614] = i[29614];
  assign o[29613] = i[29613];
  assign o[29612] = i[29612];
  assign o[29611] = i[29611];
  assign o[29610] = i[29610];
  assign o[29609] = i[29609];
  assign o[29608] = i[29608];
  assign o[29607] = i[29607];
  assign o[29606] = i[29606];
  assign o[29605] = i[29605];
  assign o[29604] = i[29604];
  assign o[29603] = i[29603];
  assign o[29602] = i[29602];
  assign o[29601] = i[29601];
  assign o[29600] = i[29600];
  assign o[29599] = i[29599];
  assign o[29598] = i[29598];
  assign o[29597] = i[29597];
  assign o[29596] = i[29596];
  assign o[29595] = i[29595];
  assign o[29594] = i[29594];
  assign o[29593] = i[29593];
  assign o[29592] = i[29592];
  assign o[29591] = i[29591];
  assign o[29590] = i[29590];
  assign o[29589] = i[29589];
  assign o[29588] = i[29588];
  assign o[29587] = i[29587];
  assign o[29586] = i[29586];
  assign o[29585] = i[29585];
  assign o[29584] = i[29584];
  assign o[29583] = i[29583];
  assign o[29582] = i[29582];
  assign o[29581] = i[29581];
  assign o[29580] = i[29580];
  assign o[29579] = i[29579];
  assign o[29578] = i[29578];
  assign o[29577] = i[29577];
  assign o[29576] = i[29576];
  assign o[29575] = i[29575];
  assign o[29574] = i[29574];
  assign o[29573] = i[29573];
  assign o[29572] = i[29572];
  assign o[29571] = i[29571];
  assign o[29570] = i[29570];
  assign o[29569] = i[29569];
  assign o[29568] = i[29568];
  assign o[29567] = i[29567];
  assign o[29566] = i[29566];
  assign o[29565] = i[29565];
  assign o[29564] = i[29564];
  assign o[29563] = i[29563];
  assign o[29562] = i[29562];
  assign o[29561] = i[29561];
  assign o[29560] = i[29560];
  assign o[29559] = i[29559];
  assign o[29558] = i[29558];
  assign o[29557] = i[29557];
  assign o[29556] = i[29556];
  assign o[29555] = i[29555];
  assign o[29554] = i[29554];
  assign o[29553] = i[29553];
  assign o[29552] = i[29552];
  assign o[29551] = i[29551];
  assign o[29550] = i[29550];
  assign o[29549] = i[29549];
  assign o[29548] = i[29548];
  assign o[29547] = i[29547];
  assign o[29546] = i[29546];
  assign o[29545] = i[29545];
  assign o[29544] = i[29544];
  assign o[29543] = i[29543];
  assign o[29542] = i[29542];
  assign o[29541] = i[29541];
  assign o[29540] = i[29540];
  assign o[29539] = i[29539];
  assign o[29538] = i[29538];
  assign o[29537] = i[29537];
  assign o[29536] = i[29536];
  assign o[29535] = i[29535];
  assign o[29534] = i[29534];
  assign o[29533] = i[29533];
  assign o[29532] = i[29532];
  assign o[29531] = i[29531];
  assign o[29530] = i[29530];
  assign o[29529] = i[29529];
  assign o[29528] = i[29528];
  assign o[29527] = i[29527];
  assign o[29526] = i[29526];
  assign o[29525] = i[29525];
  assign o[29524] = i[29524];
  assign o[29523] = i[29523];
  assign o[29522] = i[29522];
  assign o[29521] = i[29521];
  assign o[29520] = i[29520];
  assign o[29519] = i[29519];
  assign o[29518] = i[29518];
  assign o[29517] = i[29517];
  assign o[29516] = i[29516];
  assign o[29515] = i[29515];
  assign o[29514] = i[29514];
  assign o[29513] = i[29513];
  assign o[29512] = i[29512];
  assign o[29511] = i[29511];
  assign o[29510] = i[29510];
  assign o[29509] = i[29509];
  assign o[29508] = i[29508];
  assign o[29507] = i[29507];
  assign o[29506] = i[29506];
  assign o[29505] = i[29505];
  assign o[29504] = i[29504];
  assign o[29503] = i[29503];
  assign o[29502] = i[29502];
  assign o[29501] = i[29501];
  assign o[29500] = i[29500];
  assign o[29499] = i[29499];
  assign o[29498] = i[29498];
  assign o[29497] = i[29497];
  assign o[29496] = i[29496];
  assign o[29495] = i[29495];
  assign o[29494] = i[29494];
  assign o[29493] = i[29493];
  assign o[29492] = i[29492];
  assign o[29491] = i[29491];
  assign o[29490] = i[29490];
  assign o[29489] = i[29489];
  assign o[29488] = i[29488];
  assign o[29487] = i[29487];
  assign o[29486] = i[29486];
  assign o[29485] = i[29485];
  assign o[29484] = i[29484];
  assign o[29483] = i[29483];
  assign o[29482] = i[29482];
  assign o[29481] = i[29481];
  assign o[29480] = i[29480];
  assign o[29479] = i[29479];
  assign o[29478] = i[29478];
  assign o[29477] = i[29477];
  assign o[29476] = i[29476];
  assign o[29475] = i[29475];
  assign o[29474] = i[29474];
  assign o[29473] = i[29473];
  assign o[29472] = i[29472];
  assign o[29471] = i[29471];
  assign o[29470] = i[29470];
  assign o[29469] = i[29469];
  assign o[29468] = i[29468];
  assign o[29467] = i[29467];
  assign o[29466] = i[29466];
  assign o[29465] = i[29465];
  assign o[29464] = i[29464];
  assign o[29463] = i[29463];
  assign o[29462] = i[29462];
  assign o[29461] = i[29461];
  assign o[29460] = i[29460];
  assign o[29459] = i[29459];
  assign o[29458] = i[29458];
  assign o[29457] = i[29457];
  assign o[29456] = i[29456];
  assign o[29455] = i[29455];
  assign o[29454] = i[29454];
  assign o[29453] = i[29453];
  assign o[29452] = i[29452];
  assign o[29451] = i[29451];
  assign o[29450] = i[29450];
  assign o[29449] = i[29449];
  assign o[29448] = i[29448];
  assign o[29447] = i[29447];
  assign o[29446] = i[29446];
  assign o[29445] = i[29445];
  assign o[29444] = i[29444];
  assign o[29443] = i[29443];
  assign o[29442] = i[29442];
  assign o[29441] = i[29441];
  assign o[29440] = i[29440];
  assign o[29439] = i[29439];
  assign o[29438] = i[29438];
  assign o[29437] = i[29437];
  assign o[29436] = i[29436];
  assign o[29435] = i[29435];
  assign o[29434] = i[29434];
  assign o[29433] = i[29433];
  assign o[29432] = i[29432];
  assign o[29431] = i[29431];
  assign o[29430] = i[29430];
  assign o[29429] = i[29429];
  assign o[29428] = i[29428];
  assign o[29427] = i[29427];
  assign o[29426] = i[29426];
  assign o[29425] = i[29425];
  assign o[29424] = i[29424];
  assign o[29423] = i[29423];
  assign o[29422] = i[29422];
  assign o[29421] = i[29421];
  assign o[29420] = i[29420];
  assign o[29419] = i[29419];
  assign o[29418] = i[29418];
  assign o[29417] = i[29417];
  assign o[29416] = i[29416];
  assign o[29415] = i[29415];
  assign o[29414] = i[29414];
  assign o[29413] = i[29413];
  assign o[29412] = i[29412];
  assign o[29411] = i[29411];
  assign o[29410] = i[29410];
  assign o[29409] = i[29409];
  assign o[29408] = i[29408];
  assign o[29407] = i[29407];
  assign o[29406] = i[29406];
  assign o[29405] = i[29405];
  assign o[29404] = i[29404];
  assign o[29403] = i[29403];
  assign o[29402] = i[29402];
  assign o[29401] = i[29401];
  assign o[29400] = i[29400];
  assign o[29399] = i[29399];
  assign o[29398] = i[29398];
  assign o[29397] = i[29397];
  assign o[29396] = i[29396];
  assign o[29395] = i[29395];
  assign o[29394] = i[29394];
  assign o[29393] = i[29393];
  assign o[29392] = i[29392];
  assign o[29391] = i[29391];
  assign o[29390] = i[29390];
  assign o[29389] = i[29389];
  assign o[29388] = i[29388];
  assign o[29387] = i[29387];
  assign o[29386] = i[29386];
  assign o[29385] = i[29385];
  assign o[29384] = i[29384];
  assign o[29383] = i[29383];
  assign o[29382] = i[29382];
  assign o[29381] = i[29381];
  assign o[29380] = i[29380];
  assign o[29379] = i[29379];
  assign o[29378] = i[29378];
  assign o[29377] = i[29377];
  assign o[29376] = i[29376];
  assign o[29375] = i[29375];
  assign o[29374] = i[29374];
  assign o[29373] = i[29373];
  assign o[29372] = i[29372];
  assign o[29371] = i[29371];
  assign o[29370] = i[29370];
  assign o[29369] = i[29369];
  assign o[29368] = i[29368];
  assign o[29367] = i[29367];
  assign o[29366] = i[29366];
  assign o[29365] = i[29365];
  assign o[29364] = i[29364];
  assign o[29363] = i[29363];
  assign o[29362] = i[29362];
  assign o[29361] = i[29361];
  assign o[29360] = i[29360];
  assign o[29359] = i[29359];
  assign o[29358] = i[29358];
  assign o[29357] = i[29357];
  assign o[29356] = i[29356];
  assign o[29355] = i[29355];
  assign o[29354] = i[29354];
  assign o[29353] = i[29353];
  assign o[29352] = i[29352];
  assign o[29351] = i[29351];
  assign o[29350] = i[29350];
  assign o[29349] = i[29349];
  assign o[29348] = i[29348];
  assign o[29347] = i[29347];
  assign o[29346] = i[29346];
  assign o[29345] = i[29345];
  assign o[29344] = i[29344];
  assign o[29343] = i[29343];
  assign o[29342] = i[29342];
  assign o[29341] = i[29341];
  assign o[29340] = i[29340];
  assign o[29339] = i[29339];
  assign o[29338] = i[29338];
  assign o[29337] = i[29337];
  assign o[29336] = i[29336];
  assign o[29335] = i[29335];
  assign o[29334] = i[29334];
  assign o[29333] = i[29333];
  assign o[29332] = i[29332];
  assign o[29331] = i[29331];
  assign o[29330] = i[29330];
  assign o[29329] = i[29329];
  assign o[29328] = i[29328];
  assign o[29327] = i[29327];
  assign o[29326] = i[29326];
  assign o[29325] = i[29325];
  assign o[29324] = i[29324];
  assign o[29323] = i[29323];
  assign o[29322] = i[29322];
  assign o[29321] = i[29321];
  assign o[29320] = i[29320];
  assign o[29319] = i[29319];
  assign o[29318] = i[29318];
  assign o[29317] = i[29317];
  assign o[29316] = i[29316];
  assign o[29315] = i[29315];
  assign o[29314] = i[29314];
  assign o[29313] = i[29313];
  assign o[29312] = i[29312];
  assign o[29311] = i[29311];
  assign o[29310] = i[29310];
  assign o[29309] = i[29309];
  assign o[29308] = i[29308];
  assign o[29307] = i[29307];
  assign o[29306] = i[29306];
  assign o[29305] = i[29305];
  assign o[29304] = i[29304];
  assign o[29303] = i[29303];
  assign o[29302] = i[29302];
  assign o[29301] = i[29301];
  assign o[29300] = i[29300];
  assign o[29299] = i[29299];
  assign o[29298] = i[29298];
  assign o[29297] = i[29297];
  assign o[29296] = i[29296];
  assign o[29295] = i[29295];
  assign o[29294] = i[29294];
  assign o[29293] = i[29293];
  assign o[29292] = i[29292];
  assign o[29291] = i[29291];
  assign o[29290] = i[29290];
  assign o[29289] = i[29289];
  assign o[29288] = i[29288];
  assign o[29287] = i[29287];
  assign o[29286] = i[29286];
  assign o[29285] = i[29285];
  assign o[29284] = i[29284];
  assign o[29283] = i[29283];
  assign o[29282] = i[29282];
  assign o[29281] = i[29281];
  assign o[29280] = i[29280];
  assign o[29279] = i[29279];
  assign o[29278] = i[29278];
  assign o[29277] = i[29277];
  assign o[29276] = i[29276];
  assign o[29275] = i[29275];
  assign o[29274] = i[29274];
  assign o[29273] = i[29273];
  assign o[29272] = i[29272];
  assign o[29271] = i[29271];
  assign o[29270] = i[29270];
  assign o[29269] = i[29269];
  assign o[29268] = i[29268];
  assign o[29267] = i[29267];
  assign o[29266] = i[29266];
  assign o[29265] = i[29265];
  assign o[29264] = i[29264];
  assign o[29263] = i[29263];
  assign o[29262] = i[29262];
  assign o[29261] = i[29261];
  assign o[29260] = i[29260];
  assign o[29259] = i[29259];
  assign o[29258] = i[29258];
  assign o[29257] = i[29257];
  assign o[29256] = i[29256];
  assign o[29255] = i[29255];
  assign o[29254] = i[29254];
  assign o[29253] = i[29253];
  assign o[29252] = i[29252];
  assign o[29251] = i[29251];
  assign o[29250] = i[29250];
  assign o[29249] = i[29249];
  assign o[29248] = i[29248];
  assign o[29247] = i[29247];
  assign o[29246] = i[29246];
  assign o[29245] = i[29245];
  assign o[29244] = i[29244];
  assign o[29243] = i[29243];
  assign o[29242] = i[29242];
  assign o[29241] = i[29241];
  assign o[29240] = i[29240];
  assign o[29239] = i[29239];
  assign o[29238] = i[29238];
  assign o[29237] = i[29237];
  assign o[29236] = i[29236];
  assign o[29235] = i[29235];
  assign o[29234] = i[29234];
  assign o[29233] = i[29233];
  assign o[29232] = i[29232];
  assign o[29231] = i[29231];
  assign o[29230] = i[29230];
  assign o[29229] = i[29229];
  assign o[29228] = i[29228];
  assign o[29227] = i[29227];
  assign o[29226] = i[29226];
  assign o[29225] = i[29225];
  assign o[29224] = i[29224];
  assign o[29223] = i[29223];
  assign o[29222] = i[29222];
  assign o[29221] = i[29221];
  assign o[29220] = i[29220];
  assign o[29219] = i[29219];
  assign o[29218] = i[29218];
  assign o[29217] = i[29217];
  assign o[29216] = i[29216];
  assign o[29215] = i[29215];
  assign o[29214] = i[29214];
  assign o[29213] = i[29213];
  assign o[29212] = i[29212];
  assign o[29211] = i[29211];
  assign o[29210] = i[29210];
  assign o[29209] = i[29209];
  assign o[29208] = i[29208];
  assign o[29207] = i[29207];
  assign o[29206] = i[29206];
  assign o[29205] = i[29205];
  assign o[29204] = i[29204];
  assign o[29203] = i[29203];
  assign o[29202] = i[29202];
  assign o[29201] = i[29201];
  assign o[29200] = i[29200];
  assign o[29199] = i[29199];
  assign o[29198] = i[29198];
  assign o[29197] = i[29197];
  assign o[29196] = i[29196];
  assign o[29195] = i[29195];
  assign o[29194] = i[29194];
  assign o[29193] = i[29193];
  assign o[29192] = i[29192];
  assign o[29191] = i[29191];
  assign o[29190] = i[29190];
  assign o[29189] = i[29189];
  assign o[29188] = i[29188];
  assign o[29187] = i[29187];
  assign o[29186] = i[29186];
  assign o[29185] = i[29185];
  assign o[29184] = i[29184];
  assign o[29183] = i[29183];
  assign o[29182] = i[29182];
  assign o[29181] = i[29181];
  assign o[29180] = i[29180];
  assign o[29179] = i[29179];
  assign o[29178] = i[29178];
  assign o[29177] = i[29177];
  assign o[29176] = i[29176];
  assign o[29175] = i[29175];
  assign o[29174] = i[29174];
  assign o[29173] = i[29173];
  assign o[29172] = i[29172];
  assign o[29171] = i[29171];
  assign o[29170] = i[29170];
  assign o[29169] = i[29169];
  assign o[29168] = i[29168];
  assign o[29167] = i[29167];
  assign o[29166] = i[29166];
  assign o[29165] = i[29165];
  assign o[29164] = i[29164];
  assign o[29163] = i[29163];
  assign o[29162] = i[29162];
  assign o[29161] = i[29161];
  assign o[29160] = i[29160];
  assign o[29159] = i[29159];
  assign o[29158] = i[29158];
  assign o[29157] = i[29157];
  assign o[29156] = i[29156];
  assign o[29155] = i[29155];
  assign o[29154] = i[29154];
  assign o[29153] = i[29153];
  assign o[29152] = i[29152];
  assign o[29151] = i[29151];
  assign o[29150] = i[29150];
  assign o[29149] = i[29149];
  assign o[29148] = i[29148];
  assign o[29147] = i[29147];
  assign o[29146] = i[29146];
  assign o[29145] = i[29145];
  assign o[29144] = i[29144];
  assign o[29143] = i[29143];
  assign o[29142] = i[29142];
  assign o[29141] = i[29141];
  assign o[29140] = i[29140];
  assign o[29139] = i[29139];
  assign o[29138] = i[29138];
  assign o[29137] = i[29137];
  assign o[29136] = i[29136];
  assign o[29135] = i[29135];
  assign o[29134] = i[29134];
  assign o[29133] = i[29133];
  assign o[29132] = i[29132];
  assign o[29131] = i[29131];
  assign o[29130] = i[29130];
  assign o[29129] = i[29129];
  assign o[29128] = i[29128];
  assign o[29127] = i[29127];
  assign o[29126] = i[29126];
  assign o[29125] = i[29125];
  assign o[29124] = i[29124];
  assign o[29123] = i[29123];
  assign o[29122] = i[29122];
  assign o[29121] = i[29121];
  assign o[29120] = i[29120];
  assign o[29119] = i[29119];
  assign o[29118] = i[29118];
  assign o[29117] = i[29117];
  assign o[29116] = i[29116];
  assign o[29115] = i[29115];
  assign o[29114] = i[29114];
  assign o[29113] = i[29113];
  assign o[29112] = i[29112];
  assign o[29111] = i[29111];
  assign o[29110] = i[29110];
  assign o[29109] = i[29109];
  assign o[29108] = i[29108];
  assign o[29107] = i[29107];
  assign o[29106] = i[29106];
  assign o[29105] = i[29105];
  assign o[29104] = i[29104];
  assign o[29103] = i[29103];
  assign o[29102] = i[29102];
  assign o[29101] = i[29101];
  assign o[29100] = i[29100];
  assign o[29099] = i[29099];
  assign o[29098] = i[29098];
  assign o[29097] = i[29097];
  assign o[29096] = i[29096];
  assign o[29095] = i[29095];
  assign o[29094] = i[29094];
  assign o[29093] = i[29093];
  assign o[29092] = i[29092];
  assign o[29091] = i[29091];
  assign o[29090] = i[29090];
  assign o[29089] = i[29089];
  assign o[29088] = i[29088];
  assign o[29087] = i[29087];
  assign o[29086] = i[29086];
  assign o[29085] = i[29085];
  assign o[29084] = i[29084];
  assign o[29083] = i[29083];
  assign o[29082] = i[29082];
  assign o[29081] = i[29081];
  assign o[29080] = i[29080];
  assign o[29079] = i[29079];
  assign o[29078] = i[29078];
  assign o[29077] = i[29077];
  assign o[29076] = i[29076];
  assign o[29075] = i[29075];
  assign o[29074] = i[29074];
  assign o[29073] = i[29073];
  assign o[29072] = i[29072];
  assign o[29071] = i[29071];
  assign o[29070] = i[29070];
  assign o[29069] = i[29069];
  assign o[29068] = i[29068];
  assign o[29067] = i[29067];
  assign o[29066] = i[29066];
  assign o[29065] = i[29065];
  assign o[29064] = i[29064];
  assign o[29063] = i[29063];
  assign o[29062] = i[29062];
  assign o[29061] = i[29061];
  assign o[29060] = i[29060];
  assign o[29059] = i[29059];
  assign o[29058] = i[29058];
  assign o[29057] = i[29057];
  assign o[29056] = i[29056];
  assign o[29055] = i[29055];
  assign o[29054] = i[29054];
  assign o[29053] = i[29053];
  assign o[29052] = i[29052];
  assign o[29051] = i[29051];
  assign o[29050] = i[29050];
  assign o[29049] = i[29049];
  assign o[29048] = i[29048];
  assign o[29047] = i[29047];
  assign o[29046] = i[29046];
  assign o[29045] = i[29045];
  assign o[29044] = i[29044];
  assign o[29043] = i[29043];
  assign o[29042] = i[29042];
  assign o[29041] = i[29041];
  assign o[29040] = i[29040];
  assign o[29039] = i[29039];
  assign o[29038] = i[29038];
  assign o[29037] = i[29037];
  assign o[29036] = i[29036];
  assign o[29035] = i[29035];
  assign o[29034] = i[29034];
  assign o[29033] = i[29033];
  assign o[29032] = i[29032];
  assign o[29031] = i[29031];
  assign o[29030] = i[29030];
  assign o[29029] = i[29029];
  assign o[29028] = i[29028];
  assign o[29027] = i[29027];
  assign o[29026] = i[29026];
  assign o[29025] = i[29025];
  assign o[29024] = i[29024];
  assign o[29023] = i[29023];
  assign o[29022] = i[29022];
  assign o[29021] = i[29021];
  assign o[29020] = i[29020];
  assign o[29019] = i[29019];
  assign o[29018] = i[29018];
  assign o[29017] = i[29017];
  assign o[29016] = i[29016];
  assign o[29015] = i[29015];
  assign o[29014] = i[29014];
  assign o[29013] = i[29013];
  assign o[29012] = i[29012];
  assign o[29011] = i[29011];
  assign o[29010] = i[29010];
  assign o[29009] = i[29009];
  assign o[29008] = i[29008];
  assign o[29007] = i[29007];
  assign o[29006] = i[29006];
  assign o[29005] = i[29005];
  assign o[29004] = i[29004];
  assign o[29003] = i[29003];
  assign o[29002] = i[29002];
  assign o[29001] = i[29001];
  assign o[29000] = i[29000];
  assign o[28999] = i[28999];
  assign o[28998] = i[28998];
  assign o[28997] = i[28997];
  assign o[28996] = i[28996];
  assign o[28995] = i[28995];
  assign o[28994] = i[28994];
  assign o[28993] = i[28993];
  assign o[28992] = i[28992];
  assign o[28991] = i[28991];
  assign o[28990] = i[28990];
  assign o[28989] = i[28989];
  assign o[28988] = i[28988];
  assign o[28987] = i[28987];
  assign o[28986] = i[28986];
  assign o[28985] = i[28985];
  assign o[28984] = i[28984];
  assign o[28983] = i[28983];
  assign o[28982] = i[28982];
  assign o[28981] = i[28981];
  assign o[28980] = i[28980];
  assign o[28979] = i[28979];
  assign o[28978] = i[28978];
  assign o[28977] = i[28977];
  assign o[28976] = i[28976];
  assign o[28975] = i[28975];
  assign o[28974] = i[28974];
  assign o[28973] = i[28973];
  assign o[28972] = i[28972];
  assign o[28971] = i[28971];
  assign o[28970] = i[28970];
  assign o[28969] = i[28969];
  assign o[28968] = i[28968];
  assign o[28967] = i[28967];
  assign o[28966] = i[28966];
  assign o[28965] = i[28965];
  assign o[28964] = i[28964];
  assign o[28963] = i[28963];
  assign o[28962] = i[28962];
  assign o[28961] = i[28961];
  assign o[28960] = i[28960];
  assign o[28959] = i[28959];
  assign o[28958] = i[28958];
  assign o[28957] = i[28957];
  assign o[28956] = i[28956];
  assign o[28955] = i[28955];
  assign o[28954] = i[28954];
  assign o[28953] = i[28953];
  assign o[28952] = i[28952];
  assign o[28951] = i[28951];
  assign o[28950] = i[28950];
  assign o[28949] = i[28949];
  assign o[28948] = i[28948];
  assign o[28947] = i[28947];
  assign o[28946] = i[28946];
  assign o[28945] = i[28945];
  assign o[28944] = i[28944];
  assign o[28943] = i[28943];
  assign o[28942] = i[28942];
  assign o[28941] = i[28941];
  assign o[28940] = i[28940];
  assign o[28939] = i[28939];
  assign o[28938] = i[28938];
  assign o[28937] = i[28937];
  assign o[28936] = i[28936];
  assign o[28935] = i[28935];
  assign o[28934] = i[28934];
  assign o[28933] = i[28933];
  assign o[28932] = i[28932];
  assign o[28931] = i[28931];
  assign o[28930] = i[28930];
  assign o[28929] = i[28929];
  assign o[28928] = i[28928];
  assign o[28927] = i[28927];
  assign o[28926] = i[28926];
  assign o[28925] = i[28925];
  assign o[28924] = i[28924];
  assign o[28923] = i[28923];
  assign o[28922] = i[28922];
  assign o[28921] = i[28921];
  assign o[28920] = i[28920];
  assign o[28919] = i[28919];
  assign o[28918] = i[28918];
  assign o[28917] = i[28917];
  assign o[28916] = i[28916];
  assign o[28915] = i[28915];
  assign o[28914] = i[28914];
  assign o[28913] = i[28913];
  assign o[28912] = i[28912];
  assign o[28911] = i[28911];
  assign o[28910] = i[28910];
  assign o[28909] = i[28909];
  assign o[28908] = i[28908];
  assign o[28907] = i[28907];
  assign o[28906] = i[28906];
  assign o[28905] = i[28905];
  assign o[28904] = i[28904];
  assign o[28903] = i[28903];
  assign o[28902] = i[28902];
  assign o[28901] = i[28901];
  assign o[28900] = i[28900];
  assign o[28899] = i[28899];
  assign o[28898] = i[28898];
  assign o[28897] = i[28897];
  assign o[28896] = i[28896];
  assign o[28895] = i[28895];
  assign o[28894] = i[28894];
  assign o[28893] = i[28893];
  assign o[28892] = i[28892];
  assign o[28891] = i[28891];
  assign o[28890] = i[28890];
  assign o[28889] = i[28889];
  assign o[28888] = i[28888];
  assign o[28887] = i[28887];
  assign o[28886] = i[28886];
  assign o[28885] = i[28885];
  assign o[28884] = i[28884];
  assign o[28883] = i[28883];
  assign o[28882] = i[28882];
  assign o[28881] = i[28881];
  assign o[28880] = i[28880];
  assign o[28879] = i[28879];
  assign o[28878] = i[28878];
  assign o[28877] = i[28877];
  assign o[28876] = i[28876];
  assign o[28875] = i[28875];
  assign o[28874] = i[28874];
  assign o[28873] = i[28873];
  assign o[28872] = i[28872];
  assign o[28871] = i[28871];
  assign o[28870] = i[28870];
  assign o[28869] = i[28869];
  assign o[28868] = i[28868];
  assign o[28867] = i[28867];
  assign o[28866] = i[28866];
  assign o[28865] = i[28865];
  assign o[28864] = i[28864];
  assign o[28863] = i[28863];
  assign o[28862] = i[28862];
  assign o[28861] = i[28861];
  assign o[28860] = i[28860];
  assign o[28859] = i[28859];
  assign o[28858] = i[28858];
  assign o[28857] = i[28857];
  assign o[28856] = i[28856];
  assign o[28855] = i[28855];
  assign o[28854] = i[28854];
  assign o[28853] = i[28853];
  assign o[28852] = i[28852];
  assign o[28851] = i[28851];
  assign o[28850] = i[28850];
  assign o[28849] = i[28849];
  assign o[28848] = i[28848];
  assign o[28847] = i[28847];
  assign o[28846] = i[28846];
  assign o[28845] = i[28845];
  assign o[28844] = i[28844];
  assign o[28843] = i[28843];
  assign o[28842] = i[28842];
  assign o[28841] = i[28841];
  assign o[28840] = i[28840];
  assign o[28839] = i[28839];
  assign o[28838] = i[28838];
  assign o[28837] = i[28837];
  assign o[28836] = i[28836];
  assign o[28835] = i[28835];
  assign o[28834] = i[28834];
  assign o[28833] = i[28833];
  assign o[28832] = i[28832];
  assign o[28831] = i[28831];
  assign o[28830] = i[28830];
  assign o[28829] = i[28829];
  assign o[28828] = i[28828];
  assign o[28827] = i[28827];
  assign o[28826] = i[28826];
  assign o[28825] = i[28825];
  assign o[28824] = i[28824];
  assign o[28823] = i[28823];
  assign o[28822] = i[28822];
  assign o[28821] = i[28821];
  assign o[28820] = i[28820];
  assign o[28819] = i[28819];
  assign o[28818] = i[28818];
  assign o[28817] = i[28817];
  assign o[28816] = i[28816];
  assign o[28815] = i[28815];
  assign o[28814] = i[28814];
  assign o[28813] = i[28813];
  assign o[28812] = i[28812];
  assign o[28811] = i[28811];
  assign o[28810] = i[28810];
  assign o[28809] = i[28809];
  assign o[28808] = i[28808];
  assign o[28807] = i[28807];
  assign o[28806] = i[28806];
  assign o[28805] = i[28805];
  assign o[28804] = i[28804];
  assign o[28803] = i[28803];
  assign o[28802] = i[28802];
  assign o[28801] = i[28801];
  assign o[28800] = i[28800];
  assign o[28799] = i[28799];
  assign o[28798] = i[28798];
  assign o[28797] = i[28797];
  assign o[28796] = i[28796];
  assign o[28795] = i[28795];
  assign o[28794] = i[28794];
  assign o[28793] = i[28793];
  assign o[28792] = i[28792];
  assign o[28791] = i[28791];
  assign o[28790] = i[28790];
  assign o[28789] = i[28789];
  assign o[28788] = i[28788];
  assign o[28787] = i[28787];
  assign o[28786] = i[28786];
  assign o[28785] = i[28785];
  assign o[28784] = i[28784];
  assign o[28783] = i[28783];
  assign o[28782] = i[28782];
  assign o[28781] = i[28781];
  assign o[28780] = i[28780];
  assign o[28779] = i[28779];
  assign o[28778] = i[28778];
  assign o[28777] = i[28777];
  assign o[28776] = i[28776];
  assign o[28775] = i[28775];
  assign o[28774] = i[28774];
  assign o[28773] = i[28773];
  assign o[28772] = i[28772];
  assign o[28771] = i[28771];
  assign o[28770] = i[28770];
  assign o[28769] = i[28769];
  assign o[28768] = i[28768];
  assign o[28767] = i[28767];
  assign o[28766] = i[28766];
  assign o[28765] = i[28765];
  assign o[28764] = i[28764];
  assign o[28763] = i[28763];
  assign o[28762] = i[28762];
  assign o[28761] = i[28761];
  assign o[28760] = i[28760];
  assign o[28759] = i[28759];
  assign o[28758] = i[28758];
  assign o[28757] = i[28757];
  assign o[28756] = i[28756];
  assign o[28755] = i[28755];
  assign o[28754] = i[28754];
  assign o[28753] = i[28753];
  assign o[28752] = i[28752];
  assign o[28751] = i[28751];
  assign o[28750] = i[28750];
  assign o[28749] = i[28749];
  assign o[28748] = i[28748];
  assign o[28747] = i[28747];
  assign o[28746] = i[28746];
  assign o[28745] = i[28745];
  assign o[28744] = i[28744];
  assign o[28743] = i[28743];
  assign o[28742] = i[28742];
  assign o[28741] = i[28741];
  assign o[28740] = i[28740];
  assign o[28739] = i[28739];
  assign o[28738] = i[28738];
  assign o[28737] = i[28737];
  assign o[28736] = i[28736];
  assign o[28735] = i[28735];
  assign o[28734] = i[28734];
  assign o[28733] = i[28733];
  assign o[28732] = i[28732];
  assign o[28731] = i[28731];
  assign o[28730] = i[28730];
  assign o[28729] = i[28729];
  assign o[28728] = i[28728];
  assign o[28727] = i[28727];
  assign o[28726] = i[28726];
  assign o[28725] = i[28725];
  assign o[28724] = i[28724];
  assign o[28723] = i[28723];
  assign o[28722] = i[28722];
  assign o[28721] = i[28721];
  assign o[28720] = i[28720];
  assign o[28719] = i[28719];
  assign o[28718] = i[28718];
  assign o[28717] = i[28717];
  assign o[28716] = i[28716];
  assign o[28715] = i[28715];
  assign o[28714] = i[28714];
  assign o[28713] = i[28713];
  assign o[28712] = i[28712];
  assign o[28711] = i[28711];
  assign o[28710] = i[28710];
  assign o[28709] = i[28709];
  assign o[28708] = i[28708];
  assign o[28707] = i[28707];
  assign o[28706] = i[28706];
  assign o[28705] = i[28705];
  assign o[28704] = i[28704];
  assign o[28703] = i[28703];
  assign o[28702] = i[28702];
  assign o[28701] = i[28701];
  assign o[28700] = i[28700];
  assign o[28699] = i[28699];
  assign o[28698] = i[28698];
  assign o[28697] = i[28697];
  assign o[28696] = i[28696];
  assign o[28695] = i[28695];
  assign o[28694] = i[28694];
  assign o[28693] = i[28693];
  assign o[28692] = i[28692];
  assign o[28691] = i[28691];
  assign o[28690] = i[28690];
  assign o[28689] = i[28689];
  assign o[28688] = i[28688];
  assign o[28687] = i[28687];
  assign o[28686] = i[28686];
  assign o[28685] = i[28685];
  assign o[28684] = i[28684];
  assign o[28683] = i[28683];
  assign o[28682] = i[28682];
  assign o[28681] = i[28681];
  assign o[28680] = i[28680];
  assign o[28679] = i[28679];
  assign o[28678] = i[28678];
  assign o[28677] = i[28677];
  assign o[28676] = i[28676];
  assign o[28675] = i[28675];
  assign o[28674] = i[28674];
  assign o[28673] = i[28673];
  assign o[28672] = i[28672];
  assign o[28671] = i[28671];
  assign o[28670] = i[28670];
  assign o[28669] = i[28669];
  assign o[28668] = i[28668];
  assign o[28667] = i[28667];
  assign o[28666] = i[28666];
  assign o[28665] = i[28665];
  assign o[28664] = i[28664];
  assign o[28663] = i[28663];
  assign o[28662] = i[28662];
  assign o[28661] = i[28661];
  assign o[28660] = i[28660];
  assign o[28659] = i[28659];
  assign o[28658] = i[28658];
  assign o[28657] = i[28657];
  assign o[28656] = i[28656];
  assign o[28655] = i[28655];
  assign o[28654] = i[28654];
  assign o[28653] = i[28653];
  assign o[28652] = i[28652];
  assign o[28651] = i[28651];
  assign o[28650] = i[28650];
  assign o[28649] = i[28649];
  assign o[28648] = i[28648];
  assign o[28647] = i[28647];
  assign o[28646] = i[28646];
  assign o[28645] = i[28645];
  assign o[28644] = i[28644];
  assign o[28643] = i[28643];
  assign o[28642] = i[28642];
  assign o[28641] = i[28641];
  assign o[28640] = i[28640];
  assign o[28639] = i[28639];
  assign o[28638] = i[28638];
  assign o[28637] = i[28637];
  assign o[28636] = i[28636];
  assign o[28635] = i[28635];
  assign o[28634] = i[28634];
  assign o[28633] = i[28633];
  assign o[28632] = i[28632];
  assign o[28631] = i[28631];
  assign o[28630] = i[28630];
  assign o[28629] = i[28629];
  assign o[28628] = i[28628];
  assign o[28627] = i[28627];
  assign o[28626] = i[28626];
  assign o[28625] = i[28625];
  assign o[28624] = i[28624];
  assign o[28623] = i[28623];
  assign o[28622] = i[28622];
  assign o[28621] = i[28621];
  assign o[28620] = i[28620];
  assign o[28619] = i[28619];
  assign o[28618] = i[28618];
  assign o[28617] = i[28617];
  assign o[28616] = i[28616];
  assign o[28615] = i[28615];
  assign o[28614] = i[28614];
  assign o[28613] = i[28613];
  assign o[28612] = i[28612];
  assign o[28611] = i[28611];
  assign o[28610] = i[28610];
  assign o[28609] = i[28609];
  assign o[28608] = i[28608];
  assign o[28607] = i[28607];
  assign o[28606] = i[28606];
  assign o[28605] = i[28605];
  assign o[28604] = i[28604];
  assign o[28603] = i[28603];
  assign o[28602] = i[28602];
  assign o[28601] = i[28601];
  assign o[28600] = i[28600];
  assign o[28599] = i[28599];
  assign o[28598] = i[28598];
  assign o[28597] = i[28597];
  assign o[28596] = i[28596];
  assign o[28595] = i[28595];
  assign o[28594] = i[28594];
  assign o[28593] = i[28593];
  assign o[28592] = i[28592];
  assign o[28591] = i[28591];
  assign o[28590] = i[28590];
  assign o[28589] = i[28589];
  assign o[28588] = i[28588];
  assign o[28587] = i[28587];
  assign o[28586] = i[28586];
  assign o[28585] = i[28585];
  assign o[28584] = i[28584];
  assign o[28583] = i[28583];
  assign o[28582] = i[28582];
  assign o[28581] = i[28581];
  assign o[28580] = i[28580];
  assign o[28579] = i[28579];
  assign o[28578] = i[28578];
  assign o[28577] = i[28577];
  assign o[28576] = i[28576];
  assign o[28575] = i[28575];
  assign o[28574] = i[28574];
  assign o[28573] = i[28573];
  assign o[28572] = i[28572];
  assign o[28571] = i[28571];
  assign o[28570] = i[28570];
  assign o[28569] = i[28569];
  assign o[28568] = i[28568];
  assign o[28567] = i[28567];
  assign o[28566] = i[28566];
  assign o[28565] = i[28565];
  assign o[28564] = i[28564];
  assign o[28563] = i[28563];
  assign o[28562] = i[28562];
  assign o[28561] = i[28561];
  assign o[28560] = i[28560];
  assign o[28559] = i[28559];
  assign o[28558] = i[28558];
  assign o[28557] = i[28557];
  assign o[28556] = i[28556];
  assign o[28555] = i[28555];
  assign o[28554] = i[28554];
  assign o[28553] = i[28553];
  assign o[28552] = i[28552];
  assign o[28551] = i[28551];
  assign o[28550] = i[28550];
  assign o[28549] = i[28549];
  assign o[28548] = i[28548];
  assign o[28547] = i[28547];
  assign o[28546] = i[28546];
  assign o[28545] = i[28545];
  assign o[28544] = i[28544];
  assign o[28543] = i[28543];
  assign o[28542] = i[28542];
  assign o[28541] = i[28541];
  assign o[28540] = i[28540];
  assign o[28539] = i[28539];
  assign o[28538] = i[28538];
  assign o[28537] = i[28537];
  assign o[28536] = i[28536];
  assign o[28535] = i[28535];
  assign o[28534] = i[28534];
  assign o[28533] = i[28533];
  assign o[28532] = i[28532];
  assign o[28531] = i[28531];
  assign o[28530] = i[28530];
  assign o[28529] = i[28529];
  assign o[28528] = i[28528];
  assign o[28527] = i[28527];
  assign o[28526] = i[28526];
  assign o[28525] = i[28525];
  assign o[28524] = i[28524];
  assign o[28523] = i[28523];
  assign o[28522] = i[28522];
  assign o[28521] = i[28521];
  assign o[28520] = i[28520];
  assign o[28519] = i[28519];
  assign o[28518] = i[28518];
  assign o[28517] = i[28517];
  assign o[28516] = i[28516];
  assign o[28515] = i[28515];
  assign o[28514] = i[28514];
  assign o[28513] = i[28513];
  assign o[28512] = i[28512];
  assign o[28511] = i[28511];
  assign o[28510] = i[28510];
  assign o[28509] = i[28509];
  assign o[28508] = i[28508];
  assign o[28507] = i[28507];
  assign o[28506] = i[28506];
  assign o[28505] = i[28505];
  assign o[28504] = i[28504];
  assign o[28503] = i[28503];
  assign o[28502] = i[28502];
  assign o[28501] = i[28501];
  assign o[28500] = i[28500];
  assign o[28499] = i[28499];
  assign o[28498] = i[28498];
  assign o[28497] = i[28497];
  assign o[28496] = i[28496];
  assign o[28495] = i[28495];
  assign o[28494] = i[28494];
  assign o[28493] = i[28493];
  assign o[28492] = i[28492];
  assign o[28491] = i[28491];
  assign o[28490] = i[28490];
  assign o[28489] = i[28489];
  assign o[28488] = i[28488];
  assign o[28487] = i[28487];
  assign o[28486] = i[28486];
  assign o[28485] = i[28485];
  assign o[28484] = i[28484];
  assign o[28483] = i[28483];
  assign o[28482] = i[28482];
  assign o[28481] = i[28481];
  assign o[28480] = i[28480];
  assign o[28479] = i[28479];
  assign o[28478] = i[28478];
  assign o[28477] = i[28477];
  assign o[28476] = i[28476];
  assign o[28475] = i[28475];
  assign o[28474] = i[28474];
  assign o[28473] = i[28473];
  assign o[28472] = i[28472];
  assign o[28471] = i[28471];
  assign o[28470] = i[28470];
  assign o[28469] = i[28469];
  assign o[28468] = i[28468];
  assign o[28467] = i[28467];
  assign o[28466] = i[28466];
  assign o[28465] = i[28465];
  assign o[28464] = i[28464];
  assign o[28463] = i[28463];
  assign o[28462] = i[28462];
  assign o[28461] = i[28461];
  assign o[28460] = i[28460];
  assign o[28459] = i[28459];
  assign o[28458] = i[28458];
  assign o[28457] = i[28457];
  assign o[28456] = i[28456];
  assign o[28455] = i[28455];
  assign o[28454] = i[28454];
  assign o[28453] = i[28453];
  assign o[28452] = i[28452];
  assign o[28451] = i[28451];
  assign o[28450] = i[28450];
  assign o[28449] = i[28449];
  assign o[28448] = i[28448];
  assign o[28447] = i[28447];
  assign o[28446] = i[28446];
  assign o[28445] = i[28445];
  assign o[28444] = i[28444];
  assign o[28443] = i[28443];
  assign o[28442] = i[28442];
  assign o[28441] = i[28441];
  assign o[28440] = i[28440];
  assign o[28439] = i[28439];
  assign o[28438] = i[28438];
  assign o[28437] = i[28437];
  assign o[28436] = i[28436];
  assign o[28435] = i[28435];
  assign o[28434] = i[28434];
  assign o[28433] = i[28433];
  assign o[28432] = i[28432];
  assign o[28431] = i[28431];
  assign o[28430] = i[28430];
  assign o[28429] = i[28429];
  assign o[28428] = i[28428];
  assign o[28427] = i[28427];
  assign o[28426] = i[28426];
  assign o[28425] = i[28425];
  assign o[28424] = i[28424];
  assign o[28423] = i[28423];
  assign o[28422] = i[28422];
  assign o[28421] = i[28421];
  assign o[28420] = i[28420];
  assign o[28419] = i[28419];
  assign o[28418] = i[28418];
  assign o[28417] = i[28417];
  assign o[28416] = i[28416];
  assign o[28415] = i[28415];
  assign o[28414] = i[28414];
  assign o[28413] = i[28413];
  assign o[28412] = i[28412];
  assign o[28411] = i[28411];
  assign o[28410] = i[28410];
  assign o[28409] = i[28409];
  assign o[28408] = i[28408];
  assign o[28407] = i[28407];
  assign o[28406] = i[28406];
  assign o[28405] = i[28405];
  assign o[28404] = i[28404];
  assign o[28403] = i[28403];
  assign o[28402] = i[28402];
  assign o[28401] = i[28401];
  assign o[28400] = i[28400];
  assign o[28399] = i[28399];
  assign o[28398] = i[28398];
  assign o[28397] = i[28397];
  assign o[28396] = i[28396];
  assign o[28395] = i[28395];
  assign o[28394] = i[28394];
  assign o[28393] = i[28393];
  assign o[28392] = i[28392];
  assign o[28391] = i[28391];
  assign o[28390] = i[28390];
  assign o[28389] = i[28389];
  assign o[28388] = i[28388];
  assign o[28387] = i[28387];
  assign o[28386] = i[28386];
  assign o[28385] = i[28385];
  assign o[28384] = i[28384];
  assign o[28383] = i[28383];
  assign o[28382] = i[28382];
  assign o[28381] = i[28381];
  assign o[28380] = i[28380];
  assign o[28379] = i[28379];
  assign o[28378] = i[28378];
  assign o[28377] = i[28377];
  assign o[28376] = i[28376];
  assign o[28375] = i[28375];
  assign o[28374] = i[28374];
  assign o[28373] = i[28373];
  assign o[28372] = i[28372];
  assign o[28371] = i[28371];
  assign o[28370] = i[28370];
  assign o[28369] = i[28369];
  assign o[28368] = i[28368];
  assign o[28367] = i[28367];
  assign o[28366] = i[28366];
  assign o[28365] = i[28365];
  assign o[28364] = i[28364];
  assign o[28363] = i[28363];
  assign o[28362] = i[28362];
  assign o[28361] = i[28361];
  assign o[28360] = i[28360];
  assign o[28359] = i[28359];
  assign o[28358] = i[28358];
  assign o[28357] = i[28357];
  assign o[28356] = i[28356];
  assign o[28355] = i[28355];
  assign o[28354] = i[28354];
  assign o[28353] = i[28353];
  assign o[28352] = i[28352];
  assign o[28351] = i[28351];
  assign o[28350] = i[28350];
  assign o[28349] = i[28349];
  assign o[28348] = i[28348];
  assign o[28347] = i[28347];
  assign o[28346] = i[28346];
  assign o[28345] = i[28345];
  assign o[28344] = i[28344];
  assign o[28343] = i[28343];
  assign o[28342] = i[28342];
  assign o[28341] = i[28341];
  assign o[28340] = i[28340];
  assign o[28339] = i[28339];
  assign o[28338] = i[28338];
  assign o[28337] = i[28337];
  assign o[28336] = i[28336];
  assign o[28335] = i[28335];
  assign o[28334] = i[28334];
  assign o[28333] = i[28333];
  assign o[28332] = i[28332];
  assign o[28331] = i[28331];
  assign o[28330] = i[28330];
  assign o[28329] = i[28329];
  assign o[28328] = i[28328];
  assign o[28327] = i[28327];
  assign o[28326] = i[28326];
  assign o[28325] = i[28325];
  assign o[28324] = i[28324];
  assign o[28323] = i[28323];
  assign o[28322] = i[28322];
  assign o[28321] = i[28321];
  assign o[28320] = i[28320];
  assign o[28319] = i[28319];
  assign o[28318] = i[28318];
  assign o[28317] = i[28317];
  assign o[28316] = i[28316];
  assign o[28315] = i[28315];
  assign o[28314] = i[28314];
  assign o[28313] = i[28313];
  assign o[28312] = i[28312];
  assign o[28311] = i[28311];
  assign o[28310] = i[28310];
  assign o[28309] = i[28309];
  assign o[28308] = i[28308];
  assign o[28307] = i[28307];
  assign o[28306] = i[28306];
  assign o[28305] = i[28305];
  assign o[28304] = i[28304];
  assign o[28303] = i[28303];
  assign o[28302] = i[28302];
  assign o[28301] = i[28301];
  assign o[28300] = i[28300];
  assign o[28299] = i[28299];
  assign o[28298] = i[28298];
  assign o[28297] = i[28297];
  assign o[28296] = i[28296];
  assign o[28295] = i[28295];
  assign o[28294] = i[28294];
  assign o[28293] = i[28293];
  assign o[28292] = i[28292];
  assign o[28291] = i[28291];
  assign o[28290] = i[28290];
  assign o[28289] = i[28289];
  assign o[28288] = i[28288];
  assign o[28287] = i[28287];
  assign o[28286] = i[28286];
  assign o[28285] = i[28285];
  assign o[28284] = i[28284];
  assign o[28283] = i[28283];
  assign o[28282] = i[28282];
  assign o[28281] = i[28281];
  assign o[28280] = i[28280];
  assign o[28279] = i[28279];
  assign o[28278] = i[28278];
  assign o[28277] = i[28277];
  assign o[28276] = i[28276];
  assign o[28275] = i[28275];
  assign o[28274] = i[28274];
  assign o[28273] = i[28273];
  assign o[28272] = i[28272];
  assign o[28271] = i[28271];
  assign o[28270] = i[28270];
  assign o[28269] = i[28269];
  assign o[28268] = i[28268];
  assign o[28267] = i[28267];
  assign o[28266] = i[28266];
  assign o[28265] = i[28265];
  assign o[28264] = i[28264];
  assign o[28263] = i[28263];
  assign o[28262] = i[28262];
  assign o[28261] = i[28261];
  assign o[28260] = i[28260];
  assign o[28259] = i[28259];
  assign o[28258] = i[28258];
  assign o[28257] = i[28257];
  assign o[28256] = i[28256];
  assign o[28255] = i[28255];
  assign o[28254] = i[28254];
  assign o[28253] = i[28253];
  assign o[28252] = i[28252];
  assign o[28251] = i[28251];
  assign o[28250] = i[28250];
  assign o[28249] = i[28249];
  assign o[28248] = i[28248];
  assign o[28247] = i[28247];
  assign o[28246] = i[28246];
  assign o[28245] = i[28245];
  assign o[28244] = i[28244];
  assign o[28243] = i[28243];
  assign o[28242] = i[28242];
  assign o[28241] = i[28241];
  assign o[28240] = i[28240];
  assign o[28239] = i[28239];
  assign o[28238] = i[28238];
  assign o[28237] = i[28237];
  assign o[28236] = i[28236];
  assign o[28235] = i[28235];
  assign o[28234] = i[28234];
  assign o[28233] = i[28233];
  assign o[28232] = i[28232];
  assign o[28231] = i[28231];
  assign o[28230] = i[28230];
  assign o[28229] = i[28229];
  assign o[28228] = i[28228];
  assign o[28227] = i[28227];
  assign o[28226] = i[28226];
  assign o[28225] = i[28225];
  assign o[28224] = i[28224];
  assign o[28223] = i[28223];
  assign o[28222] = i[28222];
  assign o[28221] = i[28221];
  assign o[28220] = i[28220];
  assign o[28219] = i[28219];
  assign o[28218] = i[28218];
  assign o[28217] = i[28217];
  assign o[28216] = i[28216];
  assign o[28215] = i[28215];
  assign o[28214] = i[28214];
  assign o[28213] = i[28213];
  assign o[28212] = i[28212];
  assign o[28211] = i[28211];
  assign o[28210] = i[28210];
  assign o[28209] = i[28209];
  assign o[28208] = i[28208];
  assign o[28207] = i[28207];
  assign o[28206] = i[28206];
  assign o[28205] = i[28205];
  assign o[28204] = i[28204];
  assign o[28203] = i[28203];
  assign o[28202] = i[28202];
  assign o[28201] = i[28201];
  assign o[28200] = i[28200];
  assign o[28199] = i[28199];
  assign o[28198] = i[28198];
  assign o[28197] = i[28197];
  assign o[28196] = i[28196];
  assign o[28195] = i[28195];
  assign o[28194] = i[28194];
  assign o[28193] = i[28193];
  assign o[28192] = i[28192];
  assign o[28191] = i[28191];
  assign o[28190] = i[28190];
  assign o[28189] = i[28189];
  assign o[28188] = i[28188];
  assign o[28187] = i[28187];
  assign o[28186] = i[28186];
  assign o[28185] = i[28185];
  assign o[28184] = i[28184];
  assign o[28183] = i[28183];
  assign o[28182] = i[28182];
  assign o[28181] = i[28181];
  assign o[28180] = i[28180];
  assign o[28179] = i[28179];
  assign o[28178] = i[28178];
  assign o[28177] = i[28177];
  assign o[28176] = i[28176];
  assign o[28175] = i[28175];
  assign o[28174] = i[28174];
  assign o[28173] = i[28173];
  assign o[28172] = i[28172];
  assign o[28171] = i[28171];
  assign o[28170] = i[28170];
  assign o[28169] = i[28169];
  assign o[28168] = i[28168];
  assign o[28167] = i[28167];
  assign o[28166] = i[28166];
  assign o[28165] = i[28165];
  assign o[28164] = i[28164];
  assign o[28163] = i[28163];
  assign o[28162] = i[28162];
  assign o[28161] = i[28161];
  assign o[28160] = i[28160];
  assign o[28159] = i[28159];
  assign o[28158] = i[28158];
  assign o[28157] = i[28157];
  assign o[28156] = i[28156];
  assign o[28155] = i[28155];
  assign o[28154] = i[28154];
  assign o[28153] = i[28153];
  assign o[28152] = i[28152];
  assign o[28151] = i[28151];
  assign o[28150] = i[28150];
  assign o[28149] = i[28149];
  assign o[28148] = i[28148];
  assign o[28147] = i[28147];
  assign o[28146] = i[28146];
  assign o[28145] = i[28145];
  assign o[28144] = i[28144];
  assign o[28143] = i[28143];
  assign o[28142] = i[28142];
  assign o[28141] = i[28141];
  assign o[28140] = i[28140];
  assign o[28139] = i[28139];
  assign o[28138] = i[28138];
  assign o[28137] = i[28137];
  assign o[28136] = i[28136];
  assign o[28135] = i[28135];
  assign o[28134] = i[28134];
  assign o[28133] = i[28133];
  assign o[28132] = i[28132];
  assign o[28131] = i[28131];
  assign o[28130] = i[28130];
  assign o[28129] = i[28129];
  assign o[28128] = i[28128];
  assign o[28127] = i[28127];
  assign o[28126] = i[28126];
  assign o[28125] = i[28125];
  assign o[28124] = i[28124];
  assign o[28123] = i[28123];
  assign o[28122] = i[28122];
  assign o[28121] = i[28121];
  assign o[28120] = i[28120];
  assign o[28119] = i[28119];
  assign o[28118] = i[28118];
  assign o[28117] = i[28117];
  assign o[28116] = i[28116];
  assign o[28115] = i[28115];
  assign o[28114] = i[28114];
  assign o[28113] = i[28113];
  assign o[28112] = i[28112];
  assign o[28111] = i[28111];
  assign o[28110] = i[28110];
  assign o[28109] = i[28109];
  assign o[28108] = i[28108];
  assign o[28107] = i[28107];
  assign o[28106] = i[28106];
  assign o[28105] = i[28105];
  assign o[28104] = i[28104];
  assign o[28103] = i[28103];
  assign o[28102] = i[28102];
  assign o[28101] = i[28101];
  assign o[28100] = i[28100];
  assign o[28099] = i[28099];
  assign o[28098] = i[28098];
  assign o[28097] = i[28097];
  assign o[28096] = i[28096];
  assign o[28095] = i[28095];
  assign o[28094] = i[28094];
  assign o[28093] = i[28093];
  assign o[28092] = i[28092];
  assign o[28091] = i[28091];
  assign o[28090] = i[28090];
  assign o[28089] = i[28089];
  assign o[28088] = i[28088];
  assign o[28087] = i[28087];
  assign o[28086] = i[28086];
  assign o[28085] = i[28085];
  assign o[28084] = i[28084];
  assign o[28083] = i[28083];
  assign o[28082] = i[28082];
  assign o[28081] = i[28081];
  assign o[28080] = i[28080];
  assign o[28079] = i[28079];
  assign o[28078] = i[28078];
  assign o[28077] = i[28077];
  assign o[28076] = i[28076];
  assign o[28075] = i[28075];
  assign o[28074] = i[28074];
  assign o[28073] = i[28073];
  assign o[28072] = i[28072];
  assign o[28071] = i[28071];
  assign o[28070] = i[28070];
  assign o[28069] = i[28069];
  assign o[28068] = i[28068];
  assign o[28067] = i[28067];
  assign o[28066] = i[28066];
  assign o[28065] = i[28065];
  assign o[28064] = i[28064];
  assign o[28063] = i[28063];
  assign o[28062] = i[28062];
  assign o[28061] = i[28061];
  assign o[28060] = i[28060];
  assign o[28059] = i[28059];
  assign o[28058] = i[28058];
  assign o[28057] = i[28057];
  assign o[28056] = i[28056];
  assign o[28055] = i[28055];
  assign o[28054] = i[28054];
  assign o[28053] = i[28053];
  assign o[28052] = i[28052];
  assign o[28051] = i[28051];
  assign o[28050] = i[28050];
  assign o[28049] = i[28049];
  assign o[28048] = i[28048];
  assign o[28047] = i[28047];
  assign o[28046] = i[28046];
  assign o[28045] = i[28045];
  assign o[28044] = i[28044];
  assign o[28043] = i[28043];
  assign o[28042] = i[28042];
  assign o[28041] = i[28041];
  assign o[28040] = i[28040];
  assign o[28039] = i[28039];
  assign o[28038] = i[28038];
  assign o[28037] = i[28037];
  assign o[28036] = i[28036];
  assign o[28035] = i[28035];
  assign o[28034] = i[28034];
  assign o[28033] = i[28033];
  assign o[28032] = i[28032];
  assign o[28031] = i[28031];
  assign o[28030] = i[28030];
  assign o[28029] = i[28029];
  assign o[28028] = i[28028];
  assign o[28027] = i[28027];
  assign o[28026] = i[28026];
  assign o[28025] = i[28025];
  assign o[28024] = i[28024];
  assign o[28023] = i[28023];
  assign o[28022] = i[28022];
  assign o[28021] = i[28021];
  assign o[28020] = i[28020];
  assign o[28019] = i[28019];
  assign o[28018] = i[28018];
  assign o[28017] = i[28017];
  assign o[28016] = i[28016];
  assign o[28015] = i[28015];
  assign o[28014] = i[28014];
  assign o[28013] = i[28013];
  assign o[28012] = i[28012];
  assign o[28011] = i[28011];
  assign o[28010] = i[28010];
  assign o[28009] = i[28009];
  assign o[28008] = i[28008];
  assign o[28007] = i[28007];
  assign o[28006] = i[28006];
  assign o[28005] = i[28005];
  assign o[28004] = i[28004];
  assign o[28003] = i[28003];
  assign o[28002] = i[28002];
  assign o[28001] = i[28001];
  assign o[28000] = i[28000];
  assign o[27999] = i[27999];
  assign o[27998] = i[27998];
  assign o[27997] = i[27997];
  assign o[27996] = i[27996];
  assign o[27995] = i[27995];
  assign o[27994] = i[27994];
  assign o[27993] = i[27993];
  assign o[27992] = i[27992];
  assign o[27991] = i[27991];
  assign o[27990] = i[27990];
  assign o[27989] = i[27989];
  assign o[27988] = i[27988];
  assign o[27987] = i[27987];
  assign o[27986] = i[27986];
  assign o[27985] = i[27985];
  assign o[27984] = i[27984];
  assign o[27983] = i[27983];
  assign o[27982] = i[27982];
  assign o[27981] = i[27981];
  assign o[27980] = i[27980];
  assign o[27979] = i[27979];
  assign o[27978] = i[27978];
  assign o[27977] = i[27977];
  assign o[27976] = i[27976];
  assign o[27975] = i[27975];
  assign o[27974] = i[27974];
  assign o[27973] = i[27973];
  assign o[27972] = i[27972];
  assign o[27971] = i[27971];
  assign o[27970] = i[27970];
  assign o[27969] = i[27969];
  assign o[27968] = i[27968];
  assign o[27967] = i[27967];
  assign o[27966] = i[27966];
  assign o[27965] = i[27965];
  assign o[27964] = i[27964];
  assign o[27963] = i[27963];
  assign o[27962] = i[27962];
  assign o[27961] = i[27961];
  assign o[27960] = i[27960];
  assign o[27959] = i[27959];
  assign o[27958] = i[27958];
  assign o[27957] = i[27957];
  assign o[27956] = i[27956];
  assign o[27955] = i[27955];
  assign o[27954] = i[27954];
  assign o[27953] = i[27953];
  assign o[27952] = i[27952];
  assign o[27951] = i[27951];
  assign o[27950] = i[27950];
  assign o[27949] = i[27949];
  assign o[27948] = i[27948];
  assign o[27947] = i[27947];
  assign o[27946] = i[27946];
  assign o[27945] = i[27945];
  assign o[27944] = i[27944];
  assign o[27943] = i[27943];
  assign o[27942] = i[27942];
  assign o[27941] = i[27941];
  assign o[27940] = i[27940];
  assign o[27939] = i[27939];
  assign o[27938] = i[27938];
  assign o[27937] = i[27937];
  assign o[27936] = i[27936];
  assign o[27935] = i[27935];
  assign o[27934] = i[27934];
  assign o[27933] = i[27933];
  assign o[27932] = i[27932];
  assign o[27931] = i[27931];
  assign o[27930] = i[27930];
  assign o[27929] = i[27929];
  assign o[27928] = i[27928];
  assign o[27927] = i[27927];
  assign o[27926] = i[27926];
  assign o[27925] = i[27925];
  assign o[27924] = i[27924];
  assign o[27923] = i[27923];
  assign o[27922] = i[27922];
  assign o[27921] = i[27921];
  assign o[27920] = i[27920];
  assign o[27919] = i[27919];
  assign o[27918] = i[27918];
  assign o[27917] = i[27917];
  assign o[27916] = i[27916];
  assign o[27915] = i[27915];
  assign o[27914] = i[27914];
  assign o[27913] = i[27913];
  assign o[27912] = i[27912];
  assign o[27911] = i[27911];
  assign o[27910] = i[27910];
  assign o[27909] = i[27909];
  assign o[27908] = i[27908];
  assign o[27907] = i[27907];
  assign o[27906] = i[27906];
  assign o[27905] = i[27905];
  assign o[27904] = i[27904];
  assign o[27903] = i[27903];
  assign o[27902] = i[27902];
  assign o[27901] = i[27901];
  assign o[27900] = i[27900];
  assign o[27899] = i[27899];
  assign o[27898] = i[27898];
  assign o[27897] = i[27897];
  assign o[27896] = i[27896];
  assign o[27895] = i[27895];
  assign o[27894] = i[27894];
  assign o[27893] = i[27893];
  assign o[27892] = i[27892];
  assign o[27891] = i[27891];
  assign o[27890] = i[27890];
  assign o[27889] = i[27889];
  assign o[27888] = i[27888];
  assign o[27887] = i[27887];
  assign o[27886] = i[27886];
  assign o[27885] = i[27885];
  assign o[27884] = i[27884];
  assign o[27883] = i[27883];
  assign o[27882] = i[27882];
  assign o[27881] = i[27881];
  assign o[27880] = i[27880];
  assign o[27879] = i[27879];
  assign o[27878] = i[27878];
  assign o[27877] = i[27877];
  assign o[27876] = i[27876];
  assign o[27875] = i[27875];
  assign o[27874] = i[27874];
  assign o[27873] = i[27873];
  assign o[27872] = i[27872];
  assign o[27871] = i[27871];
  assign o[27870] = i[27870];
  assign o[27869] = i[27869];
  assign o[27868] = i[27868];
  assign o[27867] = i[27867];
  assign o[27866] = i[27866];
  assign o[27865] = i[27865];
  assign o[27864] = i[27864];
  assign o[27863] = i[27863];
  assign o[27862] = i[27862];
  assign o[27861] = i[27861];
  assign o[27860] = i[27860];
  assign o[27859] = i[27859];
  assign o[27858] = i[27858];
  assign o[27857] = i[27857];
  assign o[27856] = i[27856];
  assign o[27855] = i[27855];
  assign o[27854] = i[27854];
  assign o[27853] = i[27853];
  assign o[27852] = i[27852];
  assign o[27851] = i[27851];
  assign o[27850] = i[27850];
  assign o[27849] = i[27849];
  assign o[27848] = i[27848];
  assign o[27847] = i[27847];
  assign o[27846] = i[27846];
  assign o[27845] = i[27845];
  assign o[27844] = i[27844];
  assign o[27843] = i[27843];
  assign o[27842] = i[27842];
  assign o[27841] = i[27841];
  assign o[27840] = i[27840];
  assign o[27839] = i[27839];
  assign o[27838] = i[27838];
  assign o[27837] = i[27837];
  assign o[27836] = i[27836];
  assign o[27835] = i[27835];
  assign o[27834] = i[27834];
  assign o[27833] = i[27833];
  assign o[27832] = i[27832];
  assign o[27831] = i[27831];
  assign o[27830] = i[27830];
  assign o[27829] = i[27829];
  assign o[27828] = i[27828];
  assign o[27827] = i[27827];
  assign o[27826] = i[27826];
  assign o[27825] = i[27825];
  assign o[27824] = i[27824];
  assign o[27823] = i[27823];
  assign o[27822] = i[27822];
  assign o[27821] = i[27821];
  assign o[27820] = i[27820];
  assign o[27819] = i[27819];
  assign o[27818] = i[27818];
  assign o[27817] = i[27817];
  assign o[27816] = i[27816];
  assign o[27815] = i[27815];
  assign o[27814] = i[27814];
  assign o[27813] = i[27813];
  assign o[27812] = i[27812];
  assign o[27811] = i[27811];
  assign o[27810] = i[27810];
  assign o[27809] = i[27809];
  assign o[27808] = i[27808];
  assign o[27807] = i[27807];
  assign o[27806] = i[27806];
  assign o[27805] = i[27805];
  assign o[27804] = i[27804];
  assign o[27803] = i[27803];
  assign o[27802] = i[27802];
  assign o[27801] = i[27801];
  assign o[27800] = i[27800];
  assign o[27799] = i[27799];
  assign o[27798] = i[27798];
  assign o[27797] = i[27797];
  assign o[27796] = i[27796];
  assign o[27795] = i[27795];
  assign o[27794] = i[27794];
  assign o[27793] = i[27793];
  assign o[27792] = i[27792];
  assign o[27791] = i[27791];
  assign o[27790] = i[27790];
  assign o[27789] = i[27789];
  assign o[27788] = i[27788];
  assign o[27787] = i[27787];
  assign o[27786] = i[27786];
  assign o[27785] = i[27785];
  assign o[27784] = i[27784];
  assign o[27783] = i[27783];
  assign o[27782] = i[27782];
  assign o[27781] = i[27781];
  assign o[27780] = i[27780];
  assign o[27779] = i[27779];
  assign o[27778] = i[27778];
  assign o[27777] = i[27777];
  assign o[27776] = i[27776];
  assign o[27775] = i[27775];
  assign o[27774] = i[27774];
  assign o[27773] = i[27773];
  assign o[27772] = i[27772];
  assign o[27771] = i[27771];
  assign o[27770] = i[27770];
  assign o[27769] = i[27769];
  assign o[27768] = i[27768];
  assign o[27767] = i[27767];
  assign o[27766] = i[27766];
  assign o[27765] = i[27765];
  assign o[27764] = i[27764];
  assign o[27763] = i[27763];
  assign o[27762] = i[27762];
  assign o[27761] = i[27761];
  assign o[27760] = i[27760];
  assign o[27759] = i[27759];
  assign o[27758] = i[27758];
  assign o[27757] = i[27757];
  assign o[27756] = i[27756];
  assign o[27755] = i[27755];
  assign o[27754] = i[27754];
  assign o[27753] = i[27753];
  assign o[27752] = i[27752];
  assign o[27751] = i[27751];
  assign o[27750] = i[27750];
  assign o[27749] = i[27749];
  assign o[27748] = i[27748];
  assign o[27747] = i[27747];
  assign o[27746] = i[27746];
  assign o[27745] = i[27745];
  assign o[27744] = i[27744];
  assign o[27743] = i[27743];
  assign o[27742] = i[27742];
  assign o[27741] = i[27741];
  assign o[27740] = i[27740];
  assign o[27739] = i[27739];
  assign o[27738] = i[27738];
  assign o[27737] = i[27737];
  assign o[27736] = i[27736];
  assign o[27735] = i[27735];
  assign o[27734] = i[27734];
  assign o[27733] = i[27733];
  assign o[27732] = i[27732];
  assign o[27731] = i[27731];
  assign o[27730] = i[27730];
  assign o[27729] = i[27729];
  assign o[27728] = i[27728];
  assign o[27727] = i[27727];
  assign o[27726] = i[27726];
  assign o[27725] = i[27725];
  assign o[27724] = i[27724];
  assign o[27723] = i[27723];
  assign o[27722] = i[27722];
  assign o[27721] = i[27721];
  assign o[27720] = i[27720];
  assign o[27719] = i[27719];
  assign o[27718] = i[27718];
  assign o[27717] = i[27717];
  assign o[27716] = i[27716];
  assign o[27715] = i[27715];
  assign o[27714] = i[27714];
  assign o[27713] = i[27713];
  assign o[27712] = i[27712];
  assign o[27711] = i[27711];
  assign o[27710] = i[27710];
  assign o[27709] = i[27709];
  assign o[27708] = i[27708];
  assign o[27707] = i[27707];
  assign o[27706] = i[27706];
  assign o[27705] = i[27705];
  assign o[27704] = i[27704];
  assign o[27703] = i[27703];
  assign o[27702] = i[27702];
  assign o[27701] = i[27701];
  assign o[27700] = i[27700];
  assign o[27699] = i[27699];
  assign o[27698] = i[27698];
  assign o[27697] = i[27697];
  assign o[27696] = i[27696];
  assign o[27695] = i[27695];
  assign o[27694] = i[27694];
  assign o[27693] = i[27693];
  assign o[27692] = i[27692];
  assign o[27691] = i[27691];
  assign o[27690] = i[27690];
  assign o[27689] = i[27689];
  assign o[27688] = i[27688];
  assign o[27687] = i[27687];
  assign o[27686] = i[27686];
  assign o[27685] = i[27685];
  assign o[27684] = i[27684];
  assign o[27683] = i[27683];
  assign o[27682] = i[27682];
  assign o[27681] = i[27681];
  assign o[27680] = i[27680];
  assign o[27679] = i[27679];
  assign o[27678] = i[27678];
  assign o[27677] = i[27677];
  assign o[27676] = i[27676];
  assign o[27675] = i[27675];
  assign o[27674] = i[27674];
  assign o[27673] = i[27673];
  assign o[27672] = i[27672];
  assign o[27671] = i[27671];
  assign o[27670] = i[27670];
  assign o[27669] = i[27669];
  assign o[27668] = i[27668];
  assign o[27667] = i[27667];
  assign o[27666] = i[27666];
  assign o[27665] = i[27665];
  assign o[27664] = i[27664];
  assign o[27663] = i[27663];
  assign o[27662] = i[27662];
  assign o[27661] = i[27661];
  assign o[27660] = i[27660];
  assign o[27659] = i[27659];
  assign o[27658] = i[27658];
  assign o[27657] = i[27657];
  assign o[27656] = i[27656];
  assign o[27655] = i[27655];
  assign o[27654] = i[27654];
  assign o[27653] = i[27653];
  assign o[27652] = i[27652];
  assign o[27651] = i[27651];
  assign o[27650] = i[27650];
  assign o[27649] = i[27649];
  assign o[27648] = i[27648];
  assign o[27647] = i[27647];
  assign o[27646] = i[27646];
  assign o[27645] = i[27645];
  assign o[27644] = i[27644];
  assign o[27643] = i[27643];
  assign o[27642] = i[27642];
  assign o[27641] = i[27641];
  assign o[27640] = i[27640];
  assign o[27639] = i[27639];
  assign o[27638] = i[27638];
  assign o[27637] = i[27637];
  assign o[27636] = i[27636];
  assign o[27635] = i[27635];
  assign o[27634] = i[27634];
  assign o[27633] = i[27633];
  assign o[27632] = i[27632];
  assign o[27631] = i[27631];
  assign o[27630] = i[27630];
  assign o[27629] = i[27629];
  assign o[27628] = i[27628];
  assign o[27627] = i[27627];
  assign o[27626] = i[27626];
  assign o[27625] = i[27625];
  assign o[27624] = i[27624];
  assign o[27623] = i[27623];
  assign o[27622] = i[27622];
  assign o[27621] = i[27621];
  assign o[27620] = i[27620];
  assign o[27619] = i[27619];
  assign o[27618] = i[27618];
  assign o[27617] = i[27617];
  assign o[27616] = i[27616];
  assign o[27615] = i[27615];
  assign o[27614] = i[27614];
  assign o[27613] = i[27613];
  assign o[27612] = i[27612];
  assign o[27611] = i[27611];
  assign o[27610] = i[27610];
  assign o[27609] = i[27609];
  assign o[27608] = i[27608];
  assign o[27607] = i[27607];
  assign o[27606] = i[27606];
  assign o[27605] = i[27605];
  assign o[27604] = i[27604];
  assign o[27603] = i[27603];
  assign o[27602] = i[27602];
  assign o[27601] = i[27601];
  assign o[27600] = i[27600];
  assign o[27599] = i[27599];
  assign o[27598] = i[27598];
  assign o[27597] = i[27597];
  assign o[27596] = i[27596];
  assign o[27595] = i[27595];
  assign o[27594] = i[27594];
  assign o[27593] = i[27593];
  assign o[27592] = i[27592];
  assign o[27591] = i[27591];
  assign o[27590] = i[27590];
  assign o[27589] = i[27589];
  assign o[27588] = i[27588];
  assign o[27587] = i[27587];
  assign o[27586] = i[27586];
  assign o[27585] = i[27585];
  assign o[27584] = i[27584];
  assign o[27583] = i[27583];
  assign o[27582] = i[27582];
  assign o[27581] = i[27581];
  assign o[27580] = i[27580];
  assign o[27579] = i[27579];
  assign o[27578] = i[27578];
  assign o[27577] = i[27577];
  assign o[27576] = i[27576];
  assign o[27575] = i[27575];
  assign o[27574] = i[27574];
  assign o[27573] = i[27573];
  assign o[27572] = i[27572];
  assign o[27571] = i[27571];
  assign o[27570] = i[27570];
  assign o[27569] = i[27569];
  assign o[27568] = i[27568];
  assign o[27567] = i[27567];
  assign o[27566] = i[27566];
  assign o[27565] = i[27565];
  assign o[27564] = i[27564];
  assign o[27563] = i[27563];
  assign o[27562] = i[27562];
  assign o[27561] = i[27561];
  assign o[27560] = i[27560];
  assign o[27559] = i[27559];
  assign o[27558] = i[27558];
  assign o[27557] = i[27557];
  assign o[27556] = i[27556];
  assign o[27555] = i[27555];
  assign o[27554] = i[27554];
  assign o[27553] = i[27553];
  assign o[27552] = i[27552];
  assign o[27551] = i[27551];
  assign o[27550] = i[27550];
  assign o[27549] = i[27549];
  assign o[27548] = i[27548];
  assign o[27547] = i[27547];
  assign o[27546] = i[27546];
  assign o[27545] = i[27545];
  assign o[27544] = i[27544];
  assign o[27543] = i[27543];
  assign o[27542] = i[27542];
  assign o[27541] = i[27541];
  assign o[27540] = i[27540];
  assign o[27539] = i[27539];
  assign o[27538] = i[27538];
  assign o[27537] = i[27537];
  assign o[27536] = i[27536];
  assign o[27535] = i[27535];
  assign o[27534] = i[27534];
  assign o[27533] = i[27533];
  assign o[27532] = i[27532];
  assign o[27531] = i[27531];
  assign o[27530] = i[27530];
  assign o[27529] = i[27529];
  assign o[27528] = i[27528];
  assign o[27527] = i[27527];
  assign o[27526] = i[27526];
  assign o[27525] = i[27525];
  assign o[27524] = i[27524];
  assign o[27523] = i[27523];
  assign o[27522] = i[27522];
  assign o[27521] = i[27521];
  assign o[27520] = i[27520];
  assign o[27519] = i[27519];
  assign o[27518] = i[27518];
  assign o[27517] = i[27517];
  assign o[27516] = i[27516];
  assign o[27515] = i[27515];
  assign o[27514] = i[27514];
  assign o[27513] = i[27513];
  assign o[27512] = i[27512];
  assign o[27511] = i[27511];
  assign o[27510] = i[27510];
  assign o[27509] = i[27509];
  assign o[27508] = i[27508];
  assign o[27507] = i[27507];
  assign o[27506] = i[27506];
  assign o[27505] = i[27505];
  assign o[27504] = i[27504];
  assign o[27503] = i[27503];
  assign o[27502] = i[27502];
  assign o[27501] = i[27501];
  assign o[27500] = i[27500];
  assign o[27499] = i[27499];
  assign o[27498] = i[27498];
  assign o[27497] = i[27497];
  assign o[27496] = i[27496];
  assign o[27495] = i[27495];
  assign o[27494] = i[27494];
  assign o[27493] = i[27493];
  assign o[27492] = i[27492];
  assign o[27491] = i[27491];
  assign o[27490] = i[27490];
  assign o[27489] = i[27489];
  assign o[27488] = i[27488];
  assign o[27487] = i[27487];
  assign o[27486] = i[27486];
  assign o[27485] = i[27485];
  assign o[27484] = i[27484];
  assign o[27483] = i[27483];
  assign o[27482] = i[27482];
  assign o[27481] = i[27481];
  assign o[27480] = i[27480];
  assign o[27479] = i[27479];
  assign o[27478] = i[27478];
  assign o[27477] = i[27477];
  assign o[27476] = i[27476];
  assign o[27475] = i[27475];
  assign o[27474] = i[27474];
  assign o[27473] = i[27473];
  assign o[27472] = i[27472];
  assign o[27471] = i[27471];
  assign o[27470] = i[27470];
  assign o[27469] = i[27469];
  assign o[27468] = i[27468];
  assign o[27467] = i[27467];
  assign o[27466] = i[27466];
  assign o[27465] = i[27465];
  assign o[27464] = i[27464];
  assign o[27463] = i[27463];
  assign o[27462] = i[27462];
  assign o[27461] = i[27461];
  assign o[27460] = i[27460];
  assign o[27459] = i[27459];
  assign o[27458] = i[27458];
  assign o[27457] = i[27457];
  assign o[27456] = i[27456];
  assign o[27455] = i[27455];
  assign o[27454] = i[27454];
  assign o[27453] = i[27453];
  assign o[27452] = i[27452];
  assign o[27451] = i[27451];
  assign o[27450] = i[27450];
  assign o[27449] = i[27449];
  assign o[27448] = i[27448];
  assign o[27447] = i[27447];
  assign o[27446] = i[27446];
  assign o[27445] = i[27445];
  assign o[27444] = i[27444];
  assign o[27443] = i[27443];
  assign o[27442] = i[27442];
  assign o[27441] = i[27441];
  assign o[27440] = i[27440];
  assign o[27439] = i[27439];
  assign o[27438] = i[27438];
  assign o[27437] = i[27437];
  assign o[27436] = i[27436];
  assign o[27435] = i[27435];
  assign o[27434] = i[27434];
  assign o[27433] = i[27433];
  assign o[27432] = i[27432];
  assign o[27431] = i[27431];
  assign o[27430] = i[27430];
  assign o[27429] = i[27429];
  assign o[27428] = i[27428];
  assign o[27427] = i[27427];
  assign o[27426] = i[27426];
  assign o[27425] = i[27425];
  assign o[27424] = i[27424];
  assign o[27423] = i[27423];
  assign o[27422] = i[27422];
  assign o[27421] = i[27421];
  assign o[27420] = i[27420];
  assign o[27419] = i[27419];
  assign o[27418] = i[27418];
  assign o[27417] = i[27417];
  assign o[27416] = i[27416];
  assign o[27415] = i[27415];
  assign o[27414] = i[27414];
  assign o[27413] = i[27413];
  assign o[27412] = i[27412];
  assign o[27411] = i[27411];
  assign o[27410] = i[27410];
  assign o[27409] = i[27409];
  assign o[27408] = i[27408];
  assign o[27407] = i[27407];
  assign o[27406] = i[27406];
  assign o[27405] = i[27405];
  assign o[27404] = i[27404];
  assign o[27403] = i[27403];
  assign o[27402] = i[27402];
  assign o[27401] = i[27401];
  assign o[27400] = i[27400];
  assign o[27399] = i[27399];
  assign o[27398] = i[27398];
  assign o[27397] = i[27397];
  assign o[27396] = i[27396];
  assign o[27395] = i[27395];
  assign o[27394] = i[27394];
  assign o[27393] = i[27393];
  assign o[27392] = i[27392];
  assign o[27391] = i[27391];
  assign o[27390] = i[27390];
  assign o[27389] = i[27389];
  assign o[27388] = i[27388];
  assign o[27387] = i[27387];
  assign o[27386] = i[27386];
  assign o[27385] = i[27385];
  assign o[27384] = i[27384];
  assign o[27383] = i[27383];
  assign o[27382] = i[27382];
  assign o[27381] = i[27381];
  assign o[27380] = i[27380];
  assign o[27379] = i[27379];
  assign o[27378] = i[27378];
  assign o[27377] = i[27377];
  assign o[27376] = i[27376];
  assign o[27375] = i[27375];
  assign o[27374] = i[27374];
  assign o[27373] = i[27373];
  assign o[27372] = i[27372];
  assign o[27371] = i[27371];
  assign o[27370] = i[27370];
  assign o[27369] = i[27369];
  assign o[27368] = i[27368];
  assign o[27367] = i[27367];
  assign o[27366] = i[27366];
  assign o[27365] = i[27365];
  assign o[27364] = i[27364];
  assign o[27363] = i[27363];
  assign o[27362] = i[27362];
  assign o[27361] = i[27361];
  assign o[27360] = i[27360];
  assign o[27359] = i[27359];
  assign o[27358] = i[27358];
  assign o[27357] = i[27357];
  assign o[27356] = i[27356];
  assign o[27355] = i[27355];
  assign o[27354] = i[27354];
  assign o[27353] = i[27353];
  assign o[27352] = i[27352];
  assign o[27351] = i[27351];
  assign o[27350] = i[27350];
  assign o[27349] = i[27349];
  assign o[27348] = i[27348];
  assign o[27347] = i[27347];
  assign o[27346] = i[27346];
  assign o[27345] = i[27345];
  assign o[27344] = i[27344];
  assign o[27343] = i[27343];
  assign o[27342] = i[27342];
  assign o[27341] = i[27341];
  assign o[27340] = i[27340];
  assign o[27339] = i[27339];
  assign o[27338] = i[27338];
  assign o[27337] = i[27337];
  assign o[27336] = i[27336];
  assign o[27335] = i[27335];
  assign o[27334] = i[27334];
  assign o[27333] = i[27333];
  assign o[27332] = i[27332];
  assign o[27331] = i[27331];
  assign o[27330] = i[27330];
  assign o[27329] = i[27329];
  assign o[27328] = i[27328];
  assign o[27327] = i[27327];
  assign o[27326] = i[27326];
  assign o[27325] = i[27325];
  assign o[27324] = i[27324];
  assign o[27323] = i[27323];
  assign o[27322] = i[27322];
  assign o[27321] = i[27321];
  assign o[27320] = i[27320];
  assign o[27319] = i[27319];
  assign o[27318] = i[27318];
  assign o[27317] = i[27317];
  assign o[27316] = i[27316];
  assign o[27315] = i[27315];
  assign o[27314] = i[27314];
  assign o[27313] = i[27313];
  assign o[27312] = i[27312];
  assign o[27311] = i[27311];
  assign o[27310] = i[27310];
  assign o[27309] = i[27309];
  assign o[27308] = i[27308];
  assign o[27307] = i[27307];
  assign o[27306] = i[27306];
  assign o[27305] = i[27305];
  assign o[27304] = i[27304];
  assign o[27303] = i[27303];
  assign o[27302] = i[27302];
  assign o[27301] = i[27301];
  assign o[27300] = i[27300];
  assign o[27299] = i[27299];
  assign o[27298] = i[27298];
  assign o[27297] = i[27297];
  assign o[27296] = i[27296];
  assign o[27295] = i[27295];
  assign o[27294] = i[27294];
  assign o[27293] = i[27293];
  assign o[27292] = i[27292];
  assign o[27291] = i[27291];
  assign o[27290] = i[27290];
  assign o[27289] = i[27289];
  assign o[27288] = i[27288];
  assign o[27287] = i[27287];
  assign o[27286] = i[27286];
  assign o[27285] = i[27285];
  assign o[27284] = i[27284];
  assign o[27283] = i[27283];
  assign o[27282] = i[27282];
  assign o[27281] = i[27281];
  assign o[27280] = i[27280];
  assign o[27279] = i[27279];
  assign o[27278] = i[27278];
  assign o[27277] = i[27277];
  assign o[27276] = i[27276];
  assign o[27275] = i[27275];
  assign o[27274] = i[27274];
  assign o[27273] = i[27273];
  assign o[27272] = i[27272];
  assign o[27271] = i[27271];
  assign o[27270] = i[27270];
  assign o[27269] = i[27269];
  assign o[27268] = i[27268];
  assign o[27267] = i[27267];
  assign o[27266] = i[27266];
  assign o[27265] = i[27265];
  assign o[27264] = i[27264];
  assign o[27263] = i[27263];
  assign o[27262] = i[27262];
  assign o[27261] = i[27261];
  assign o[27260] = i[27260];
  assign o[27259] = i[27259];
  assign o[27258] = i[27258];
  assign o[27257] = i[27257];
  assign o[27256] = i[27256];
  assign o[27255] = i[27255];
  assign o[27254] = i[27254];
  assign o[27253] = i[27253];
  assign o[27252] = i[27252];
  assign o[27251] = i[27251];
  assign o[27250] = i[27250];
  assign o[27249] = i[27249];
  assign o[27248] = i[27248];
  assign o[27247] = i[27247];
  assign o[27246] = i[27246];
  assign o[27245] = i[27245];
  assign o[27244] = i[27244];
  assign o[27243] = i[27243];
  assign o[27242] = i[27242];
  assign o[27241] = i[27241];
  assign o[27240] = i[27240];
  assign o[27239] = i[27239];
  assign o[27238] = i[27238];
  assign o[27237] = i[27237];
  assign o[27236] = i[27236];
  assign o[27235] = i[27235];
  assign o[27234] = i[27234];
  assign o[27233] = i[27233];
  assign o[27232] = i[27232];
  assign o[27231] = i[27231];
  assign o[27230] = i[27230];
  assign o[27229] = i[27229];
  assign o[27228] = i[27228];
  assign o[27227] = i[27227];
  assign o[27226] = i[27226];
  assign o[27225] = i[27225];
  assign o[27224] = i[27224];
  assign o[27223] = i[27223];
  assign o[27222] = i[27222];
  assign o[27221] = i[27221];
  assign o[27220] = i[27220];
  assign o[27219] = i[27219];
  assign o[27218] = i[27218];
  assign o[27217] = i[27217];
  assign o[27216] = i[27216];
  assign o[27215] = i[27215];
  assign o[27214] = i[27214];
  assign o[27213] = i[27213];
  assign o[27212] = i[27212];
  assign o[27211] = i[27211];
  assign o[27210] = i[27210];
  assign o[27209] = i[27209];
  assign o[27208] = i[27208];
  assign o[27207] = i[27207];
  assign o[27206] = i[27206];
  assign o[27205] = i[27205];
  assign o[27204] = i[27204];
  assign o[27203] = i[27203];
  assign o[27202] = i[27202];
  assign o[27201] = i[27201];
  assign o[27200] = i[27200];
  assign o[27199] = i[27199];
  assign o[27198] = i[27198];
  assign o[27197] = i[27197];
  assign o[27196] = i[27196];
  assign o[27195] = i[27195];
  assign o[27194] = i[27194];
  assign o[27193] = i[27193];
  assign o[27192] = i[27192];
  assign o[27191] = i[27191];
  assign o[27190] = i[27190];
  assign o[27189] = i[27189];
  assign o[27188] = i[27188];
  assign o[27187] = i[27187];
  assign o[27186] = i[27186];
  assign o[27185] = i[27185];
  assign o[27184] = i[27184];
  assign o[27183] = i[27183];
  assign o[27182] = i[27182];
  assign o[27181] = i[27181];
  assign o[27180] = i[27180];
  assign o[27179] = i[27179];
  assign o[27178] = i[27178];
  assign o[27177] = i[27177];
  assign o[27176] = i[27176];
  assign o[27175] = i[27175];
  assign o[27174] = i[27174];
  assign o[27173] = i[27173];
  assign o[27172] = i[27172];
  assign o[27171] = i[27171];
  assign o[27170] = i[27170];
  assign o[27169] = i[27169];
  assign o[27168] = i[27168];
  assign o[27167] = i[27167];
  assign o[27166] = i[27166];
  assign o[27165] = i[27165];
  assign o[27164] = i[27164];
  assign o[27163] = i[27163];
  assign o[27162] = i[27162];
  assign o[27161] = i[27161];
  assign o[27160] = i[27160];
  assign o[27159] = i[27159];
  assign o[27158] = i[27158];
  assign o[27157] = i[27157];
  assign o[27156] = i[27156];
  assign o[27155] = i[27155];
  assign o[27154] = i[27154];
  assign o[27153] = i[27153];
  assign o[27152] = i[27152];
  assign o[27151] = i[27151];
  assign o[27150] = i[27150];
  assign o[27149] = i[27149];
  assign o[27148] = i[27148];
  assign o[27147] = i[27147];
  assign o[27146] = i[27146];
  assign o[27145] = i[27145];
  assign o[27144] = i[27144];
  assign o[27143] = i[27143];
  assign o[27142] = i[27142];
  assign o[27141] = i[27141];
  assign o[27140] = i[27140];
  assign o[27139] = i[27139];
  assign o[27138] = i[27138];
  assign o[27137] = i[27137];
  assign o[27136] = i[27136];
  assign o[27135] = i[27135];
  assign o[27134] = i[27134];
  assign o[27133] = i[27133];
  assign o[27132] = i[27132];
  assign o[27131] = i[27131];
  assign o[27130] = i[27130];
  assign o[27129] = i[27129];
  assign o[27128] = i[27128];
  assign o[27127] = i[27127];
  assign o[27126] = i[27126];
  assign o[27125] = i[27125];
  assign o[27124] = i[27124];
  assign o[27123] = i[27123];
  assign o[27122] = i[27122];
  assign o[27121] = i[27121];
  assign o[27120] = i[27120];
  assign o[27119] = i[27119];
  assign o[27118] = i[27118];
  assign o[27117] = i[27117];
  assign o[27116] = i[27116];
  assign o[27115] = i[27115];
  assign o[27114] = i[27114];
  assign o[27113] = i[27113];
  assign o[27112] = i[27112];
  assign o[27111] = i[27111];
  assign o[27110] = i[27110];
  assign o[27109] = i[27109];
  assign o[27108] = i[27108];
  assign o[27107] = i[27107];
  assign o[27106] = i[27106];
  assign o[27105] = i[27105];
  assign o[27104] = i[27104];
  assign o[27103] = i[27103];
  assign o[27102] = i[27102];
  assign o[27101] = i[27101];
  assign o[27100] = i[27100];
  assign o[27099] = i[27099];
  assign o[27098] = i[27098];
  assign o[27097] = i[27097];
  assign o[27096] = i[27096];
  assign o[27095] = i[27095];
  assign o[27094] = i[27094];
  assign o[27093] = i[27093];
  assign o[27092] = i[27092];
  assign o[27091] = i[27091];
  assign o[27090] = i[27090];
  assign o[27089] = i[27089];
  assign o[27088] = i[27088];
  assign o[27087] = i[27087];
  assign o[27086] = i[27086];
  assign o[27085] = i[27085];
  assign o[27084] = i[27084];
  assign o[27083] = i[27083];
  assign o[27082] = i[27082];
  assign o[27081] = i[27081];
  assign o[27080] = i[27080];
  assign o[27079] = i[27079];
  assign o[27078] = i[27078];
  assign o[27077] = i[27077];
  assign o[27076] = i[27076];
  assign o[27075] = i[27075];
  assign o[27074] = i[27074];
  assign o[27073] = i[27073];
  assign o[27072] = i[27072];
  assign o[27071] = i[27071];
  assign o[27070] = i[27070];
  assign o[27069] = i[27069];
  assign o[27068] = i[27068];
  assign o[27067] = i[27067];
  assign o[27066] = i[27066];
  assign o[27065] = i[27065];
  assign o[27064] = i[27064];
  assign o[27063] = i[27063];
  assign o[27062] = i[27062];
  assign o[27061] = i[27061];
  assign o[27060] = i[27060];
  assign o[27059] = i[27059];
  assign o[27058] = i[27058];
  assign o[27057] = i[27057];
  assign o[27056] = i[27056];
  assign o[27055] = i[27055];
  assign o[27054] = i[27054];
  assign o[27053] = i[27053];
  assign o[27052] = i[27052];
  assign o[27051] = i[27051];
  assign o[27050] = i[27050];
  assign o[27049] = i[27049];
  assign o[27048] = i[27048];
  assign o[27047] = i[27047];
  assign o[27046] = i[27046];
  assign o[27045] = i[27045];
  assign o[27044] = i[27044];
  assign o[27043] = i[27043];
  assign o[27042] = i[27042];
  assign o[27041] = i[27041];
  assign o[27040] = i[27040];
  assign o[27039] = i[27039];
  assign o[27038] = i[27038];
  assign o[27037] = i[27037];
  assign o[27036] = i[27036];
  assign o[27035] = i[27035];
  assign o[27034] = i[27034];
  assign o[27033] = i[27033];
  assign o[27032] = i[27032];
  assign o[27031] = i[27031];
  assign o[27030] = i[27030];
  assign o[27029] = i[27029];
  assign o[27028] = i[27028];
  assign o[27027] = i[27027];
  assign o[27026] = i[27026];
  assign o[27025] = i[27025];
  assign o[27024] = i[27024];
  assign o[27023] = i[27023];
  assign o[27022] = i[27022];
  assign o[27021] = i[27021];
  assign o[27020] = i[27020];
  assign o[27019] = i[27019];
  assign o[27018] = i[27018];
  assign o[27017] = i[27017];
  assign o[27016] = i[27016];
  assign o[27015] = i[27015];
  assign o[27014] = i[27014];
  assign o[27013] = i[27013];
  assign o[27012] = i[27012];
  assign o[27011] = i[27011];
  assign o[27010] = i[27010];
  assign o[27009] = i[27009];
  assign o[27008] = i[27008];
  assign o[27007] = i[27007];
  assign o[27006] = i[27006];
  assign o[27005] = i[27005];
  assign o[27004] = i[27004];
  assign o[27003] = i[27003];
  assign o[27002] = i[27002];
  assign o[27001] = i[27001];
  assign o[27000] = i[27000];
  assign o[26999] = i[26999];
  assign o[26998] = i[26998];
  assign o[26997] = i[26997];
  assign o[26996] = i[26996];
  assign o[26995] = i[26995];
  assign o[26994] = i[26994];
  assign o[26993] = i[26993];
  assign o[26992] = i[26992];
  assign o[26991] = i[26991];
  assign o[26990] = i[26990];
  assign o[26989] = i[26989];
  assign o[26988] = i[26988];
  assign o[26987] = i[26987];
  assign o[26986] = i[26986];
  assign o[26985] = i[26985];
  assign o[26984] = i[26984];
  assign o[26983] = i[26983];
  assign o[26982] = i[26982];
  assign o[26981] = i[26981];
  assign o[26980] = i[26980];
  assign o[26979] = i[26979];
  assign o[26978] = i[26978];
  assign o[26977] = i[26977];
  assign o[26976] = i[26976];
  assign o[26975] = i[26975];
  assign o[26974] = i[26974];
  assign o[26973] = i[26973];
  assign o[26972] = i[26972];
  assign o[26971] = i[26971];
  assign o[26970] = i[26970];
  assign o[26969] = i[26969];
  assign o[26968] = i[26968];
  assign o[26967] = i[26967];
  assign o[26966] = i[26966];
  assign o[26965] = i[26965];
  assign o[26964] = i[26964];
  assign o[26963] = i[26963];
  assign o[26962] = i[26962];
  assign o[26961] = i[26961];
  assign o[26960] = i[26960];
  assign o[26959] = i[26959];
  assign o[26958] = i[26958];
  assign o[26957] = i[26957];
  assign o[26956] = i[26956];
  assign o[26955] = i[26955];
  assign o[26954] = i[26954];
  assign o[26953] = i[26953];
  assign o[26952] = i[26952];
  assign o[26951] = i[26951];
  assign o[26950] = i[26950];
  assign o[26949] = i[26949];
  assign o[26948] = i[26948];
  assign o[26947] = i[26947];
  assign o[26946] = i[26946];
  assign o[26945] = i[26945];
  assign o[26944] = i[26944];
  assign o[26943] = i[26943];
  assign o[26942] = i[26942];
  assign o[26941] = i[26941];
  assign o[26940] = i[26940];
  assign o[26939] = i[26939];
  assign o[26938] = i[26938];
  assign o[26937] = i[26937];
  assign o[26936] = i[26936];
  assign o[26935] = i[26935];
  assign o[26934] = i[26934];
  assign o[26933] = i[26933];
  assign o[26932] = i[26932];
  assign o[26931] = i[26931];
  assign o[26930] = i[26930];
  assign o[26929] = i[26929];
  assign o[26928] = i[26928];
  assign o[26927] = i[26927];
  assign o[26926] = i[26926];
  assign o[26925] = i[26925];
  assign o[26924] = i[26924];
  assign o[26923] = i[26923];
  assign o[26922] = i[26922];
  assign o[26921] = i[26921];
  assign o[26920] = i[26920];
  assign o[26919] = i[26919];
  assign o[26918] = i[26918];
  assign o[26917] = i[26917];
  assign o[26916] = i[26916];
  assign o[26915] = i[26915];
  assign o[26914] = i[26914];
  assign o[26913] = i[26913];
  assign o[26912] = i[26912];
  assign o[26911] = i[26911];
  assign o[26910] = i[26910];
  assign o[26909] = i[26909];
  assign o[26908] = i[26908];
  assign o[26907] = i[26907];
  assign o[26906] = i[26906];
  assign o[26905] = i[26905];
  assign o[26904] = i[26904];
  assign o[26903] = i[26903];
  assign o[26902] = i[26902];
  assign o[26901] = i[26901];
  assign o[26900] = i[26900];
  assign o[26899] = i[26899];
  assign o[26898] = i[26898];
  assign o[26897] = i[26897];
  assign o[26896] = i[26896];
  assign o[26895] = i[26895];
  assign o[26894] = i[26894];
  assign o[26893] = i[26893];
  assign o[26892] = i[26892];
  assign o[26891] = i[26891];
  assign o[26890] = i[26890];
  assign o[26889] = i[26889];
  assign o[26888] = i[26888];
  assign o[26887] = i[26887];
  assign o[26886] = i[26886];
  assign o[26885] = i[26885];
  assign o[26884] = i[26884];
  assign o[26883] = i[26883];
  assign o[26882] = i[26882];
  assign o[26881] = i[26881];
  assign o[26880] = i[26880];
  assign o[26879] = i[26879];
  assign o[26878] = i[26878];
  assign o[26877] = i[26877];
  assign o[26876] = i[26876];
  assign o[26875] = i[26875];
  assign o[26874] = i[26874];
  assign o[26873] = i[26873];
  assign o[26872] = i[26872];
  assign o[26871] = i[26871];
  assign o[26870] = i[26870];
  assign o[26869] = i[26869];
  assign o[26868] = i[26868];
  assign o[26867] = i[26867];
  assign o[26866] = i[26866];
  assign o[26865] = i[26865];
  assign o[26864] = i[26864];
  assign o[26863] = i[26863];
  assign o[26862] = i[26862];
  assign o[26861] = i[26861];
  assign o[26860] = i[26860];
  assign o[26859] = i[26859];
  assign o[26858] = i[26858];
  assign o[26857] = i[26857];
  assign o[26856] = i[26856];
  assign o[26855] = i[26855];
  assign o[26854] = i[26854];
  assign o[26853] = i[26853];
  assign o[26852] = i[26852];
  assign o[26851] = i[26851];
  assign o[26850] = i[26850];
  assign o[26849] = i[26849];
  assign o[26848] = i[26848];
  assign o[26847] = i[26847];
  assign o[26846] = i[26846];
  assign o[26845] = i[26845];
  assign o[26844] = i[26844];
  assign o[26843] = i[26843];
  assign o[26842] = i[26842];
  assign o[26841] = i[26841];
  assign o[26840] = i[26840];
  assign o[26839] = i[26839];
  assign o[26838] = i[26838];
  assign o[26837] = i[26837];
  assign o[26836] = i[26836];
  assign o[26835] = i[26835];
  assign o[26834] = i[26834];
  assign o[26833] = i[26833];
  assign o[26832] = i[26832];
  assign o[26831] = i[26831];
  assign o[26830] = i[26830];
  assign o[26829] = i[26829];
  assign o[26828] = i[26828];
  assign o[26827] = i[26827];
  assign o[26826] = i[26826];
  assign o[26825] = i[26825];
  assign o[26824] = i[26824];
  assign o[26823] = i[26823];
  assign o[26822] = i[26822];
  assign o[26821] = i[26821];
  assign o[26820] = i[26820];
  assign o[26819] = i[26819];
  assign o[26818] = i[26818];
  assign o[26817] = i[26817];
  assign o[26816] = i[26816];
  assign o[26815] = i[26815];
  assign o[26814] = i[26814];
  assign o[26813] = i[26813];
  assign o[26812] = i[26812];
  assign o[26811] = i[26811];
  assign o[26810] = i[26810];
  assign o[26809] = i[26809];
  assign o[26808] = i[26808];
  assign o[26807] = i[26807];
  assign o[26806] = i[26806];
  assign o[26805] = i[26805];
  assign o[26804] = i[26804];
  assign o[26803] = i[26803];
  assign o[26802] = i[26802];
  assign o[26801] = i[26801];
  assign o[26800] = i[26800];
  assign o[26799] = i[26799];
  assign o[26798] = i[26798];
  assign o[26797] = i[26797];
  assign o[26796] = i[26796];
  assign o[26795] = i[26795];
  assign o[26794] = i[26794];
  assign o[26793] = i[26793];
  assign o[26792] = i[26792];
  assign o[26791] = i[26791];
  assign o[26790] = i[26790];
  assign o[26789] = i[26789];
  assign o[26788] = i[26788];
  assign o[26787] = i[26787];
  assign o[26786] = i[26786];
  assign o[26785] = i[26785];
  assign o[26784] = i[26784];
  assign o[26783] = i[26783];
  assign o[26782] = i[26782];
  assign o[26781] = i[26781];
  assign o[26780] = i[26780];
  assign o[26779] = i[26779];
  assign o[26778] = i[26778];
  assign o[26777] = i[26777];
  assign o[26776] = i[26776];
  assign o[26775] = i[26775];
  assign o[26774] = i[26774];
  assign o[26773] = i[26773];
  assign o[26772] = i[26772];
  assign o[26771] = i[26771];
  assign o[26770] = i[26770];
  assign o[26769] = i[26769];
  assign o[26768] = i[26768];
  assign o[26767] = i[26767];
  assign o[26766] = i[26766];
  assign o[26765] = i[26765];
  assign o[26764] = i[26764];
  assign o[26763] = i[26763];
  assign o[26762] = i[26762];
  assign o[26761] = i[26761];
  assign o[26760] = i[26760];
  assign o[26759] = i[26759];
  assign o[26758] = i[26758];
  assign o[26757] = i[26757];
  assign o[26756] = i[26756];
  assign o[26755] = i[26755];
  assign o[26754] = i[26754];
  assign o[26753] = i[26753];
  assign o[26752] = i[26752];
  assign o[26751] = i[26751];
  assign o[26750] = i[26750];
  assign o[26749] = i[26749];
  assign o[26748] = i[26748];
  assign o[26747] = i[26747];
  assign o[26746] = i[26746];
  assign o[26745] = i[26745];
  assign o[26744] = i[26744];
  assign o[26743] = i[26743];
  assign o[26742] = i[26742];
  assign o[26741] = i[26741];
  assign o[26740] = i[26740];
  assign o[26739] = i[26739];
  assign o[26738] = i[26738];
  assign o[26737] = i[26737];
  assign o[26736] = i[26736];
  assign o[26735] = i[26735];
  assign o[26734] = i[26734];
  assign o[26733] = i[26733];
  assign o[26732] = i[26732];
  assign o[26731] = i[26731];
  assign o[26730] = i[26730];
  assign o[26729] = i[26729];
  assign o[26728] = i[26728];
  assign o[26727] = i[26727];
  assign o[26726] = i[26726];
  assign o[26725] = i[26725];
  assign o[26724] = i[26724];
  assign o[26723] = i[26723];
  assign o[26722] = i[26722];
  assign o[26721] = i[26721];
  assign o[26720] = i[26720];
  assign o[26719] = i[26719];
  assign o[26718] = i[26718];
  assign o[26717] = i[26717];
  assign o[26716] = i[26716];
  assign o[26715] = i[26715];
  assign o[26714] = i[26714];
  assign o[26713] = i[26713];
  assign o[26712] = i[26712];
  assign o[26711] = i[26711];
  assign o[26710] = i[26710];
  assign o[26709] = i[26709];
  assign o[26708] = i[26708];
  assign o[26707] = i[26707];
  assign o[26706] = i[26706];
  assign o[26705] = i[26705];
  assign o[26704] = i[26704];
  assign o[26703] = i[26703];
  assign o[26702] = i[26702];
  assign o[26701] = i[26701];
  assign o[26700] = i[26700];
  assign o[26699] = i[26699];
  assign o[26698] = i[26698];
  assign o[26697] = i[26697];
  assign o[26696] = i[26696];
  assign o[26695] = i[26695];
  assign o[26694] = i[26694];
  assign o[26693] = i[26693];
  assign o[26692] = i[26692];
  assign o[26691] = i[26691];
  assign o[26690] = i[26690];
  assign o[26689] = i[26689];
  assign o[26688] = i[26688];
  assign o[26687] = i[26687];
  assign o[26686] = i[26686];
  assign o[26685] = i[26685];
  assign o[26684] = i[26684];
  assign o[26683] = i[26683];
  assign o[26682] = i[26682];
  assign o[26681] = i[26681];
  assign o[26680] = i[26680];
  assign o[26679] = i[26679];
  assign o[26678] = i[26678];
  assign o[26677] = i[26677];
  assign o[26676] = i[26676];
  assign o[26675] = i[26675];
  assign o[26674] = i[26674];
  assign o[26673] = i[26673];
  assign o[26672] = i[26672];
  assign o[26671] = i[26671];
  assign o[26670] = i[26670];
  assign o[26669] = i[26669];
  assign o[26668] = i[26668];
  assign o[26667] = i[26667];
  assign o[26666] = i[26666];
  assign o[26665] = i[26665];
  assign o[26664] = i[26664];
  assign o[26663] = i[26663];
  assign o[26662] = i[26662];
  assign o[26661] = i[26661];
  assign o[26660] = i[26660];
  assign o[26659] = i[26659];
  assign o[26658] = i[26658];
  assign o[26657] = i[26657];
  assign o[26656] = i[26656];
  assign o[26655] = i[26655];
  assign o[26654] = i[26654];
  assign o[26653] = i[26653];
  assign o[26652] = i[26652];
  assign o[26651] = i[26651];
  assign o[26650] = i[26650];
  assign o[26649] = i[26649];
  assign o[26648] = i[26648];
  assign o[26647] = i[26647];
  assign o[26646] = i[26646];
  assign o[26645] = i[26645];
  assign o[26644] = i[26644];
  assign o[26643] = i[26643];
  assign o[26642] = i[26642];
  assign o[26641] = i[26641];
  assign o[26640] = i[26640];
  assign o[26639] = i[26639];
  assign o[26638] = i[26638];
  assign o[26637] = i[26637];
  assign o[26636] = i[26636];
  assign o[26635] = i[26635];
  assign o[26634] = i[26634];
  assign o[26633] = i[26633];
  assign o[26632] = i[26632];
  assign o[26631] = i[26631];
  assign o[26630] = i[26630];
  assign o[26629] = i[26629];
  assign o[26628] = i[26628];
  assign o[26627] = i[26627];
  assign o[26626] = i[26626];
  assign o[26625] = i[26625];
  assign o[26624] = i[26624];
  assign o[26623] = i[26623];
  assign o[26622] = i[26622];
  assign o[26621] = i[26621];
  assign o[26620] = i[26620];
  assign o[26619] = i[26619];
  assign o[26618] = i[26618];
  assign o[26617] = i[26617];
  assign o[26616] = i[26616];
  assign o[26615] = i[26615];
  assign o[26614] = i[26614];
  assign o[26613] = i[26613];
  assign o[26612] = i[26612];
  assign o[26611] = i[26611];
  assign o[26610] = i[26610];
  assign o[26609] = i[26609];
  assign o[26608] = i[26608];
  assign o[26607] = i[26607];
  assign o[26606] = i[26606];
  assign o[26605] = i[26605];
  assign o[26604] = i[26604];
  assign o[26603] = i[26603];
  assign o[26602] = i[26602];
  assign o[26601] = i[26601];
  assign o[26600] = i[26600];
  assign o[26599] = i[26599];
  assign o[26598] = i[26598];
  assign o[26597] = i[26597];
  assign o[26596] = i[26596];
  assign o[26595] = i[26595];
  assign o[26594] = i[26594];
  assign o[26593] = i[26593];
  assign o[26592] = i[26592];
  assign o[26591] = i[26591];
  assign o[26590] = i[26590];
  assign o[26589] = i[26589];
  assign o[26588] = i[26588];
  assign o[26587] = i[26587];
  assign o[26586] = i[26586];
  assign o[26585] = i[26585];
  assign o[26584] = i[26584];
  assign o[26583] = i[26583];
  assign o[26582] = i[26582];
  assign o[26581] = i[26581];
  assign o[26580] = i[26580];
  assign o[26579] = i[26579];
  assign o[26578] = i[26578];
  assign o[26577] = i[26577];
  assign o[26576] = i[26576];
  assign o[26575] = i[26575];
  assign o[26574] = i[26574];
  assign o[26573] = i[26573];
  assign o[26572] = i[26572];
  assign o[26571] = i[26571];
  assign o[26570] = i[26570];
  assign o[26569] = i[26569];
  assign o[26568] = i[26568];
  assign o[26567] = i[26567];
  assign o[26566] = i[26566];
  assign o[26565] = i[26565];
  assign o[26564] = i[26564];
  assign o[26563] = i[26563];
  assign o[26562] = i[26562];
  assign o[26561] = i[26561];
  assign o[26560] = i[26560];
  assign o[26559] = i[26559];
  assign o[26558] = i[26558];
  assign o[26557] = i[26557];
  assign o[26556] = i[26556];
  assign o[26555] = i[26555];
  assign o[26554] = i[26554];
  assign o[26553] = i[26553];
  assign o[26552] = i[26552];
  assign o[26551] = i[26551];
  assign o[26550] = i[26550];
  assign o[26549] = i[26549];
  assign o[26548] = i[26548];
  assign o[26547] = i[26547];
  assign o[26546] = i[26546];
  assign o[26545] = i[26545];
  assign o[26544] = i[26544];
  assign o[26543] = i[26543];
  assign o[26542] = i[26542];
  assign o[26541] = i[26541];
  assign o[26540] = i[26540];
  assign o[26539] = i[26539];
  assign o[26538] = i[26538];
  assign o[26537] = i[26537];
  assign o[26536] = i[26536];
  assign o[26535] = i[26535];
  assign o[26534] = i[26534];
  assign o[26533] = i[26533];
  assign o[26532] = i[26532];
  assign o[26531] = i[26531];
  assign o[26530] = i[26530];
  assign o[26529] = i[26529];
  assign o[26528] = i[26528];
  assign o[26527] = i[26527];
  assign o[26526] = i[26526];
  assign o[26525] = i[26525];
  assign o[26524] = i[26524];
  assign o[26523] = i[26523];
  assign o[26522] = i[26522];
  assign o[26521] = i[26521];
  assign o[26520] = i[26520];
  assign o[26519] = i[26519];
  assign o[26518] = i[26518];
  assign o[26517] = i[26517];
  assign o[26516] = i[26516];
  assign o[26515] = i[26515];
  assign o[26514] = i[26514];
  assign o[26513] = i[26513];
  assign o[26512] = i[26512];
  assign o[26511] = i[26511];
  assign o[26510] = i[26510];
  assign o[26509] = i[26509];
  assign o[26508] = i[26508];
  assign o[26507] = i[26507];
  assign o[26506] = i[26506];
  assign o[26505] = i[26505];
  assign o[26504] = i[26504];
  assign o[26503] = i[26503];
  assign o[26502] = i[26502];
  assign o[26501] = i[26501];
  assign o[26500] = i[26500];
  assign o[26499] = i[26499];
  assign o[26498] = i[26498];
  assign o[26497] = i[26497];
  assign o[26496] = i[26496];
  assign o[26495] = i[26495];
  assign o[26494] = i[26494];
  assign o[26493] = i[26493];
  assign o[26492] = i[26492];
  assign o[26491] = i[26491];
  assign o[26490] = i[26490];
  assign o[26489] = i[26489];
  assign o[26488] = i[26488];
  assign o[26487] = i[26487];
  assign o[26486] = i[26486];
  assign o[26485] = i[26485];
  assign o[26484] = i[26484];
  assign o[26483] = i[26483];
  assign o[26482] = i[26482];
  assign o[26481] = i[26481];
  assign o[26480] = i[26480];
  assign o[26479] = i[26479];
  assign o[26478] = i[26478];
  assign o[26477] = i[26477];
  assign o[26476] = i[26476];
  assign o[26475] = i[26475];
  assign o[26474] = i[26474];
  assign o[26473] = i[26473];
  assign o[26472] = i[26472];
  assign o[26471] = i[26471];
  assign o[26470] = i[26470];
  assign o[26469] = i[26469];
  assign o[26468] = i[26468];
  assign o[26467] = i[26467];
  assign o[26466] = i[26466];
  assign o[26465] = i[26465];
  assign o[26464] = i[26464];
  assign o[26463] = i[26463];
  assign o[26462] = i[26462];
  assign o[26461] = i[26461];
  assign o[26460] = i[26460];
  assign o[26459] = i[26459];
  assign o[26458] = i[26458];
  assign o[26457] = i[26457];
  assign o[26456] = i[26456];
  assign o[26455] = i[26455];
  assign o[26454] = i[26454];
  assign o[26453] = i[26453];
  assign o[26452] = i[26452];
  assign o[26451] = i[26451];
  assign o[26450] = i[26450];
  assign o[26449] = i[26449];
  assign o[26448] = i[26448];
  assign o[26447] = i[26447];
  assign o[26446] = i[26446];
  assign o[26445] = i[26445];
  assign o[26444] = i[26444];
  assign o[26443] = i[26443];
  assign o[26442] = i[26442];
  assign o[26441] = i[26441];
  assign o[26440] = i[26440];
  assign o[26439] = i[26439];
  assign o[26438] = i[26438];
  assign o[26437] = i[26437];
  assign o[26436] = i[26436];
  assign o[26435] = i[26435];
  assign o[26434] = i[26434];
  assign o[26433] = i[26433];
  assign o[26432] = i[26432];
  assign o[26431] = i[26431];
  assign o[26430] = i[26430];
  assign o[26429] = i[26429];
  assign o[26428] = i[26428];
  assign o[26427] = i[26427];
  assign o[26426] = i[26426];
  assign o[26425] = i[26425];
  assign o[26424] = i[26424];
  assign o[26423] = i[26423];
  assign o[26422] = i[26422];
  assign o[26421] = i[26421];
  assign o[26420] = i[26420];
  assign o[26419] = i[26419];
  assign o[26418] = i[26418];
  assign o[26417] = i[26417];
  assign o[26416] = i[26416];
  assign o[26415] = i[26415];
  assign o[26414] = i[26414];
  assign o[26413] = i[26413];
  assign o[26412] = i[26412];
  assign o[26411] = i[26411];
  assign o[26410] = i[26410];
  assign o[26409] = i[26409];
  assign o[26408] = i[26408];
  assign o[26407] = i[26407];
  assign o[26406] = i[26406];
  assign o[26405] = i[26405];
  assign o[26404] = i[26404];
  assign o[26403] = i[26403];
  assign o[26402] = i[26402];
  assign o[26401] = i[26401];
  assign o[26400] = i[26400];
  assign o[26399] = i[26399];
  assign o[26398] = i[26398];
  assign o[26397] = i[26397];
  assign o[26396] = i[26396];
  assign o[26395] = i[26395];
  assign o[26394] = i[26394];
  assign o[26393] = i[26393];
  assign o[26392] = i[26392];
  assign o[26391] = i[26391];
  assign o[26390] = i[26390];
  assign o[26389] = i[26389];
  assign o[26388] = i[26388];
  assign o[26387] = i[26387];
  assign o[26386] = i[26386];
  assign o[26385] = i[26385];
  assign o[26384] = i[26384];
  assign o[26383] = i[26383];
  assign o[26382] = i[26382];
  assign o[26381] = i[26381];
  assign o[26380] = i[26380];
  assign o[26379] = i[26379];
  assign o[26378] = i[26378];
  assign o[26377] = i[26377];
  assign o[26376] = i[26376];
  assign o[26375] = i[26375];
  assign o[26374] = i[26374];
  assign o[26373] = i[26373];
  assign o[26372] = i[26372];
  assign o[26371] = i[26371];
  assign o[26370] = i[26370];
  assign o[26369] = i[26369];
  assign o[26368] = i[26368];
  assign o[26367] = i[26367];
  assign o[26366] = i[26366];
  assign o[26365] = i[26365];
  assign o[26364] = i[26364];
  assign o[26363] = i[26363];
  assign o[26362] = i[26362];
  assign o[26361] = i[26361];
  assign o[26360] = i[26360];
  assign o[26359] = i[26359];
  assign o[26358] = i[26358];
  assign o[26357] = i[26357];
  assign o[26356] = i[26356];
  assign o[26355] = i[26355];
  assign o[26354] = i[26354];
  assign o[26353] = i[26353];
  assign o[26352] = i[26352];
  assign o[26351] = i[26351];
  assign o[26350] = i[26350];
  assign o[26349] = i[26349];
  assign o[26348] = i[26348];
  assign o[26347] = i[26347];
  assign o[26346] = i[26346];
  assign o[26345] = i[26345];
  assign o[26344] = i[26344];
  assign o[26343] = i[26343];
  assign o[26342] = i[26342];
  assign o[26341] = i[26341];
  assign o[26340] = i[26340];
  assign o[26339] = i[26339];
  assign o[26338] = i[26338];
  assign o[26337] = i[26337];
  assign o[26336] = i[26336];
  assign o[26335] = i[26335];
  assign o[26334] = i[26334];
  assign o[26333] = i[26333];
  assign o[26332] = i[26332];
  assign o[26331] = i[26331];
  assign o[26330] = i[26330];
  assign o[26329] = i[26329];
  assign o[26328] = i[26328];
  assign o[26327] = i[26327];
  assign o[26326] = i[26326];
  assign o[26325] = i[26325];
  assign o[26324] = i[26324];
  assign o[26323] = i[26323];
  assign o[26322] = i[26322];
  assign o[26321] = i[26321];
  assign o[26320] = i[26320];
  assign o[26319] = i[26319];
  assign o[26318] = i[26318];
  assign o[26317] = i[26317];
  assign o[26316] = i[26316];
  assign o[26315] = i[26315];
  assign o[26314] = i[26314];
  assign o[26313] = i[26313];
  assign o[26312] = i[26312];
  assign o[26311] = i[26311];
  assign o[26310] = i[26310];
  assign o[26309] = i[26309];
  assign o[26308] = i[26308];
  assign o[26307] = i[26307];
  assign o[26306] = i[26306];
  assign o[26305] = i[26305];
  assign o[26304] = i[26304];
  assign o[26303] = i[26303];
  assign o[26302] = i[26302];
  assign o[26301] = i[26301];
  assign o[26300] = i[26300];
  assign o[26299] = i[26299];
  assign o[26298] = i[26298];
  assign o[26297] = i[26297];
  assign o[26296] = i[26296];
  assign o[26295] = i[26295];
  assign o[26294] = i[26294];
  assign o[26293] = i[26293];
  assign o[26292] = i[26292];
  assign o[26291] = i[26291];
  assign o[26290] = i[26290];
  assign o[26289] = i[26289];
  assign o[26288] = i[26288];
  assign o[26287] = i[26287];
  assign o[26286] = i[26286];
  assign o[26285] = i[26285];
  assign o[26284] = i[26284];
  assign o[26283] = i[26283];
  assign o[26282] = i[26282];
  assign o[26281] = i[26281];
  assign o[26280] = i[26280];
  assign o[26279] = i[26279];
  assign o[26278] = i[26278];
  assign o[26277] = i[26277];
  assign o[26276] = i[26276];
  assign o[26275] = i[26275];
  assign o[26274] = i[26274];
  assign o[26273] = i[26273];
  assign o[26272] = i[26272];
  assign o[26271] = i[26271];
  assign o[26270] = i[26270];
  assign o[26269] = i[26269];
  assign o[26268] = i[26268];
  assign o[26267] = i[26267];
  assign o[26266] = i[26266];
  assign o[26265] = i[26265];
  assign o[26264] = i[26264];
  assign o[26263] = i[26263];
  assign o[26262] = i[26262];
  assign o[26261] = i[26261];
  assign o[26260] = i[26260];
  assign o[26259] = i[26259];
  assign o[26258] = i[26258];
  assign o[26257] = i[26257];
  assign o[26256] = i[26256];
  assign o[26255] = i[26255];
  assign o[26254] = i[26254];
  assign o[26253] = i[26253];
  assign o[26252] = i[26252];
  assign o[26251] = i[26251];
  assign o[26250] = i[26250];
  assign o[26249] = i[26249];
  assign o[26248] = i[26248];
  assign o[26247] = i[26247];
  assign o[26246] = i[26246];
  assign o[26245] = i[26245];
  assign o[26244] = i[26244];
  assign o[26243] = i[26243];
  assign o[26242] = i[26242];
  assign o[26241] = i[26241];
  assign o[26240] = i[26240];
  assign o[26239] = i[26239];
  assign o[26238] = i[26238];
  assign o[26237] = i[26237];
  assign o[26236] = i[26236];
  assign o[26235] = i[26235];
  assign o[26234] = i[26234];
  assign o[26233] = i[26233];
  assign o[26232] = i[26232];
  assign o[26231] = i[26231];
  assign o[26230] = i[26230];
  assign o[26229] = i[26229];
  assign o[26228] = i[26228];
  assign o[26227] = i[26227];
  assign o[26226] = i[26226];
  assign o[26225] = i[26225];
  assign o[26224] = i[26224];
  assign o[26223] = i[26223];
  assign o[26222] = i[26222];
  assign o[26221] = i[26221];
  assign o[26220] = i[26220];
  assign o[26219] = i[26219];
  assign o[26218] = i[26218];
  assign o[26217] = i[26217];
  assign o[26216] = i[26216];
  assign o[26215] = i[26215];
  assign o[26214] = i[26214];
  assign o[26213] = i[26213];
  assign o[26212] = i[26212];
  assign o[26211] = i[26211];
  assign o[26210] = i[26210];
  assign o[26209] = i[26209];
  assign o[26208] = i[26208];
  assign o[26207] = i[26207];
  assign o[26206] = i[26206];
  assign o[26205] = i[26205];
  assign o[26204] = i[26204];
  assign o[26203] = i[26203];
  assign o[26202] = i[26202];
  assign o[26201] = i[26201];
  assign o[26200] = i[26200];
  assign o[26199] = i[26199];
  assign o[26198] = i[26198];
  assign o[26197] = i[26197];
  assign o[26196] = i[26196];
  assign o[26195] = i[26195];
  assign o[26194] = i[26194];
  assign o[26193] = i[26193];
  assign o[26192] = i[26192];
  assign o[26191] = i[26191];
  assign o[26190] = i[26190];
  assign o[26189] = i[26189];
  assign o[26188] = i[26188];
  assign o[26187] = i[26187];
  assign o[26186] = i[26186];
  assign o[26185] = i[26185];
  assign o[26184] = i[26184];
  assign o[26183] = i[26183];
  assign o[26182] = i[26182];
  assign o[26181] = i[26181];
  assign o[26180] = i[26180];
  assign o[26179] = i[26179];
  assign o[26178] = i[26178];
  assign o[26177] = i[26177];
  assign o[26176] = i[26176];
  assign o[26175] = i[26175];
  assign o[26174] = i[26174];
  assign o[26173] = i[26173];
  assign o[26172] = i[26172];
  assign o[26171] = i[26171];
  assign o[26170] = i[26170];
  assign o[26169] = i[26169];
  assign o[26168] = i[26168];
  assign o[26167] = i[26167];
  assign o[26166] = i[26166];
  assign o[26165] = i[26165];
  assign o[26164] = i[26164];
  assign o[26163] = i[26163];
  assign o[26162] = i[26162];
  assign o[26161] = i[26161];
  assign o[26160] = i[26160];
  assign o[26159] = i[26159];
  assign o[26158] = i[26158];
  assign o[26157] = i[26157];
  assign o[26156] = i[26156];
  assign o[26155] = i[26155];
  assign o[26154] = i[26154];
  assign o[26153] = i[26153];
  assign o[26152] = i[26152];
  assign o[26151] = i[26151];
  assign o[26150] = i[26150];
  assign o[26149] = i[26149];
  assign o[26148] = i[26148];
  assign o[26147] = i[26147];
  assign o[26146] = i[26146];
  assign o[26145] = i[26145];
  assign o[26144] = i[26144];
  assign o[26143] = i[26143];
  assign o[26142] = i[26142];
  assign o[26141] = i[26141];
  assign o[26140] = i[26140];
  assign o[26139] = i[26139];
  assign o[26138] = i[26138];
  assign o[26137] = i[26137];
  assign o[26136] = i[26136];
  assign o[26135] = i[26135];
  assign o[26134] = i[26134];
  assign o[26133] = i[26133];
  assign o[26132] = i[26132];
  assign o[26131] = i[26131];
  assign o[26130] = i[26130];
  assign o[26129] = i[26129];
  assign o[26128] = i[26128];
  assign o[26127] = i[26127];
  assign o[26126] = i[26126];
  assign o[26125] = i[26125];
  assign o[26124] = i[26124];
  assign o[26123] = i[26123];
  assign o[26122] = i[26122];
  assign o[26121] = i[26121];
  assign o[26120] = i[26120];
  assign o[26119] = i[26119];
  assign o[26118] = i[26118];
  assign o[26117] = i[26117];
  assign o[26116] = i[26116];
  assign o[26115] = i[26115];
  assign o[26114] = i[26114];
  assign o[26113] = i[26113];
  assign o[26112] = i[26112];
  assign o[26111] = i[26111];
  assign o[26110] = i[26110];
  assign o[26109] = i[26109];
  assign o[26108] = i[26108];
  assign o[26107] = i[26107];
  assign o[26106] = i[26106];
  assign o[26105] = i[26105];
  assign o[26104] = i[26104];
  assign o[26103] = i[26103];
  assign o[26102] = i[26102];
  assign o[26101] = i[26101];
  assign o[26100] = i[26100];
  assign o[26099] = i[26099];
  assign o[26098] = i[26098];
  assign o[26097] = i[26097];
  assign o[26096] = i[26096];
  assign o[26095] = i[26095];
  assign o[26094] = i[26094];
  assign o[26093] = i[26093];
  assign o[26092] = i[26092];
  assign o[26091] = i[26091];
  assign o[26090] = i[26090];
  assign o[26089] = i[26089];
  assign o[26088] = i[26088];
  assign o[26087] = i[26087];
  assign o[26086] = i[26086];
  assign o[26085] = i[26085];
  assign o[26084] = i[26084];
  assign o[26083] = i[26083];
  assign o[26082] = i[26082];
  assign o[26081] = i[26081];
  assign o[26080] = i[26080];
  assign o[26079] = i[26079];
  assign o[26078] = i[26078];
  assign o[26077] = i[26077];
  assign o[26076] = i[26076];
  assign o[26075] = i[26075];
  assign o[26074] = i[26074];
  assign o[26073] = i[26073];
  assign o[26072] = i[26072];
  assign o[26071] = i[26071];
  assign o[26070] = i[26070];
  assign o[26069] = i[26069];
  assign o[26068] = i[26068];
  assign o[26067] = i[26067];
  assign o[26066] = i[26066];
  assign o[26065] = i[26065];
  assign o[26064] = i[26064];
  assign o[26063] = i[26063];
  assign o[26062] = i[26062];
  assign o[26061] = i[26061];
  assign o[26060] = i[26060];
  assign o[26059] = i[26059];
  assign o[26058] = i[26058];
  assign o[26057] = i[26057];
  assign o[26056] = i[26056];
  assign o[26055] = i[26055];
  assign o[26054] = i[26054];
  assign o[26053] = i[26053];
  assign o[26052] = i[26052];
  assign o[26051] = i[26051];
  assign o[26050] = i[26050];
  assign o[26049] = i[26049];
  assign o[26048] = i[26048];
  assign o[26047] = i[26047];
  assign o[26046] = i[26046];
  assign o[26045] = i[26045];
  assign o[26044] = i[26044];
  assign o[26043] = i[26043];
  assign o[26042] = i[26042];
  assign o[26041] = i[26041];
  assign o[26040] = i[26040];
  assign o[26039] = i[26039];
  assign o[26038] = i[26038];
  assign o[26037] = i[26037];
  assign o[26036] = i[26036];
  assign o[26035] = i[26035];
  assign o[26034] = i[26034];
  assign o[26033] = i[26033];
  assign o[26032] = i[26032];
  assign o[26031] = i[26031];
  assign o[26030] = i[26030];
  assign o[26029] = i[26029];
  assign o[26028] = i[26028];
  assign o[26027] = i[26027];
  assign o[26026] = i[26026];
  assign o[26025] = i[26025];
  assign o[26024] = i[26024];
  assign o[26023] = i[26023];
  assign o[26022] = i[26022];
  assign o[26021] = i[26021];
  assign o[26020] = i[26020];
  assign o[26019] = i[26019];
  assign o[26018] = i[26018];
  assign o[26017] = i[26017];
  assign o[26016] = i[26016];
  assign o[26015] = i[26015];
  assign o[26014] = i[26014];
  assign o[26013] = i[26013];
  assign o[26012] = i[26012];
  assign o[26011] = i[26011];
  assign o[26010] = i[26010];
  assign o[26009] = i[26009];
  assign o[26008] = i[26008];
  assign o[26007] = i[26007];
  assign o[26006] = i[26006];
  assign o[26005] = i[26005];
  assign o[26004] = i[26004];
  assign o[26003] = i[26003];
  assign o[26002] = i[26002];
  assign o[26001] = i[26001];
  assign o[26000] = i[26000];
  assign o[25999] = i[25999];
  assign o[25998] = i[25998];
  assign o[25997] = i[25997];
  assign o[25996] = i[25996];
  assign o[25995] = i[25995];
  assign o[25994] = i[25994];
  assign o[25993] = i[25993];
  assign o[25992] = i[25992];
  assign o[25991] = i[25991];
  assign o[25990] = i[25990];
  assign o[25989] = i[25989];
  assign o[25988] = i[25988];
  assign o[25987] = i[25987];
  assign o[25986] = i[25986];
  assign o[25985] = i[25985];
  assign o[25984] = i[25984];
  assign o[25983] = i[25983];
  assign o[25982] = i[25982];
  assign o[25981] = i[25981];
  assign o[25980] = i[25980];
  assign o[25979] = i[25979];
  assign o[25978] = i[25978];
  assign o[25977] = i[25977];
  assign o[25976] = i[25976];
  assign o[25975] = i[25975];
  assign o[25974] = i[25974];
  assign o[25973] = i[25973];
  assign o[25972] = i[25972];
  assign o[25971] = i[25971];
  assign o[25970] = i[25970];
  assign o[25969] = i[25969];
  assign o[25968] = i[25968];
  assign o[25967] = i[25967];
  assign o[25966] = i[25966];
  assign o[25965] = i[25965];
  assign o[25964] = i[25964];
  assign o[25963] = i[25963];
  assign o[25962] = i[25962];
  assign o[25961] = i[25961];
  assign o[25960] = i[25960];
  assign o[25959] = i[25959];
  assign o[25958] = i[25958];
  assign o[25957] = i[25957];
  assign o[25956] = i[25956];
  assign o[25955] = i[25955];
  assign o[25954] = i[25954];
  assign o[25953] = i[25953];
  assign o[25952] = i[25952];
  assign o[25951] = i[25951];
  assign o[25950] = i[25950];
  assign o[25949] = i[25949];
  assign o[25948] = i[25948];
  assign o[25947] = i[25947];
  assign o[25946] = i[25946];
  assign o[25945] = i[25945];
  assign o[25944] = i[25944];
  assign o[25943] = i[25943];
  assign o[25942] = i[25942];
  assign o[25941] = i[25941];
  assign o[25940] = i[25940];
  assign o[25939] = i[25939];
  assign o[25938] = i[25938];
  assign o[25937] = i[25937];
  assign o[25936] = i[25936];
  assign o[25935] = i[25935];
  assign o[25934] = i[25934];
  assign o[25933] = i[25933];
  assign o[25932] = i[25932];
  assign o[25931] = i[25931];
  assign o[25930] = i[25930];
  assign o[25929] = i[25929];
  assign o[25928] = i[25928];
  assign o[25927] = i[25927];
  assign o[25926] = i[25926];
  assign o[25925] = i[25925];
  assign o[25924] = i[25924];
  assign o[25923] = i[25923];
  assign o[25922] = i[25922];
  assign o[25921] = i[25921];
  assign o[25920] = i[25920];
  assign o[25919] = i[25919];
  assign o[25918] = i[25918];
  assign o[25917] = i[25917];
  assign o[25916] = i[25916];
  assign o[25915] = i[25915];
  assign o[25914] = i[25914];
  assign o[25913] = i[25913];
  assign o[25912] = i[25912];
  assign o[25911] = i[25911];
  assign o[25910] = i[25910];
  assign o[25909] = i[25909];
  assign o[25908] = i[25908];
  assign o[25907] = i[25907];
  assign o[25906] = i[25906];
  assign o[25905] = i[25905];
  assign o[25904] = i[25904];
  assign o[25903] = i[25903];
  assign o[25902] = i[25902];
  assign o[25901] = i[25901];
  assign o[25900] = i[25900];
  assign o[25899] = i[25899];
  assign o[25898] = i[25898];
  assign o[25897] = i[25897];
  assign o[25896] = i[25896];
  assign o[25895] = i[25895];
  assign o[25894] = i[25894];
  assign o[25893] = i[25893];
  assign o[25892] = i[25892];
  assign o[25891] = i[25891];
  assign o[25890] = i[25890];
  assign o[25889] = i[25889];
  assign o[25888] = i[25888];
  assign o[25887] = i[25887];
  assign o[25886] = i[25886];
  assign o[25885] = i[25885];
  assign o[25884] = i[25884];
  assign o[25883] = i[25883];
  assign o[25882] = i[25882];
  assign o[25881] = i[25881];
  assign o[25880] = i[25880];
  assign o[25879] = i[25879];
  assign o[25878] = i[25878];
  assign o[25877] = i[25877];
  assign o[25876] = i[25876];
  assign o[25875] = i[25875];
  assign o[25874] = i[25874];
  assign o[25873] = i[25873];
  assign o[25872] = i[25872];
  assign o[25871] = i[25871];
  assign o[25870] = i[25870];
  assign o[25869] = i[25869];
  assign o[25868] = i[25868];
  assign o[25867] = i[25867];
  assign o[25866] = i[25866];
  assign o[25865] = i[25865];
  assign o[25864] = i[25864];
  assign o[25863] = i[25863];
  assign o[25862] = i[25862];
  assign o[25861] = i[25861];
  assign o[25860] = i[25860];
  assign o[25859] = i[25859];
  assign o[25858] = i[25858];
  assign o[25857] = i[25857];
  assign o[25856] = i[25856];
  assign o[25855] = i[25855];
  assign o[25854] = i[25854];
  assign o[25853] = i[25853];
  assign o[25852] = i[25852];
  assign o[25851] = i[25851];
  assign o[25850] = i[25850];
  assign o[25849] = i[25849];
  assign o[25848] = i[25848];
  assign o[25847] = i[25847];
  assign o[25846] = i[25846];
  assign o[25845] = i[25845];
  assign o[25844] = i[25844];
  assign o[25843] = i[25843];
  assign o[25842] = i[25842];
  assign o[25841] = i[25841];
  assign o[25840] = i[25840];
  assign o[25839] = i[25839];
  assign o[25838] = i[25838];
  assign o[25837] = i[25837];
  assign o[25836] = i[25836];
  assign o[25835] = i[25835];
  assign o[25834] = i[25834];
  assign o[25833] = i[25833];
  assign o[25832] = i[25832];
  assign o[25831] = i[25831];
  assign o[25830] = i[25830];
  assign o[25829] = i[25829];
  assign o[25828] = i[25828];
  assign o[25827] = i[25827];
  assign o[25826] = i[25826];
  assign o[25825] = i[25825];
  assign o[25824] = i[25824];
  assign o[25823] = i[25823];
  assign o[25822] = i[25822];
  assign o[25821] = i[25821];
  assign o[25820] = i[25820];
  assign o[25819] = i[25819];
  assign o[25818] = i[25818];
  assign o[25817] = i[25817];
  assign o[25816] = i[25816];
  assign o[25815] = i[25815];
  assign o[25814] = i[25814];
  assign o[25813] = i[25813];
  assign o[25812] = i[25812];
  assign o[25811] = i[25811];
  assign o[25810] = i[25810];
  assign o[25809] = i[25809];
  assign o[25808] = i[25808];
  assign o[25807] = i[25807];
  assign o[25806] = i[25806];
  assign o[25805] = i[25805];
  assign o[25804] = i[25804];
  assign o[25803] = i[25803];
  assign o[25802] = i[25802];
  assign o[25801] = i[25801];
  assign o[25800] = i[25800];
  assign o[25799] = i[25799];
  assign o[25798] = i[25798];
  assign o[25797] = i[25797];
  assign o[25796] = i[25796];
  assign o[25795] = i[25795];
  assign o[25794] = i[25794];
  assign o[25793] = i[25793];
  assign o[25792] = i[25792];
  assign o[25791] = i[25791];
  assign o[25790] = i[25790];
  assign o[25789] = i[25789];
  assign o[25788] = i[25788];
  assign o[25787] = i[25787];
  assign o[25786] = i[25786];
  assign o[25785] = i[25785];
  assign o[25784] = i[25784];
  assign o[25783] = i[25783];
  assign o[25782] = i[25782];
  assign o[25781] = i[25781];
  assign o[25780] = i[25780];
  assign o[25779] = i[25779];
  assign o[25778] = i[25778];
  assign o[25777] = i[25777];
  assign o[25776] = i[25776];
  assign o[25775] = i[25775];
  assign o[25774] = i[25774];
  assign o[25773] = i[25773];
  assign o[25772] = i[25772];
  assign o[25771] = i[25771];
  assign o[25770] = i[25770];
  assign o[25769] = i[25769];
  assign o[25768] = i[25768];
  assign o[25767] = i[25767];
  assign o[25766] = i[25766];
  assign o[25765] = i[25765];
  assign o[25764] = i[25764];
  assign o[25763] = i[25763];
  assign o[25762] = i[25762];
  assign o[25761] = i[25761];
  assign o[25760] = i[25760];
  assign o[25759] = i[25759];
  assign o[25758] = i[25758];
  assign o[25757] = i[25757];
  assign o[25756] = i[25756];
  assign o[25755] = i[25755];
  assign o[25754] = i[25754];
  assign o[25753] = i[25753];
  assign o[25752] = i[25752];
  assign o[25751] = i[25751];
  assign o[25750] = i[25750];
  assign o[25749] = i[25749];
  assign o[25748] = i[25748];
  assign o[25747] = i[25747];
  assign o[25746] = i[25746];
  assign o[25745] = i[25745];
  assign o[25744] = i[25744];
  assign o[25743] = i[25743];
  assign o[25742] = i[25742];
  assign o[25741] = i[25741];
  assign o[25740] = i[25740];
  assign o[25739] = i[25739];
  assign o[25738] = i[25738];
  assign o[25737] = i[25737];
  assign o[25736] = i[25736];
  assign o[25735] = i[25735];
  assign o[25734] = i[25734];
  assign o[25733] = i[25733];
  assign o[25732] = i[25732];
  assign o[25731] = i[25731];
  assign o[25730] = i[25730];
  assign o[25729] = i[25729];
  assign o[25728] = i[25728];
  assign o[25727] = i[25727];
  assign o[25726] = i[25726];
  assign o[25725] = i[25725];
  assign o[25724] = i[25724];
  assign o[25723] = i[25723];
  assign o[25722] = i[25722];
  assign o[25721] = i[25721];
  assign o[25720] = i[25720];
  assign o[25719] = i[25719];
  assign o[25718] = i[25718];
  assign o[25717] = i[25717];
  assign o[25716] = i[25716];
  assign o[25715] = i[25715];
  assign o[25714] = i[25714];
  assign o[25713] = i[25713];
  assign o[25712] = i[25712];
  assign o[25711] = i[25711];
  assign o[25710] = i[25710];
  assign o[25709] = i[25709];
  assign o[25708] = i[25708];
  assign o[25707] = i[25707];
  assign o[25706] = i[25706];
  assign o[25705] = i[25705];
  assign o[25704] = i[25704];
  assign o[25703] = i[25703];
  assign o[25702] = i[25702];
  assign o[25701] = i[25701];
  assign o[25700] = i[25700];
  assign o[25699] = i[25699];
  assign o[25698] = i[25698];
  assign o[25697] = i[25697];
  assign o[25696] = i[25696];
  assign o[25695] = i[25695];
  assign o[25694] = i[25694];
  assign o[25693] = i[25693];
  assign o[25692] = i[25692];
  assign o[25691] = i[25691];
  assign o[25690] = i[25690];
  assign o[25689] = i[25689];
  assign o[25688] = i[25688];
  assign o[25687] = i[25687];
  assign o[25686] = i[25686];
  assign o[25685] = i[25685];
  assign o[25684] = i[25684];
  assign o[25683] = i[25683];
  assign o[25682] = i[25682];
  assign o[25681] = i[25681];
  assign o[25680] = i[25680];
  assign o[25679] = i[25679];
  assign o[25678] = i[25678];
  assign o[25677] = i[25677];
  assign o[25676] = i[25676];
  assign o[25675] = i[25675];
  assign o[25674] = i[25674];
  assign o[25673] = i[25673];
  assign o[25672] = i[25672];
  assign o[25671] = i[25671];
  assign o[25670] = i[25670];
  assign o[25669] = i[25669];
  assign o[25668] = i[25668];
  assign o[25667] = i[25667];
  assign o[25666] = i[25666];
  assign o[25665] = i[25665];
  assign o[25664] = i[25664];
  assign o[25663] = i[25663];
  assign o[25662] = i[25662];
  assign o[25661] = i[25661];
  assign o[25660] = i[25660];
  assign o[25659] = i[25659];
  assign o[25658] = i[25658];
  assign o[25657] = i[25657];
  assign o[25656] = i[25656];
  assign o[25655] = i[25655];
  assign o[25654] = i[25654];
  assign o[25653] = i[25653];
  assign o[25652] = i[25652];
  assign o[25651] = i[25651];
  assign o[25650] = i[25650];
  assign o[25649] = i[25649];
  assign o[25648] = i[25648];
  assign o[25647] = i[25647];
  assign o[25646] = i[25646];
  assign o[25645] = i[25645];
  assign o[25644] = i[25644];
  assign o[25643] = i[25643];
  assign o[25642] = i[25642];
  assign o[25641] = i[25641];
  assign o[25640] = i[25640];
  assign o[25639] = i[25639];
  assign o[25638] = i[25638];
  assign o[25637] = i[25637];
  assign o[25636] = i[25636];
  assign o[25635] = i[25635];
  assign o[25634] = i[25634];
  assign o[25633] = i[25633];
  assign o[25632] = i[25632];
  assign o[25631] = i[25631];
  assign o[25630] = i[25630];
  assign o[25629] = i[25629];
  assign o[25628] = i[25628];
  assign o[25627] = i[25627];
  assign o[25626] = i[25626];
  assign o[25625] = i[25625];
  assign o[25624] = i[25624];
  assign o[25623] = i[25623];
  assign o[25622] = i[25622];
  assign o[25621] = i[25621];
  assign o[25620] = i[25620];
  assign o[25619] = i[25619];
  assign o[25618] = i[25618];
  assign o[25617] = i[25617];
  assign o[25616] = i[25616];
  assign o[25615] = i[25615];
  assign o[25614] = i[25614];
  assign o[25613] = i[25613];
  assign o[25612] = i[25612];
  assign o[25611] = i[25611];
  assign o[25610] = i[25610];
  assign o[25609] = i[25609];
  assign o[25608] = i[25608];
  assign o[25607] = i[25607];
  assign o[25606] = i[25606];
  assign o[25605] = i[25605];
  assign o[25604] = i[25604];
  assign o[25603] = i[25603];
  assign o[25602] = i[25602];
  assign o[25601] = i[25601];
  assign o[25600] = i[25600];
  assign o[25599] = i[25599];
  assign o[25598] = i[25598];
  assign o[25597] = i[25597];
  assign o[25596] = i[25596];
  assign o[25595] = i[25595];
  assign o[25594] = i[25594];
  assign o[25593] = i[25593];
  assign o[25592] = i[25592];
  assign o[25591] = i[25591];
  assign o[25590] = i[25590];
  assign o[25589] = i[25589];
  assign o[25588] = i[25588];
  assign o[25587] = i[25587];
  assign o[25586] = i[25586];
  assign o[25585] = i[25585];
  assign o[25584] = i[25584];
  assign o[25583] = i[25583];
  assign o[25582] = i[25582];
  assign o[25581] = i[25581];
  assign o[25580] = i[25580];
  assign o[25579] = i[25579];
  assign o[25578] = i[25578];
  assign o[25577] = i[25577];
  assign o[25576] = i[25576];
  assign o[25575] = i[25575];
  assign o[25574] = i[25574];
  assign o[25573] = i[25573];
  assign o[25572] = i[25572];
  assign o[25571] = i[25571];
  assign o[25570] = i[25570];
  assign o[25569] = i[25569];
  assign o[25568] = i[25568];
  assign o[25567] = i[25567];
  assign o[25566] = i[25566];
  assign o[25565] = i[25565];
  assign o[25564] = i[25564];
  assign o[25563] = i[25563];
  assign o[25562] = i[25562];
  assign o[25561] = i[25561];
  assign o[25560] = i[25560];
  assign o[25559] = i[25559];
  assign o[25558] = i[25558];
  assign o[25557] = i[25557];
  assign o[25556] = i[25556];
  assign o[25555] = i[25555];
  assign o[25554] = i[25554];
  assign o[25553] = i[25553];
  assign o[25552] = i[25552];
  assign o[25551] = i[25551];
  assign o[25550] = i[25550];
  assign o[25549] = i[25549];
  assign o[25548] = i[25548];
  assign o[25547] = i[25547];
  assign o[25546] = i[25546];
  assign o[25545] = i[25545];
  assign o[25544] = i[25544];
  assign o[25543] = i[25543];
  assign o[25542] = i[25542];
  assign o[25541] = i[25541];
  assign o[25540] = i[25540];
  assign o[25539] = i[25539];
  assign o[25538] = i[25538];
  assign o[25537] = i[25537];
  assign o[25536] = i[25536];
  assign o[25535] = i[25535];
  assign o[25534] = i[25534];
  assign o[25533] = i[25533];
  assign o[25532] = i[25532];
  assign o[25531] = i[25531];
  assign o[25530] = i[25530];
  assign o[25529] = i[25529];
  assign o[25528] = i[25528];
  assign o[25527] = i[25527];
  assign o[25526] = i[25526];
  assign o[25525] = i[25525];
  assign o[25524] = i[25524];
  assign o[25523] = i[25523];
  assign o[25522] = i[25522];
  assign o[25521] = i[25521];
  assign o[25520] = i[25520];
  assign o[25519] = i[25519];
  assign o[25518] = i[25518];
  assign o[25517] = i[25517];
  assign o[25516] = i[25516];
  assign o[25515] = i[25515];
  assign o[25514] = i[25514];
  assign o[25513] = i[25513];
  assign o[25512] = i[25512];
  assign o[25511] = i[25511];
  assign o[25510] = i[25510];
  assign o[25509] = i[25509];
  assign o[25508] = i[25508];
  assign o[25507] = i[25507];
  assign o[25506] = i[25506];
  assign o[25505] = i[25505];
  assign o[25504] = i[25504];
  assign o[25503] = i[25503];
  assign o[25502] = i[25502];
  assign o[25501] = i[25501];
  assign o[25500] = i[25500];
  assign o[25499] = i[25499];
  assign o[25498] = i[25498];
  assign o[25497] = i[25497];
  assign o[25496] = i[25496];
  assign o[25495] = i[25495];
  assign o[25494] = i[25494];
  assign o[25493] = i[25493];
  assign o[25492] = i[25492];
  assign o[25491] = i[25491];
  assign o[25490] = i[25490];
  assign o[25489] = i[25489];
  assign o[25488] = i[25488];
  assign o[25487] = i[25487];
  assign o[25486] = i[25486];
  assign o[25485] = i[25485];
  assign o[25484] = i[25484];
  assign o[25483] = i[25483];
  assign o[25482] = i[25482];
  assign o[25481] = i[25481];
  assign o[25480] = i[25480];
  assign o[25479] = i[25479];
  assign o[25478] = i[25478];
  assign o[25477] = i[25477];
  assign o[25476] = i[25476];
  assign o[25475] = i[25475];
  assign o[25474] = i[25474];
  assign o[25473] = i[25473];
  assign o[25472] = i[25472];
  assign o[25471] = i[25471];
  assign o[25470] = i[25470];
  assign o[25469] = i[25469];
  assign o[25468] = i[25468];
  assign o[25467] = i[25467];
  assign o[25466] = i[25466];
  assign o[25465] = i[25465];
  assign o[25464] = i[25464];
  assign o[25463] = i[25463];
  assign o[25462] = i[25462];
  assign o[25461] = i[25461];
  assign o[25460] = i[25460];
  assign o[25459] = i[25459];
  assign o[25458] = i[25458];
  assign o[25457] = i[25457];
  assign o[25456] = i[25456];
  assign o[25455] = i[25455];
  assign o[25454] = i[25454];
  assign o[25453] = i[25453];
  assign o[25452] = i[25452];
  assign o[25451] = i[25451];
  assign o[25450] = i[25450];
  assign o[25449] = i[25449];
  assign o[25448] = i[25448];
  assign o[25447] = i[25447];
  assign o[25446] = i[25446];
  assign o[25445] = i[25445];
  assign o[25444] = i[25444];
  assign o[25443] = i[25443];
  assign o[25442] = i[25442];
  assign o[25441] = i[25441];
  assign o[25440] = i[25440];
  assign o[25439] = i[25439];
  assign o[25438] = i[25438];
  assign o[25437] = i[25437];
  assign o[25436] = i[25436];
  assign o[25435] = i[25435];
  assign o[25434] = i[25434];
  assign o[25433] = i[25433];
  assign o[25432] = i[25432];
  assign o[25431] = i[25431];
  assign o[25430] = i[25430];
  assign o[25429] = i[25429];
  assign o[25428] = i[25428];
  assign o[25427] = i[25427];
  assign o[25426] = i[25426];
  assign o[25425] = i[25425];
  assign o[25424] = i[25424];
  assign o[25423] = i[25423];
  assign o[25422] = i[25422];
  assign o[25421] = i[25421];
  assign o[25420] = i[25420];
  assign o[25419] = i[25419];
  assign o[25418] = i[25418];
  assign o[25417] = i[25417];
  assign o[25416] = i[25416];
  assign o[25415] = i[25415];
  assign o[25414] = i[25414];
  assign o[25413] = i[25413];
  assign o[25412] = i[25412];
  assign o[25411] = i[25411];
  assign o[25410] = i[25410];
  assign o[25409] = i[25409];
  assign o[25408] = i[25408];
  assign o[25407] = i[25407];
  assign o[25406] = i[25406];
  assign o[25405] = i[25405];
  assign o[25404] = i[25404];
  assign o[25403] = i[25403];
  assign o[25402] = i[25402];
  assign o[25401] = i[25401];
  assign o[25400] = i[25400];
  assign o[25399] = i[25399];
  assign o[25398] = i[25398];
  assign o[25397] = i[25397];
  assign o[25396] = i[25396];
  assign o[25395] = i[25395];
  assign o[25394] = i[25394];
  assign o[25393] = i[25393];
  assign o[25392] = i[25392];
  assign o[25391] = i[25391];
  assign o[25390] = i[25390];
  assign o[25389] = i[25389];
  assign o[25388] = i[25388];
  assign o[25387] = i[25387];
  assign o[25386] = i[25386];
  assign o[25385] = i[25385];
  assign o[25384] = i[25384];
  assign o[25383] = i[25383];
  assign o[25382] = i[25382];
  assign o[25381] = i[25381];
  assign o[25380] = i[25380];
  assign o[25379] = i[25379];
  assign o[25378] = i[25378];
  assign o[25377] = i[25377];
  assign o[25376] = i[25376];
  assign o[25375] = i[25375];
  assign o[25374] = i[25374];
  assign o[25373] = i[25373];
  assign o[25372] = i[25372];
  assign o[25371] = i[25371];
  assign o[25370] = i[25370];
  assign o[25369] = i[25369];
  assign o[25368] = i[25368];
  assign o[25367] = i[25367];
  assign o[25366] = i[25366];
  assign o[25365] = i[25365];
  assign o[25364] = i[25364];
  assign o[25363] = i[25363];
  assign o[25362] = i[25362];
  assign o[25361] = i[25361];
  assign o[25360] = i[25360];
  assign o[25359] = i[25359];
  assign o[25358] = i[25358];
  assign o[25357] = i[25357];
  assign o[25356] = i[25356];
  assign o[25355] = i[25355];
  assign o[25354] = i[25354];
  assign o[25353] = i[25353];
  assign o[25352] = i[25352];
  assign o[25351] = i[25351];
  assign o[25350] = i[25350];
  assign o[25349] = i[25349];
  assign o[25348] = i[25348];
  assign o[25347] = i[25347];
  assign o[25346] = i[25346];
  assign o[25345] = i[25345];
  assign o[25344] = i[25344];
  assign o[25343] = i[25343];
  assign o[25342] = i[25342];
  assign o[25341] = i[25341];
  assign o[25340] = i[25340];
  assign o[25339] = i[25339];
  assign o[25338] = i[25338];
  assign o[25337] = i[25337];
  assign o[25336] = i[25336];
  assign o[25335] = i[25335];
  assign o[25334] = i[25334];
  assign o[25333] = i[25333];
  assign o[25332] = i[25332];
  assign o[25331] = i[25331];
  assign o[25330] = i[25330];
  assign o[25329] = i[25329];
  assign o[25328] = i[25328];
  assign o[25327] = i[25327];
  assign o[25326] = i[25326];
  assign o[25325] = i[25325];
  assign o[25324] = i[25324];
  assign o[25323] = i[25323];
  assign o[25322] = i[25322];
  assign o[25321] = i[25321];
  assign o[25320] = i[25320];
  assign o[25319] = i[25319];
  assign o[25318] = i[25318];
  assign o[25317] = i[25317];
  assign o[25316] = i[25316];
  assign o[25315] = i[25315];
  assign o[25314] = i[25314];
  assign o[25313] = i[25313];
  assign o[25312] = i[25312];
  assign o[25311] = i[25311];
  assign o[25310] = i[25310];
  assign o[25309] = i[25309];
  assign o[25308] = i[25308];
  assign o[25307] = i[25307];
  assign o[25306] = i[25306];
  assign o[25305] = i[25305];
  assign o[25304] = i[25304];
  assign o[25303] = i[25303];
  assign o[25302] = i[25302];
  assign o[25301] = i[25301];
  assign o[25300] = i[25300];
  assign o[25299] = i[25299];
  assign o[25298] = i[25298];
  assign o[25297] = i[25297];
  assign o[25296] = i[25296];
  assign o[25295] = i[25295];
  assign o[25294] = i[25294];
  assign o[25293] = i[25293];
  assign o[25292] = i[25292];
  assign o[25291] = i[25291];
  assign o[25290] = i[25290];
  assign o[25289] = i[25289];
  assign o[25288] = i[25288];
  assign o[25287] = i[25287];
  assign o[25286] = i[25286];
  assign o[25285] = i[25285];
  assign o[25284] = i[25284];
  assign o[25283] = i[25283];
  assign o[25282] = i[25282];
  assign o[25281] = i[25281];
  assign o[25280] = i[25280];
  assign o[25279] = i[25279];
  assign o[25278] = i[25278];
  assign o[25277] = i[25277];
  assign o[25276] = i[25276];
  assign o[25275] = i[25275];
  assign o[25274] = i[25274];
  assign o[25273] = i[25273];
  assign o[25272] = i[25272];
  assign o[25271] = i[25271];
  assign o[25270] = i[25270];
  assign o[25269] = i[25269];
  assign o[25268] = i[25268];
  assign o[25267] = i[25267];
  assign o[25266] = i[25266];
  assign o[25265] = i[25265];
  assign o[25264] = i[25264];
  assign o[25263] = i[25263];
  assign o[25262] = i[25262];
  assign o[25261] = i[25261];
  assign o[25260] = i[25260];
  assign o[25259] = i[25259];
  assign o[25258] = i[25258];
  assign o[25257] = i[25257];
  assign o[25256] = i[25256];
  assign o[25255] = i[25255];
  assign o[25254] = i[25254];
  assign o[25253] = i[25253];
  assign o[25252] = i[25252];
  assign o[25251] = i[25251];
  assign o[25250] = i[25250];
  assign o[25249] = i[25249];
  assign o[25248] = i[25248];
  assign o[25247] = i[25247];
  assign o[25246] = i[25246];
  assign o[25245] = i[25245];
  assign o[25244] = i[25244];
  assign o[25243] = i[25243];
  assign o[25242] = i[25242];
  assign o[25241] = i[25241];
  assign o[25240] = i[25240];
  assign o[25239] = i[25239];
  assign o[25238] = i[25238];
  assign o[25237] = i[25237];
  assign o[25236] = i[25236];
  assign o[25235] = i[25235];
  assign o[25234] = i[25234];
  assign o[25233] = i[25233];
  assign o[25232] = i[25232];
  assign o[25231] = i[25231];
  assign o[25230] = i[25230];
  assign o[25229] = i[25229];
  assign o[25228] = i[25228];
  assign o[25227] = i[25227];
  assign o[25226] = i[25226];
  assign o[25225] = i[25225];
  assign o[25224] = i[25224];
  assign o[25223] = i[25223];
  assign o[25222] = i[25222];
  assign o[25221] = i[25221];
  assign o[25220] = i[25220];
  assign o[25219] = i[25219];
  assign o[25218] = i[25218];
  assign o[25217] = i[25217];
  assign o[25216] = i[25216];
  assign o[25215] = i[25215];
  assign o[25214] = i[25214];
  assign o[25213] = i[25213];
  assign o[25212] = i[25212];
  assign o[25211] = i[25211];
  assign o[25210] = i[25210];
  assign o[25209] = i[25209];
  assign o[25208] = i[25208];
  assign o[25207] = i[25207];
  assign o[25206] = i[25206];
  assign o[25205] = i[25205];
  assign o[25204] = i[25204];
  assign o[25203] = i[25203];
  assign o[25202] = i[25202];
  assign o[25201] = i[25201];
  assign o[25200] = i[25200];
  assign o[25199] = i[25199];
  assign o[25198] = i[25198];
  assign o[25197] = i[25197];
  assign o[25196] = i[25196];
  assign o[25195] = i[25195];
  assign o[25194] = i[25194];
  assign o[25193] = i[25193];
  assign o[25192] = i[25192];
  assign o[25191] = i[25191];
  assign o[25190] = i[25190];
  assign o[25189] = i[25189];
  assign o[25188] = i[25188];
  assign o[25187] = i[25187];
  assign o[25186] = i[25186];
  assign o[25185] = i[25185];
  assign o[25184] = i[25184];
  assign o[25183] = i[25183];
  assign o[25182] = i[25182];
  assign o[25181] = i[25181];
  assign o[25180] = i[25180];
  assign o[25179] = i[25179];
  assign o[25178] = i[25178];
  assign o[25177] = i[25177];
  assign o[25176] = i[25176];
  assign o[25175] = i[25175];
  assign o[25174] = i[25174];
  assign o[25173] = i[25173];
  assign o[25172] = i[25172];
  assign o[25171] = i[25171];
  assign o[25170] = i[25170];
  assign o[25169] = i[25169];
  assign o[25168] = i[25168];
  assign o[25167] = i[25167];
  assign o[25166] = i[25166];
  assign o[25165] = i[25165];
  assign o[25164] = i[25164];
  assign o[25163] = i[25163];
  assign o[25162] = i[25162];
  assign o[25161] = i[25161];
  assign o[25160] = i[25160];
  assign o[25159] = i[25159];
  assign o[25158] = i[25158];
  assign o[25157] = i[25157];
  assign o[25156] = i[25156];
  assign o[25155] = i[25155];
  assign o[25154] = i[25154];
  assign o[25153] = i[25153];
  assign o[25152] = i[25152];
  assign o[25151] = i[25151];
  assign o[25150] = i[25150];
  assign o[25149] = i[25149];
  assign o[25148] = i[25148];
  assign o[25147] = i[25147];
  assign o[25146] = i[25146];
  assign o[25145] = i[25145];
  assign o[25144] = i[25144];
  assign o[25143] = i[25143];
  assign o[25142] = i[25142];
  assign o[25141] = i[25141];
  assign o[25140] = i[25140];
  assign o[25139] = i[25139];
  assign o[25138] = i[25138];
  assign o[25137] = i[25137];
  assign o[25136] = i[25136];
  assign o[25135] = i[25135];
  assign o[25134] = i[25134];
  assign o[25133] = i[25133];
  assign o[25132] = i[25132];
  assign o[25131] = i[25131];
  assign o[25130] = i[25130];
  assign o[25129] = i[25129];
  assign o[25128] = i[25128];
  assign o[25127] = i[25127];
  assign o[25126] = i[25126];
  assign o[25125] = i[25125];
  assign o[25124] = i[25124];
  assign o[25123] = i[25123];
  assign o[25122] = i[25122];
  assign o[25121] = i[25121];
  assign o[25120] = i[25120];
  assign o[25119] = i[25119];
  assign o[25118] = i[25118];
  assign o[25117] = i[25117];
  assign o[25116] = i[25116];
  assign o[25115] = i[25115];
  assign o[25114] = i[25114];
  assign o[25113] = i[25113];
  assign o[25112] = i[25112];
  assign o[25111] = i[25111];
  assign o[25110] = i[25110];
  assign o[25109] = i[25109];
  assign o[25108] = i[25108];
  assign o[25107] = i[25107];
  assign o[25106] = i[25106];
  assign o[25105] = i[25105];
  assign o[25104] = i[25104];
  assign o[25103] = i[25103];
  assign o[25102] = i[25102];
  assign o[25101] = i[25101];
  assign o[25100] = i[25100];
  assign o[25099] = i[25099];
  assign o[25098] = i[25098];
  assign o[25097] = i[25097];
  assign o[25096] = i[25096];
  assign o[25095] = i[25095];
  assign o[25094] = i[25094];
  assign o[25093] = i[25093];
  assign o[25092] = i[25092];
  assign o[25091] = i[25091];
  assign o[25090] = i[25090];
  assign o[25089] = i[25089];
  assign o[25088] = i[25088];
  assign o[25087] = i[25087];
  assign o[25086] = i[25086];
  assign o[25085] = i[25085];
  assign o[25084] = i[25084];
  assign o[25083] = i[25083];
  assign o[25082] = i[25082];
  assign o[25081] = i[25081];
  assign o[25080] = i[25080];
  assign o[25079] = i[25079];
  assign o[25078] = i[25078];
  assign o[25077] = i[25077];
  assign o[25076] = i[25076];
  assign o[25075] = i[25075];
  assign o[25074] = i[25074];
  assign o[25073] = i[25073];
  assign o[25072] = i[25072];
  assign o[25071] = i[25071];
  assign o[25070] = i[25070];
  assign o[25069] = i[25069];
  assign o[25068] = i[25068];
  assign o[25067] = i[25067];
  assign o[25066] = i[25066];
  assign o[25065] = i[25065];
  assign o[25064] = i[25064];
  assign o[25063] = i[25063];
  assign o[25062] = i[25062];
  assign o[25061] = i[25061];
  assign o[25060] = i[25060];
  assign o[25059] = i[25059];
  assign o[25058] = i[25058];
  assign o[25057] = i[25057];
  assign o[25056] = i[25056];
  assign o[25055] = i[25055];
  assign o[25054] = i[25054];
  assign o[25053] = i[25053];
  assign o[25052] = i[25052];
  assign o[25051] = i[25051];
  assign o[25050] = i[25050];
  assign o[25049] = i[25049];
  assign o[25048] = i[25048];
  assign o[25047] = i[25047];
  assign o[25046] = i[25046];
  assign o[25045] = i[25045];
  assign o[25044] = i[25044];
  assign o[25043] = i[25043];
  assign o[25042] = i[25042];
  assign o[25041] = i[25041];
  assign o[25040] = i[25040];
  assign o[25039] = i[25039];
  assign o[25038] = i[25038];
  assign o[25037] = i[25037];
  assign o[25036] = i[25036];
  assign o[25035] = i[25035];
  assign o[25034] = i[25034];
  assign o[25033] = i[25033];
  assign o[25032] = i[25032];
  assign o[25031] = i[25031];
  assign o[25030] = i[25030];
  assign o[25029] = i[25029];
  assign o[25028] = i[25028];
  assign o[25027] = i[25027];
  assign o[25026] = i[25026];
  assign o[25025] = i[25025];
  assign o[25024] = i[25024];
  assign o[25023] = i[25023];
  assign o[25022] = i[25022];
  assign o[25021] = i[25021];
  assign o[25020] = i[25020];
  assign o[25019] = i[25019];
  assign o[25018] = i[25018];
  assign o[25017] = i[25017];
  assign o[25016] = i[25016];
  assign o[25015] = i[25015];
  assign o[25014] = i[25014];
  assign o[25013] = i[25013];
  assign o[25012] = i[25012];
  assign o[25011] = i[25011];
  assign o[25010] = i[25010];
  assign o[25009] = i[25009];
  assign o[25008] = i[25008];
  assign o[25007] = i[25007];
  assign o[25006] = i[25006];
  assign o[25005] = i[25005];
  assign o[25004] = i[25004];
  assign o[25003] = i[25003];
  assign o[25002] = i[25002];
  assign o[25001] = i[25001];
  assign o[25000] = i[25000];
  assign o[24999] = i[24999];
  assign o[24998] = i[24998];
  assign o[24997] = i[24997];
  assign o[24996] = i[24996];
  assign o[24995] = i[24995];
  assign o[24994] = i[24994];
  assign o[24993] = i[24993];
  assign o[24992] = i[24992];
  assign o[24991] = i[24991];
  assign o[24990] = i[24990];
  assign o[24989] = i[24989];
  assign o[24988] = i[24988];
  assign o[24987] = i[24987];
  assign o[24986] = i[24986];
  assign o[24985] = i[24985];
  assign o[24984] = i[24984];
  assign o[24983] = i[24983];
  assign o[24982] = i[24982];
  assign o[24981] = i[24981];
  assign o[24980] = i[24980];
  assign o[24979] = i[24979];
  assign o[24978] = i[24978];
  assign o[24977] = i[24977];
  assign o[24976] = i[24976];
  assign o[24975] = i[24975];
  assign o[24974] = i[24974];
  assign o[24973] = i[24973];
  assign o[24972] = i[24972];
  assign o[24971] = i[24971];
  assign o[24970] = i[24970];
  assign o[24969] = i[24969];
  assign o[24968] = i[24968];
  assign o[24967] = i[24967];
  assign o[24966] = i[24966];
  assign o[24965] = i[24965];
  assign o[24964] = i[24964];
  assign o[24963] = i[24963];
  assign o[24962] = i[24962];
  assign o[24961] = i[24961];
  assign o[24960] = i[24960];
  assign o[24959] = i[24959];
  assign o[24958] = i[24958];
  assign o[24957] = i[24957];
  assign o[24956] = i[24956];
  assign o[24955] = i[24955];
  assign o[24954] = i[24954];
  assign o[24953] = i[24953];
  assign o[24952] = i[24952];
  assign o[24951] = i[24951];
  assign o[24950] = i[24950];
  assign o[24949] = i[24949];
  assign o[24948] = i[24948];
  assign o[24947] = i[24947];
  assign o[24946] = i[24946];
  assign o[24945] = i[24945];
  assign o[24944] = i[24944];
  assign o[24943] = i[24943];
  assign o[24942] = i[24942];
  assign o[24941] = i[24941];
  assign o[24940] = i[24940];
  assign o[24939] = i[24939];
  assign o[24938] = i[24938];
  assign o[24937] = i[24937];
  assign o[24936] = i[24936];
  assign o[24935] = i[24935];
  assign o[24934] = i[24934];
  assign o[24933] = i[24933];
  assign o[24932] = i[24932];
  assign o[24931] = i[24931];
  assign o[24930] = i[24930];
  assign o[24929] = i[24929];
  assign o[24928] = i[24928];
  assign o[24927] = i[24927];
  assign o[24926] = i[24926];
  assign o[24925] = i[24925];
  assign o[24924] = i[24924];
  assign o[24923] = i[24923];
  assign o[24922] = i[24922];
  assign o[24921] = i[24921];
  assign o[24920] = i[24920];
  assign o[24919] = i[24919];
  assign o[24918] = i[24918];
  assign o[24917] = i[24917];
  assign o[24916] = i[24916];
  assign o[24915] = i[24915];
  assign o[24914] = i[24914];
  assign o[24913] = i[24913];
  assign o[24912] = i[24912];
  assign o[24911] = i[24911];
  assign o[24910] = i[24910];
  assign o[24909] = i[24909];
  assign o[24908] = i[24908];
  assign o[24907] = i[24907];
  assign o[24906] = i[24906];
  assign o[24905] = i[24905];
  assign o[24904] = i[24904];
  assign o[24903] = i[24903];
  assign o[24902] = i[24902];
  assign o[24901] = i[24901];
  assign o[24900] = i[24900];
  assign o[24899] = i[24899];
  assign o[24898] = i[24898];
  assign o[24897] = i[24897];
  assign o[24896] = i[24896];
  assign o[24895] = i[24895];
  assign o[24894] = i[24894];
  assign o[24893] = i[24893];
  assign o[24892] = i[24892];
  assign o[24891] = i[24891];
  assign o[24890] = i[24890];
  assign o[24889] = i[24889];
  assign o[24888] = i[24888];
  assign o[24887] = i[24887];
  assign o[24886] = i[24886];
  assign o[24885] = i[24885];
  assign o[24884] = i[24884];
  assign o[24883] = i[24883];
  assign o[24882] = i[24882];
  assign o[24881] = i[24881];
  assign o[24880] = i[24880];
  assign o[24879] = i[24879];
  assign o[24878] = i[24878];
  assign o[24877] = i[24877];
  assign o[24876] = i[24876];
  assign o[24875] = i[24875];
  assign o[24874] = i[24874];
  assign o[24873] = i[24873];
  assign o[24872] = i[24872];
  assign o[24871] = i[24871];
  assign o[24870] = i[24870];
  assign o[24869] = i[24869];
  assign o[24868] = i[24868];
  assign o[24867] = i[24867];
  assign o[24866] = i[24866];
  assign o[24865] = i[24865];
  assign o[24864] = i[24864];
  assign o[24863] = i[24863];
  assign o[24862] = i[24862];
  assign o[24861] = i[24861];
  assign o[24860] = i[24860];
  assign o[24859] = i[24859];
  assign o[24858] = i[24858];
  assign o[24857] = i[24857];
  assign o[24856] = i[24856];
  assign o[24855] = i[24855];
  assign o[24854] = i[24854];
  assign o[24853] = i[24853];
  assign o[24852] = i[24852];
  assign o[24851] = i[24851];
  assign o[24850] = i[24850];
  assign o[24849] = i[24849];
  assign o[24848] = i[24848];
  assign o[24847] = i[24847];
  assign o[24846] = i[24846];
  assign o[24845] = i[24845];
  assign o[24844] = i[24844];
  assign o[24843] = i[24843];
  assign o[24842] = i[24842];
  assign o[24841] = i[24841];
  assign o[24840] = i[24840];
  assign o[24839] = i[24839];
  assign o[24838] = i[24838];
  assign o[24837] = i[24837];
  assign o[24836] = i[24836];
  assign o[24835] = i[24835];
  assign o[24834] = i[24834];
  assign o[24833] = i[24833];
  assign o[24832] = i[24832];
  assign o[24831] = i[24831];
  assign o[24830] = i[24830];
  assign o[24829] = i[24829];
  assign o[24828] = i[24828];
  assign o[24827] = i[24827];
  assign o[24826] = i[24826];
  assign o[24825] = i[24825];
  assign o[24824] = i[24824];
  assign o[24823] = i[24823];
  assign o[24822] = i[24822];
  assign o[24821] = i[24821];
  assign o[24820] = i[24820];
  assign o[24819] = i[24819];
  assign o[24818] = i[24818];
  assign o[24817] = i[24817];
  assign o[24816] = i[24816];
  assign o[24815] = i[24815];
  assign o[24814] = i[24814];
  assign o[24813] = i[24813];
  assign o[24812] = i[24812];
  assign o[24811] = i[24811];
  assign o[24810] = i[24810];
  assign o[24809] = i[24809];
  assign o[24808] = i[24808];
  assign o[24807] = i[24807];
  assign o[24806] = i[24806];
  assign o[24805] = i[24805];
  assign o[24804] = i[24804];
  assign o[24803] = i[24803];
  assign o[24802] = i[24802];
  assign o[24801] = i[24801];
  assign o[24800] = i[24800];
  assign o[24799] = i[24799];
  assign o[24798] = i[24798];
  assign o[24797] = i[24797];
  assign o[24796] = i[24796];
  assign o[24795] = i[24795];
  assign o[24794] = i[24794];
  assign o[24793] = i[24793];
  assign o[24792] = i[24792];
  assign o[24791] = i[24791];
  assign o[24790] = i[24790];
  assign o[24789] = i[24789];
  assign o[24788] = i[24788];
  assign o[24787] = i[24787];
  assign o[24786] = i[24786];
  assign o[24785] = i[24785];
  assign o[24784] = i[24784];
  assign o[24783] = i[24783];
  assign o[24782] = i[24782];
  assign o[24781] = i[24781];
  assign o[24780] = i[24780];
  assign o[24779] = i[24779];
  assign o[24778] = i[24778];
  assign o[24777] = i[24777];
  assign o[24776] = i[24776];
  assign o[24775] = i[24775];
  assign o[24774] = i[24774];
  assign o[24773] = i[24773];
  assign o[24772] = i[24772];
  assign o[24771] = i[24771];
  assign o[24770] = i[24770];
  assign o[24769] = i[24769];
  assign o[24768] = i[24768];
  assign o[24767] = i[24767];
  assign o[24766] = i[24766];
  assign o[24765] = i[24765];
  assign o[24764] = i[24764];
  assign o[24763] = i[24763];
  assign o[24762] = i[24762];
  assign o[24761] = i[24761];
  assign o[24760] = i[24760];
  assign o[24759] = i[24759];
  assign o[24758] = i[24758];
  assign o[24757] = i[24757];
  assign o[24756] = i[24756];
  assign o[24755] = i[24755];
  assign o[24754] = i[24754];
  assign o[24753] = i[24753];
  assign o[24752] = i[24752];
  assign o[24751] = i[24751];
  assign o[24750] = i[24750];
  assign o[24749] = i[24749];
  assign o[24748] = i[24748];
  assign o[24747] = i[24747];
  assign o[24746] = i[24746];
  assign o[24745] = i[24745];
  assign o[24744] = i[24744];
  assign o[24743] = i[24743];
  assign o[24742] = i[24742];
  assign o[24741] = i[24741];
  assign o[24740] = i[24740];
  assign o[24739] = i[24739];
  assign o[24738] = i[24738];
  assign o[24737] = i[24737];
  assign o[24736] = i[24736];
  assign o[24735] = i[24735];
  assign o[24734] = i[24734];
  assign o[24733] = i[24733];
  assign o[24732] = i[24732];
  assign o[24731] = i[24731];
  assign o[24730] = i[24730];
  assign o[24729] = i[24729];
  assign o[24728] = i[24728];
  assign o[24727] = i[24727];
  assign o[24726] = i[24726];
  assign o[24725] = i[24725];
  assign o[24724] = i[24724];
  assign o[24723] = i[24723];
  assign o[24722] = i[24722];
  assign o[24721] = i[24721];
  assign o[24720] = i[24720];
  assign o[24719] = i[24719];
  assign o[24718] = i[24718];
  assign o[24717] = i[24717];
  assign o[24716] = i[24716];
  assign o[24715] = i[24715];
  assign o[24714] = i[24714];
  assign o[24713] = i[24713];
  assign o[24712] = i[24712];
  assign o[24711] = i[24711];
  assign o[24710] = i[24710];
  assign o[24709] = i[24709];
  assign o[24708] = i[24708];
  assign o[24707] = i[24707];
  assign o[24706] = i[24706];
  assign o[24705] = i[24705];
  assign o[24704] = i[24704];
  assign o[24703] = i[24703];
  assign o[24702] = i[24702];
  assign o[24701] = i[24701];
  assign o[24700] = i[24700];
  assign o[24699] = i[24699];
  assign o[24698] = i[24698];
  assign o[24697] = i[24697];
  assign o[24696] = i[24696];
  assign o[24695] = i[24695];
  assign o[24694] = i[24694];
  assign o[24693] = i[24693];
  assign o[24692] = i[24692];
  assign o[24691] = i[24691];
  assign o[24690] = i[24690];
  assign o[24689] = i[24689];
  assign o[24688] = i[24688];
  assign o[24687] = i[24687];
  assign o[24686] = i[24686];
  assign o[24685] = i[24685];
  assign o[24684] = i[24684];
  assign o[24683] = i[24683];
  assign o[24682] = i[24682];
  assign o[24681] = i[24681];
  assign o[24680] = i[24680];
  assign o[24679] = i[24679];
  assign o[24678] = i[24678];
  assign o[24677] = i[24677];
  assign o[24676] = i[24676];
  assign o[24675] = i[24675];
  assign o[24674] = i[24674];
  assign o[24673] = i[24673];
  assign o[24672] = i[24672];
  assign o[24671] = i[24671];
  assign o[24670] = i[24670];
  assign o[24669] = i[24669];
  assign o[24668] = i[24668];
  assign o[24667] = i[24667];
  assign o[24666] = i[24666];
  assign o[24665] = i[24665];
  assign o[24664] = i[24664];
  assign o[24663] = i[24663];
  assign o[24662] = i[24662];
  assign o[24661] = i[24661];
  assign o[24660] = i[24660];
  assign o[24659] = i[24659];
  assign o[24658] = i[24658];
  assign o[24657] = i[24657];
  assign o[24656] = i[24656];
  assign o[24655] = i[24655];
  assign o[24654] = i[24654];
  assign o[24653] = i[24653];
  assign o[24652] = i[24652];
  assign o[24651] = i[24651];
  assign o[24650] = i[24650];
  assign o[24649] = i[24649];
  assign o[24648] = i[24648];
  assign o[24647] = i[24647];
  assign o[24646] = i[24646];
  assign o[24645] = i[24645];
  assign o[24644] = i[24644];
  assign o[24643] = i[24643];
  assign o[24642] = i[24642];
  assign o[24641] = i[24641];
  assign o[24640] = i[24640];
  assign o[24639] = i[24639];
  assign o[24638] = i[24638];
  assign o[24637] = i[24637];
  assign o[24636] = i[24636];
  assign o[24635] = i[24635];
  assign o[24634] = i[24634];
  assign o[24633] = i[24633];
  assign o[24632] = i[24632];
  assign o[24631] = i[24631];
  assign o[24630] = i[24630];
  assign o[24629] = i[24629];
  assign o[24628] = i[24628];
  assign o[24627] = i[24627];
  assign o[24626] = i[24626];
  assign o[24625] = i[24625];
  assign o[24624] = i[24624];
  assign o[24623] = i[24623];
  assign o[24622] = i[24622];
  assign o[24621] = i[24621];
  assign o[24620] = i[24620];
  assign o[24619] = i[24619];
  assign o[24618] = i[24618];
  assign o[24617] = i[24617];
  assign o[24616] = i[24616];
  assign o[24615] = i[24615];
  assign o[24614] = i[24614];
  assign o[24613] = i[24613];
  assign o[24612] = i[24612];
  assign o[24611] = i[24611];
  assign o[24610] = i[24610];
  assign o[24609] = i[24609];
  assign o[24608] = i[24608];
  assign o[24607] = i[24607];
  assign o[24606] = i[24606];
  assign o[24605] = i[24605];
  assign o[24604] = i[24604];
  assign o[24603] = i[24603];
  assign o[24602] = i[24602];
  assign o[24601] = i[24601];
  assign o[24600] = i[24600];
  assign o[24599] = i[24599];
  assign o[24598] = i[24598];
  assign o[24597] = i[24597];
  assign o[24596] = i[24596];
  assign o[24595] = i[24595];
  assign o[24594] = i[24594];
  assign o[24593] = i[24593];
  assign o[24592] = i[24592];
  assign o[24591] = i[24591];
  assign o[24590] = i[24590];
  assign o[24589] = i[24589];
  assign o[24588] = i[24588];
  assign o[24587] = i[24587];
  assign o[24586] = i[24586];
  assign o[24585] = i[24585];
  assign o[24584] = i[24584];
  assign o[24583] = i[24583];
  assign o[24582] = i[24582];
  assign o[24581] = i[24581];
  assign o[24580] = i[24580];
  assign o[24579] = i[24579];
  assign o[24578] = i[24578];
  assign o[24577] = i[24577];
  assign o[24576] = i[24576];
  assign o[24575] = i[24575];
  assign o[24574] = i[24574];
  assign o[24573] = i[24573];
  assign o[24572] = i[24572];
  assign o[24571] = i[24571];
  assign o[24570] = i[24570];
  assign o[24569] = i[24569];
  assign o[24568] = i[24568];
  assign o[24567] = i[24567];
  assign o[24566] = i[24566];
  assign o[24565] = i[24565];
  assign o[24564] = i[24564];
  assign o[24563] = i[24563];
  assign o[24562] = i[24562];
  assign o[24561] = i[24561];
  assign o[24560] = i[24560];
  assign o[24559] = i[24559];
  assign o[24558] = i[24558];
  assign o[24557] = i[24557];
  assign o[24556] = i[24556];
  assign o[24555] = i[24555];
  assign o[24554] = i[24554];
  assign o[24553] = i[24553];
  assign o[24552] = i[24552];
  assign o[24551] = i[24551];
  assign o[24550] = i[24550];
  assign o[24549] = i[24549];
  assign o[24548] = i[24548];
  assign o[24547] = i[24547];
  assign o[24546] = i[24546];
  assign o[24545] = i[24545];
  assign o[24544] = i[24544];
  assign o[24543] = i[24543];
  assign o[24542] = i[24542];
  assign o[24541] = i[24541];
  assign o[24540] = i[24540];
  assign o[24539] = i[24539];
  assign o[24538] = i[24538];
  assign o[24537] = i[24537];
  assign o[24536] = i[24536];
  assign o[24535] = i[24535];
  assign o[24534] = i[24534];
  assign o[24533] = i[24533];
  assign o[24532] = i[24532];
  assign o[24531] = i[24531];
  assign o[24530] = i[24530];
  assign o[24529] = i[24529];
  assign o[24528] = i[24528];
  assign o[24527] = i[24527];
  assign o[24526] = i[24526];
  assign o[24525] = i[24525];
  assign o[24524] = i[24524];
  assign o[24523] = i[24523];
  assign o[24522] = i[24522];
  assign o[24521] = i[24521];
  assign o[24520] = i[24520];
  assign o[24519] = i[24519];
  assign o[24518] = i[24518];
  assign o[24517] = i[24517];
  assign o[24516] = i[24516];
  assign o[24515] = i[24515];
  assign o[24514] = i[24514];
  assign o[24513] = i[24513];
  assign o[24512] = i[24512];
  assign o[24511] = i[24511];
  assign o[24510] = i[24510];
  assign o[24509] = i[24509];
  assign o[24508] = i[24508];
  assign o[24507] = i[24507];
  assign o[24506] = i[24506];
  assign o[24505] = i[24505];
  assign o[24504] = i[24504];
  assign o[24503] = i[24503];
  assign o[24502] = i[24502];
  assign o[24501] = i[24501];
  assign o[24500] = i[24500];
  assign o[24499] = i[24499];
  assign o[24498] = i[24498];
  assign o[24497] = i[24497];
  assign o[24496] = i[24496];
  assign o[24495] = i[24495];
  assign o[24494] = i[24494];
  assign o[24493] = i[24493];
  assign o[24492] = i[24492];
  assign o[24491] = i[24491];
  assign o[24490] = i[24490];
  assign o[24489] = i[24489];
  assign o[24488] = i[24488];
  assign o[24487] = i[24487];
  assign o[24486] = i[24486];
  assign o[24485] = i[24485];
  assign o[24484] = i[24484];
  assign o[24483] = i[24483];
  assign o[24482] = i[24482];
  assign o[24481] = i[24481];
  assign o[24480] = i[24480];
  assign o[24479] = i[24479];
  assign o[24478] = i[24478];
  assign o[24477] = i[24477];
  assign o[24476] = i[24476];
  assign o[24475] = i[24475];
  assign o[24474] = i[24474];
  assign o[24473] = i[24473];
  assign o[24472] = i[24472];
  assign o[24471] = i[24471];
  assign o[24470] = i[24470];
  assign o[24469] = i[24469];
  assign o[24468] = i[24468];
  assign o[24467] = i[24467];
  assign o[24466] = i[24466];
  assign o[24465] = i[24465];
  assign o[24464] = i[24464];
  assign o[24463] = i[24463];
  assign o[24462] = i[24462];
  assign o[24461] = i[24461];
  assign o[24460] = i[24460];
  assign o[24459] = i[24459];
  assign o[24458] = i[24458];
  assign o[24457] = i[24457];
  assign o[24456] = i[24456];
  assign o[24455] = i[24455];
  assign o[24454] = i[24454];
  assign o[24453] = i[24453];
  assign o[24452] = i[24452];
  assign o[24451] = i[24451];
  assign o[24450] = i[24450];
  assign o[24449] = i[24449];
  assign o[24448] = i[24448];
  assign o[24447] = i[24447];
  assign o[24446] = i[24446];
  assign o[24445] = i[24445];
  assign o[24444] = i[24444];
  assign o[24443] = i[24443];
  assign o[24442] = i[24442];
  assign o[24441] = i[24441];
  assign o[24440] = i[24440];
  assign o[24439] = i[24439];
  assign o[24438] = i[24438];
  assign o[24437] = i[24437];
  assign o[24436] = i[24436];
  assign o[24435] = i[24435];
  assign o[24434] = i[24434];
  assign o[24433] = i[24433];
  assign o[24432] = i[24432];
  assign o[24431] = i[24431];
  assign o[24430] = i[24430];
  assign o[24429] = i[24429];
  assign o[24428] = i[24428];
  assign o[24427] = i[24427];
  assign o[24426] = i[24426];
  assign o[24425] = i[24425];
  assign o[24424] = i[24424];
  assign o[24423] = i[24423];
  assign o[24422] = i[24422];
  assign o[24421] = i[24421];
  assign o[24420] = i[24420];
  assign o[24419] = i[24419];
  assign o[24418] = i[24418];
  assign o[24417] = i[24417];
  assign o[24416] = i[24416];
  assign o[24415] = i[24415];
  assign o[24414] = i[24414];
  assign o[24413] = i[24413];
  assign o[24412] = i[24412];
  assign o[24411] = i[24411];
  assign o[24410] = i[24410];
  assign o[24409] = i[24409];
  assign o[24408] = i[24408];
  assign o[24407] = i[24407];
  assign o[24406] = i[24406];
  assign o[24405] = i[24405];
  assign o[24404] = i[24404];
  assign o[24403] = i[24403];
  assign o[24402] = i[24402];
  assign o[24401] = i[24401];
  assign o[24400] = i[24400];
  assign o[24399] = i[24399];
  assign o[24398] = i[24398];
  assign o[24397] = i[24397];
  assign o[24396] = i[24396];
  assign o[24395] = i[24395];
  assign o[24394] = i[24394];
  assign o[24393] = i[24393];
  assign o[24392] = i[24392];
  assign o[24391] = i[24391];
  assign o[24390] = i[24390];
  assign o[24389] = i[24389];
  assign o[24388] = i[24388];
  assign o[24387] = i[24387];
  assign o[24386] = i[24386];
  assign o[24385] = i[24385];
  assign o[24384] = i[24384];
  assign o[24383] = i[24383];
  assign o[24382] = i[24382];
  assign o[24381] = i[24381];
  assign o[24380] = i[24380];
  assign o[24379] = i[24379];
  assign o[24378] = i[24378];
  assign o[24377] = i[24377];
  assign o[24376] = i[24376];
  assign o[24375] = i[24375];
  assign o[24374] = i[24374];
  assign o[24373] = i[24373];
  assign o[24372] = i[24372];
  assign o[24371] = i[24371];
  assign o[24370] = i[24370];
  assign o[24369] = i[24369];
  assign o[24368] = i[24368];
  assign o[24367] = i[24367];
  assign o[24366] = i[24366];
  assign o[24365] = i[24365];
  assign o[24364] = i[24364];
  assign o[24363] = i[24363];
  assign o[24362] = i[24362];
  assign o[24361] = i[24361];
  assign o[24360] = i[24360];
  assign o[24359] = i[24359];
  assign o[24358] = i[24358];
  assign o[24357] = i[24357];
  assign o[24356] = i[24356];
  assign o[24355] = i[24355];
  assign o[24354] = i[24354];
  assign o[24353] = i[24353];
  assign o[24352] = i[24352];
  assign o[24351] = i[24351];
  assign o[24350] = i[24350];
  assign o[24349] = i[24349];
  assign o[24348] = i[24348];
  assign o[24347] = i[24347];
  assign o[24346] = i[24346];
  assign o[24345] = i[24345];
  assign o[24344] = i[24344];
  assign o[24343] = i[24343];
  assign o[24342] = i[24342];
  assign o[24341] = i[24341];
  assign o[24340] = i[24340];
  assign o[24339] = i[24339];
  assign o[24338] = i[24338];
  assign o[24337] = i[24337];
  assign o[24336] = i[24336];
  assign o[24335] = i[24335];
  assign o[24334] = i[24334];
  assign o[24333] = i[24333];
  assign o[24332] = i[24332];
  assign o[24331] = i[24331];
  assign o[24330] = i[24330];
  assign o[24329] = i[24329];
  assign o[24328] = i[24328];
  assign o[24327] = i[24327];
  assign o[24326] = i[24326];
  assign o[24325] = i[24325];
  assign o[24324] = i[24324];
  assign o[24323] = i[24323];
  assign o[24322] = i[24322];
  assign o[24321] = i[24321];
  assign o[24320] = i[24320];
  assign o[24319] = i[24319];
  assign o[24318] = i[24318];
  assign o[24317] = i[24317];
  assign o[24316] = i[24316];
  assign o[24315] = i[24315];
  assign o[24314] = i[24314];
  assign o[24313] = i[24313];
  assign o[24312] = i[24312];
  assign o[24311] = i[24311];
  assign o[24310] = i[24310];
  assign o[24309] = i[24309];
  assign o[24308] = i[24308];
  assign o[24307] = i[24307];
  assign o[24306] = i[24306];
  assign o[24305] = i[24305];
  assign o[24304] = i[24304];
  assign o[24303] = i[24303];
  assign o[24302] = i[24302];
  assign o[24301] = i[24301];
  assign o[24300] = i[24300];
  assign o[24299] = i[24299];
  assign o[24298] = i[24298];
  assign o[24297] = i[24297];
  assign o[24296] = i[24296];
  assign o[24295] = i[24295];
  assign o[24294] = i[24294];
  assign o[24293] = i[24293];
  assign o[24292] = i[24292];
  assign o[24291] = i[24291];
  assign o[24290] = i[24290];
  assign o[24289] = i[24289];
  assign o[24288] = i[24288];
  assign o[24287] = i[24287];
  assign o[24286] = i[24286];
  assign o[24285] = i[24285];
  assign o[24284] = i[24284];
  assign o[24283] = i[24283];
  assign o[24282] = i[24282];
  assign o[24281] = i[24281];
  assign o[24280] = i[24280];
  assign o[24279] = i[24279];
  assign o[24278] = i[24278];
  assign o[24277] = i[24277];
  assign o[24276] = i[24276];
  assign o[24275] = i[24275];
  assign o[24274] = i[24274];
  assign o[24273] = i[24273];
  assign o[24272] = i[24272];
  assign o[24271] = i[24271];
  assign o[24270] = i[24270];
  assign o[24269] = i[24269];
  assign o[24268] = i[24268];
  assign o[24267] = i[24267];
  assign o[24266] = i[24266];
  assign o[24265] = i[24265];
  assign o[24264] = i[24264];
  assign o[24263] = i[24263];
  assign o[24262] = i[24262];
  assign o[24261] = i[24261];
  assign o[24260] = i[24260];
  assign o[24259] = i[24259];
  assign o[24258] = i[24258];
  assign o[24257] = i[24257];
  assign o[24256] = i[24256];
  assign o[24255] = i[24255];
  assign o[24254] = i[24254];
  assign o[24253] = i[24253];
  assign o[24252] = i[24252];
  assign o[24251] = i[24251];
  assign o[24250] = i[24250];
  assign o[24249] = i[24249];
  assign o[24248] = i[24248];
  assign o[24247] = i[24247];
  assign o[24246] = i[24246];
  assign o[24245] = i[24245];
  assign o[24244] = i[24244];
  assign o[24243] = i[24243];
  assign o[24242] = i[24242];
  assign o[24241] = i[24241];
  assign o[24240] = i[24240];
  assign o[24239] = i[24239];
  assign o[24238] = i[24238];
  assign o[24237] = i[24237];
  assign o[24236] = i[24236];
  assign o[24235] = i[24235];
  assign o[24234] = i[24234];
  assign o[24233] = i[24233];
  assign o[24232] = i[24232];
  assign o[24231] = i[24231];
  assign o[24230] = i[24230];
  assign o[24229] = i[24229];
  assign o[24228] = i[24228];
  assign o[24227] = i[24227];
  assign o[24226] = i[24226];
  assign o[24225] = i[24225];
  assign o[24224] = i[24224];
  assign o[24223] = i[24223];
  assign o[24222] = i[24222];
  assign o[24221] = i[24221];
  assign o[24220] = i[24220];
  assign o[24219] = i[24219];
  assign o[24218] = i[24218];
  assign o[24217] = i[24217];
  assign o[24216] = i[24216];
  assign o[24215] = i[24215];
  assign o[24214] = i[24214];
  assign o[24213] = i[24213];
  assign o[24212] = i[24212];
  assign o[24211] = i[24211];
  assign o[24210] = i[24210];
  assign o[24209] = i[24209];
  assign o[24208] = i[24208];
  assign o[24207] = i[24207];
  assign o[24206] = i[24206];
  assign o[24205] = i[24205];
  assign o[24204] = i[24204];
  assign o[24203] = i[24203];
  assign o[24202] = i[24202];
  assign o[24201] = i[24201];
  assign o[24200] = i[24200];
  assign o[24199] = i[24199];
  assign o[24198] = i[24198];
  assign o[24197] = i[24197];
  assign o[24196] = i[24196];
  assign o[24195] = i[24195];
  assign o[24194] = i[24194];
  assign o[24193] = i[24193];
  assign o[24192] = i[24192];
  assign o[24191] = i[24191];
  assign o[24190] = i[24190];
  assign o[24189] = i[24189];
  assign o[24188] = i[24188];
  assign o[24187] = i[24187];
  assign o[24186] = i[24186];
  assign o[24185] = i[24185];
  assign o[24184] = i[24184];
  assign o[24183] = i[24183];
  assign o[24182] = i[24182];
  assign o[24181] = i[24181];
  assign o[24180] = i[24180];
  assign o[24179] = i[24179];
  assign o[24178] = i[24178];
  assign o[24177] = i[24177];
  assign o[24176] = i[24176];
  assign o[24175] = i[24175];
  assign o[24174] = i[24174];
  assign o[24173] = i[24173];
  assign o[24172] = i[24172];
  assign o[24171] = i[24171];
  assign o[24170] = i[24170];
  assign o[24169] = i[24169];
  assign o[24168] = i[24168];
  assign o[24167] = i[24167];
  assign o[24166] = i[24166];
  assign o[24165] = i[24165];
  assign o[24164] = i[24164];
  assign o[24163] = i[24163];
  assign o[24162] = i[24162];
  assign o[24161] = i[24161];
  assign o[24160] = i[24160];
  assign o[24159] = i[24159];
  assign o[24158] = i[24158];
  assign o[24157] = i[24157];
  assign o[24156] = i[24156];
  assign o[24155] = i[24155];
  assign o[24154] = i[24154];
  assign o[24153] = i[24153];
  assign o[24152] = i[24152];
  assign o[24151] = i[24151];
  assign o[24150] = i[24150];
  assign o[24149] = i[24149];
  assign o[24148] = i[24148];
  assign o[24147] = i[24147];
  assign o[24146] = i[24146];
  assign o[24145] = i[24145];
  assign o[24144] = i[24144];
  assign o[24143] = i[24143];
  assign o[24142] = i[24142];
  assign o[24141] = i[24141];
  assign o[24140] = i[24140];
  assign o[24139] = i[24139];
  assign o[24138] = i[24138];
  assign o[24137] = i[24137];
  assign o[24136] = i[24136];
  assign o[24135] = i[24135];
  assign o[24134] = i[24134];
  assign o[24133] = i[24133];
  assign o[24132] = i[24132];
  assign o[24131] = i[24131];
  assign o[24130] = i[24130];
  assign o[24129] = i[24129];
  assign o[24128] = i[24128];
  assign o[24127] = i[24127];
  assign o[24126] = i[24126];
  assign o[24125] = i[24125];
  assign o[24124] = i[24124];
  assign o[24123] = i[24123];
  assign o[24122] = i[24122];
  assign o[24121] = i[24121];
  assign o[24120] = i[24120];
  assign o[24119] = i[24119];
  assign o[24118] = i[24118];
  assign o[24117] = i[24117];
  assign o[24116] = i[24116];
  assign o[24115] = i[24115];
  assign o[24114] = i[24114];
  assign o[24113] = i[24113];
  assign o[24112] = i[24112];
  assign o[24111] = i[24111];
  assign o[24110] = i[24110];
  assign o[24109] = i[24109];
  assign o[24108] = i[24108];
  assign o[24107] = i[24107];
  assign o[24106] = i[24106];
  assign o[24105] = i[24105];
  assign o[24104] = i[24104];
  assign o[24103] = i[24103];
  assign o[24102] = i[24102];
  assign o[24101] = i[24101];
  assign o[24100] = i[24100];
  assign o[24099] = i[24099];
  assign o[24098] = i[24098];
  assign o[24097] = i[24097];
  assign o[24096] = i[24096];
  assign o[24095] = i[24095];
  assign o[24094] = i[24094];
  assign o[24093] = i[24093];
  assign o[24092] = i[24092];
  assign o[24091] = i[24091];
  assign o[24090] = i[24090];
  assign o[24089] = i[24089];
  assign o[24088] = i[24088];
  assign o[24087] = i[24087];
  assign o[24086] = i[24086];
  assign o[24085] = i[24085];
  assign o[24084] = i[24084];
  assign o[24083] = i[24083];
  assign o[24082] = i[24082];
  assign o[24081] = i[24081];
  assign o[24080] = i[24080];
  assign o[24079] = i[24079];
  assign o[24078] = i[24078];
  assign o[24077] = i[24077];
  assign o[24076] = i[24076];
  assign o[24075] = i[24075];
  assign o[24074] = i[24074];
  assign o[24073] = i[24073];
  assign o[24072] = i[24072];
  assign o[24071] = i[24071];
  assign o[24070] = i[24070];
  assign o[24069] = i[24069];
  assign o[24068] = i[24068];
  assign o[24067] = i[24067];
  assign o[24066] = i[24066];
  assign o[24065] = i[24065];
  assign o[24064] = i[24064];
  assign o[24063] = i[24063];
  assign o[24062] = i[24062];
  assign o[24061] = i[24061];
  assign o[24060] = i[24060];
  assign o[24059] = i[24059];
  assign o[24058] = i[24058];
  assign o[24057] = i[24057];
  assign o[24056] = i[24056];
  assign o[24055] = i[24055];
  assign o[24054] = i[24054];
  assign o[24053] = i[24053];
  assign o[24052] = i[24052];
  assign o[24051] = i[24051];
  assign o[24050] = i[24050];
  assign o[24049] = i[24049];
  assign o[24048] = i[24048];
  assign o[24047] = i[24047];
  assign o[24046] = i[24046];
  assign o[24045] = i[24045];
  assign o[24044] = i[24044];
  assign o[24043] = i[24043];
  assign o[24042] = i[24042];
  assign o[24041] = i[24041];
  assign o[24040] = i[24040];
  assign o[24039] = i[24039];
  assign o[24038] = i[24038];
  assign o[24037] = i[24037];
  assign o[24036] = i[24036];
  assign o[24035] = i[24035];
  assign o[24034] = i[24034];
  assign o[24033] = i[24033];
  assign o[24032] = i[24032];
  assign o[24031] = i[24031];
  assign o[24030] = i[24030];
  assign o[24029] = i[24029];
  assign o[24028] = i[24028];
  assign o[24027] = i[24027];
  assign o[24026] = i[24026];
  assign o[24025] = i[24025];
  assign o[24024] = i[24024];
  assign o[24023] = i[24023];
  assign o[24022] = i[24022];
  assign o[24021] = i[24021];
  assign o[24020] = i[24020];
  assign o[24019] = i[24019];
  assign o[24018] = i[24018];
  assign o[24017] = i[24017];
  assign o[24016] = i[24016];
  assign o[24015] = i[24015];
  assign o[24014] = i[24014];
  assign o[24013] = i[24013];
  assign o[24012] = i[24012];
  assign o[24011] = i[24011];
  assign o[24010] = i[24010];
  assign o[24009] = i[24009];
  assign o[24008] = i[24008];
  assign o[24007] = i[24007];
  assign o[24006] = i[24006];
  assign o[24005] = i[24005];
  assign o[24004] = i[24004];
  assign o[24003] = i[24003];
  assign o[24002] = i[24002];
  assign o[24001] = i[24001];
  assign o[24000] = i[24000];
  assign o[23999] = i[23999];
  assign o[23998] = i[23998];
  assign o[23997] = i[23997];
  assign o[23996] = i[23996];
  assign o[23995] = i[23995];
  assign o[23994] = i[23994];
  assign o[23993] = i[23993];
  assign o[23992] = i[23992];
  assign o[23991] = i[23991];
  assign o[23990] = i[23990];
  assign o[23989] = i[23989];
  assign o[23988] = i[23988];
  assign o[23987] = i[23987];
  assign o[23986] = i[23986];
  assign o[23985] = i[23985];
  assign o[23984] = i[23984];
  assign o[23983] = i[23983];
  assign o[23982] = i[23982];
  assign o[23981] = i[23981];
  assign o[23980] = i[23980];
  assign o[23979] = i[23979];
  assign o[23978] = i[23978];
  assign o[23977] = i[23977];
  assign o[23976] = i[23976];
  assign o[23975] = i[23975];
  assign o[23974] = i[23974];
  assign o[23973] = i[23973];
  assign o[23972] = i[23972];
  assign o[23971] = i[23971];
  assign o[23970] = i[23970];
  assign o[23969] = i[23969];
  assign o[23968] = i[23968];
  assign o[23967] = i[23967];
  assign o[23966] = i[23966];
  assign o[23965] = i[23965];
  assign o[23964] = i[23964];
  assign o[23963] = i[23963];
  assign o[23962] = i[23962];
  assign o[23961] = i[23961];
  assign o[23960] = i[23960];
  assign o[23959] = i[23959];
  assign o[23958] = i[23958];
  assign o[23957] = i[23957];
  assign o[23956] = i[23956];
  assign o[23955] = i[23955];
  assign o[23954] = i[23954];
  assign o[23953] = i[23953];
  assign o[23952] = i[23952];
  assign o[23951] = i[23951];
  assign o[23950] = i[23950];
  assign o[23949] = i[23949];
  assign o[23948] = i[23948];
  assign o[23947] = i[23947];
  assign o[23946] = i[23946];
  assign o[23945] = i[23945];
  assign o[23944] = i[23944];
  assign o[23943] = i[23943];
  assign o[23942] = i[23942];
  assign o[23941] = i[23941];
  assign o[23940] = i[23940];
  assign o[23939] = i[23939];
  assign o[23938] = i[23938];
  assign o[23937] = i[23937];
  assign o[23936] = i[23936];
  assign o[23935] = i[23935];
  assign o[23934] = i[23934];
  assign o[23933] = i[23933];
  assign o[23932] = i[23932];
  assign o[23931] = i[23931];
  assign o[23930] = i[23930];
  assign o[23929] = i[23929];
  assign o[23928] = i[23928];
  assign o[23927] = i[23927];
  assign o[23926] = i[23926];
  assign o[23925] = i[23925];
  assign o[23924] = i[23924];
  assign o[23923] = i[23923];
  assign o[23922] = i[23922];
  assign o[23921] = i[23921];
  assign o[23920] = i[23920];
  assign o[23919] = i[23919];
  assign o[23918] = i[23918];
  assign o[23917] = i[23917];
  assign o[23916] = i[23916];
  assign o[23915] = i[23915];
  assign o[23914] = i[23914];
  assign o[23913] = i[23913];
  assign o[23912] = i[23912];
  assign o[23911] = i[23911];
  assign o[23910] = i[23910];
  assign o[23909] = i[23909];
  assign o[23908] = i[23908];
  assign o[23907] = i[23907];
  assign o[23906] = i[23906];
  assign o[23905] = i[23905];
  assign o[23904] = i[23904];
  assign o[23903] = i[23903];
  assign o[23902] = i[23902];
  assign o[23901] = i[23901];
  assign o[23900] = i[23900];
  assign o[23899] = i[23899];
  assign o[23898] = i[23898];
  assign o[23897] = i[23897];
  assign o[23896] = i[23896];
  assign o[23895] = i[23895];
  assign o[23894] = i[23894];
  assign o[23893] = i[23893];
  assign o[23892] = i[23892];
  assign o[23891] = i[23891];
  assign o[23890] = i[23890];
  assign o[23889] = i[23889];
  assign o[23888] = i[23888];
  assign o[23887] = i[23887];
  assign o[23886] = i[23886];
  assign o[23885] = i[23885];
  assign o[23884] = i[23884];
  assign o[23883] = i[23883];
  assign o[23882] = i[23882];
  assign o[23881] = i[23881];
  assign o[23880] = i[23880];
  assign o[23879] = i[23879];
  assign o[23878] = i[23878];
  assign o[23877] = i[23877];
  assign o[23876] = i[23876];
  assign o[23875] = i[23875];
  assign o[23874] = i[23874];
  assign o[23873] = i[23873];
  assign o[23872] = i[23872];
  assign o[23871] = i[23871];
  assign o[23870] = i[23870];
  assign o[23869] = i[23869];
  assign o[23868] = i[23868];
  assign o[23867] = i[23867];
  assign o[23866] = i[23866];
  assign o[23865] = i[23865];
  assign o[23864] = i[23864];
  assign o[23863] = i[23863];
  assign o[23862] = i[23862];
  assign o[23861] = i[23861];
  assign o[23860] = i[23860];
  assign o[23859] = i[23859];
  assign o[23858] = i[23858];
  assign o[23857] = i[23857];
  assign o[23856] = i[23856];
  assign o[23855] = i[23855];
  assign o[23854] = i[23854];
  assign o[23853] = i[23853];
  assign o[23852] = i[23852];
  assign o[23851] = i[23851];
  assign o[23850] = i[23850];
  assign o[23849] = i[23849];
  assign o[23848] = i[23848];
  assign o[23847] = i[23847];
  assign o[23846] = i[23846];
  assign o[23845] = i[23845];
  assign o[23844] = i[23844];
  assign o[23843] = i[23843];
  assign o[23842] = i[23842];
  assign o[23841] = i[23841];
  assign o[23840] = i[23840];
  assign o[23839] = i[23839];
  assign o[23838] = i[23838];
  assign o[23837] = i[23837];
  assign o[23836] = i[23836];
  assign o[23835] = i[23835];
  assign o[23834] = i[23834];
  assign o[23833] = i[23833];
  assign o[23832] = i[23832];
  assign o[23831] = i[23831];
  assign o[23830] = i[23830];
  assign o[23829] = i[23829];
  assign o[23828] = i[23828];
  assign o[23827] = i[23827];
  assign o[23826] = i[23826];
  assign o[23825] = i[23825];
  assign o[23824] = i[23824];
  assign o[23823] = i[23823];
  assign o[23822] = i[23822];
  assign o[23821] = i[23821];
  assign o[23820] = i[23820];
  assign o[23819] = i[23819];
  assign o[23818] = i[23818];
  assign o[23817] = i[23817];
  assign o[23816] = i[23816];
  assign o[23815] = i[23815];
  assign o[23814] = i[23814];
  assign o[23813] = i[23813];
  assign o[23812] = i[23812];
  assign o[23811] = i[23811];
  assign o[23810] = i[23810];
  assign o[23809] = i[23809];
  assign o[23808] = i[23808];
  assign o[23807] = i[23807];
  assign o[23806] = i[23806];
  assign o[23805] = i[23805];
  assign o[23804] = i[23804];
  assign o[23803] = i[23803];
  assign o[23802] = i[23802];
  assign o[23801] = i[23801];
  assign o[23800] = i[23800];
  assign o[23799] = i[23799];
  assign o[23798] = i[23798];
  assign o[23797] = i[23797];
  assign o[23796] = i[23796];
  assign o[23795] = i[23795];
  assign o[23794] = i[23794];
  assign o[23793] = i[23793];
  assign o[23792] = i[23792];
  assign o[23791] = i[23791];
  assign o[23790] = i[23790];
  assign o[23789] = i[23789];
  assign o[23788] = i[23788];
  assign o[23787] = i[23787];
  assign o[23786] = i[23786];
  assign o[23785] = i[23785];
  assign o[23784] = i[23784];
  assign o[23783] = i[23783];
  assign o[23782] = i[23782];
  assign o[23781] = i[23781];
  assign o[23780] = i[23780];
  assign o[23779] = i[23779];
  assign o[23778] = i[23778];
  assign o[23777] = i[23777];
  assign o[23776] = i[23776];
  assign o[23775] = i[23775];
  assign o[23774] = i[23774];
  assign o[23773] = i[23773];
  assign o[23772] = i[23772];
  assign o[23771] = i[23771];
  assign o[23770] = i[23770];
  assign o[23769] = i[23769];
  assign o[23768] = i[23768];
  assign o[23767] = i[23767];
  assign o[23766] = i[23766];
  assign o[23765] = i[23765];
  assign o[23764] = i[23764];
  assign o[23763] = i[23763];
  assign o[23762] = i[23762];
  assign o[23761] = i[23761];
  assign o[23760] = i[23760];
  assign o[23759] = i[23759];
  assign o[23758] = i[23758];
  assign o[23757] = i[23757];
  assign o[23756] = i[23756];
  assign o[23755] = i[23755];
  assign o[23754] = i[23754];
  assign o[23753] = i[23753];
  assign o[23752] = i[23752];
  assign o[23751] = i[23751];
  assign o[23750] = i[23750];
  assign o[23749] = i[23749];
  assign o[23748] = i[23748];
  assign o[23747] = i[23747];
  assign o[23746] = i[23746];
  assign o[23745] = i[23745];
  assign o[23744] = i[23744];
  assign o[23743] = i[23743];
  assign o[23742] = i[23742];
  assign o[23741] = i[23741];
  assign o[23740] = i[23740];
  assign o[23739] = i[23739];
  assign o[23738] = i[23738];
  assign o[23737] = i[23737];
  assign o[23736] = i[23736];
  assign o[23735] = i[23735];
  assign o[23734] = i[23734];
  assign o[23733] = i[23733];
  assign o[23732] = i[23732];
  assign o[23731] = i[23731];
  assign o[23730] = i[23730];
  assign o[23729] = i[23729];
  assign o[23728] = i[23728];
  assign o[23727] = i[23727];
  assign o[23726] = i[23726];
  assign o[23725] = i[23725];
  assign o[23724] = i[23724];
  assign o[23723] = i[23723];
  assign o[23722] = i[23722];
  assign o[23721] = i[23721];
  assign o[23720] = i[23720];
  assign o[23719] = i[23719];
  assign o[23718] = i[23718];
  assign o[23717] = i[23717];
  assign o[23716] = i[23716];
  assign o[23715] = i[23715];
  assign o[23714] = i[23714];
  assign o[23713] = i[23713];
  assign o[23712] = i[23712];
  assign o[23711] = i[23711];
  assign o[23710] = i[23710];
  assign o[23709] = i[23709];
  assign o[23708] = i[23708];
  assign o[23707] = i[23707];
  assign o[23706] = i[23706];
  assign o[23705] = i[23705];
  assign o[23704] = i[23704];
  assign o[23703] = i[23703];
  assign o[23702] = i[23702];
  assign o[23701] = i[23701];
  assign o[23700] = i[23700];
  assign o[23699] = i[23699];
  assign o[23698] = i[23698];
  assign o[23697] = i[23697];
  assign o[23696] = i[23696];
  assign o[23695] = i[23695];
  assign o[23694] = i[23694];
  assign o[23693] = i[23693];
  assign o[23692] = i[23692];
  assign o[23691] = i[23691];
  assign o[23690] = i[23690];
  assign o[23689] = i[23689];
  assign o[23688] = i[23688];
  assign o[23687] = i[23687];
  assign o[23686] = i[23686];
  assign o[23685] = i[23685];
  assign o[23684] = i[23684];
  assign o[23683] = i[23683];
  assign o[23682] = i[23682];
  assign o[23681] = i[23681];
  assign o[23680] = i[23680];
  assign o[23679] = i[23679];
  assign o[23678] = i[23678];
  assign o[23677] = i[23677];
  assign o[23676] = i[23676];
  assign o[23675] = i[23675];
  assign o[23674] = i[23674];
  assign o[23673] = i[23673];
  assign o[23672] = i[23672];
  assign o[23671] = i[23671];
  assign o[23670] = i[23670];
  assign o[23669] = i[23669];
  assign o[23668] = i[23668];
  assign o[23667] = i[23667];
  assign o[23666] = i[23666];
  assign o[23665] = i[23665];
  assign o[23664] = i[23664];
  assign o[23663] = i[23663];
  assign o[23662] = i[23662];
  assign o[23661] = i[23661];
  assign o[23660] = i[23660];
  assign o[23659] = i[23659];
  assign o[23658] = i[23658];
  assign o[23657] = i[23657];
  assign o[23656] = i[23656];
  assign o[23655] = i[23655];
  assign o[23654] = i[23654];
  assign o[23653] = i[23653];
  assign o[23652] = i[23652];
  assign o[23651] = i[23651];
  assign o[23650] = i[23650];
  assign o[23649] = i[23649];
  assign o[23648] = i[23648];
  assign o[23647] = i[23647];
  assign o[23646] = i[23646];
  assign o[23645] = i[23645];
  assign o[23644] = i[23644];
  assign o[23643] = i[23643];
  assign o[23642] = i[23642];
  assign o[23641] = i[23641];
  assign o[23640] = i[23640];
  assign o[23639] = i[23639];
  assign o[23638] = i[23638];
  assign o[23637] = i[23637];
  assign o[23636] = i[23636];
  assign o[23635] = i[23635];
  assign o[23634] = i[23634];
  assign o[23633] = i[23633];
  assign o[23632] = i[23632];
  assign o[23631] = i[23631];
  assign o[23630] = i[23630];
  assign o[23629] = i[23629];
  assign o[23628] = i[23628];
  assign o[23627] = i[23627];
  assign o[23626] = i[23626];
  assign o[23625] = i[23625];
  assign o[23624] = i[23624];
  assign o[23623] = i[23623];
  assign o[23622] = i[23622];
  assign o[23621] = i[23621];
  assign o[23620] = i[23620];
  assign o[23619] = i[23619];
  assign o[23618] = i[23618];
  assign o[23617] = i[23617];
  assign o[23616] = i[23616];
  assign o[23615] = i[23615];
  assign o[23614] = i[23614];
  assign o[23613] = i[23613];
  assign o[23612] = i[23612];
  assign o[23611] = i[23611];
  assign o[23610] = i[23610];
  assign o[23609] = i[23609];
  assign o[23608] = i[23608];
  assign o[23607] = i[23607];
  assign o[23606] = i[23606];
  assign o[23605] = i[23605];
  assign o[23604] = i[23604];
  assign o[23603] = i[23603];
  assign o[23602] = i[23602];
  assign o[23601] = i[23601];
  assign o[23600] = i[23600];
  assign o[23599] = i[23599];
  assign o[23598] = i[23598];
  assign o[23597] = i[23597];
  assign o[23596] = i[23596];
  assign o[23595] = i[23595];
  assign o[23594] = i[23594];
  assign o[23593] = i[23593];
  assign o[23592] = i[23592];
  assign o[23591] = i[23591];
  assign o[23590] = i[23590];
  assign o[23589] = i[23589];
  assign o[23588] = i[23588];
  assign o[23587] = i[23587];
  assign o[23586] = i[23586];
  assign o[23585] = i[23585];
  assign o[23584] = i[23584];
  assign o[23583] = i[23583];
  assign o[23582] = i[23582];
  assign o[23581] = i[23581];
  assign o[23580] = i[23580];
  assign o[23579] = i[23579];
  assign o[23578] = i[23578];
  assign o[23577] = i[23577];
  assign o[23576] = i[23576];
  assign o[23575] = i[23575];
  assign o[23574] = i[23574];
  assign o[23573] = i[23573];
  assign o[23572] = i[23572];
  assign o[23571] = i[23571];
  assign o[23570] = i[23570];
  assign o[23569] = i[23569];
  assign o[23568] = i[23568];
  assign o[23567] = i[23567];
  assign o[23566] = i[23566];
  assign o[23565] = i[23565];
  assign o[23564] = i[23564];
  assign o[23563] = i[23563];
  assign o[23562] = i[23562];
  assign o[23561] = i[23561];
  assign o[23560] = i[23560];
  assign o[23559] = i[23559];
  assign o[23558] = i[23558];
  assign o[23557] = i[23557];
  assign o[23556] = i[23556];
  assign o[23555] = i[23555];
  assign o[23554] = i[23554];
  assign o[23553] = i[23553];
  assign o[23552] = i[23552];
  assign o[23551] = i[23551];
  assign o[23550] = i[23550];
  assign o[23549] = i[23549];
  assign o[23548] = i[23548];
  assign o[23547] = i[23547];
  assign o[23546] = i[23546];
  assign o[23545] = i[23545];
  assign o[23544] = i[23544];
  assign o[23543] = i[23543];
  assign o[23542] = i[23542];
  assign o[23541] = i[23541];
  assign o[23540] = i[23540];
  assign o[23539] = i[23539];
  assign o[23538] = i[23538];
  assign o[23537] = i[23537];
  assign o[23536] = i[23536];
  assign o[23535] = i[23535];
  assign o[23534] = i[23534];
  assign o[23533] = i[23533];
  assign o[23532] = i[23532];
  assign o[23531] = i[23531];
  assign o[23530] = i[23530];
  assign o[23529] = i[23529];
  assign o[23528] = i[23528];
  assign o[23527] = i[23527];
  assign o[23526] = i[23526];
  assign o[23525] = i[23525];
  assign o[23524] = i[23524];
  assign o[23523] = i[23523];
  assign o[23522] = i[23522];
  assign o[23521] = i[23521];
  assign o[23520] = i[23520];
  assign o[23519] = i[23519];
  assign o[23518] = i[23518];
  assign o[23517] = i[23517];
  assign o[23516] = i[23516];
  assign o[23515] = i[23515];
  assign o[23514] = i[23514];
  assign o[23513] = i[23513];
  assign o[23512] = i[23512];
  assign o[23511] = i[23511];
  assign o[23510] = i[23510];
  assign o[23509] = i[23509];
  assign o[23508] = i[23508];
  assign o[23507] = i[23507];
  assign o[23506] = i[23506];
  assign o[23505] = i[23505];
  assign o[23504] = i[23504];
  assign o[23503] = i[23503];
  assign o[23502] = i[23502];
  assign o[23501] = i[23501];
  assign o[23500] = i[23500];
  assign o[23499] = i[23499];
  assign o[23498] = i[23498];
  assign o[23497] = i[23497];
  assign o[23496] = i[23496];
  assign o[23495] = i[23495];
  assign o[23494] = i[23494];
  assign o[23493] = i[23493];
  assign o[23492] = i[23492];
  assign o[23491] = i[23491];
  assign o[23490] = i[23490];
  assign o[23489] = i[23489];
  assign o[23488] = i[23488];
  assign o[23487] = i[23487];
  assign o[23486] = i[23486];
  assign o[23485] = i[23485];
  assign o[23484] = i[23484];
  assign o[23483] = i[23483];
  assign o[23482] = i[23482];
  assign o[23481] = i[23481];
  assign o[23480] = i[23480];
  assign o[23479] = i[23479];
  assign o[23478] = i[23478];
  assign o[23477] = i[23477];
  assign o[23476] = i[23476];
  assign o[23475] = i[23475];
  assign o[23474] = i[23474];
  assign o[23473] = i[23473];
  assign o[23472] = i[23472];
  assign o[23471] = i[23471];
  assign o[23470] = i[23470];
  assign o[23469] = i[23469];
  assign o[23468] = i[23468];
  assign o[23467] = i[23467];
  assign o[23466] = i[23466];
  assign o[23465] = i[23465];
  assign o[23464] = i[23464];
  assign o[23463] = i[23463];
  assign o[23462] = i[23462];
  assign o[23461] = i[23461];
  assign o[23460] = i[23460];
  assign o[23459] = i[23459];
  assign o[23458] = i[23458];
  assign o[23457] = i[23457];
  assign o[23456] = i[23456];
  assign o[23455] = i[23455];
  assign o[23454] = i[23454];
  assign o[23453] = i[23453];
  assign o[23452] = i[23452];
  assign o[23451] = i[23451];
  assign o[23450] = i[23450];
  assign o[23449] = i[23449];
  assign o[23448] = i[23448];
  assign o[23447] = i[23447];
  assign o[23446] = i[23446];
  assign o[23445] = i[23445];
  assign o[23444] = i[23444];
  assign o[23443] = i[23443];
  assign o[23442] = i[23442];
  assign o[23441] = i[23441];
  assign o[23440] = i[23440];
  assign o[23439] = i[23439];
  assign o[23438] = i[23438];
  assign o[23437] = i[23437];
  assign o[23436] = i[23436];
  assign o[23435] = i[23435];
  assign o[23434] = i[23434];
  assign o[23433] = i[23433];
  assign o[23432] = i[23432];
  assign o[23431] = i[23431];
  assign o[23430] = i[23430];
  assign o[23429] = i[23429];
  assign o[23428] = i[23428];
  assign o[23427] = i[23427];
  assign o[23426] = i[23426];
  assign o[23425] = i[23425];
  assign o[23424] = i[23424];
  assign o[23423] = i[23423];
  assign o[23422] = i[23422];
  assign o[23421] = i[23421];
  assign o[23420] = i[23420];
  assign o[23419] = i[23419];
  assign o[23418] = i[23418];
  assign o[23417] = i[23417];
  assign o[23416] = i[23416];
  assign o[23415] = i[23415];
  assign o[23414] = i[23414];
  assign o[23413] = i[23413];
  assign o[23412] = i[23412];
  assign o[23411] = i[23411];
  assign o[23410] = i[23410];
  assign o[23409] = i[23409];
  assign o[23408] = i[23408];
  assign o[23407] = i[23407];
  assign o[23406] = i[23406];
  assign o[23405] = i[23405];
  assign o[23404] = i[23404];
  assign o[23403] = i[23403];
  assign o[23402] = i[23402];
  assign o[23401] = i[23401];
  assign o[23400] = i[23400];
  assign o[23399] = i[23399];
  assign o[23398] = i[23398];
  assign o[23397] = i[23397];
  assign o[23396] = i[23396];
  assign o[23395] = i[23395];
  assign o[23394] = i[23394];
  assign o[23393] = i[23393];
  assign o[23392] = i[23392];
  assign o[23391] = i[23391];
  assign o[23390] = i[23390];
  assign o[23389] = i[23389];
  assign o[23388] = i[23388];
  assign o[23387] = i[23387];
  assign o[23386] = i[23386];
  assign o[23385] = i[23385];
  assign o[23384] = i[23384];
  assign o[23383] = i[23383];
  assign o[23382] = i[23382];
  assign o[23381] = i[23381];
  assign o[23380] = i[23380];
  assign o[23379] = i[23379];
  assign o[23378] = i[23378];
  assign o[23377] = i[23377];
  assign o[23376] = i[23376];
  assign o[23375] = i[23375];
  assign o[23374] = i[23374];
  assign o[23373] = i[23373];
  assign o[23372] = i[23372];
  assign o[23371] = i[23371];
  assign o[23370] = i[23370];
  assign o[23369] = i[23369];
  assign o[23368] = i[23368];
  assign o[23367] = i[23367];
  assign o[23366] = i[23366];
  assign o[23365] = i[23365];
  assign o[23364] = i[23364];
  assign o[23363] = i[23363];
  assign o[23362] = i[23362];
  assign o[23361] = i[23361];
  assign o[23360] = i[23360];
  assign o[23359] = i[23359];
  assign o[23358] = i[23358];
  assign o[23357] = i[23357];
  assign o[23356] = i[23356];
  assign o[23355] = i[23355];
  assign o[23354] = i[23354];
  assign o[23353] = i[23353];
  assign o[23352] = i[23352];
  assign o[23351] = i[23351];
  assign o[23350] = i[23350];
  assign o[23349] = i[23349];
  assign o[23348] = i[23348];
  assign o[23347] = i[23347];
  assign o[23346] = i[23346];
  assign o[23345] = i[23345];
  assign o[23344] = i[23344];
  assign o[23343] = i[23343];
  assign o[23342] = i[23342];
  assign o[23341] = i[23341];
  assign o[23340] = i[23340];
  assign o[23339] = i[23339];
  assign o[23338] = i[23338];
  assign o[23337] = i[23337];
  assign o[23336] = i[23336];
  assign o[23335] = i[23335];
  assign o[23334] = i[23334];
  assign o[23333] = i[23333];
  assign o[23332] = i[23332];
  assign o[23331] = i[23331];
  assign o[23330] = i[23330];
  assign o[23329] = i[23329];
  assign o[23328] = i[23328];
  assign o[23327] = i[23327];
  assign o[23326] = i[23326];
  assign o[23325] = i[23325];
  assign o[23324] = i[23324];
  assign o[23323] = i[23323];
  assign o[23322] = i[23322];
  assign o[23321] = i[23321];
  assign o[23320] = i[23320];
  assign o[23319] = i[23319];
  assign o[23318] = i[23318];
  assign o[23317] = i[23317];
  assign o[23316] = i[23316];
  assign o[23315] = i[23315];
  assign o[23314] = i[23314];
  assign o[23313] = i[23313];
  assign o[23312] = i[23312];
  assign o[23311] = i[23311];
  assign o[23310] = i[23310];
  assign o[23309] = i[23309];
  assign o[23308] = i[23308];
  assign o[23307] = i[23307];
  assign o[23306] = i[23306];
  assign o[23305] = i[23305];
  assign o[23304] = i[23304];
  assign o[23303] = i[23303];
  assign o[23302] = i[23302];
  assign o[23301] = i[23301];
  assign o[23300] = i[23300];
  assign o[23299] = i[23299];
  assign o[23298] = i[23298];
  assign o[23297] = i[23297];
  assign o[23296] = i[23296];
  assign o[23295] = i[23295];
  assign o[23294] = i[23294];
  assign o[23293] = i[23293];
  assign o[23292] = i[23292];
  assign o[23291] = i[23291];
  assign o[23290] = i[23290];
  assign o[23289] = i[23289];
  assign o[23288] = i[23288];
  assign o[23287] = i[23287];
  assign o[23286] = i[23286];
  assign o[23285] = i[23285];
  assign o[23284] = i[23284];
  assign o[23283] = i[23283];
  assign o[23282] = i[23282];
  assign o[23281] = i[23281];
  assign o[23280] = i[23280];
  assign o[23279] = i[23279];
  assign o[23278] = i[23278];
  assign o[23277] = i[23277];
  assign o[23276] = i[23276];
  assign o[23275] = i[23275];
  assign o[23274] = i[23274];
  assign o[23273] = i[23273];
  assign o[23272] = i[23272];
  assign o[23271] = i[23271];
  assign o[23270] = i[23270];
  assign o[23269] = i[23269];
  assign o[23268] = i[23268];
  assign o[23267] = i[23267];
  assign o[23266] = i[23266];
  assign o[23265] = i[23265];
  assign o[23264] = i[23264];
  assign o[23263] = i[23263];
  assign o[23262] = i[23262];
  assign o[23261] = i[23261];
  assign o[23260] = i[23260];
  assign o[23259] = i[23259];
  assign o[23258] = i[23258];
  assign o[23257] = i[23257];
  assign o[23256] = i[23256];
  assign o[23255] = i[23255];
  assign o[23254] = i[23254];
  assign o[23253] = i[23253];
  assign o[23252] = i[23252];
  assign o[23251] = i[23251];
  assign o[23250] = i[23250];
  assign o[23249] = i[23249];
  assign o[23248] = i[23248];
  assign o[23247] = i[23247];
  assign o[23246] = i[23246];
  assign o[23245] = i[23245];
  assign o[23244] = i[23244];
  assign o[23243] = i[23243];
  assign o[23242] = i[23242];
  assign o[23241] = i[23241];
  assign o[23240] = i[23240];
  assign o[23239] = i[23239];
  assign o[23238] = i[23238];
  assign o[23237] = i[23237];
  assign o[23236] = i[23236];
  assign o[23235] = i[23235];
  assign o[23234] = i[23234];
  assign o[23233] = i[23233];
  assign o[23232] = i[23232];
  assign o[23231] = i[23231];
  assign o[23230] = i[23230];
  assign o[23229] = i[23229];
  assign o[23228] = i[23228];
  assign o[23227] = i[23227];
  assign o[23226] = i[23226];
  assign o[23225] = i[23225];
  assign o[23224] = i[23224];
  assign o[23223] = i[23223];
  assign o[23222] = i[23222];
  assign o[23221] = i[23221];
  assign o[23220] = i[23220];
  assign o[23219] = i[23219];
  assign o[23218] = i[23218];
  assign o[23217] = i[23217];
  assign o[23216] = i[23216];
  assign o[23215] = i[23215];
  assign o[23214] = i[23214];
  assign o[23213] = i[23213];
  assign o[23212] = i[23212];
  assign o[23211] = i[23211];
  assign o[23210] = i[23210];
  assign o[23209] = i[23209];
  assign o[23208] = i[23208];
  assign o[23207] = i[23207];
  assign o[23206] = i[23206];
  assign o[23205] = i[23205];
  assign o[23204] = i[23204];
  assign o[23203] = i[23203];
  assign o[23202] = i[23202];
  assign o[23201] = i[23201];
  assign o[23200] = i[23200];
  assign o[23199] = i[23199];
  assign o[23198] = i[23198];
  assign o[23197] = i[23197];
  assign o[23196] = i[23196];
  assign o[23195] = i[23195];
  assign o[23194] = i[23194];
  assign o[23193] = i[23193];
  assign o[23192] = i[23192];
  assign o[23191] = i[23191];
  assign o[23190] = i[23190];
  assign o[23189] = i[23189];
  assign o[23188] = i[23188];
  assign o[23187] = i[23187];
  assign o[23186] = i[23186];
  assign o[23185] = i[23185];
  assign o[23184] = i[23184];
  assign o[23183] = i[23183];
  assign o[23182] = i[23182];
  assign o[23181] = i[23181];
  assign o[23180] = i[23180];
  assign o[23179] = i[23179];
  assign o[23178] = i[23178];
  assign o[23177] = i[23177];
  assign o[23176] = i[23176];
  assign o[23175] = i[23175];
  assign o[23174] = i[23174];
  assign o[23173] = i[23173];
  assign o[23172] = i[23172];
  assign o[23171] = i[23171];
  assign o[23170] = i[23170];
  assign o[23169] = i[23169];
  assign o[23168] = i[23168];
  assign o[23167] = i[23167];
  assign o[23166] = i[23166];
  assign o[23165] = i[23165];
  assign o[23164] = i[23164];
  assign o[23163] = i[23163];
  assign o[23162] = i[23162];
  assign o[23161] = i[23161];
  assign o[23160] = i[23160];
  assign o[23159] = i[23159];
  assign o[23158] = i[23158];
  assign o[23157] = i[23157];
  assign o[23156] = i[23156];
  assign o[23155] = i[23155];
  assign o[23154] = i[23154];
  assign o[23153] = i[23153];
  assign o[23152] = i[23152];
  assign o[23151] = i[23151];
  assign o[23150] = i[23150];
  assign o[23149] = i[23149];
  assign o[23148] = i[23148];
  assign o[23147] = i[23147];
  assign o[23146] = i[23146];
  assign o[23145] = i[23145];
  assign o[23144] = i[23144];
  assign o[23143] = i[23143];
  assign o[23142] = i[23142];
  assign o[23141] = i[23141];
  assign o[23140] = i[23140];
  assign o[23139] = i[23139];
  assign o[23138] = i[23138];
  assign o[23137] = i[23137];
  assign o[23136] = i[23136];
  assign o[23135] = i[23135];
  assign o[23134] = i[23134];
  assign o[23133] = i[23133];
  assign o[23132] = i[23132];
  assign o[23131] = i[23131];
  assign o[23130] = i[23130];
  assign o[23129] = i[23129];
  assign o[23128] = i[23128];
  assign o[23127] = i[23127];
  assign o[23126] = i[23126];
  assign o[23125] = i[23125];
  assign o[23124] = i[23124];
  assign o[23123] = i[23123];
  assign o[23122] = i[23122];
  assign o[23121] = i[23121];
  assign o[23120] = i[23120];
  assign o[23119] = i[23119];
  assign o[23118] = i[23118];
  assign o[23117] = i[23117];
  assign o[23116] = i[23116];
  assign o[23115] = i[23115];
  assign o[23114] = i[23114];
  assign o[23113] = i[23113];
  assign o[23112] = i[23112];
  assign o[23111] = i[23111];
  assign o[23110] = i[23110];
  assign o[23109] = i[23109];
  assign o[23108] = i[23108];
  assign o[23107] = i[23107];
  assign o[23106] = i[23106];
  assign o[23105] = i[23105];
  assign o[23104] = i[23104];
  assign o[23103] = i[23103];
  assign o[23102] = i[23102];
  assign o[23101] = i[23101];
  assign o[23100] = i[23100];
  assign o[23099] = i[23099];
  assign o[23098] = i[23098];
  assign o[23097] = i[23097];
  assign o[23096] = i[23096];
  assign o[23095] = i[23095];
  assign o[23094] = i[23094];
  assign o[23093] = i[23093];
  assign o[23092] = i[23092];
  assign o[23091] = i[23091];
  assign o[23090] = i[23090];
  assign o[23089] = i[23089];
  assign o[23088] = i[23088];
  assign o[23087] = i[23087];
  assign o[23086] = i[23086];
  assign o[23085] = i[23085];
  assign o[23084] = i[23084];
  assign o[23083] = i[23083];
  assign o[23082] = i[23082];
  assign o[23081] = i[23081];
  assign o[23080] = i[23080];
  assign o[23079] = i[23079];
  assign o[23078] = i[23078];
  assign o[23077] = i[23077];
  assign o[23076] = i[23076];
  assign o[23075] = i[23075];
  assign o[23074] = i[23074];
  assign o[23073] = i[23073];
  assign o[23072] = i[23072];
  assign o[23071] = i[23071];
  assign o[23070] = i[23070];
  assign o[23069] = i[23069];
  assign o[23068] = i[23068];
  assign o[23067] = i[23067];
  assign o[23066] = i[23066];
  assign o[23065] = i[23065];
  assign o[23064] = i[23064];
  assign o[23063] = i[23063];
  assign o[23062] = i[23062];
  assign o[23061] = i[23061];
  assign o[23060] = i[23060];
  assign o[23059] = i[23059];
  assign o[23058] = i[23058];
  assign o[23057] = i[23057];
  assign o[23056] = i[23056];
  assign o[23055] = i[23055];
  assign o[23054] = i[23054];
  assign o[23053] = i[23053];
  assign o[23052] = i[23052];
  assign o[23051] = i[23051];
  assign o[23050] = i[23050];
  assign o[23049] = i[23049];
  assign o[23048] = i[23048];
  assign o[23047] = i[23047];
  assign o[23046] = i[23046];
  assign o[23045] = i[23045];
  assign o[23044] = i[23044];
  assign o[23043] = i[23043];
  assign o[23042] = i[23042];
  assign o[23041] = i[23041];
  assign o[23040] = i[23040];
  assign o[23039] = i[23039];
  assign o[23038] = i[23038];
  assign o[23037] = i[23037];
  assign o[23036] = i[23036];
  assign o[23035] = i[23035];
  assign o[23034] = i[23034];
  assign o[23033] = i[23033];
  assign o[23032] = i[23032];
  assign o[23031] = i[23031];
  assign o[23030] = i[23030];
  assign o[23029] = i[23029];
  assign o[23028] = i[23028];
  assign o[23027] = i[23027];
  assign o[23026] = i[23026];
  assign o[23025] = i[23025];
  assign o[23024] = i[23024];
  assign o[23023] = i[23023];
  assign o[23022] = i[23022];
  assign o[23021] = i[23021];
  assign o[23020] = i[23020];
  assign o[23019] = i[23019];
  assign o[23018] = i[23018];
  assign o[23017] = i[23017];
  assign o[23016] = i[23016];
  assign o[23015] = i[23015];
  assign o[23014] = i[23014];
  assign o[23013] = i[23013];
  assign o[23012] = i[23012];
  assign o[23011] = i[23011];
  assign o[23010] = i[23010];
  assign o[23009] = i[23009];
  assign o[23008] = i[23008];
  assign o[23007] = i[23007];
  assign o[23006] = i[23006];
  assign o[23005] = i[23005];
  assign o[23004] = i[23004];
  assign o[23003] = i[23003];
  assign o[23002] = i[23002];
  assign o[23001] = i[23001];
  assign o[23000] = i[23000];
  assign o[22999] = i[22999];
  assign o[22998] = i[22998];
  assign o[22997] = i[22997];
  assign o[22996] = i[22996];
  assign o[22995] = i[22995];
  assign o[22994] = i[22994];
  assign o[22993] = i[22993];
  assign o[22992] = i[22992];
  assign o[22991] = i[22991];
  assign o[22990] = i[22990];
  assign o[22989] = i[22989];
  assign o[22988] = i[22988];
  assign o[22987] = i[22987];
  assign o[22986] = i[22986];
  assign o[22985] = i[22985];
  assign o[22984] = i[22984];
  assign o[22983] = i[22983];
  assign o[22982] = i[22982];
  assign o[22981] = i[22981];
  assign o[22980] = i[22980];
  assign o[22979] = i[22979];
  assign o[22978] = i[22978];
  assign o[22977] = i[22977];
  assign o[22976] = i[22976];
  assign o[22975] = i[22975];
  assign o[22974] = i[22974];
  assign o[22973] = i[22973];
  assign o[22972] = i[22972];
  assign o[22971] = i[22971];
  assign o[22970] = i[22970];
  assign o[22969] = i[22969];
  assign o[22968] = i[22968];
  assign o[22967] = i[22967];
  assign o[22966] = i[22966];
  assign o[22965] = i[22965];
  assign o[22964] = i[22964];
  assign o[22963] = i[22963];
  assign o[22962] = i[22962];
  assign o[22961] = i[22961];
  assign o[22960] = i[22960];
  assign o[22959] = i[22959];
  assign o[22958] = i[22958];
  assign o[22957] = i[22957];
  assign o[22956] = i[22956];
  assign o[22955] = i[22955];
  assign o[22954] = i[22954];
  assign o[22953] = i[22953];
  assign o[22952] = i[22952];
  assign o[22951] = i[22951];
  assign o[22950] = i[22950];
  assign o[22949] = i[22949];
  assign o[22948] = i[22948];
  assign o[22947] = i[22947];
  assign o[22946] = i[22946];
  assign o[22945] = i[22945];
  assign o[22944] = i[22944];
  assign o[22943] = i[22943];
  assign o[22942] = i[22942];
  assign o[22941] = i[22941];
  assign o[22940] = i[22940];
  assign o[22939] = i[22939];
  assign o[22938] = i[22938];
  assign o[22937] = i[22937];
  assign o[22936] = i[22936];
  assign o[22935] = i[22935];
  assign o[22934] = i[22934];
  assign o[22933] = i[22933];
  assign o[22932] = i[22932];
  assign o[22931] = i[22931];
  assign o[22930] = i[22930];
  assign o[22929] = i[22929];
  assign o[22928] = i[22928];
  assign o[22927] = i[22927];
  assign o[22926] = i[22926];
  assign o[22925] = i[22925];
  assign o[22924] = i[22924];
  assign o[22923] = i[22923];
  assign o[22922] = i[22922];
  assign o[22921] = i[22921];
  assign o[22920] = i[22920];
  assign o[22919] = i[22919];
  assign o[22918] = i[22918];
  assign o[22917] = i[22917];
  assign o[22916] = i[22916];
  assign o[22915] = i[22915];
  assign o[22914] = i[22914];
  assign o[22913] = i[22913];
  assign o[22912] = i[22912];
  assign o[22911] = i[22911];
  assign o[22910] = i[22910];
  assign o[22909] = i[22909];
  assign o[22908] = i[22908];
  assign o[22907] = i[22907];
  assign o[22906] = i[22906];
  assign o[22905] = i[22905];
  assign o[22904] = i[22904];
  assign o[22903] = i[22903];
  assign o[22902] = i[22902];
  assign o[22901] = i[22901];
  assign o[22900] = i[22900];
  assign o[22899] = i[22899];
  assign o[22898] = i[22898];
  assign o[22897] = i[22897];
  assign o[22896] = i[22896];
  assign o[22895] = i[22895];
  assign o[22894] = i[22894];
  assign o[22893] = i[22893];
  assign o[22892] = i[22892];
  assign o[22891] = i[22891];
  assign o[22890] = i[22890];
  assign o[22889] = i[22889];
  assign o[22888] = i[22888];
  assign o[22887] = i[22887];
  assign o[22886] = i[22886];
  assign o[22885] = i[22885];
  assign o[22884] = i[22884];
  assign o[22883] = i[22883];
  assign o[22882] = i[22882];
  assign o[22881] = i[22881];
  assign o[22880] = i[22880];
  assign o[22879] = i[22879];
  assign o[22878] = i[22878];
  assign o[22877] = i[22877];
  assign o[22876] = i[22876];
  assign o[22875] = i[22875];
  assign o[22874] = i[22874];
  assign o[22873] = i[22873];
  assign o[22872] = i[22872];
  assign o[22871] = i[22871];
  assign o[22870] = i[22870];
  assign o[22869] = i[22869];
  assign o[22868] = i[22868];
  assign o[22867] = i[22867];
  assign o[22866] = i[22866];
  assign o[22865] = i[22865];
  assign o[22864] = i[22864];
  assign o[22863] = i[22863];
  assign o[22862] = i[22862];
  assign o[22861] = i[22861];
  assign o[22860] = i[22860];
  assign o[22859] = i[22859];
  assign o[22858] = i[22858];
  assign o[22857] = i[22857];
  assign o[22856] = i[22856];
  assign o[22855] = i[22855];
  assign o[22854] = i[22854];
  assign o[22853] = i[22853];
  assign o[22852] = i[22852];
  assign o[22851] = i[22851];
  assign o[22850] = i[22850];
  assign o[22849] = i[22849];
  assign o[22848] = i[22848];
  assign o[22847] = i[22847];
  assign o[22846] = i[22846];
  assign o[22845] = i[22845];
  assign o[22844] = i[22844];
  assign o[22843] = i[22843];
  assign o[22842] = i[22842];
  assign o[22841] = i[22841];
  assign o[22840] = i[22840];
  assign o[22839] = i[22839];
  assign o[22838] = i[22838];
  assign o[22837] = i[22837];
  assign o[22836] = i[22836];
  assign o[22835] = i[22835];
  assign o[22834] = i[22834];
  assign o[22833] = i[22833];
  assign o[22832] = i[22832];
  assign o[22831] = i[22831];
  assign o[22830] = i[22830];
  assign o[22829] = i[22829];
  assign o[22828] = i[22828];
  assign o[22827] = i[22827];
  assign o[22826] = i[22826];
  assign o[22825] = i[22825];
  assign o[22824] = i[22824];
  assign o[22823] = i[22823];
  assign o[22822] = i[22822];
  assign o[22821] = i[22821];
  assign o[22820] = i[22820];
  assign o[22819] = i[22819];
  assign o[22818] = i[22818];
  assign o[22817] = i[22817];
  assign o[22816] = i[22816];
  assign o[22815] = i[22815];
  assign o[22814] = i[22814];
  assign o[22813] = i[22813];
  assign o[22812] = i[22812];
  assign o[22811] = i[22811];
  assign o[22810] = i[22810];
  assign o[22809] = i[22809];
  assign o[22808] = i[22808];
  assign o[22807] = i[22807];
  assign o[22806] = i[22806];
  assign o[22805] = i[22805];
  assign o[22804] = i[22804];
  assign o[22803] = i[22803];
  assign o[22802] = i[22802];
  assign o[22801] = i[22801];
  assign o[22800] = i[22800];
  assign o[22799] = i[22799];
  assign o[22798] = i[22798];
  assign o[22797] = i[22797];
  assign o[22796] = i[22796];
  assign o[22795] = i[22795];
  assign o[22794] = i[22794];
  assign o[22793] = i[22793];
  assign o[22792] = i[22792];
  assign o[22791] = i[22791];
  assign o[22790] = i[22790];
  assign o[22789] = i[22789];
  assign o[22788] = i[22788];
  assign o[22787] = i[22787];
  assign o[22786] = i[22786];
  assign o[22785] = i[22785];
  assign o[22784] = i[22784];
  assign o[22783] = i[22783];
  assign o[22782] = i[22782];
  assign o[22781] = i[22781];
  assign o[22780] = i[22780];
  assign o[22779] = i[22779];
  assign o[22778] = i[22778];
  assign o[22777] = i[22777];
  assign o[22776] = i[22776];
  assign o[22775] = i[22775];
  assign o[22774] = i[22774];
  assign o[22773] = i[22773];
  assign o[22772] = i[22772];
  assign o[22771] = i[22771];
  assign o[22770] = i[22770];
  assign o[22769] = i[22769];
  assign o[22768] = i[22768];
  assign o[22767] = i[22767];
  assign o[22766] = i[22766];
  assign o[22765] = i[22765];
  assign o[22764] = i[22764];
  assign o[22763] = i[22763];
  assign o[22762] = i[22762];
  assign o[22761] = i[22761];
  assign o[22760] = i[22760];
  assign o[22759] = i[22759];
  assign o[22758] = i[22758];
  assign o[22757] = i[22757];
  assign o[22756] = i[22756];
  assign o[22755] = i[22755];
  assign o[22754] = i[22754];
  assign o[22753] = i[22753];
  assign o[22752] = i[22752];
  assign o[22751] = i[22751];
  assign o[22750] = i[22750];
  assign o[22749] = i[22749];
  assign o[22748] = i[22748];
  assign o[22747] = i[22747];
  assign o[22746] = i[22746];
  assign o[22745] = i[22745];
  assign o[22744] = i[22744];
  assign o[22743] = i[22743];
  assign o[22742] = i[22742];
  assign o[22741] = i[22741];
  assign o[22740] = i[22740];
  assign o[22739] = i[22739];
  assign o[22738] = i[22738];
  assign o[22737] = i[22737];
  assign o[22736] = i[22736];
  assign o[22735] = i[22735];
  assign o[22734] = i[22734];
  assign o[22733] = i[22733];
  assign o[22732] = i[22732];
  assign o[22731] = i[22731];
  assign o[22730] = i[22730];
  assign o[22729] = i[22729];
  assign o[22728] = i[22728];
  assign o[22727] = i[22727];
  assign o[22726] = i[22726];
  assign o[22725] = i[22725];
  assign o[22724] = i[22724];
  assign o[22723] = i[22723];
  assign o[22722] = i[22722];
  assign o[22721] = i[22721];
  assign o[22720] = i[22720];
  assign o[22719] = i[22719];
  assign o[22718] = i[22718];
  assign o[22717] = i[22717];
  assign o[22716] = i[22716];
  assign o[22715] = i[22715];
  assign o[22714] = i[22714];
  assign o[22713] = i[22713];
  assign o[22712] = i[22712];
  assign o[22711] = i[22711];
  assign o[22710] = i[22710];
  assign o[22709] = i[22709];
  assign o[22708] = i[22708];
  assign o[22707] = i[22707];
  assign o[22706] = i[22706];
  assign o[22705] = i[22705];
  assign o[22704] = i[22704];
  assign o[22703] = i[22703];
  assign o[22702] = i[22702];
  assign o[22701] = i[22701];
  assign o[22700] = i[22700];
  assign o[22699] = i[22699];
  assign o[22698] = i[22698];
  assign o[22697] = i[22697];
  assign o[22696] = i[22696];
  assign o[22695] = i[22695];
  assign o[22694] = i[22694];
  assign o[22693] = i[22693];
  assign o[22692] = i[22692];
  assign o[22691] = i[22691];
  assign o[22690] = i[22690];
  assign o[22689] = i[22689];
  assign o[22688] = i[22688];
  assign o[22687] = i[22687];
  assign o[22686] = i[22686];
  assign o[22685] = i[22685];
  assign o[22684] = i[22684];
  assign o[22683] = i[22683];
  assign o[22682] = i[22682];
  assign o[22681] = i[22681];
  assign o[22680] = i[22680];
  assign o[22679] = i[22679];
  assign o[22678] = i[22678];
  assign o[22677] = i[22677];
  assign o[22676] = i[22676];
  assign o[22675] = i[22675];
  assign o[22674] = i[22674];
  assign o[22673] = i[22673];
  assign o[22672] = i[22672];
  assign o[22671] = i[22671];
  assign o[22670] = i[22670];
  assign o[22669] = i[22669];
  assign o[22668] = i[22668];
  assign o[22667] = i[22667];
  assign o[22666] = i[22666];
  assign o[22665] = i[22665];
  assign o[22664] = i[22664];
  assign o[22663] = i[22663];
  assign o[22662] = i[22662];
  assign o[22661] = i[22661];
  assign o[22660] = i[22660];
  assign o[22659] = i[22659];
  assign o[22658] = i[22658];
  assign o[22657] = i[22657];
  assign o[22656] = i[22656];
  assign o[22655] = i[22655];
  assign o[22654] = i[22654];
  assign o[22653] = i[22653];
  assign o[22652] = i[22652];
  assign o[22651] = i[22651];
  assign o[22650] = i[22650];
  assign o[22649] = i[22649];
  assign o[22648] = i[22648];
  assign o[22647] = i[22647];
  assign o[22646] = i[22646];
  assign o[22645] = i[22645];
  assign o[22644] = i[22644];
  assign o[22643] = i[22643];
  assign o[22642] = i[22642];
  assign o[22641] = i[22641];
  assign o[22640] = i[22640];
  assign o[22639] = i[22639];
  assign o[22638] = i[22638];
  assign o[22637] = i[22637];
  assign o[22636] = i[22636];
  assign o[22635] = i[22635];
  assign o[22634] = i[22634];
  assign o[22633] = i[22633];
  assign o[22632] = i[22632];
  assign o[22631] = i[22631];
  assign o[22630] = i[22630];
  assign o[22629] = i[22629];
  assign o[22628] = i[22628];
  assign o[22627] = i[22627];
  assign o[22626] = i[22626];
  assign o[22625] = i[22625];
  assign o[22624] = i[22624];
  assign o[22623] = i[22623];
  assign o[22622] = i[22622];
  assign o[22621] = i[22621];
  assign o[22620] = i[22620];
  assign o[22619] = i[22619];
  assign o[22618] = i[22618];
  assign o[22617] = i[22617];
  assign o[22616] = i[22616];
  assign o[22615] = i[22615];
  assign o[22614] = i[22614];
  assign o[22613] = i[22613];
  assign o[22612] = i[22612];
  assign o[22611] = i[22611];
  assign o[22610] = i[22610];
  assign o[22609] = i[22609];
  assign o[22608] = i[22608];
  assign o[22607] = i[22607];
  assign o[22606] = i[22606];
  assign o[22605] = i[22605];
  assign o[22604] = i[22604];
  assign o[22603] = i[22603];
  assign o[22602] = i[22602];
  assign o[22601] = i[22601];
  assign o[22600] = i[22600];
  assign o[22599] = i[22599];
  assign o[22598] = i[22598];
  assign o[22597] = i[22597];
  assign o[22596] = i[22596];
  assign o[22595] = i[22595];
  assign o[22594] = i[22594];
  assign o[22593] = i[22593];
  assign o[22592] = i[22592];
  assign o[22591] = i[22591];
  assign o[22590] = i[22590];
  assign o[22589] = i[22589];
  assign o[22588] = i[22588];
  assign o[22587] = i[22587];
  assign o[22586] = i[22586];
  assign o[22585] = i[22585];
  assign o[22584] = i[22584];
  assign o[22583] = i[22583];
  assign o[22582] = i[22582];
  assign o[22581] = i[22581];
  assign o[22580] = i[22580];
  assign o[22579] = i[22579];
  assign o[22578] = i[22578];
  assign o[22577] = i[22577];
  assign o[22576] = i[22576];
  assign o[22575] = i[22575];
  assign o[22574] = i[22574];
  assign o[22573] = i[22573];
  assign o[22572] = i[22572];
  assign o[22571] = i[22571];
  assign o[22570] = i[22570];
  assign o[22569] = i[22569];
  assign o[22568] = i[22568];
  assign o[22567] = i[22567];
  assign o[22566] = i[22566];
  assign o[22565] = i[22565];
  assign o[22564] = i[22564];
  assign o[22563] = i[22563];
  assign o[22562] = i[22562];
  assign o[22561] = i[22561];
  assign o[22560] = i[22560];
  assign o[22559] = i[22559];
  assign o[22558] = i[22558];
  assign o[22557] = i[22557];
  assign o[22556] = i[22556];
  assign o[22555] = i[22555];
  assign o[22554] = i[22554];
  assign o[22553] = i[22553];
  assign o[22552] = i[22552];
  assign o[22551] = i[22551];
  assign o[22550] = i[22550];
  assign o[22549] = i[22549];
  assign o[22548] = i[22548];
  assign o[22547] = i[22547];
  assign o[22546] = i[22546];
  assign o[22545] = i[22545];
  assign o[22544] = i[22544];
  assign o[22543] = i[22543];
  assign o[22542] = i[22542];
  assign o[22541] = i[22541];
  assign o[22540] = i[22540];
  assign o[22539] = i[22539];
  assign o[22538] = i[22538];
  assign o[22537] = i[22537];
  assign o[22536] = i[22536];
  assign o[22535] = i[22535];
  assign o[22534] = i[22534];
  assign o[22533] = i[22533];
  assign o[22532] = i[22532];
  assign o[22531] = i[22531];
  assign o[22530] = i[22530];
  assign o[22529] = i[22529];
  assign o[22528] = i[22528];
  assign o[22527] = i[22527];
  assign o[22526] = i[22526];
  assign o[22525] = i[22525];
  assign o[22524] = i[22524];
  assign o[22523] = i[22523];
  assign o[22522] = i[22522];
  assign o[22521] = i[22521];
  assign o[22520] = i[22520];
  assign o[22519] = i[22519];
  assign o[22518] = i[22518];
  assign o[22517] = i[22517];
  assign o[22516] = i[22516];
  assign o[22515] = i[22515];
  assign o[22514] = i[22514];
  assign o[22513] = i[22513];
  assign o[22512] = i[22512];
  assign o[22511] = i[22511];
  assign o[22510] = i[22510];
  assign o[22509] = i[22509];
  assign o[22508] = i[22508];
  assign o[22507] = i[22507];
  assign o[22506] = i[22506];
  assign o[22505] = i[22505];
  assign o[22504] = i[22504];
  assign o[22503] = i[22503];
  assign o[22502] = i[22502];
  assign o[22501] = i[22501];
  assign o[22500] = i[22500];
  assign o[22499] = i[22499];
  assign o[22498] = i[22498];
  assign o[22497] = i[22497];
  assign o[22496] = i[22496];
  assign o[22495] = i[22495];
  assign o[22494] = i[22494];
  assign o[22493] = i[22493];
  assign o[22492] = i[22492];
  assign o[22491] = i[22491];
  assign o[22490] = i[22490];
  assign o[22489] = i[22489];
  assign o[22488] = i[22488];
  assign o[22487] = i[22487];
  assign o[22486] = i[22486];
  assign o[22485] = i[22485];
  assign o[22484] = i[22484];
  assign o[22483] = i[22483];
  assign o[22482] = i[22482];
  assign o[22481] = i[22481];
  assign o[22480] = i[22480];
  assign o[22479] = i[22479];
  assign o[22478] = i[22478];
  assign o[22477] = i[22477];
  assign o[22476] = i[22476];
  assign o[22475] = i[22475];
  assign o[22474] = i[22474];
  assign o[22473] = i[22473];
  assign o[22472] = i[22472];
  assign o[22471] = i[22471];
  assign o[22470] = i[22470];
  assign o[22469] = i[22469];
  assign o[22468] = i[22468];
  assign o[22467] = i[22467];
  assign o[22466] = i[22466];
  assign o[22465] = i[22465];
  assign o[22464] = i[22464];
  assign o[22463] = i[22463];
  assign o[22462] = i[22462];
  assign o[22461] = i[22461];
  assign o[22460] = i[22460];
  assign o[22459] = i[22459];
  assign o[22458] = i[22458];
  assign o[22457] = i[22457];
  assign o[22456] = i[22456];
  assign o[22455] = i[22455];
  assign o[22454] = i[22454];
  assign o[22453] = i[22453];
  assign o[22452] = i[22452];
  assign o[22451] = i[22451];
  assign o[22450] = i[22450];
  assign o[22449] = i[22449];
  assign o[22448] = i[22448];
  assign o[22447] = i[22447];
  assign o[22446] = i[22446];
  assign o[22445] = i[22445];
  assign o[22444] = i[22444];
  assign o[22443] = i[22443];
  assign o[22442] = i[22442];
  assign o[22441] = i[22441];
  assign o[22440] = i[22440];
  assign o[22439] = i[22439];
  assign o[22438] = i[22438];
  assign o[22437] = i[22437];
  assign o[22436] = i[22436];
  assign o[22435] = i[22435];
  assign o[22434] = i[22434];
  assign o[22433] = i[22433];
  assign o[22432] = i[22432];
  assign o[22431] = i[22431];
  assign o[22430] = i[22430];
  assign o[22429] = i[22429];
  assign o[22428] = i[22428];
  assign o[22427] = i[22427];
  assign o[22426] = i[22426];
  assign o[22425] = i[22425];
  assign o[22424] = i[22424];
  assign o[22423] = i[22423];
  assign o[22422] = i[22422];
  assign o[22421] = i[22421];
  assign o[22420] = i[22420];
  assign o[22419] = i[22419];
  assign o[22418] = i[22418];
  assign o[22417] = i[22417];
  assign o[22416] = i[22416];
  assign o[22415] = i[22415];
  assign o[22414] = i[22414];
  assign o[22413] = i[22413];
  assign o[22412] = i[22412];
  assign o[22411] = i[22411];
  assign o[22410] = i[22410];
  assign o[22409] = i[22409];
  assign o[22408] = i[22408];
  assign o[22407] = i[22407];
  assign o[22406] = i[22406];
  assign o[22405] = i[22405];
  assign o[22404] = i[22404];
  assign o[22403] = i[22403];
  assign o[22402] = i[22402];
  assign o[22401] = i[22401];
  assign o[22400] = i[22400];
  assign o[22399] = i[22399];
  assign o[22398] = i[22398];
  assign o[22397] = i[22397];
  assign o[22396] = i[22396];
  assign o[22395] = i[22395];
  assign o[22394] = i[22394];
  assign o[22393] = i[22393];
  assign o[22392] = i[22392];
  assign o[22391] = i[22391];
  assign o[22390] = i[22390];
  assign o[22389] = i[22389];
  assign o[22388] = i[22388];
  assign o[22387] = i[22387];
  assign o[22386] = i[22386];
  assign o[22385] = i[22385];
  assign o[22384] = i[22384];
  assign o[22383] = i[22383];
  assign o[22382] = i[22382];
  assign o[22381] = i[22381];
  assign o[22380] = i[22380];
  assign o[22379] = i[22379];
  assign o[22378] = i[22378];
  assign o[22377] = i[22377];
  assign o[22376] = i[22376];
  assign o[22375] = i[22375];
  assign o[22374] = i[22374];
  assign o[22373] = i[22373];
  assign o[22372] = i[22372];
  assign o[22371] = i[22371];
  assign o[22370] = i[22370];
  assign o[22369] = i[22369];
  assign o[22368] = i[22368];
  assign o[22367] = i[22367];
  assign o[22366] = i[22366];
  assign o[22365] = i[22365];
  assign o[22364] = i[22364];
  assign o[22363] = i[22363];
  assign o[22362] = i[22362];
  assign o[22361] = i[22361];
  assign o[22360] = i[22360];
  assign o[22359] = i[22359];
  assign o[22358] = i[22358];
  assign o[22357] = i[22357];
  assign o[22356] = i[22356];
  assign o[22355] = i[22355];
  assign o[22354] = i[22354];
  assign o[22353] = i[22353];
  assign o[22352] = i[22352];
  assign o[22351] = i[22351];
  assign o[22350] = i[22350];
  assign o[22349] = i[22349];
  assign o[22348] = i[22348];
  assign o[22347] = i[22347];
  assign o[22346] = i[22346];
  assign o[22345] = i[22345];
  assign o[22344] = i[22344];
  assign o[22343] = i[22343];
  assign o[22342] = i[22342];
  assign o[22341] = i[22341];
  assign o[22340] = i[22340];
  assign o[22339] = i[22339];
  assign o[22338] = i[22338];
  assign o[22337] = i[22337];
  assign o[22336] = i[22336];
  assign o[22335] = i[22335];
  assign o[22334] = i[22334];
  assign o[22333] = i[22333];
  assign o[22332] = i[22332];
  assign o[22331] = i[22331];
  assign o[22330] = i[22330];
  assign o[22329] = i[22329];
  assign o[22328] = i[22328];
  assign o[22327] = i[22327];
  assign o[22326] = i[22326];
  assign o[22325] = i[22325];
  assign o[22324] = i[22324];
  assign o[22323] = i[22323];
  assign o[22322] = i[22322];
  assign o[22321] = i[22321];
  assign o[22320] = i[22320];
  assign o[22319] = i[22319];
  assign o[22318] = i[22318];
  assign o[22317] = i[22317];
  assign o[22316] = i[22316];
  assign o[22315] = i[22315];
  assign o[22314] = i[22314];
  assign o[22313] = i[22313];
  assign o[22312] = i[22312];
  assign o[22311] = i[22311];
  assign o[22310] = i[22310];
  assign o[22309] = i[22309];
  assign o[22308] = i[22308];
  assign o[22307] = i[22307];
  assign o[22306] = i[22306];
  assign o[22305] = i[22305];
  assign o[22304] = i[22304];
  assign o[22303] = i[22303];
  assign o[22302] = i[22302];
  assign o[22301] = i[22301];
  assign o[22300] = i[22300];
  assign o[22299] = i[22299];
  assign o[22298] = i[22298];
  assign o[22297] = i[22297];
  assign o[22296] = i[22296];
  assign o[22295] = i[22295];
  assign o[22294] = i[22294];
  assign o[22293] = i[22293];
  assign o[22292] = i[22292];
  assign o[22291] = i[22291];
  assign o[22290] = i[22290];
  assign o[22289] = i[22289];
  assign o[22288] = i[22288];
  assign o[22287] = i[22287];
  assign o[22286] = i[22286];
  assign o[22285] = i[22285];
  assign o[22284] = i[22284];
  assign o[22283] = i[22283];
  assign o[22282] = i[22282];
  assign o[22281] = i[22281];
  assign o[22280] = i[22280];
  assign o[22279] = i[22279];
  assign o[22278] = i[22278];
  assign o[22277] = i[22277];
  assign o[22276] = i[22276];
  assign o[22275] = i[22275];
  assign o[22274] = i[22274];
  assign o[22273] = i[22273];
  assign o[22272] = i[22272];
  assign o[22271] = i[22271];
  assign o[22270] = i[22270];
  assign o[22269] = i[22269];
  assign o[22268] = i[22268];
  assign o[22267] = i[22267];
  assign o[22266] = i[22266];
  assign o[22265] = i[22265];
  assign o[22264] = i[22264];
  assign o[22263] = i[22263];
  assign o[22262] = i[22262];
  assign o[22261] = i[22261];
  assign o[22260] = i[22260];
  assign o[22259] = i[22259];
  assign o[22258] = i[22258];
  assign o[22257] = i[22257];
  assign o[22256] = i[22256];
  assign o[22255] = i[22255];
  assign o[22254] = i[22254];
  assign o[22253] = i[22253];
  assign o[22252] = i[22252];
  assign o[22251] = i[22251];
  assign o[22250] = i[22250];
  assign o[22249] = i[22249];
  assign o[22248] = i[22248];
  assign o[22247] = i[22247];
  assign o[22246] = i[22246];
  assign o[22245] = i[22245];
  assign o[22244] = i[22244];
  assign o[22243] = i[22243];
  assign o[22242] = i[22242];
  assign o[22241] = i[22241];
  assign o[22240] = i[22240];
  assign o[22239] = i[22239];
  assign o[22238] = i[22238];
  assign o[22237] = i[22237];
  assign o[22236] = i[22236];
  assign o[22235] = i[22235];
  assign o[22234] = i[22234];
  assign o[22233] = i[22233];
  assign o[22232] = i[22232];
  assign o[22231] = i[22231];
  assign o[22230] = i[22230];
  assign o[22229] = i[22229];
  assign o[22228] = i[22228];
  assign o[22227] = i[22227];
  assign o[22226] = i[22226];
  assign o[22225] = i[22225];
  assign o[22224] = i[22224];
  assign o[22223] = i[22223];
  assign o[22222] = i[22222];
  assign o[22221] = i[22221];
  assign o[22220] = i[22220];
  assign o[22219] = i[22219];
  assign o[22218] = i[22218];
  assign o[22217] = i[22217];
  assign o[22216] = i[22216];
  assign o[22215] = i[22215];
  assign o[22214] = i[22214];
  assign o[22213] = i[22213];
  assign o[22212] = i[22212];
  assign o[22211] = i[22211];
  assign o[22210] = i[22210];
  assign o[22209] = i[22209];
  assign o[22208] = i[22208];
  assign o[22207] = i[22207];
  assign o[22206] = i[22206];
  assign o[22205] = i[22205];
  assign o[22204] = i[22204];
  assign o[22203] = i[22203];
  assign o[22202] = i[22202];
  assign o[22201] = i[22201];
  assign o[22200] = i[22200];
  assign o[22199] = i[22199];
  assign o[22198] = i[22198];
  assign o[22197] = i[22197];
  assign o[22196] = i[22196];
  assign o[22195] = i[22195];
  assign o[22194] = i[22194];
  assign o[22193] = i[22193];
  assign o[22192] = i[22192];
  assign o[22191] = i[22191];
  assign o[22190] = i[22190];
  assign o[22189] = i[22189];
  assign o[22188] = i[22188];
  assign o[22187] = i[22187];
  assign o[22186] = i[22186];
  assign o[22185] = i[22185];
  assign o[22184] = i[22184];
  assign o[22183] = i[22183];
  assign o[22182] = i[22182];
  assign o[22181] = i[22181];
  assign o[22180] = i[22180];
  assign o[22179] = i[22179];
  assign o[22178] = i[22178];
  assign o[22177] = i[22177];
  assign o[22176] = i[22176];
  assign o[22175] = i[22175];
  assign o[22174] = i[22174];
  assign o[22173] = i[22173];
  assign o[22172] = i[22172];
  assign o[22171] = i[22171];
  assign o[22170] = i[22170];
  assign o[22169] = i[22169];
  assign o[22168] = i[22168];
  assign o[22167] = i[22167];
  assign o[22166] = i[22166];
  assign o[22165] = i[22165];
  assign o[22164] = i[22164];
  assign o[22163] = i[22163];
  assign o[22162] = i[22162];
  assign o[22161] = i[22161];
  assign o[22160] = i[22160];
  assign o[22159] = i[22159];
  assign o[22158] = i[22158];
  assign o[22157] = i[22157];
  assign o[22156] = i[22156];
  assign o[22155] = i[22155];
  assign o[22154] = i[22154];
  assign o[22153] = i[22153];
  assign o[22152] = i[22152];
  assign o[22151] = i[22151];
  assign o[22150] = i[22150];
  assign o[22149] = i[22149];
  assign o[22148] = i[22148];
  assign o[22147] = i[22147];
  assign o[22146] = i[22146];
  assign o[22145] = i[22145];
  assign o[22144] = i[22144];
  assign o[22143] = i[22143];
  assign o[22142] = i[22142];
  assign o[22141] = i[22141];
  assign o[22140] = i[22140];
  assign o[22139] = i[22139];
  assign o[22138] = i[22138];
  assign o[22137] = i[22137];
  assign o[22136] = i[22136];
  assign o[22135] = i[22135];
  assign o[22134] = i[22134];
  assign o[22133] = i[22133];
  assign o[22132] = i[22132];
  assign o[22131] = i[22131];
  assign o[22130] = i[22130];
  assign o[22129] = i[22129];
  assign o[22128] = i[22128];
  assign o[22127] = i[22127];
  assign o[22126] = i[22126];
  assign o[22125] = i[22125];
  assign o[22124] = i[22124];
  assign o[22123] = i[22123];
  assign o[22122] = i[22122];
  assign o[22121] = i[22121];
  assign o[22120] = i[22120];
  assign o[22119] = i[22119];
  assign o[22118] = i[22118];
  assign o[22117] = i[22117];
  assign o[22116] = i[22116];
  assign o[22115] = i[22115];
  assign o[22114] = i[22114];
  assign o[22113] = i[22113];
  assign o[22112] = i[22112];
  assign o[22111] = i[22111];
  assign o[22110] = i[22110];
  assign o[22109] = i[22109];
  assign o[22108] = i[22108];
  assign o[22107] = i[22107];
  assign o[22106] = i[22106];
  assign o[22105] = i[22105];
  assign o[22104] = i[22104];
  assign o[22103] = i[22103];
  assign o[22102] = i[22102];
  assign o[22101] = i[22101];
  assign o[22100] = i[22100];
  assign o[22099] = i[22099];
  assign o[22098] = i[22098];
  assign o[22097] = i[22097];
  assign o[22096] = i[22096];
  assign o[22095] = i[22095];
  assign o[22094] = i[22094];
  assign o[22093] = i[22093];
  assign o[22092] = i[22092];
  assign o[22091] = i[22091];
  assign o[22090] = i[22090];
  assign o[22089] = i[22089];
  assign o[22088] = i[22088];
  assign o[22087] = i[22087];
  assign o[22086] = i[22086];
  assign o[22085] = i[22085];
  assign o[22084] = i[22084];
  assign o[22083] = i[22083];
  assign o[22082] = i[22082];
  assign o[22081] = i[22081];
  assign o[22080] = i[22080];
  assign o[22079] = i[22079];
  assign o[22078] = i[22078];
  assign o[22077] = i[22077];
  assign o[22076] = i[22076];
  assign o[22075] = i[22075];
  assign o[22074] = i[22074];
  assign o[22073] = i[22073];
  assign o[22072] = i[22072];
  assign o[22071] = i[22071];
  assign o[22070] = i[22070];
  assign o[22069] = i[22069];
  assign o[22068] = i[22068];
  assign o[22067] = i[22067];
  assign o[22066] = i[22066];
  assign o[22065] = i[22065];
  assign o[22064] = i[22064];
  assign o[22063] = i[22063];
  assign o[22062] = i[22062];
  assign o[22061] = i[22061];
  assign o[22060] = i[22060];
  assign o[22059] = i[22059];
  assign o[22058] = i[22058];
  assign o[22057] = i[22057];
  assign o[22056] = i[22056];
  assign o[22055] = i[22055];
  assign o[22054] = i[22054];
  assign o[22053] = i[22053];
  assign o[22052] = i[22052];
  assign o[22051] = i[22051];
  assign o[22050] = i[22050];
  assign o[22049] = i[22049];
  assign o[22048] = i[22048];
  assign o[22047] = i[22047];
  assign o[22046] = i[22046];
  assign o[22045] = i[22045];
  assign o[22044] = i[22044];
  assign o[22043] = i[22043];
  assign o[22042] = i[22042];
  assign o[22041] = i[22041];
  assign o[22040] = i[22040];
  assign o[22039] = i[22039];
  assign o[22038] = i[22038];
  assign o[22037] = i[22037];
  assign o[22036] = i[22036];
  assign o[22035] = i[22035];
  assign o[22034] = i[22034];
  assign o[22033] = i[22033];
  assign o[22032] = i[22032];
  assign o[22031] = i[22031];
  assign o[22030] = i[22030];
  assign o[22029] = i[22029];
  assign o[22028] = i[22028];
  assign o[22027] = i[22027];
  assign o[22026] = i[22026];
  assign o[22025] = i[22025];
  assign o[22024] = i[22024];
  assign o[22023] = i[22023];
  assign o[22022] = i[22022];
  assign o[22021] = i[22021];
  assign o[22020] = i[22020];
  assign o[22019] = i[22019];
  assign o[22018] = i[22018];
  assign o[22017] = i[22017];
  assign o[22016] = i[22016];
  assign o[22015] = i[22015];
  assign o[22014] = i[22014];
  assign o[22013] = i[22013];
  assign o[22012] = i[22012];
  assign o[22011] = i[22011];
  assign o[22010] = i[22010];
  assign o[22009] = i[22009];
  assign o[22008] = i[22008];
  assign o[22007] = i[22007];
  assign o[22006] = i[22006];
  assign o[22005] = i[22005];
  assign o[22004] = i[22004];
  assign o[22003] = i[22003];
  assign o[22002] = i[22002];
  assign o[22001] = i[22001];
  assign o[22000] = i[22000];
  assign o[21999] = i[21999];
  assign o[21998] = i[21998];
  assign o[21997] = i[21997];
  assign o[21996] = i[21996];
  assign o[21995] = i[21995];
  assign o[21994] = i[21994];
  assign o[21993] = i[21993];
  assign o[21992] = i[21992];
  assign o[21991] = i[21991];
  assign o[21990] = i[21990];
  assign o[21989] = i[21989];
  assign o[21988] = i[21988];
  assign o[21987] = i[21987];
  assign o[21986] = i[21986];
  assign o[21985] = i[21985];
  assign o[21984] = i[21984];
  assign o[21983] = i[21983];
  assign o[21982] = i[21982];
  assign o[21981] = i[21981];
  assign o[21980] = i[21980];
  assign o[21979] = i[21979];
  assign o[21978] = i[21978];
  assign o[21977] = i[21977];
  assign o[21976] = i[21976];
  assign o[21975] = i[21975];
  assign o[21974] = i[21974];
  assign o[21973] = i[21973];
  assign o[21972] = i[21972];
  assign o[21971] = i[21971];
  assign o[21970] = i[21970];
  assign o[21969] = i[21969];
  assign o[21968] = i[21968];
  assign o[21967] = i[21967];
  assign o[21966] = i[21966];
  assign o[21965] = i[21965];
  assign o[21964] = i[21964];
  assign o[21963] = i[21963];
  assign o[21962] = i[21962];
  assign o[21961] = i[21961];
  assign o[21960] = i[21960];
  assign o[21959] = i[21959];
  assign o[21958] = i[21958];
  assign o[21957] = i[21957];
  assign o[21956] = i[21956];
  assign o[21955] = i[21955];
  assign o[21954] = i[21954];
  assign o[21953] = i[21953];
  assign o[21952] = i[21952];
  assign o[21951] = i[21951];
  assign o[21950] = i[21950];
  assign o[21949] = i[21949];
  assign o[21948] = i[21948];
  assign o[21947] = i[21947];
  assign o[21946] = i[21946];
  assign o[21945] = i[21945];
  assign o[21944] = i[21944];
  assign o[21943] = i[21943];
  assign o[21942] = i[21942];
  assign o[21941] = i[21941];
  assign o[21940] = i[21940];
  assign o[21939] = i[21939];
  assign o[21938] = i[21938];
  assign o[21937] = i[21937];
  assign o[21936] = i[21936];
  assign o[21935] = i[21935];
  assign o[21934] = i[21934];
  assign o[21933] = i[21933];
  assign o[21932] = i[21932];
  assign o[21931] = i[21931];
  assign o[21930] = i[21930];
  assign o[21929] = i[21929];
  assign o[21928] = i[21928];
  assign o[21927] = i[21927];
  assign o[21926] = i[21926];
  assign o[21925] = i[21925];
  assign o[21924] = i[21924];
  assign o[21923] = i[21923];
  assign o[21922] = i[21922];
  assign o[21921] = i[21921];
  assign o[21920] = i[21920];
  assign o[21919] = i[21919];
  assign o[21918] = i[21918];
  assign o[21917] = i[21917];
  assign o[21916] = i[21916];
  assign o[21915] = i[21915];
  assign o[21914] = i[21914];
  assign o[21913] = i[21913];
  assign o[21912] = i[21912];
  assign o[21911] = i[21911];
  assign o[21910] = i[21910];
  assign o[21909] = i[21909];
  assign o[21908] = i[21908];
  assign o[21907] = i[21907];
  assign o[21906] = i[21906];
  assign o[21905] = i[21905];
  assign o[21904] = i[21904];
  assign o[21903] = i[21903];
  assign o[21902] = i[21902];
  assign o[21901] = i[21901];
  assign o[21900] = i[21900];
  assign o[21899] = i[21899];
  assign o[21898] = i[21898];
  assign o[21897] = i[21897];
  assign o[21896] = i[21896];
  assign o[21895] = i[21895];
  assign o[21894] = i[21894];
  assign o[21893] = i[21893];
  assign o[21892] = i[21892];
  assign o[21891] = i[21891];
  assign o[21890] = i[21890];
  assign o[21889] = i[21889];
  assign o[21888] = i[21888];
  assign o[21887] = i[21887];
  assign o[21886] = i[21886];
  assign o[21885] = i[21885];
  assign o[21884] = i[21884];
  assign o[21883] = i[21883];
  assign o[21882] = i[21882];
  assign o[21881] = i[21881];
  assign o[21880] = i[21880];
  assign o[21879] = i[21879];
  assign o[21878] = i[21878];
  assign o[21877] = i[21877];
  assign o[21876] = i[21876];
  assign o[21875] = i[21875];
  assign o[21874] = i[21874];
  assign o[21873] = i[21873];
  assign o[21872] = i[21872];
  assign o[21871] = i[21871];
  assign o[21870] = i[21870];
  assign o[21869] = i[21869];
  assign o[21868] = i[21868];
  assign o[21867] = i[21867];
  assign o[21866] = i[21866];
  assign o[21865] = i[21865];
  assign o[21864] = i[21864];
  assign o[21863] = i[21863];
  assign o[21862] = i[21862];
  assign o[21861] = i[21861];
  assign o[21860] = i[21860];
  assign o[21859] = i[21859];
  assign o[21858] = i[21858];
  assign o[21857] = i[21857];
  assign o[21856] = i[21856];
  assign o[21855] = i[21855];
  assign o[21854] = i[21854];
  assign o[21853] = i[21853];
  assign o[21852] = i[21852];
  assign o[21851] = i[21851];
  assign o[21850] = i[21850];
  assign o[21849] = i[21849];
  assign o[21848] = i[21848];
  assign o[21847] = i[21847];
  assign o[21846] = i[21846];
  assign o[21845] = i[21845];
  assign o[21844] = i[21844];
  assign o[21843] = i[21843];
  assign o[21842] = i[21842];
  assign o[21841] = i[21841];
  assign o[21840] = i[21840];
  assign o[21839] = i[21839];
  assign o[21838] = i[21838];
  assign o[21837] = i[21837];
  assign o[21836] = i[21836];
  assign o[21835] = i[21835];
  assign o[21834] = i[21834];
  assign o[21833] = i[21833];
  assign o[21832] = i[21832];
  assign o[21831] = i[21831];
  assign o[21830] = i[21830];
  assign o[21829] = i[21829];
  assign o[21828] = i[21828];
  assign o[21827] = i[21827];
  assign o[21826] = i[21826];
  assign o[21825] = i[21825];
  assign o[21824] = i[21824];
  assign o[21823] = i[21823];
  assign o[21822] = i[21822];
  assign o[21821] = i[21821];
  assign o[21820] = i[21820];
  assign o[21819] = i[21819];
  assign o[21818] = i[21818];
  assign o[21817] = i[21817];
  assign o[21816] = i[21816];
  assign o[21815] = i[21815];
  assign o[21814] = i[21814];
  assign o[21813] = i[21813];
  assign o[21812] = i[21812];
  assign o[21811] = i[21811];
  assign o[21810] = i[21810];
  assign o[21809] = i[21809];
  assign o[21808] = i[21808];
  assign o[21807] = i[21807];
  assign o[21806] = i[21806];
  assign o[21805] = i[21805];
  assign o[21804] = i[21804];
  assign o[21803] = i[21803];
  assign o[21802] = i[21802];
  assign o[21801] = i[21801];
  assign o[21800] = i[21800];
  assign o[21799] = i[21799];
  assign o[21798] = i[21798];
  assign o[21797] = i[21797];
  assign o[21796] = i[21796];
  assign o[21795] = i[21795];
  assign o[21794] = i[21794];
  assign o[21793] = i[21793];
  assign o[21792] = i[21792];
  assign o[21791] = i[21791];
  assign o[21790] = i[21790];
  assign o[21789] = i[21789];
  assign o[21788] = i[21788];
  assign o[21787] = i[21787];
  assign o[21786] = i[21786];
  assign o[21785] = i[21785];
  assign o[21784] = i[21784];
  assign o[21783] = i[21783];
  assign o[21782] = i[21782];
  assign o[21781] = i[21781];
  assign o[21780] = i[21780];
  assign o[21779] = i[21779];
  assign o[21778] = i[21778];
  assign o[21777] = i[21777];
  assign o[21776] = i[21776];
  assign o[21775] = i[21775];
  assign o[21774] = i[21774];
  assign o[21773] = i[21773];
  assign o[21772] = i[21772];
  assign o[21771] = i[21771];
  assign o[21770] = i[21770];
  assign o[21769] = i[21769];
  assign o[21768] = i[21768];
  assign o[21767] = i[21767];
  assign o[21766] = i[21766];
  assign o[21765] = i[21765];
  assign o[21764] = i[21764];
  assign o[21763] = i[21763];
  assign o[21762] = i[21762];
  assign o[21761] = i[21761];
  assign o[21760] = i[21760];
  assign o[21759] = i[21759];
  assign o[21758] = i[21758];
  assign o[21757] = i[21757];
  assign o[21756] = i[21756];
  assign o[21755] = i[21755];
  assign o[21754] = i[21754];
  assign o[21753] = i[21753];
  assign o[21752] = i[21752];
  assign o[21751] = i[21751];
  assign o[21750] = i[21750];
  assign o[21749] = i[21749];
  assign o[21748] = i[21748];
  assign o[21747] = i[21747];
  assign o[21746] = i[21746];
  assign o[21745] = i[21745];
  assign o[21744] = i[21744];
  assign o[21743] = i[21743];
  assign o[21742] = i[21742];
  assign o[21741] = i[21741];
  assign o[21740] = i[21740];
  assign o[21739] = i[21739];
  assign o[21738] = i[21738];
  assign o[21737] = i[21737];
  assign o[21736] = i[21736];
  assign o[21735] = i[21735];
  assign o[21734] = i[21734];
  assign o[21733] = i[21733];
  assign o[21732] = i[21732];
  assign o[21731] = i[21731];
  assign o[21730] = i[21730];
  assign o[21729] = i[21729];
  assign o[21728] = i[21728];
  assign o[21727] = i[21727];
  assign o[21726] = i[21726];
  assign o[21725] = i[21725];
  assign o[21724] = i[21724];
  assign o[21723] = i[21723];
  assign o[21722] = i[21722];
  assign o[21721] = i[21721];
  assign o[21720] = i[21720];
  assign o[21719] = i[21719];
  assign o[21718] = i[21718];
  assign o[21717] = i[21717];
  assign o[21716] = i[21716];
  assign o[21715] = i[21715];
  assign o[21714] = i[21714];
  assign o[21713] = i[21713];
  assign o[21712] = i[21712];
  assign o[21711] = i[21711];
  assign o[21710] = i[21710];
  assign o[21709] = i[21709];
  assign o[21708] = i[21708];
  assign o[21707] = i[21707];
  assign o[21706] = i[21706];
  assign o[21705] = i[21705];
  assign o[21704] = i[21704];
  assign o[21703] = i[21703];
  assign o[21702] = i[21702];
  assign o[21701] = i[21701];
  assign o[21700] = i[21700];
  assign o[21699] = i[21699];
  assign o[21698] = i[21698];
  assign o[21697] = i[21697];
  assign o[21696] = i[21696];
  assign o[21695] = i[21695];
  assign o[21694] = i[21694];
  assign o[21693] = i[21693];
  assign o[21692] = i[21692];
  assign o[21691] = i[21691];
  assign o[21690] = i[21690];
  assign o[21689] = i[21689];
  assign o[21688] = i[21688];
  assign o[21687] = i[21687];
  assign o[21686] = i[21686];
  assign o[21685] = i[21685];
  assign o[21684] = i[21684];
  assign o[21683] = i[21683];
  assign o[21682] = i[21682];
  assign o[21681] = i[21681];
  assign o[21680] = i[21680];
  assign o[21679] = i[21679];
  assign o[21678] = i[21678];
  assign o[21677] = i[21677];
  assign o[21676] = i[21676];
  assign o[21675] = i[21675];
  assign o[21674] = i[21674];
  assign o[21673] = i[21673];
  assign o[21672] = i[21672];
  assign o[21671] = i[21671];
  assign o[21670] = i[21670];
  assign o[21669] = i[21669];
  assign o[21668] = i[21668];
  assign o[21667] = i[21667];
  assign o[21666] = i[21666];
  assign o[21665] = i[21665];
  assign o[21664] = i[21664];
  assign o[21663] = i[21663];
  assign o[21662] = i[21662];
  assign o[21661] = i[21661];
  assign o[21660] = i[21660];
  assign o[21659] = i[21659];
  assign o[21658] = i[21658];
  assign o[21657] = i[21657];
  assign o[21656] = i[21656];
  assign o[21655] = i[21655];
  assign o[21654] = i[21654];
  assign o[21653] = i[21653];
  assign o[21652] = i[21652];
  assign o[21651] = i[21651];
  assign o[21650] = i[21650];
  assign o[21649] = i[21649];
  assign o[21648] = i[21648];
  assign o[21647] = i[21647];
  assign o[21646] = i[21646];
  assign o[21645] = i[21645];
  assign o[21644] = i[21644];
  assign o[21643] = i[21643];
  assign o[21642] = i[21642];
  assign o[21641] = i[21641];
  assign o[21640] = i[21640];
  assign o[21639] = i[21639];
  assign o[21638] = i[21638];
  assign o[21637] = i[21637];
  assign o[21636] = i[21636];
  assign o[21635] = i[21635];
  assign o[21634] = i[21634];
  assign o[21633] = i[21633];
  assign o[21632] = i[21632];
  assign o[21631] = i[21631];
  assign o[21630] = i[21630];
  assign o[21629] = i[21629];
  assign o[21628] = i[21628];
  assign o[21627] = i[21627];
  assign o[21626] = i[21626];
  assign o[21625] = i[21625];
  assign o[21624] = i[21624];
  assign o[21623] = i[21623];
  assign o[21622] = i[21622];
  assign o[21621] = i[21621];
  assign o[21620] = i[21620];
  assign o[21619] = i[21619];
  assign o[21618] = i[21618];
  assign o[21617] = i[21617];
  assign o[21616] = i[21616];
  assign o[21615] = i[21615];
  assign o[21614] = i[21614];
  assign o[21613] = i[21613];
  assign o[21612] = i[21612];
  assign o[21611] = i[21611];
  assign o[21610] = i[21610];
  assign o[21609] = i[21609];
  assign o[21608] = i[21608];
  assign o[21607] = i[21607];
  assign o[21606] = i[21606];
  assign o[21605] = i[21605];
  assign o[21604] = i[21604];
  assign o[21603] = i[21603];
  assign o[21602] = i[21602];
  assign o[21601] = i[21601];
  assign o[21600] = i[21600];
  assign o[21599] = i[21599];
  assign o[21598] = i[21598];
  assign o[21597] = i[21597];
  assign o[21596] = i[21596];
  assign o[21595] = i[21595];
  assign o[21594] = i[21594];
  assign o[21593] = i[21593];
  assign o[21592] = i[21592];
  assign o[21591] = i[21591];
  assign o[21590] = i[21590];
  assign o[21589] = i[21589];
  assign o[21588] = i[21588];
  assign o[21587] = i[21587];
  assign o[21586] = i[21586];
  assign o[21585] = i[21585];
  assign o[21584] = i[21584];
  assign o[21583] = i[21583];
  assign o[21582] = i[21582];
  assign o[21581] = i[21581];
  assign o[21580] = i[21580];
  assign o[21579] = i[21579];
  assign o[21578] = i[21578];
  assign o[21577] = i[21577];
  assign o[21576] = i[21576];
  assign o[21575] = i[21575];
  assign o[21574] = i[21574];
  assign o[21573] = i[21573];
  assign o[21572] = i[21572];
  assign o[21571] = i[21571];
  assign o[21570] = i[21570];
  assign o[21569] = i[21569];
  assign o[21568] = i[21568];
  assign o[21567] = i[21567];
  assign o[21566] = i[21566];
  assign o[21565] = i[21565];
  assign o[21564] = i[21564];
  assign o[21563] = i[21563];
  assign o[21562] = i[21562];
  assign o[21561] = i[21561];
  assign o[21560] = i[21560];
  assign o[21559] = i[21559];
  assign o[21558] = i[21558];
  assign o[21557] = i[21557];
  assign o[21556] = i[21556];
  assign o[21555] = i[21555];
  assign o[21554] = i[21554];
  assign o[21553] = i[21553];
  assign o[21552] = i[21552];
  assign o[21551] = i[21551];
  assign o[21550] = i[21550];
  assign o[21549] = i[21549];
  assign o[21548] = i[21548];
  assign o[21547] = i[21547];
  assign o[21546] = i[21546];
  assign o[21545] = i[21545];
  assign o[21544] = i[21544];
  assign o[21543] = i[21543];
  assign o[21542] = i[21542];
  assign o[21541] = i[21541];
  assign o[21540] = i[21540];
  assign o[21539] = i[21539];
  assign o[21538] = i[21538];
  assign o[21537] = i[21537];
  assign o[21536] = i[21536];
  assign o[21535] = i[21535];
  assign o[21534] = i[21534];
  assign o[21533] = i[21533];
  assign o[21532] = i[21532];
  assign o[21531] = i[21531];
  assign o[21530] = i[21530];
  assign o[21529] = i[21529];
  assign o[21528] = i[21528];
  assign o[21527] = i[21527];
  assign o[21526] = i[21526];
  assign o[21525] = i[21525];
  assign o[21524] = i[21524];
  assign o[21523] = i[21523];
  assign o[21522] = i[21522];
  assign o[21521] = i[21521];
  assign o[21520] = i[21520];
  assign o[21519] = i[21519];
  assign o[21518] = i[21518];
  assign o[21517] = i[21517];
  assign o[21516] = i[21516];
  assign o[21515] = i[21515];
  assign o[21514] = i[21514];
  assign o[21513] = i[21513];
  assign o[21512] = i[21512];
  assign o[21511] = i[21511];
  assign o[21510] = i[21510];
  assign o[21509] = i[21509];
  assign o[21508] = i[21508];
  assign o[21507] = i[21507];
  assign o[21506] = i[21506];
  assign o[21505] = i[21505];
  assign o[21504] = i[21504];
  assign o[21503] = i[21503];
  assign o[21502] = i[21502];
  assign o[21501] = i[21501];
  assign o[21500] = i[21500];
  assign o[21499] = i[21499];
  assign o[21498] = i[21498];
  assign o[21497] = i[21497];
  assign o[21496] = i[21496];
  assign o[21495] = i[21495];
  assign o[21494] = i[21494];
  assign o[21493] = i[21493];
  assign o[21492] = i[21492];
  assign o[21491] = i[21491];
  assign o[21490] = i[21490];
  assign o[21489] = i[21489];
  assign o[21488] = i[21488];
  assign o[21487] = i[21487];
  assign o[21486] = i[21486];
  assign o[21485] = i[21485];
  assign o[21484] = i[21484];
  assign o[21483] = i[21483];
  assign o[21482] = i[21482];
  assign o[21481] = i[21481];
  assign o[21480] = i[21480];
  assign o[21479] = i[21479];
  assign o[21478] = i[21478];
  assign o[21477] = i[21477];
  assign o[21476] = i[21476];
  assign o[21475] = i[21475];
  assign o[21474] = i[21474];
  assign o[21473] = i[21473];
  assign o[21472] = i[21472];
  assign o[21471] = i[21471];
  assign o[21470] = i[21470];
  assign o[21469] = i[21469];
  assign o[21468] = i[21468];
  assign o[21467] = i[21467];
  assign o[21466] = i[21466];
  assign o[21465] = i[21465];
  assign o[21464] = i[21464];
  assign o[21463] = i[21463];
  assign o[21462] = i[21462];
  assign o[21461] = i[21461];
  assign o[21460] = i[21460];
  assign o[21459] = i[21459];
  assign o[21458] = i[21458];
  assign o[21457] = i[21457];
  assign o[21456] = i[21456];
  assign o[21455] = i[21455];
  assign o[21454] = i[21454];
  assign o[21453] = i[21453];
  assign o[21452] = i[21452];
  assign o[21451] = i[21451];
  assign o[21450] = i[21450];
  assign o[21449] = i[21449];
  assign o[21448] = i[21448];
  assign o[21447] = i[21447];
  assign o[21446] = i[21446];
  assign o[21445] = i[21445];
  assign o[21444] = i[21444];
  assign o[21443] = i[21443];
  assign o[21442] = i[21442];
  assign o[21441] = i[21441];
  assign o[21440] = i[21440];
  assign o[21439] = i[21439];
  assign o[21438] = i[21438];
  assign o[21437] = i[21437];
  assign o[21436] = i[21436];
  assign o[21435] = i[21435];
  assign o[21434] = i[21434];
  assign o[21433] = i[21433];
  assign o[21432] = i[21432];
  assign o[21431] = i[21431];
  assign o[21430] = i[21430];
  assign o[21429] = i[21429];
  assign o[21428] = i[21428];
  assign o[21427] = i[21427];
  assign o[21426] = i[21426];
  assign o[21425] = i[21425];
  assign o[21424] = i[21424];
  assign o[21423] = i[21423];
  assign o[21422] = i[21422];
  assign o[21421] = i[21421];
  assign o[21420] = i[21420];
  assign o[21419] = i[21419];
  assign o[21418] = i[21418];
  assign o[21417] = i[21417];
  assign o[21416] = i[21416];
  assign o[21415] = i[21415];
  assign o[21414] = i[21414];
  assign o[21413] = i[21413];
  assign o[21412] = i[21412];
  assign o[21411] = i[21411];
  assign o[21410] = i[21410];
  assign o[21409] = i[21409];
  assign o[21408] = i[21408];
  assign o[21407] = i[21407];
  assign o[21406] = i[21406];
  assign o[21405] = i[21405];
  assign o[21404] = i[21404];
  assign o[21403] = i[21403];
  assign o[21402] = i[21402];
  assign o[21401] = i[21401];
  assign o[21400] = i[21400];
  assign o[21399] = i[21399];
  assign o[21398] = i[21398];
  assign o[21397] = i[21397];
  assign o[21396] = i[21396];
  assign o[21395] = i[21395];
  assign o[21394] = i[21394];
  assign o[21393] = i[21393];
  assign o[21392] = i[21392];
  assign o[21391] = i[21391];
  assign o[21390] = i[21390];
  assign o[21389] = i[21389];
  assign o[21388] = i[21388];
  assign o[21387] = i[21387];
  assign o[21386] = i[21386];
  assign o[21385] = i[21385];
  assign o[21384] = i[21384];
  assign o[21383] = i[21383];
  assign o[21382] = i[21382];
  assign o[21381] = i[21381];
  assign o[21380] = i[21380];
  assign o[21379] = i[21379];
  assign o[21378] = i[21378];
  assign o[21377] = i[21377];
  assign o[21376] = i[21376];
  assign o[21375] = i[21375];
  assign o[21374] = i[21374];
  assign o[21373] = i[21373];
  assign o[21372] = i[21372];
  assign o[21371] = i[21371];
  assign o[21370] = i[21370];
  assign o[21369] = i[21369];
  assign o[21368] = i[21368];
  assign o[21367] = i[21367];
  assign o[21366] = i[21366];
  assign o[21365] = i[21365];
  assign o[21364] = i[21364];
  assign o[21363] = i[21363];
  assign o[21362] = i[21362];
  assign o[21361] = i[21361];
  assign o[21360] = i[21360];
  assign o[21359] = i[21359];
  assign o[21358] = i[21358];
  assign o[21357] = i[21357];
  assign o[21356] = i[21356];
  assign o[21355] = i[21355];
  assign o[21354] = i[21354];
  assign o[21353] = i[21353];
  assign o[21352] = i[21352];
  assign o[21351] = i[21351];
  assign o[21350] = i[21350];
  assign o[21349] = i[21349];
  assign o[21348] = i[21348];
  assign o[21347] = i[21347];
  assign o[21346] = i[21346];
  assign o[21345] = i[21345];
  assign o[21344] = i[21344];
  assign o[21343] = i[21343];
  assign o[21342] = i[21342];
  assign o[21341] = i[21341];
  assign o[21340] = i[21340];
  assign o[21339] = i[21339];
  assign o[21338] = i[21338];
  assign o[21337] = i[21337];
  assign o[21336] = i[21336];
  assign o[21335] = i[21335];
  assign o[21334] = i[21334];
  assign o[21333] = i[21333];
  assign o[21332] = i[21332];
  assign o[21331] = i[21331];
  assign o[21330] = i[21330];
  assign o[21329] = i[21329];
  assign o[21328] = i[21328];
  assign o[21327] = i[21327];
  assign o[21326] = i[21326];
  assign o[21325] = i[21325];
  assign o[21324] = i[21324];
  assign o[21323] = i[21323];
  assign o[21322] = i[21322];
  assign o[21321] = i[21321];
  assign o[21320] = i[21320];
  assign o[21319] = i[21319];
  assign o[21318] = i[21318];
  assign o[21317] = i[21317];
  assign o[21316] = i[21316];
  assign o[21315] = i[21315];
  assign o[21314] = i[21314];
  assign o[21313] = i[21313];
  assign o[21312] = i[21312];
  assign o[21311] = i[21311];
  assign o[21310] = i[21310];
  assign o[21309] = i[21309];
  assign o[21308] = i[21308];
  assign o[21307] = i[21307];
  assign o[21306] = i[21306];
  assign o[21305] = i[21305];
  assign o[21304] = i[21304];
  assign o[21303] = i[21303];
  assign o[21302] = i[21302];
  assign o[21301] = i[21301];
  assign o[21300] = i[21300];
  assign o[21299] = i[21299];
  assign o[21298] = i[21298];
  assign o[21297] = i[21297];
  assign o[21296] = i[21296];
  assign o[21295] = i[21295];
  assign o[21294] = i[21294];
  assign o[21293] = i[21293];
  assign o[21292] = i[21292];
  assign o[21291] = i[21291];
  assign o[21290] = i[21290];
  assign o[21289] = i[21289];
  assign o[21288] = i[21288];
  assign o[21287] = i[21287];
  assign o[21286] = i[21286];
  assign o[21285] = i[21285];
  assign o[21284] = i[21284];
  assign o[21283] = i[21283];
  assign o[21282] = i[21282];
  assign o[21281] = i[21281];
  assign o[21280] = i[21280];
  assign o[21279] = i[21279];
  assign o[21278] = i[21278];
  assign o[21277] = i[21277];
  assign o[21276] = i[21276];
  assign o[21275] = i[21275];
  assign o[21274] = i[21274];
  assign o[21273] = i[21273];
  assign o[21272] = i[21272];
  assign o[21271] = i[21271];
  assign o[21270] = i[21270];
  assign o[21269] = i[21269];
  assign o[21268] = i[21268];
  assign o[21267] = i[21267];
  assign o[21266] = i[21266];
  assign o[21265] = i[21265];
  assign o[21264] = i[21264];
  assign o[21263] = i[21263];
  assign o[21262] = i[21262];
  assign o[21261] = i[21261];
  assign o[21260] = i[21260];
  assign o[21259] = i[21259];
  assign o[21258] = i[21258];
  assign o[21257] = i[21257];
  assign o[21256] = i[21256];
  assign o[21255] = i[21255];
  assign o[21254] = i[21254];
  assign o[21253] = i[21253];
  assign o[21252] = i[21252];
  assign o[21251] = i[21251];
  assign o[21250] = i[21250];
  assign o[21249] = i[21249];
  assign o[21248] = i[21248];
  assign o[21247] = i[21247];
  assign o[21246] = i[21246];
  assign o[21245] = i[21245];
  assign o[21244] = i[21244];
  assign o[21243] = i[21243];
  assign o[21242] = i[21242];
  assign o[21241] = i[21241];
  assign o[21240] = i[21240];
  assign o[21239] = i[21239];
  assign o[21238] = i[21238];
  assign o[21237] = i[21237];
  assign o[21236] = i[21236];
  assign o[21235] = i[21235];
  assign o[21234] = i[21234];
  assign o[21233] = i[21233];
  assign o[21232] = i[21232];
  assign o[21231] = i[21231];
  assign o[21230] = i[21230];
  assign o[21229] = i[21229];
  assign o[21228] = i[21228];
  assign o[21227] = i[21227];
  assign o[21226] = i[21226];
  assign o[21225] = i[21225];
  assign o[21224] = i[21224];
  assign o[21223] = i[21223];
  assign o[21222] = i[21222];
  assign o[21221] = i[21221];
  assign o[21220] = i[21220];
  assign o[21219] = i[21219];
  assign o[21218] = i[21218];
  assign o[21217] = i[21217];
  assign o[21216] = i[21216];
  assign o[21215] = i[21215];
  assign o[21214] = i[21214];
  assign o[21213] = i[21213];
  assign o[21212] = i[21212];
  assign o[21211] = i[21211];
  assign o[21210] = i[21210];
  assign o[21209] = i[21209];
  assign o[21208] = i[21208];
  assign o[21207] = i[21207];
  assign o[21206] = i[21206];
  assign o[21205] = i[21205];
  assign o[21204] = i[21204];
  assign o[21203] = i[21203];
  assign o[21202] = i[21202];
  assign o[21201] = i[21201];
  assign o[21200] = i[21200];
  assign o[21199] = i[21199];
  assign o[21198] = i[21198];
  assign o[21197] = i[21197];
  assign o[21196] = i[21196];
  assign o[21195] = i[21195];
  assign o[21194] = i[21194];
  assign o[21193] = i[21193];
  assign o[21192] = i[21192];
  assign o[21191] = i[21191];
  assign o[21190] = i[21190];
  assign o[21189] = i[21189];
  assign o[21188] = i[21188];
  assign o[21187] = i[21187];
  assign o[21186] = i[21186];
  assign o[21185] = i[21185];
  assign o[21184] = i[21184];
  assign o[21183] = i[21183];
  assign o[21182] = i[21182];
  assign o[21181] = i[21181];
  assign o[21180] = i[21180];
  assign o[21179] = i[21179];
  assign o[21178] = i[21178];
  assign o[21177] = i[21177];
  assign o[21176] = i[21176];
  assign o[21175] = i[21175];
  assign o[21174] = i[21174];
  assign o[21173] = i[21173];
  assign o[21172] = i[21172];
  assign o[21171] = i[21171];
  assign o[21170] = i[21170];
  assign o[21169] = i[21169];
  assign o[21168] = i[21168];
  assign o[21167] = i[21167];
  assign o[21166] = i[21166];
  assign o[21165] = i[21165];
  assign o[21164] = i[21164];
  assign o[21163] = i[21163];
  assign o[21162] = i[21162];
  assign o[21161] = i[21161];
  assign o[21160] = i[21160];
  assign o[21159] = i[21159];
  assign o[21158] = i[21158];
  assign o[21157] = i[21157];
  assign o[21156] = i[21156];
  assign o[21155] = i[21155];
  assign o[21154] = i[21154];
  assign o[21153] = i[21153];
  assign o[21152] = i[21152];
  assign o[21151] = i[21151];
  assign o[21150] = i[21150];
  assign o[21149] = i[21149];
  assign o[21148] = i[21148];
  assign o[21147] = i[21147];
  assign o[21146] = i[21146];
  assign o[21145] = i[21145];
  assign o[21144] = i[21144];
  assign o[21143] = i[21143];
  assign o[21142] = i[21142];
  assign o[21141] = i[21141];
  assign o[21140] = i[21140];
  assign o[21139] = i[21139];
  assign o[21138] = i[21138];
  assign o[21137] = i[21137];
  assign o[21136] = i[21136];
  assign o[21135] = i[21135];
  assign o[21134] = i[21134];
  assign o[21133] = i[21133];
  assign o[21132] = i[21132];
  assign o[21131] = i[21131];
  assign o[21130] = i[21130];
  assign o[21129] = i[21129];
  assign o[21128] = i[21128];
  assign o[21127] = i[21127];
  assign o[21126] = i[21126];
  assign o[21125] = i[21125];
  assign o[21124] = i[21124];
  assign o[21123] = i[21123];
  assign o[21122] = i[21122];
  assign o[21121] = i[21121];
  assign o[21120] = i[21120];
  assign o[21119] = i[21119];
  assign o[21118] = i[21118];
  assign o[21117] = i[21117];
  assign o[21116] = i[21116];
  assign o[21115] = i[21115];
  assign o[21114] = i[21114];
  assign o[21113] = i[21113];
  assign o[21112] = i[21112];
  assign o[21111] = i[21111];
  assign o[21110] = i[21110];
  assign o[21109] = i[21109];
  assign o[21108] = i[21108];
  assign o[21107] = i[21107];
  assign o[21106] = i[21106];
  assign o[21105] = i[21105];
  assign o[21104] = i[21104];
  assign o[21103] = i[21103];
  assign o[21102] = i[21102];
  assign o[21101] = i[21101];
  assign o[21100] = i[21100];
  assign o[21099] = i[21099];
  assign o[21098] = i[21098];
  assign o[21097] = i[21097];
  assign o[21096] = i[21096];
  assign o[21095] = i[21095];
  assign o[21094] = i[21094];
  assign o[21093] = i[21093];
  assign o[21092] = i[21092];
  assign o[21091] = i[21091];
  assign o[21090] = i[21090];
  assign o[21089] = i[21089];
  assign o[21088] = i[21088];
  assign o[21087] = i[21087];
  assign o[21086] = i[21086];
  assign o[21085] = i[21085];
  assign o[21084] = i[21084];
  assign o[21083] = i[21083];
  assign o[21082] = i[21082];
  assign o[21081] = i[21081];
  assign o[21080] = i[21080];
  assign o[21079] = i[21079];
  assign o[21078] = i[21078];
  assign o[21077] = i[21077];
  assign o[21076] = i[21076];
  assign o[21075] = i[21075];
  assign o[21074] = i[21074];
  assign o[21073] = i[21073];
  assign o[21072] = i[21072];
  assign o[21071] = i[21071];
  assign o[21070] = i[21070];
  assign o[21069] = i[21069];
  assign o[21068] = i[21068];
  assign o[21067] = i[21067];
  assign o[21066] = i[21066];
  assign o[21065] = i[21065];
  assign o[21064] = i[21064];
  assign o[21063] = i[21063];
  assign o[21062] = i[21062];
  assign o[21061] = i[21061];
  assign o[21060] = i[21060];
  assign o[21059] = i[21059];
  assign o[21058] = i[21058];
  assign o[21057] = i[21057];
  assign o[21056] = i[21056];
  assign o[21055] = i[21055];
  assign o[21054] = i[21054];
  assign o[21053] = i[21053];
  assign o[21052] = i[21052];
  assign o[21051] = i[21051];
  assign o[21050] = i[21050];
  assign o[21049] = i[21049];
  assign o[21048] = i[21048];
  assign o[21047] = i[21047];
  assign o[21046] = i[21046];
  assign o[21045] = i[21045];
  assign o[21044] = i[21044];
  assign o[21043] = i[21043];
  assign o[21042] = i[21042];
  assign o[21041] = i[21041];
  assign o[21040] = i[21040];
  assign o[21039] = i[21039];
  assign o[21038] = i[21038];
  assign o[21037] = i[21037];
  assign o[21036] = i[21036];
  assign o[21035] = i[21035];
  assign o[21034] = i[21034];
  assign o[21033] = i[21033];
  assign o[21032] = i[21032];
  assign o[21031] = i[21031];
  assign o[21030] = i[21030];
  assign o[21029] = i[21029];
  assign o[21028] = i[21028];
  assign o[21027] = i[21027];
  assign o[21026] = i[21026];
  assign o[21025] = i[21025];
  assign o[21024] = i[21024];
  assign o[21023] = i[21023];
  assign o[21022] = i[21022];
  assign o[21021] = i[21021];
  assign o[21020] = i[21020];
  assign o[21019] = i[21019];
  assign o[21018] = i[21018];
  assign o[21017] = i[21017];
  assign o[21016] = i[21016];
  assign o[21015] = i[21015];
  assign o[21014] = i[21014];
  assign o[21013] = i[21013];
  assign o[21012] = i[21012];
  assign o[21011] = i[21011];
  assign o[21010] = i[21010];
  assign o[21009] = i[21009];
  assign o[21008] = i[21008];
  assign o[21007] = i[21007];
  assign o[21006] = i[21006];
  assign o[21005] = i[21005];
  assign o[21004] = i[21004];
  assign o[21003] = i[21003];
  assign o[21002] = i[21002];
  assign o[21001] = i[21001];
  assign o[21000] = i[21000];
  assign o[20999] = i[20999];
  assign o[20998] = i[20998];
  assign o[20997] = i[20997];
  assign o[20996] = i[20996];
  assign o[20995] = i[20995];
  assign o[20994] = i[20994];
  assign o[20993] = i[20993];
  assign o[20992] = i[20992];
  assign o[20991] = i[20991];
  assign o[20990] = i[20990];
  assign o[20989] = i[20989];
  assign o[20988] = i[20988];
  assign o[20987] = i[20987];
  assign o[20986] = i[20986];
  assign o[20985] = i[20985];
  assign o[20984] = i[20984];
  assign o[20983] = i[20983];
  assign o[20982] = i[20982];
  assign o[20981] = i[20981];
  assign o[20980] = i[20980];
  assign o[20979] = i[20979];
  assign o[20978] = i[20978];
  assign o[20977] = i[20977];
  assign o[20976] = i[20976];
  assign o[20975] = i[20975];
  assign o[20974] = i[20974];
  assign o[20973] = i[20973];
  assign o[20972] = i[20972];
  assign o[20971] = i[20971];
  assign o[20970] = i[20970];
  assign o[20969] = i[20969];
  assign o[20968] = i[20968];
  assign o[20967] = i[20967];
  assign o[20966] = i[20966];
  assign o[20965] = i[20965];
  assign o[20964] = i[20964];
  assign o[20963] = i[20963];
  assign o[20962] = i[20962];
  assign o[20961] = i[20961];
  assign o[20960] = i[20960];
  assign o[20959] = i[20959];
  assign o[20958] = i[20958];
  assign o[20957] = i[20957];
  assign o[20956] = i[20956];
  assign o[20955] = i[20955];
  assign o[20954] = i[20954];
  assign o[20953] = i[20953];
  assign o[20952] = i[20952];
  assign o[20951] = i[20951];
  assign o[20950] = i[20950];
  assign o[20949] = i[20949];
  assign o[20948] = i[20948];
  assign o[20947] = i[20947];
  assign o[20946] = i[20946];
  assign o[20945] = i[20945];
  assign o[20944] = i[20944];
  assign o[20943] = i[20943];
  assign o[20942] = i[20942];
  assign o[20941] = i[20941];
  assign o[20940] = i[20940];
  assign o[20939] = i[20939];
  assign o[20938] = i[20938];
  assign o[20937] = i[20937];
  assign o[20936] = i[20936];
  assign o[20935] = i[20935];
  assign o[20934] = i[20934];
  assign o[20933] = i[20933];
  assign o[20932] = i[20932];
  assign o[20931] = i[20931];
  assign o[20930] = i[20930];
  assign o[20929] = i[20929];
  assign o[20928] = i[20928];
  assign o[20927] = i[20927];
  assign o[20926] = i[20926];
  assign o[20925] = i[20925];
  assign o[20924] = i[20924];
  assign o[20923] = i[20923];
  assign o[20922] = i[20922];
  assign o[20921] = i[20921];
  assign o[20920] = i[20920];
  assign o[20919] = i[20919];
  assign o[20918] = i[20918];
  assign o[20917] = i[20917];
  assign o[20916] = i[20916];
  assign o[20915] = i[20915];
  assign o[20914] = i[20914];
  assign o[20913] = i[20913];
  assign o[20912] = i[20912];
  assign o[20911] = i[20911];
  assign o[20910] = i[20910];
  assign o[20909] = i[20909];
  assign o[20908] = i[20908];
  assign o[20907] = i[20907];
  assign o[20906] = i[20906];
  assign o[20905] = i[20905];
  assign o[20904] = i[20904];
  assign o[20903] = i[20903];
  assign o[20902] = i[20902];
  assign o[20901] = i[20901];
  assign o[20900] = i[20900];
  assign o[20899] = i[20899];
  assign o[20898] = i[20898];
  assign o[20897] = i[20897];
  assign o[20896] = i[20896];
  assign o[20895] = i[20895];
  assign o[20894] = i[20894];
  assign o[20893] = i[20893];
  assign o[20892] = i[20892];
  assign o[20891] = i[20891];
  assign o[20890] = i[20890];
  assign o[20889] = i[20889];
  assign o[20888] = i[20888];
  assign o[20887] = i[20887];
  assign o[20886] = i[20886];
  assign o[20885] = i[20885];
  assign o[20884] = i[20884];
  assign o[20883] = i[20883];
  assign o[20882] = i[20882];
  assign o[20881] = i[20881];
  assign o[20880] = i[20880];
  assign o[20879] = i[20879];
  assign o[20878] = i[20878];
  assign o[20877] = i[20877];
  assign o[20876] = i[20876];
  assign o[20875] = i[20875];
  assign o[20874] = i[20874];
  assign o[20873] = i[20873];
  assign o[20872] = i[20872];
  assign o[20871] = i[20871];
  assign o[20870] = i[20870];
  assign o[20869] = i[20869];
  assign o[20868] = i[20868];
  assign o[20867] = i[20867];
  assign o[20866] = i[20866];
  assign o[20865] = i[20865];
  assign o[20864] = i[20864];
  assign o[20863] = i[20863];
  assign o[20862] = i[20862];
  assign o[20861] = i[20861];
  assign o[20860] = i[20860];
  assign o[20859] = i[20859];
  assign o[20858] = i[20858];
  assign o[20857] = i[20857];
  assign o[20856] = i[20856];
  assign o[20855] = i[20855];
  assign o[20854] = i[20854];
  assign o[20853] = i[20853];
  assign o[20852] = i[20852];
  assign o[20851] = i[20851];
  assign o[20850] = i[20850];
  assign o[20849] = i[20849];
  assign o[20848] = i[20848];
  assign o[20847] = i[20847];
  assign o[20846] = i[20846];
  assign o[20845] = i[20845];
  assign o[20844] = i[20844];
  assign o[20843] = i[20843];
  assign o[20842] = i[20842];
  assign o[20841] = i[20841];
  assign o[20840] = i[20840];
  assign o[20839] = i[20839];
  assign o[20838] = i[20838];
  assign o[20837] = i[20837];
  assign o[20836] = i[20836];
  assign o[20835] = i[20835];
  assign o[20834] = i[20834];
  assign o[20833] = i[20833];
  assign o[20832] = i[20832];
  assign o[20831] = i[20831];
  assign o[20830] = i[20830];
  assign o[20829] = i[20829];
  assign o[20828] = i[20828];
  assign o[20827] = i[20827];
  assign o[20826] = i[20826];
  assign o[20825] = i[20825];
  assign o[20824] = i[20824];
  assign o[20823] = i[20823];
  assign o[20822] = i[20822];
  assign o[20821] = i[20821];
  assign o[20820] = i[20820];
  assign o[20819] = i[20819];
  assign o[20818] = i[20818];
  assign o[20817] = i[20817];
  assign o[20816] = i[20816];
  assign o[20815] = i[20815];
  assign o[20814] = i[20814];
  assign o[20813] = i[20813];
  assign o[20812] = i[20812];
  assign o[20811] = i[20811];
  assign o[20810] = i[20810];
  assign o[20809] = i[20809];
  assign o[20808] = i[20808];
  assign o[20807] = i[20807];
  assign o[20806] = i[20806];
  assign o[20805] = i[20805];
  assign o[20804] = i[20804];
  assign o[20803] = i[20803];
  assign o[20802] = i[20802];
  assign o[20801] = i[20801];
  assign o[20800] = i[20800];
  assign o[20799] = i[20799];
  assign o[20798] = i[20798];
  assign o[20797] = i[20797];
  assign o[20796] = i[20796];
  assign o[20795] = i[20795];
  assign o[20794] = i[20794];
  assign o[20793] = i[20793];
  assign o[20792] = i[20792];
  assign o[20791] = i[20791];
  assign o[20790] = i[20790];
  assign o[20789] = i[20789];
  assign o[20788] = i[20788];
  assign o[20787] = i[20787];
  assign o[20786] = i[20786];
  assign o[20785] = i[20785];
  assign o[20784] = i[20784];
  assign o[20783] = i[20783];
  assign o[20782] = i[20782];
  assign o[20781] = i[20781];
  assign o[20780] = i[20780];
  assign o[20779] = i[20779];
  assign o[20778] = i[20778];
  assign o[20777] = i[20777];
  assign o[20776] = i[20776];
  assign o[20775] = i[20775];
  assign o[20774] = i[20774];
  assign o[20773] = i[20773];
  assign o[20772] = i[20772];
  assign o[20771] = i[20771];
  assign o[20770] = i[20770];
  assign o[20769] = i[20769];
  assign o[20768] = i[20768];
  assign o[20767] = i[20767];
  assign o[20766] = i[20766];
  assign o[20765] = i[20765];
  assign o[20764] = i[20764];
  assign o[20763] = i[20763];
  assign o[20762] = i[20762];
  assign o[20761] = i[20761];
  assign o[20760] = i[20760];
  assign o[20759] = i[20759];
  assign o[20758] = i[20758];
  assign o[20757] = i[20757];
  assign o[20756] = i[20756];
  assign o[20755] = i[20755];
  assign o[20754] = i[20754];
  assign o[20753] = i[20753];
  assign o[20752] = i[20752];
  assign o[20751] = i[20751];
  assign o[20750] = i[20750];
  assign o[20749] = i[20749];
  assign o[20748] = i[20748];
  assign o[20747] = i[20747];
  assign o[20746] = i[20746];
  assign o[20745] = i[20745];
  assign o[20744] = i[20744];
  assign o[20743] = i[20743];
  assign o[20742] = i[20742];
  assign o[20741] = i[20741];
  assign o[20740] = i[20740];
  assign o[20739] = i[20739];
  assign o[20738] = i[20738];
  assign o[20737] = i[20737];
  assign o[20736] = i[20736];
  assign o[20735] = i[20735];
  assign o[20734] = i[20734];
  assign o[20733] = i[20733];
  assign o[20732] = i[20732];
  assign o[20731] = i[20731];
  assign o[20730] = i[20730];
  assign o[20729] = i[20729];
  assign o[20728] = i[20728];
  assign o[20727] = i[20727];
  assign o[20726] = i[20726];
  assign o[20725] = i[20725];
  assign o[20724] = i[20724];
  assign o[20723] = i[20723];
  assign o[20722] = i[20722];
  assign o[20721] = i[20721];
  assign o[20720] = i[20720];
  assign o[20719] = i[20719];
  assign o[20718] = i[20718];
  assign o[20717] = i[20717];
  assign o[20716] = i[20716];
  assign o[20715] = i[20715];
  assign o[20714] = i[20714];
  assign o[20713] = i[20713];
  assign o[20712] = i[20712];
  assign o[20711] = i[20711];
  assign o[20710] = i[20710];
  assign o[20709] = i[20709];
  assign o[20708] = i[20708];
  assign o[20707] = i[20707];
  assign o[20706] = i[20706];
  assign o[20705] = i[20705];
  assign o[20704] = i[20704];
  assign o[20703] = i[20703];
  assign o[20702] = i[20702];
  assign o[20701] = i[20701];
  assign o[20700] = i[20700];
  assign o[20699] = i[20699];
  assign o[20698] = i[20698];
  assign o[20697] = i[20697];
  assign o[20696] = i[20696];
  assign o[20695] = i[20695];
  assign o[20694] = i[20694];
  assign o[20693] = i[20693];
  assign o[20692] = i[20692];
  assign o[20691] = i[20691];
  assign o[20690] = i[20690];
  assign o[20689] = i[20689];
  assign o[20688] = i[20688];
  assign o[20687] = i[20687];
  assign o[20686] = i[20686];
  assign o[20685] = i[20685];
  assign o[20684] = i[20684];
  assign o[20683] = i[20683];
  assign o[20682] = i[20682];
  assign o[20681] = i[20681];
  assign o[20680] = i[20680];
  assign o[20679] = i[20679];
  assign o[20678] = i[20678];
  assign o[20677] = i[20677];
  assign o[20676] = i[20676];
  assign o[20675] = i[20675];
  assign o[20674] = i[20674];
  assign o[20673] = i[20673];
  assign o[20672] = i[20672];
  assign o[20671] = i[20671];
  assign o[20670] = i[20670];
  assign o[20669] = i[20669];
  assign o[20668] = i[20668];
  assign o[20667] = i[20667];
  assign o[20666] = i[20666];
  assign o[20665] = i[20665];
  assign o[20664] = i[20664];
  assign o[20663] = i[20663];
  assign o[20662] = i[20662];
  assign o[20661] = i[20661];
  assign o[20660] = i[20660];
  assign o[20659] = i[20659];
  assign o[20658] = i[20658];
  assign o[20657] = i[20657];
  assign o[20656] = i[20656];
  assign o[20655] = i[20655];
  assign o[20654] = i[20654];
  assign o[20653] = i[20653];
  assign o[20652] = i[20652];
  assign o[20651] = i[20651];
  assign o[20650] = i[20650];
  assign o[20649] = i[20649];
  assign o[20648] = i[20648];
  assign o[20647] = i[20647];
  assign o[20646] = i[20646];
  assign o[20645] = i[20645];
  assign o[20644] = i[20644];
  assign o[20643] = i[20643];
  assign o[20642] = i[20642];
  assign o[20641] = i[20641];
  assign o[20640] = i[20640];
  assign o[20639] = i[20639];
  assign o[20638] = i[20638];
  assign o[20637] = i[20637];
  assign o[20636] = i[20636];
  assign o[20635] = i[20635];
  assign o[20634] = i[20634];
  assign o[20633] = i[20633];
  assign o[20632] = i[20632];
  assign o[20631] = i[20631];
  assign o[20630] = i[20630];
  assign o[20629] = i[20629];
  assign o[20628] = i[20628];
  assign o[20627] = i[20627];
  assign o[20626] = i[20626];
  assign o[20625] = i[20625];
  assign o[20624] = i[20624];
  assign o[20623] = i[20623];
  assign o[20622] = i[20622];
  assign o[20621] = i[20621];
  assign o[20620] = i[20620];
  assign o[20619] = i[20619];
  assign o[20618] = i[20618];
  assign o[20617] = i[20617];
  assign o[20616] = i[20616];
  assign o[20615] = i[20615];
  assign o[20614] = i[20614];
  assign o[20613] = i[20613];
  assign o[20612] = i[20612];
  assign o[20611] = i[20611];
  assign o[20610] = i[20610];
  assign o[20609] = i[20609];
  assign o[20608] = i[20608];
  assign o[20607] = i[20607];
  assign o[20606] = i[20606];
  assign o[20605] = i[20605];
  assign o[20604] = i[20604];
  assign o[20603] = i[20603];
  assign o[20602] = i[20602];
  assign o[20601] = i[20601];
  assign o[20600] = i[20600];
  assign o[20599] = i[20599];
  assign o[20598] = i[20598];
  assign o[20597] = i[20597];
  assign o[20596] = i[20596];
  assign o[20595] = i[20595];
  assign o[20594] = i[20594];
  assign o[20593] = i[20593];
  assign o[20592] = i[20592];
  assign o[20591] = i[20591];
  assign o[20590] = i[20590];
  assign o[20589] = i[20589];
  assign o[20588] = i[20588];
  assign o[20587] = i[20587];
  assign o[20586] = i[20586];
  assign o[20585] = i[20585];
  assign o[20584] = i[20584];
  assign o[20583] = i[20583];
  assign o[20582] = i[20582];
  assign o[20581] = i[20581];
  assign o[20580] = i[20580];
  assign o[20579] = i[20579];
  assign o[20578] = i[20578];
  assign o[20577] = i[20577];
  assign o[20576] = i[20576];
  assign o[20575] = i[20575];
  assign o[20574] = i[20574];
  assign o[20573] = i[20573];
  assign o[20572] = i[20572];
  assign o[20571] = i[20571];
  assign o[20570] = i[20570];
  assign o[20569] = i[20569];
  assign o[20568] = i[20568];
  assign o[20567] = i[20567];
  assign o[20566] = i[20566];
  assign o[20565] = i[20565];
  assign o[20564] = i[20564];
  assign o[20563] = i[20563];
  assign o[20562] = i[20562];
  assign o[20561] = i[20561];
  assign o[20560] = i[20560];
  assign o[20559] = i[20559];
  assign o[20558] = i[20558];
  assign o[20557] = i[20557];
  assign o[20556] = i[20556];
  assign o[20555] = i[20555];
  assign o[20554] = i[20554];
  assign o[20553] = i[20553];
  assign o[20552] = i[20552];
  assign o[20551] = i[20551];
  assign o[20550] = i[20550];
  assign o[20549] = i[20549];
  assign o[20548] = i[20548];
  assign o[20547] = i[20547];
  assign o[20546] = i[20546];
  assign o[20545] = i[20545];
  assign o[20544] = i[20544];
  assign o[20543] = i[20543];
  assign o[20542] = i[20542];
  assign o[20541] = i[20541];
  assign o[20540] = i[20540];
  assign o[20539] = i[20539];
  assign o[20538] = i[20538];
  assign o[20537] = i[20537];
  assign o[20536] = i[20536];
  assign o[20535] = i[20535];
  assign o[20534] = i[20534];
  assign o[20533] = i[20533];
  assign o[20532] = i[20532];
  assign o[20531] = i[20531];
  assign o[20530] = i[20530];
  assign o[20529] = i[20529];
  assign o[20528] = i[20528];
  assign o[20527] = i[20527];
  assign o[20526] = i[20526];
  assign o[20525] = i[20525];
  assign o[20524] = i[20524];
  assign o[20523] = i[20523];
  assign o[20522] = i[20522];
  assign o[20521] = i[20521];
  assign o[20520] = i[20520];
  assign o[20519] = i[20519];
  assign o[20518] = i[20518];
  assign o[20517] = i[20517];
  assign o[20516] = i[20516];
  assign o[20515] = i[20515];
  assign o[20514] = i[20514];
  assign o[20513] = i[20513];
  assign o[20512] = i[20512];
  assign o[20511] = i[20511];
  assign o[20510] = i[20510];
  assign o[20509] = i[20509];
  assign o[20508] = i[20508];
  assign o[20507] = i[20507];
  assign o[20506] = i[20506];
  assign o[20505] = i[20505];
  assign o[20504] = i[20504];
  assign o[20503] = i[20503];
  assign o[20502] = i[20502];
  assign o[20501] = i[20501];
  assign o[20500] = i[20500];
  assign o[20499] = i[20499];
  assign o[20498] = i[20498];
  assign o[20497] = i[20497];
  assign o[20496] = i[20496];
  assign o[20495] = i[20495];
  assign o[20494] = i[20494];
  assign o[20493] = i[20493];
  assign o[20492] = i[20492];
  assign o[20491] = i[20491];
  assign o[20490] = i[20490];
  assign o[20489] = i[20489];
  assign o[20488] = i[20488];
  assign o[20487] = i[20487];
  assign o[20486] = i[20486];
  assign o[20485] = i[20485];
  assign o[20484] = i[20484];
  assign o[20483] = i[20483];
  assign o[20482] = i[20482];
  assign o[20481] = i[20481];
  assign o[20480] = i[20480];
  assign o[20479] = i[20479];
  assign o[20478] = i[20478];
  assign o[20477] = i[20477];
  assign o[20476] = i[20476];
  assign o[20475] = i[20475];
  assign o[20474] = i[20474];
  assign o[20473] = i[20473];
  assign o[20472] = i[20472];
  assign o[20471] = i[20471];
  assign o[20470] = i[20470];
  assign o[20469] = i[20469];
  assign o[20468] = i[20468];
  assign o[20467] = i[20467];
  assign o[20466] = i[20466];
  assign o[20465] = i[20465];
  assign o[20464] = i[20464];
  assign o[20463] = i[20463];
  assign o[20462] = i[20462];
  assign o[20461] = i[20461];
  assign o[20460] = i[20460];
  assign o[20459] = i[20459];
  assign o[20458] = i[20458];
  assign o[20457] = i[20457];
  assign o[20456] = i[20456];
  assign o[20455] = i[20455];
  assign o[20454] = i[20454];
  assign o[20453] = i[20453];
  assign o[20452] = i[20452];
  assign o[20451] = i[20451];
  assign o[20450] = i[20450];
  assign o[20449] = i[20449];
  assign o[20448] = i[20448];
  assign o[20447] = i[20447];
  assign o[20446] = i[20446];
  assign o[20445] = i[20445];
  assign o[20444] = i[20444];
  assign o[20443] = i[20443];
  assign o[20442] = i[20442];
  assign o[20441] = i[20441];
  assign o[20440] = i[20440];
  assign o[20439] = i[20439];
  assign o[20438] = i[20438];
  assign o[20437] = i[20437];
  assign o[20436] = i[20436];
  assign o[20435] = i[20435];
  assign o[20434] = i[20434];
  assign o[20433] = i[20433];
  assign o[20432] = i[20432];
  assign o[20431] = i[20431];
  assign o[20430] = i[20430];
  assign o[20429] = i[20429];
  assign o[20428] = i[20428];
  assign o[20427] = i[20427];
  assign o[20426] = i[20426];
  assign o[20425] = i[20425];
  assign o[20424] = i[20424];
  assign o[20423] = i[20423];
  assign o[20422] = i[20422];
  assign o[20421] = i[20421];
  assign o[20420] = i[20420];
  assign o[20419] = i[20419];
  assign o[20418] = i[20418];
  assign o[20417] = i[20417];
  assign o[20416] = i[20416];
  assign o[20415] = i[20415];
  assign o[20414] = i[20414];
  assign o[20413] = i[20413];
  assign o[20412] = i[20412];
  assign o[20411] = i[20411];
  assign o[20410] = i[20410];
  assign o[20409] = i[20409];
  assign o[20408] = i[20408];
  assign o[20407] = i[20407];
  assign o[20406] = i[20406];
  assign o[20405] = i[20405];
  assign o[20404] = i[20404];
  assign o[20403] = i[20403];
  assign o[20402] = i[20402];
  assign o[20401] = i[20401];
  assign o[20400] = i[20400];
  assign o[20399] = i[20399];
  assign o[20398] = i[20398];
  assign o[20397] = i[20397];
  assign o[20396] = i[20396];
  assign o[20395] = i[20395];
  assign o[20394] = i[20394];
  assign o[20393] = i[20393];
  assign o[20392] = i[20392];
  assign o[20391] = i[20391];
  assign o[20390] = i[20390];
  assign o[20389] = i[20389];
  assign o[20388] = i[20388];
  assign o[20387] = i[20387];
  assign o[20386] = i[20386];
  assign o[20385] = i[20385];
  assign o[20384] = i[20384];
  assign o[20383] = i[20383];
  assign o[20382] = i[20382];
  assign o[20381] = i[20381];
  assign o[20380] = i[20380];
  assign o[20379] = i[20379];
  assign o[20378] = i[20378];
  assign o[20377] = i[20377];
  assign o[20376] = i[20376];
  assign o[20375] = i[20375];
  assign o[20374] = i[20374];
  assign o[20373] = i[20373];
  assign o[20372] = i[20372];
  assign o[20371] = i[20371];
  assign o[20370] = i[20370];
  assign o[20369] = i[20369];
  assign o[20368] = i[20368];
  assign o[20367] = i[20367];
  assign o[20366] = i[20366];
  assign o[20365] = i[20365];
  assign o[20364] = i[20364];
  assign o[20363] = i[20363];
  assign o[20362] = i[20362];
  assign o[20361] = i[20361];
  assign o[20360] = i[20360];
  assign o[20359] = i[20359];
  assign o[20358] = i[20358];
  assign o[20357] = i[20357];
  assign o[20356] = i[20356];
  assign o[20355] = i[20355];
  assign o[20354] = i[20354];
  assign o[20353] = i[20353];
  assign o[20352] = i[20352];
  assign o[20351] = i[20351];
  assign o[20350] = i[20350];
  assign o[20349] = i[20349];
  assign o[20348] = i[20348];
  assign o[20347] = i[20347];
  assign o[20346] = i[20346];
  assign o[20345] = i[20345];
  assign o[20344] = i[20344];
  assign o[20343] = i[20343];
  assign o[20342] = i[20342];
  assign o[20341] = i[20341];
  assign o[20340] = i[20340];
  assign o[20339] = i[20339];
  assign o[20338] = i[20338];
  assign o[20337] = i[20337];
  assign o[20336] = i[20336];
  assign o[20335] = i[20335];
  assign o[20334] = i[20334];
  assign o[20333] = i[20333];
  assign o[20332] = i[20332];
  assign o[20331] = i[20331];
  assign o[20330] = i[20330];
  assign o[20329] = i[20329];
  assign o[20328] = i[20328];
  assign o[20327] = i[20327];
  assign o[20326] = i[20326];
  assign o[20325] = i[20325];
  assign o[20324] = i[20324];
  assign o[20323] = i[20323];
  assign o[20322] = i[20322];
  assign o[20321] = i[20321];
  assign o[20320] = i[20320];
  assign o[20319] = i[20319];
  assign o[20318] = i[20318];
  assign o[20317] = i[20317];
  assign o[20316] = i[20316];
  assign o[20315] = i[20315];
  assign o[20314] = i[20314];
  assign o[20313] = i[20313];
  assign o[20312] = i[20312];
  assign o[20311] = i[20311];
  assign o[20310] = i[20310];
  assign o[20309] = i[20309];
  assign o[20308] = i[20308];
  assign o[20307] = i[20307];
  assign o[20306] = i[20306];
  assign o[20305] = i[20305];
  assign o[20304] = i[20304];
  assign o[20303] = i[20303];
  assign o[20302] = i[20302];
  assign o[20301] = i[20301];
  assign o[20300] = i[20300];
  assign o[20299] = i[20299];
  assign o[20298] = i[20298];
  assign o[20297] = i[20297];
  assign o[20296] = i[20296];
  assign o[20295] = i[20295];
  assign o[20294] = i[20294];
  assign o[20293] = i[20293];
  assign o[20292] = i[20292];
  assign o[20291] = i[20291];
  assign o[20290] = i[20290];
  assign o[20289] = i[20289];
  assign o[20288] = i[20288];
  assign o[20287] = i[20287];
  assign o[20286] = i[20286];
  assign o[20285] = i[20285];
  assign o[20284] = i[20284];
  assign o[20283] = i[20283];
  assign o[20282] = i[20282];
  assign o[20281] = i[20281];
  assign o[20280] = i[20280];
  assign o[20279] = i[20279];
  assign o[20278] = i[20278];
  assign o[20277] = i[20277];
  assign o[20276] = i[20276];
  assign o[20275] = i[20275];
  assign o[20274] = i[20274];
  assign o[20273] = i[20273];
  assign o[20272] = i[20272];
  assign o[20271] = i[20271];
  assign o[20270] = i[20270];
  assign o[20269] = i[20269];
  assign o[20268] = i[20268];
  assign o[20267] = i[20267];
  assign o[20266] = i[20266];
  assign o[20265] = i[20265];
  assign o[20264] = i[20264];
  assign o[20263] = i[20263];
  assign o[20262] = i[20262];
  assign o[20261] = i[20261];
  assign o[20260] = i[20260];
  assign o[20259] = i[20259];
  assign o[20258] = i[20258];
  assign o[20257] = i[20257];
  assign o[20256] = i[20256];
  assign o[20255] = i[20255];
  assign o[20254] = i[20254];
  assign o[20253] = i[20253];
  assign o[20252] = i[20252];
  assign o[20251] = i[20251];
  assign o[20250] = i[20250];
  assign o[20249] = i[20249];
  assign o[20248] = i[20248];
  assign o[20247] = i[20247];
  assign o[20246] = i[20246];
  assign o[20245] = i[20245];
  assign o[20244] = i[20244];
  assign o[20243] = i[20243];
  assign o[20242] = i[20242];
  assign o[20241] = i[20241];
  assign o[20240] = i[20240];
  assign o[20239] = i[20239];
  assign o[20238] = i[20238];
  assign o[20237] = i[20237];
  assign o[20236] = i[20236];
  assign o[20235] = i[20235];
  assign o[20234] = i[20234];
  assign o[20233] = i[20233];
  assign o[20232] = i[20232];
  assign o[20231] = i[20231];
  assign o[20230] = i[20230];
  assign o[20229] = i[20229];
  assign o[20228] = i[20228];
  assign o[20227] = i[20227];
  assign o[20226] = i[20226];
  assign o[20225] = i[20225];
  assign o[20224] = i[20224];
  assign o[20223] = i[20223];
  assign o[20222] = i[20222];
  assign o[20221] = i[20221];
  assign o[20220] = i[20220];
  assign o[20219] = i[20219];
  assign o[20218] = i[20218];
  assign o[20217] = i[20217];
  assign o[20216] = i[20216];
  assign o[20215] = i[20215];
  assign o[20214] = i[20214];
  assign o[20213] = i[20213];
  assign o[20212] = i[20212];
  assign o[20211] = i[20211];
  assign o[20210] = i[20210];
  assign o[20209] = i[20209];
  assign o[20208] = i[20208];
  assign o[20207] = i[20207];
  assign o[20206] = i[20206];
  assign o[20205] = i[20205];
  assign o[20204] = i[20204];
  assign o[20203] = i[20203];
  assign o[20202] = i[20202];
  assign o[20201] = i[20201];
  assign o[20200] = i[20200];
  assign o[20199] = i[20199];
  assign o[20198] = i[20198];
  assign o[20197] = i[20197];
  assign o[20196] = i[20196];
  assign o[20195] = i[20195];
  assign o[20194] = i[20194];
  assign o[20193] = i[20193];
  assign o[20192] = i[20192];
  assign o[20191] = i[20191];
  assign o[20190] = i[20190];
  assign o[20189] = i[20189];
  assign o[20188] = i[20188];
  assign o[20187] = i[20187];
  assign o[20186] = i[20186];
  assign o[20185] = i[20185];
  assign o[20184] = i[20184];
  assign o[20183] = i[20183];
  assign o[20182] = i[20182];
  assign o[20181] = i[20181];
  assign o[20180] = i[20180];
  assign o[20179] = i[20179];
  assign o[20178] = i[20178];
  assign o[20177] = i[20177];
  assign o[20176] = i[20176];
  assign o[20175] = i[20175];
  assign o[20174] = i[20174];
  assign o[20173] = i[20173];
  assign o[20172] = i[20172];
  assign o[20171] = i[20171];
  assign o[20170] = i[20170];
  assign o[20169] = i[20169];
  assign o[20168] = i[20168];
  assign o[20167] = i[20167];
  assign o[20166] = i[20166];
  assign o[20165] = i[20165];
  assign o[20164] = i[20164];
  assign o[20163] = i[20163];
  assign o[20162] = i[20162];
  assign o[20161] = i[20161];
  assign o[20160] = i[20160];
  assign o[20159] = i[20159];
  assign o[20158] = i[20158];
  assign o[20157] = i[20157];
  assign o[20156] = i[20156];
  assign o[20155] = i[20155];
  assign o[20154] = i[20154];
  assign o[20153] = i[20153];
  assign o[20152] = i[20152];
  assign o[20151] = i[20151];
  assign o[20150] = i[20150];
  assign o[20149] = i[20149];
  assign o[20148] = i[20148];
  assign o[20147] = i[20147];
  assign o[20146] = i[20146];
  assign o[20145] = i[20145];
  assign o[20144] = i[20144];
  assign o[20143] = i[20143];
  assign o[20142] = i[20142];
  assign o[20141] = i[20141];
  assign o[20140] = i[20140];
  assign o[20139] = i[20139];
  assign o[20138] = i[20138];
  assign o[20137] = i[20137];
  assign o[20136] = i[20136];
  assign o[20135] = i[20135];
  assign o[20134] = i[20134];
  assign o[20133] = i[20133];
  assign o[20132] = i[20132];
  assign o[20131] = i[20131];
  assign o[20130] = i[20130];
  assign o[20129] = i[20129];
  assign o[20128] = i[20128];
  assign o[20127] = i[20127];
  assign o[20126] = i[20126];
  assign o[20125] = i[20125];
  assign o[20124] = i[20124];
  assign o[20123] = i[20123];
  assign o[20122] = i[20122];
  assign o[20121] = i[20121];
  assign o[20120] = i[20120];
  assign o[20119] = i[20119];
  assign o[20118] = i[20118];
  assign o[20117] = i[20117];
  assign o[20116] = i[20116];
  assign o[20115] = i[20115];
  assign o[20114] = i[20114];
  assign o[20113] = i[20113];
  assign o[20112] = i[20112];
  assign o[20111] = i[20111];
  assign o[20110] = i[20110];
  assign o[20109] = i[20109];
  assign o[20108] = i[20108];
  assign o[20107] = i[20107];
  assign o[20106] = i[20106];
  assign o[20105] = i[20105];
  assign o[20104] = i[20104];
  assign o[20103] = i[20103];
  assign o[20102] = i[20102];
  assign o[20101] = i[20101];
  assign o[20100] = i[20100];
  assign o[20099] = i[20099];
  assign o[20098] = i[20098];
  assign o[20097] = i[20097];
  assign o[20096] = i[20096];
  assign o[20095] = i[20095];
  assign o[20094] = i[20094];
  assign o[20093] = i[20093];
  assign o[20092] = i[20092];
  assign o[20091] = i[20091];
  assign o[20090] = i[20090];
  assign o[20089] = i[20089];
  assign o[20088] = i[20088];
  assign o[20087] = i[20087];
  assign o[20086] = i[20086];
  assign o[20085] = i[20085];
  assign o[20084] = i[20084];
  assign o[20083] = i[20083];
  assign o[20082] = i[20082];
  assign o[20081] = i[20081];
  assign o[20080] = i[20080];
  assign o[20079] = i[20079];
  assign o[20078] = i[20078];
  assign o[20077] = i[20077];
  assign o[20076] = i[20076];
  assign o[20075] = i[20075];
  assign o[20074] = i[20074];
  assign o[20073] = i[20073];
  assign o[20072] = i[20072];
  assign o[20071] = i[20071];
  assign o[20070] = i[20070];
  assign o[20069] = i[20069];
  assign o[20068] = i[20068];
  assign o[20067] = i[20067];
  assign o[20066] = i[20066];
  assign o[20065] = i[20065];
  assign o[20064] = i[20064];
  assign o[20063] = i[20063];
  assign o[20062] = i[20062];
  assign o[20061] = i[20061];
  assign o[20060] = i[20060];
  assign o[20059] = i[20059];
  assign o[20058] = i[20058];
  assign o[20057] = i[20057];
  assign o[20056] = i[20056];
  assign o[20055] = i[20055];
  assign o[20054] = i[20054];
  assign o[20053] = i[20053];
  assign o[20052] = i[20052];
  assign o[20051] = i[20051];
  assign o[20050] = i[20050];
  assign o[20049] = i[20049];
  assign o[20048] = i[20048];
  assign o[20047] = i[20047];
  assign o[20046] = i[20046];
  assign o[20045] = i[20045];
  assign o[20044] = i[20044];
  assign o[20043] = i[20043];
  assign o[20042] = i[20042];
  assign o[20041] = i[20041];
  assign o[20040] = i[20040];
  assign o[20039] = i[20039];
  assign o[20038] = i[20038];
  assign o[20037] = i[20037];
  assign o[20036] = i[20036];
  assign o[20035] = i[20035];
  assign o[20034] = i[20034];
  assign o[20033] = i[20033];
  assign o[20032] = i[20032];
  assign o[20031] = i[20031];
  assign o[20030] = i[20030];
  assign o[20029] = i[20029];
  assign o[20028] = i[20028];
  assign o[20027] = i[20027];
  assign o[20026] = i[20026];
  assign o[20025] = i[20025];
  assign o[20024] = i[20024];
  assign o[20023] = i[20023];
  assign o[20022] = i[20022];
  assign o[20021] = i[20021];
  assign o[20020] = i[20020];
  assign o[20019] = i[20019];
  assign o[20018] = i[20018];
  assign o[20017] = i[20017];
  assign o[20016] = i[20016];
  assign o[20015] = i[20015];
  assign o[20014] = i[20014];
  assign o[20013] = i[20013];
  assign o[20012] = i[20012];
  assign o[20011] = i[20011];
  assign o[20010] = i[20010];
  assign o[20009] = i[20009];
  assign o[20008] = i[20008];
  assign o[20007] = i[20007];
  assign o[20006] = i[20006];
  assign o[20005] = i[20005];
  assign o[20004] = i[20004];
  assign o[20003] = i[20003];
  assign o[20002] = i[20002];
  assign o[20001] = i[20001];
  assign o[20000] = i[20000];
  assign o[19999] = i[19999];
  assign o[19998] = i[19998];
  assign o[19997] = i[19997];
  assign o[19996] = i[19996];
  assign o[19995] = i[19995];
  assign o[19994] = i[19994];
  assign o[19993] = i[19993];
  assign o[19992] = i[19992];
  assign o[19991] = i[19991];
  assign o[19990] = i[19990];
  assign o[19989] = i[19989];
  assign o[19988] = i[19988];
  assign o[19987] = i[19987];
  assign o[19986] = i[19986];
  assign o[19985] = i[19985];
  assign o[19984] = i[19984];
  assign o[19983] = i[19983];
  assign o[19982] = i[19982];
  assign o[19981] = i[19981];
  assign o[19980] = i[19980];
  assign o[19979] = i[19979];
  assign o[19978] = i[19978];
  assign o[19977] = i[19977];
  assign o[19976] = i[19976];
  assign o[19975] = i[19975];
  assign o[19974] = i[19974];
  assign o[19973] = i[19973];
  assign o[19972] = i[19972];
  assign o[19971] = i[19971];
  assign o[19970] = i[19970];
  assign o[19969] = i[19969];
  assign o[19968] = i[19968];
  assign o[19967] = i[19967];
  assign o[19966] = i[19966];
  assign o[19965] = i[19965];
  assign o[19964] = i[19964];
  assign o[19963] = i[19963];
  assign o[19962] = i[19962];
  assign o[19961] = i[19961];
  assign o[19960] = i[19960];
  assign o[19959] = i[19959];
  assign o[19958] = i[19958];
  assign o[19957] = i[19957];
  assign o[19956] = i[19956];
  assign o[19955] = i[19955];
  assign o[19954] = i[19954];
  assign o[19953] = i[19953];
  assign o[19952] = i[19952];
  assign o[19951] = i[19951];
  assign o[19950] = i[19950];
  assign o[19949] = i[19949];
  assign o[19948] = i[19948];
  assign o[19947] = i[19947];
  assign o[19946] = i[19946];
  assign o[19945] = i[19945];
  assign o[19944] = i[19944];
  assign o[19943] = i[19943];
  assign o[19942] = i[19942];
  assign o[19941] = i[19941];
  assign o[19940] = i[19940];
  assign o[19939] = i[19939];
  assign o[19938] = i[19938];
  assign o[19937] = i[19937];
  assign o[19936] = i[19936];
  assign o[19935] = i[19935];
  assign o[19934] = i[19934];
  assign o[19933] = i[19933];
  assign o[19932] = i[19932];
  assign o[19931] = i[19931];
  assign o[19930] = i[19930];
  assign o[19929] = i[19929];
  assign o[19928] = i[19928];
  assign o[19927] = i[19927];
  assign o[19926] = i[19926];
  assign o[19925] = i[19925];
  assign o[19924] = i[19924];
  assign o[19923] = i[19923];
  assign o[19922] = i[19922];
  assign o[19921] = i[19921];
  assign o[19920] = i[19920];
  assign o[19919] = i[19919];
  assign o[19918] = i[19918];
  assign o[19917] = i[19917];
  assign o[19916] = i[19916];
  assign o[19915] = i[19915];
  assign o[19914] = i[19914];
  assign o[19913] = i[19913];
  assign o[19912] = i[19912];
  assign o[19911] = i[19911];
  assign o[19910] = i[19910];
  assign o[19909] = i[19909];
  assign o[19908] = i[19908];
  assign o[19907] = i[19907];
  assign o[19906] = i[19906];
  assign o[19905] = i[19905];
  assign o[19904] = i[19904];
  assign o[19903] = i[19903];
  assign o[19902] = i[19902];
  assign o[19901] = i[19901];
  assign o[19900] = i[19900];
  assign o[19899] = i[19899];
  assign o[19898] = i[19898];
  assign o[19897] = i[19897];
  assign o[19896] = i[19896];
  assign o[19895] = i[19895];
  assign o[19894] = i[19894];
  assign o[19893] = i[19893];
  assign o[19892] = i[19892];
  assign o[19891] = i[19891];
  assign o[19890] = i[19890];
  assign o[19889] = i[19889];
  assign o[19888] = i[19888];
  assign o[19887] = i[19887];
  assign o[19886] = i[19886];
  assign o[19885] = i[19885];
  assign o[19884] = i[19884];
  assign o[19883] = i[19883];
  assign o[19882] = i[19882];
  assign o[19881] = i[19881];
  assign o[19880] = i[19880];
  assign o[19879] = i[19879];
  assign o[19878] = i[19878];
  assign o[19877] = i[19877];
  assign o[19876] = i[19876];
  assign o[19875] = i[19875];
  assign o[19874] = i[19874];
  assign o[19873] = i[19873];
  assign o[19872] = i[19872];
  assign o[19871] = i[19871];
  assign o[19870] = i[19870];
  assign o[19869] = i[19869];
  assign o[19868] = i[19868];
  assign o[19867] = i[19867];
  assign o[19866] = i[19866];
  assign o[19865] = i[19865];
  assign o[19864] = i[19864];
  assign o[19863] = i[19863];
  assign o[19862] = i[19862];
  assign o[19861] = i[19861];
  assign o[19860] = i[19860];
  assign o[19859] = i[19859];
  assign o[19858] = i[19858];
  assign o[19857] = i[19857];
  assign o[19856] = i[19856];
  assign o[19855] = i[19855];
  assign o[19854] = i[19854];
  assign o[19853] = i[19853];
  assign o[19852] = i[19852];
  assign o[19851] = i[19851];
  assign o[19850] = i[19850];
  assign o[19849] = i[19849];
  assign o[19848] = i[19848];
  assign o[19847] = i[19847];
  assign o[19846] = i[19846];
  assign o[19845] = i[19845];
  assign o[19844] = i[19844];
  assign o[19843] = i[19843];
  assign o[19842] = i[19842];
  assign o[19841] = i[19841];
  assign o[19840] = i[19840];
  assign o[19839] = i[19839];
  assign o[19838] = i[19838];
  assign o[19837] = i[19837];
  assign o[19836] = i[19836];
  assign o[19835] = i[19835];
  assign o[19834] = i[19834];
  assign o[19833] = i[19833];
  assign o[19832] = i[19832];
  assign o[19831] = i[19831];
  assign o[19830] = i[19830];
  assign o[19829] = i[19829];
  assign o[19828] = i[19828];
  assign o[19827] = i[19827];
  assign o[19826] = i[19826];
  assign o[19825] = i[19825];
  assign o[19824] = i[19824];
  assign o[19823] = i[19823];
  assign o[19822] = i[19822];
  assign o[19821] = i[19821];
  assign o[19820] = i[19820];
  assign o[19819] = i[19819];
  assign o[19818] = i[19818];
  assign o[19817] = i[19817];
  assign o[19816] = i[19816];
  assign o[19815] = i[19815];
  assign o[19814] = i[19814];
  assign o[19813] = i[19813];
  assign o[19812] = i[19812];
  assign o[19811] = i[19811];
  assign o[19810] = i[19810];
  assign o[19809] = i[19809];
  assign o[19808] = i[19808];
  assign o[19807] = i[19807];
  assign o[19806] = i[19806];
  assign o[19805] = i[19805];
  assign o[19804] = i[19804];
  assign o[19803] = i[19803];
  assign o[19802] = i[19802];
  assign o[19801] = i[19801];
  assign o[19800] = i[19800];
  assign o[19799] = i[19799];
  assign o[19798] = i[19798];
  assign o[19797] = i[19797];
  assign o[19796] = i[19796];
  assign o[19795] = i[19795];
  assign o[19794] = i[19794];
  assign o[19793] = i[19793];
  assign o[19792] = i[19792];
  assign o[19791] = i[19791];
  assign o[19790] = i[19790];
  assign o[19789] = i[19789];
  assign o[19788] = i[19788];
  assign o[19787] = i[19787];
  assign o[19786] = i[19786];
  assign o[19785] = i[19785];
  assign o[19784] = i[19784];
  assign o[19783] = i[19783];
  assign o[19782] = i[19782];
  assign o[19781] = i[19781];
  assign o[19780] = i[19780];
  assign o[19779] = i[19779];
  assign o[19778] = i[19778];
  assign o[19777] = i[19777];
  assign o[19776] = i[19776];
  assign o[19775] = i[19775];
  assign o[19774] = i[19774];
  assign o[19773] = i[19773];
  assign o[19772] = i[19772];
  assign o[19771] = i[19771];
  assign o[19770] = i[19770];
  assign o[19769] = i[19769];
  assign o[19768] = i[19768];
  assign o[19767] = i[19767];
  assign o[19766] = i[19766];
  assign o[19765] = i[19765];
  assign o[19764] = i[19764];
  assign o[19763] = i[19763];
  assign o[19762] = i[19762];
  assign o[19761] = i[19761];
  assign o[19760] = i[19760];
  assign o[19759] = i[19759];
  assign o[19758] = i[19758];
  assign o[19757] = i[19757];
  assign o[19756] = i[19756];
  assign o[19755] = i[19755];
  assign o[19754] = i[19754];
  assign o[19753] = i[19753];
  assign o[19752] = i[19752];
  assign o[19751] = i[19751];
  assign o[19750] = i[19750];
  assign o[19749] = i[19749];
  assign o[19748] = i[19748];
  assign o[19747] = i[19747];
  assign o[19746] = i[19746];
  assign o[19745] = i[19745];
  assign o[19744] = i[19744];
  assign o[19743] = i[19743];
  assign o[19742] = i[19742];
  assign o[19741] = i[19741];
  assign o[19740] = i[19740];
  assign o[19739] = i[19739];
  assign o[19738] = i[19738];
  assign o[19737] = i[19737];
  assign o[19736] = i[19736];
  assign o[19735] = i[19735];
  assign o[19734] = i[19734];
  assign o[19733] = i[19733];
  assign o[19732] = i[19732];
  assign o[19731] = i[19731];
  assign o[19730] = i[19730];
  assign o[19729] = i[19729];
  assign o[19728] = i[19728];
  assign o[19727] = i[19727];
  assign o[19726] = i[19726];
  assign o[19725] = i[19725];
  assign o[19724] = i[19724];
  assign o[19723] = i[19723];
  assign o[19722] = i[19722];
  assign o[19721] = i[19721];
  assign o[19720] = i[19720];
  assign o[19719] = i[19719];
  assign o[19718] = i[19718];
  assign o[19717] = i[19717];
  assign o[19716] = i[19716];
  assign o[19715] = i[19715];
  assign o[19714] = i[19714];
  assign o[19713] = i[19713];
  assign o[19712] = i[19712];
  assign o[19711] = i[19711];
  assign o[19710] = i[19710];
  assign o[19709] = i[19709];
  assign o[19708] = i[19708];
  assign o[19707] = i[19707];
  assign o[19706] = i[19706];
  assign o[19705] = i[19705];
  assign o[19704] = i[19704];
  assign o[19703] = i[19703];
  assign o[19702] = i[19702];
  assign o[19701] = i[19701];
  assign o[19700] = i[19700];
  assign o[19699] = i[19699];
  assign o[19698] = i[19698];
  assign o[19697] = i[19697];
  assign o[19696] = i[19696];
  assign o[19695] = i[19695];
  assign o[19694] = i[19694];
  assign o[19693] = i[19693];
  assign o[19692] = i[19692];
  assign o[19691] = i[19691];
  assign o[19690] = i[19690];
  assign o[19689] = i[19689];
  assign o[19688] = i[19688];
  assign o[19687] = i[19687];
  assign o[19686] = i[19686];
  assign o[19685] = i[19685];
  assign o[19684] = i[19684];
  assign o[19683] = i[19683];
  assign o[19682] = i[19682];
  assign o[19681] = i[19681];
  assign o[19680] = i[19680];
  assign o[19679] = i[19679];
  assign o[19678] = i[19678];
  assign o[19677] = i[19677];
  assign o[19676] = i[19676];
  assign o[19675] = i[19675];
  assign o[19674] = i[19674];
  assign o[19673] = i[19673];
  assign o[19672] = i[19672];
  assign o[19671] = i[19671];
  assign o[19670] = i[19670];
  assign o[19669] = i[19669];
  assign o[19668] = i[19668];
  assign o[19667] = i[19667];
  assign o[19666] = i[19666];
  assign o[19665] = i[19665];
  assign o[19664] = i[19664];
  assign o[19663] = i[19663];
  assign o[19662] = i[19662];
  assign o[19661] = i[19661];
  assign o[19660] = i[19660];
  assign o[19659] = i[19659];
  assign o[19658] = i[19658];
  assign o[19657] = i[19657];
  assign o[19656] = i[19656];
  assign o[19655] = i[19655];
  assign o[19654] = i[19654];
  assign o[19653] = i[19653];
  assign o[19652] = i[19652];
  assign o[19651] = i[19651];
  assign o[19650] = i[19650];
  assign o[19649] = i[19649];
  assign o[19648] = i[19648];
  assign o[19647] = i[19647];
  assign o[19646] = i[19646];
  assign o[19645] = i[19645];
  assign o[19644] = i[19644];
  assign o[19643] = i[19643];
  assign o[19642] = i[19642];
  assign o[19641] = i[19641];
  assign o[19640] = i[19640];
  assign o[19639] = i[19639];
  assign o[19638] = i[19638];
  assign o[19637] = i[19637];
  assign o[19636] = i[19636];
  assign o[19635] = i[19635];
  assign o[19634] = i[19634];
  assign o[19633] = i[19633];
  assign o[19632] = i[19632];
  assign o[19631] = i[19631];
  assign o[19630] = i[19630];
  assign o[19629] = i[19629];
  assign o[19628] = i[19628];
  assign o[19627] = i[19627];
  assign o[19626] = i[19626];
  assign o[19625] = i[19625];
  assign o[19624] = i[19624];
  assign o[19623] = i[19623];
  assign o[19622] = i[19622];
  assign o[19621] = i[19621];
  assign o[19620] = i[19620];
  assign o[19619] = i[19619];
  assign o[19618] = i[19618];
  assign o[19617] = i[19617];
  assign o[19616] = i[19616];
  assign o[19615] = i[19615];
  assign o[19614] = i[19614];
  assign o[19613] = i[19613];
  assign o[19612] = i[19612];
  assign o[19611] = i[19611];
  assign o[19610] = i[19610];
  assign o[19609] = i[19609];
  assign o[19608] = i[19608];
  assign o[19607] = i[19607];
  assign o[19606] = i[19606];
  assign o[19605] = i[19605];
  assign o[19604] = i[19604];
  assign o[19603] = i[19603];
  assign o[19602] = i[19602];
  assign o[19601] = i[19601];
  assign o[19600] = i[19600];
  assign o[19599] = i[19599];
  assign o[19598] = i[19598];
  assign o[19597] = i[19597];
  assign o[19596] = i[19596];
  assign o[19595] = i[19595];
  assign o[19594] = i[19594];
  assign o[19593] = i[19593];
  assign o[19592] = i[19592];
  assign o[19591] = i[19591];
  assign o[19590] = i[19590];
  assign o[19589] = i[19589];
  assign o[19588] = i[19588];
  assign o[19587] = i[19587];
  assign o[19586] = i[19586];
  assign o[19585] = i[19585];
  assign o[19584] = i[19584];
  assign o[19583] = i[19583];
  assign o[19582] = i[19582];
  assign o[19581] = i[19581];
  assign o[19580] = i[19580];
  assign o[19579] = i[19579];
  assign o[19578] = i[19578];
  assign o[19577] = i[19577];
  assign o[19576] = i[19576];
  assign o[19575] = i[19575];
  assign o[19574] = i[19574];
  assign o[19573] = i[19573];
  assign o[19572] = i[19572];
  assign o[19571] = i[19571];
  assign o[19570] = i[19570];
  assign o[19569] = i[19569];
  assign o[19568] = i[19568];
  assign o[19567] = i[19567];
  assign o[19566] = i[19566];
  assign o[19565] = i[19565];
  assign o[19564] = i[19564];
  assign o[19563] = i[19563];
  assign o[19562] = i[19562];
  assign o[19561] = i[19561];
  assign o[19560] = i[19560];
  assign o[19559] = i[19559];
  assign o[19558] = i[19558];
  assign o[19557] = i[19557];
  assign o[19556] = i[19556];
  assign o[19555] = i[19555];
  assign o[19554] = i[19554];
  assign o[19553] = i[19553];
  assign o[19552] = i[19552];
  assign o[19551] = i[19551];
  assign o[19550] = i[19550];
  assign o[19549] = i[19549];
  assign o[19548] = i[19548];
  assign o[19547] = i[19547];
  assign o[19546] = i[19546];
  assign o[19545] = i[19545];
  assign o[19544] = i[19544];
  assign o[19543] = i[19543];
  assign o[19542] = i[19542];
  assign o[19541] = i[19541];
  assign o[19540] = i[19540];
  assign o[19539] = i[19539];
  assign o[19538] = i[19538];
  assign o[19537] = i[19537];
  assign o[19536] = i[19536];
  assign o[19535] = i[19535];
  assign o[19534] = i[19534];
  assign o[19533] = i[19533];
  assign o[19532] = i[19532];
  assign o[19531] = i[19531];
  assign o[19530] = i[19530];
  assign o[19529] = i[19529];
  assign o[19528] = i[19528];
  assign o[19527] = i[19527];
  assign o[19526] = i[19526];
  assign o[19525] = i[19525];
  assign o[19524] = i[19524];
  assign o[19523] = i[19523];
  assign o[19522] = i[19522];
  assign o[19521] = i[19521];
  assign o[19520] = i[19520];
  assign o[19519] = i[19519];
  assign o[19518] = i[19518];
  assign o[19517] = i[19517];
  assign o[19516] = i[19516];
  assign o[19515] = i[19515];
  assign o[19514] = i[19514];
  assign o[19513] = i[19513];
  assign o[19512] = i[19512];
  assign o[19511] = i[19511];
  assign o[19510] = i[19510];
  assign o[19509] = i[19509];
  assign o[19508] = i[19508];
  assign o[19507] = i[19507];
  assign o[19506] = i[19506];
  assign o[19505] = i[19505];
  assign o[19504] = i[19504];
  assign o[19503] = i[19503];
  assign o[19502] = i[19502];
  assign o[19501] = i[19501];
  assign o[19500] = i[19500];
  assign o[19499] = i[19499];
  assign o[19498] = i[19498];
  assign o[19497] = i[19497];
  assign o[19496] = i[19496];
  assign o[19495] = i[19495];
  assign o[19494] = i[19494];
  assign o[19493] = i[19493];
  assign o[19492] = i[19492];
  assign o[19491] = i[19491];
  assign o[19490] = i[19490];
  assign o[19489] = i[19489];
  assign o[19488] = i[19488];
  assign o[19487] = i[19487];
  assign o[19486] = i[19486];
  assign o[19485] = i[19485];
  assign o[19484] = i[19484];
  assign o[19483] = i[19483];
  assign o[19482] = i[19482];
  assign o[19481] = i[19481];
  assign o[19480] = i[19480];
  assign o[19479] = i[19479];
  assign o[19478] = i[19478];
  assign o[19477] = i[19477];
  assign o[19476] = i[19476];
  assign o[19475] = i[19475];
  assign o[19474] = i[19474];
  assign o[19473] = i[19473];
  assign o[19472] = i[19472];
  assign o[19471] = i[19471];
  assign o[19470] = i[19470];
  assign o[19469] = i[19469];
  assign o[19468] = i[19468];
  assign o[19467] = i[19467];
  assign o[19466] = i[19466];
  assign o[19465] = i[19465];
  assign o[19464] = i[19464];
  assign o[19463] = i[19463];
  assign o[19462] = i[19462];
  assign o[19461] = i[19461];
  assign o[19460] = i[19460];
  assign o[19459] = i[19459];
  assign o[19458] = i[19458];
  assign o[19457] = i[19457];
  assign o[19456] = i[19456];
  assign o[19455] = i[19455];
  assign o[19454] = i[19454];
  assign o[19453] = i[19453];
  assign o[19452] = i[19452];
  assign o[19451] = i[19451];
  assign o[19450] = i[19450];
  assign o[19449] = i[19449];
  assign o[19448] = i[19448];
  assign o[19447] = i[19447];
  assign o[19446] = i[19446];
  assign o[19445] = i[19445];
  assign o[19444] = i[19444];
  assign o[19443] = i[19443];
  assign o[19442] = i[19442];
  assign o[19441] = i[19441];
  assign o[19440] = i[19440];
  assign o[19439] = i[19439];
  assign o[19438] = i[19438];
  assign o[19437] = i[19437];
  assign o[19436] = i[19436];
  assign o[19435] = i[19435];
  assign o[19434] = i[19434];
  assign o[19433] = i[19433];
  assign o[19432] = i[19432];
  assign o[19431] = i[19431];
  assign o[19430] = i[19430];
  assign o[19429] = i[19429];
  assign o[19428] = i[19428];
  assign o[19427] = i[19427];
  assign o[19426] = i[19426];
  assign o[19425] = i[19425];
  assign o[19424] = i[19424];
  assign o[19423] = i[19423];
  assign o[19422] = i[19422];
  assign o[19421] = i[19421];
  assign o[19420] = i[19420];
  assign o[19419] = i[19419];
  assign o[19418] = i[19418];
  assign o[19417] = i[19417];
  assign o[19416] = i[19416];
  assign o[19415] = i[19415];
  assign o[19414] = i[19414];
  assign o[19413] = i[19413];
  assign o[19412] = i[19412];
  assign o[19411] = i[19411];
  assign o[19410] = i[19410];
  assign o[19409] = i[19409];
  assign o[19408] = i[19408];
  assign o[19407] = i[19407];
  assign o[19406] = i[19406];
  assign o[19405] = i[19405];
  assign o[19404] = i[19404];
  assign o[19403] = i[19403];
  assign o[19402] = i[19402];
  assign o[19401] = i[19401];
  assign o[19400] = i[19400];
  assign o[19399] = i[19399];
  assign o[19398] = i[19398];
  assign o[19397] = i[19397];
  assign o[19396] = i[19396];
  assign o[19395] = i[19395];
  assign o[19394] = i[19394];
  assign o[19393] = i[19393];
  assign o[19392] = i[19392];
  assign o[19391] = i[19391];
  assign o[19390] = i[19390];
  assign o[19389] = i[19389];
  assign o[19388] = i[19388];
  assign o[19387] = i[19387];
  assign o[19386] = i[19386];
  assign o[19385] = i[19385];
  assign o[19384] = i[19384];
  assign o[19383] = i[19383];
  assign o[19382] = i[19382];
  assign o[19381] = i[19381];
  assign o[19380] = i[19380];
  assign o[19379] = i[19379];
  assign o[19378] = i[19378];
  assign o[19377] = i[19377];
  assign o[19376] = i[19376];
  assign o[19375] = i[19375];
  assign o[19374] = i[19374];
  assign o[19373] = i[19373];
  assign o[19372] = i[19372];
  assign o[19371] = i[19371];
  assign o[19370] = i[19370];
  assign o[19369] = i[19369];
  assign o[19368] = i[19368];
  assign o[19367] = i[19367];
  assign o[19366] = i[19366];
  assign o[19365] = i[19365];
  assign o[19364] = i[19364];
  assign o[19363] = i[19363];
  assign o[19362] = i[19362];
  assign o[19361] = i[19361];
  assign o[19360] = i[19360];
  assign o[19359] = i[19359];
  assign o[19358] = i[19358];
  assign o[19357] = i[19357];
  assign o[19356] = i[19356];
  assign o[19355] = i[19355];
  assign o[19354] = i[19354];
  assign o[19353] = i[19353];
  assign o[19352] = i[19352];
  assign o[19351] = i[19351];
  assign o[19350] = i[19350];
  assign o[19349] = i[19349];
  assign o[19348] = i[19348];
  assign o[19347] = i[19347];
  assign o[19346] = i[19346];
  assign o[19345] = i[19345];
  assign o[19344] = i[19344];
  assign o[19343] = i[19343];
  assign o[19342] = i[19342];
  assign o[19341] = i[19341];
  assign o[19340] = i[19340];
  assign o[19339] = i[19339];
  assign o[19338] = i[19338];
  assign o[19337] = i[19337];
  assign o[19336] = i[19336];
  assign o[19335] = i[19335];
  assign o[19334] = i[19334];
  assign o[19333] = i[19333];
  assign o[19332] = i[19332];
  assign o[19331] = i[19331];
  assign o[19330] = i[19330];
  assign o[19329] = i[19329];
  assign o[19328] = i[19328];
  assign o[19327] = i[19327];
  assign o[19326] = i[19326];
  assign o[19325] = i[19325];
  assign o[19324] = i[19324];
  assign o[19323] = i[19323];
  assign o[19322] = i[19322];
  assign o[19321] = i[19321];
  assign o[19320] = i[19320];
  assign o[19319] = i[19319];
  assign o[19318] = i[19318];
  assign o[19317] = i[19317];
  assign o[19316] = i[19316];
  assign o[19315] = i[19315];
  assign o[19314] = i[19314];
  assign o[19313] = i[19313];
  assign o[19312] = i[19312];
  assign o[19311] = i[19311];
  assign o[19310] = i[19310];
  assign o[19309] = i[19309];
  assign o[19308] = i[19308];
  assign o[19307] = i[19307];
  assign o[19306] = i[19306];
  assign o[19305] = i[19305];
  assign o[19304] = i[19304];
  assign o[19303] = i[19303];
  assign o[19302] = i[19302];
  assign o[19301] = i[19301];
  assign o[19300] = i[19300];
  assign o[19299] = i[19299];
  assign o[19298] = i[19298];
  assign o[19297] = i[19297];
  assign o[19296] = i[19296];
  assign o[19295] = i[19295];
  assign o[19294] = i[19294];
  assign o[19293] = i[19293];
  assign o[19292] = i[19292];
  assign o[19291] = i[19291];
  assign o[19290] = i[19290];
  assign o[19289] = i[19289];
  assign o[19288] = i[19288];
  assign o[19287] = i[19287];
  assign o[19286] = i[19286];
  assign o[19285] = i[19285];
  assign o[19284] = i[19284];
  assign o[19283] = i[19283];
  assign o[19282] = i[19282];
  assign o[19281] = i[19281];
  assign o[19280] = i[19280];
  assign o[19279] = i[19279];
  assign o[19278] = i[19278];
  assign o[19277] = i[19277];
  assign o[19276] = i[19276];
  assign o[19275] = i[19275];
  assign o[19274] = i[19274];
  assign o[19273] = i[19273];
  assign o[19272] = i[19272];
  assign o[19271] = i[19271];
  assign o[19270] = i[19270];
  assign o[19269] = i[19269];
  assign o[19268] = i[19268];
  assign o[19267] = i[19267];
  assign o[19266] = i[19266];
  assign o[19265] = i[19265];
  assign o[19264] = i[19264];
  assign o[19263] = i[19263];
  assign o[19262] = i[19262];
  assign o[19261] = i[19261];
  assign o[19260] = i[19260];
  assign o[19259] = i[19259];
  assign o[19258] = i[19258];
  assign o[19257] = i[19257];
  assign o[19256] = i[19256];
  assign o[19255] = i[19255];
  assign o[19254] = i[19254];
  assign o[19253] = i[19253];
  assign o[19252] = i[19252];
  assign o[19251] = i[19251];
  assign o[19250] = i[19250];
  assign o[19249] = i[19249];
  assign o[19248] = i[19248];
  assign o[19247] = i[19247];
  assign o[19246] = i[19246];
  assign o[19245] = i[19245];
  assign o[19244] = i[19244];
  assign o[19243] = i[19243];
  assign o[19242] = i[19242];
  assign o[19241] = i[19241];
  assign o[19240] = i[19240];
  assign o[19239] = i[19239];
  assign o[19238] = i[19238];
  assign o[19237] = i[19237];
  assign o[19236] = i[19236];
  assign o[19235] = i[19235];
  assign o[19234] = i[19234];
  assign o[19233] = i[19233];
  assign o[19232] = i[19232];
  assign o[19231] = i[19231];
  assign o[19230] = i[19230];
  assign o[19229] = i[19229];
  assign o[19228] = i[19228];
  assign o[19227] = i[19227];
  assign o[19226] = i[19226];
  assign o[19225] = i[19225];
  assign o[19224] = i[19224];
  assign o[19223] = i[19223];
  assign o[19222] = i[19222];
  assign o[19221] = i[19221];
  assign o[19220] = i[19220];
  assign o[19219] = i[19219];
  assign o[19218] = i[19218];
  assign o[19217] = i[19217];
  assign o[19216] = i[19216];
  assign o[19215] = i[19215];
  assign o[19214] = i[19214];
  assign o[19213] = i[19213];
  assign o[19212] = i[19212];
  assign o[19211] = i[19211];
  assign o[19210] = i[19210];
  assign o[19209] = i[19209];
  assign o[19208] = i[19208];
  assign o[19207] = i[19207];
  assign o[19206] = i[19206];
  assign o[19205] = i[19205];
  assign o[19204] = i[19204];
  assign o[19203] = i[19203];
  assign o[19202] = i[19202];
  assign o[19201] = i[19201];
  assign o[19200] = i[19200];
  assign o[19199] = i[19199];
  assign o[19198] = i[19198];
  assign o[19197] = i[19197];
  assign o[19196] = i[19196];
  assign o[19195] = i[19195];
  assign o[19194] = i[19194];
  assign o[19193] = i[19193];
  assign o[19192] = i[19192];
  assign o[19191] = i[19191];
  assign o[19190] = i[19190];
  assign o[19189] = i[19189];
  assign o[19188] = i[19188];
  assign o[19187] = i[19187];
  assign o[19186] = i[19186];
  assign o[19185] = i[19185];
  assign o[19184] = i[19184];
  assign o[19183] = i[19183];
  assign o[19182] = i[19182];
  assign o[19181] = i[19181];
  assign o[19180] = i[19180];
  assign o[19179] = i[19179];
  assign o[19178] = i[19178];
  assign o[19177] = i[19177];
  assign o[19176] = i[19176];
  assign o[19175] = i[19175];
  assign o[19174] = i[19174];
  assign o[19173] = i[19173];
  assign o[19172] = i[19172];
  assign o[19171] = i[19171];
  assign o[19170] = i[19170];
  assign o[19169] = i[19169];
  assign o[19168] = i[19168];
  assign o[19167] = i[19167];
  assign o[19166] = i[19166];
  assign o[19165] = i[19165];
  assign o[19164] = i[19164];
  assign o[19163] = i[19163];
  assign o[19162] = i[19162];
  assign o[19161] = i[19161];
  assign o[19160] = i[19160];
  assign o[19159] = i[19159];
  assign o[19158] = i[19158];
  assign o[19157] = i[19157];
  assign o[19156] = i[19156];
  assign o[19155] = i[19155];
  assign o[19154] = i[19154];
  assign o[19153] = i[19153];
  assign o[19152] = i[19152];
  assign o[19151] = i[19151];
  assign o[19150] = i[19150];
  assign o[19149] = i[19149];
  assign o[19148] = i[19148];
  assign o[19147] = i[19147];
  assign o[19146] = i[19146];
  assign o[19145] = i[19145];
  assign o[19144] = i[19144];
  assign o[19143] = i[19143];
  assign o[19142] = i[19142];
  assign o[19141] = i[19141];
  assign o[19140] = i[19140];
  assign o[19139] = i[19139];
  assign o[19138] = i[19138];
  assign o[19137] = i[19137];
  assign o[19136] = i[19136];
  assign o[19135] = i[19135];
  assign o[19134] = i[19134];
  assign o[19133] = i[19133];
  assign o[19132] = i[19132];
  assign o[19131] = i[19131];
  assign o[19130] = i[19130];
  assign o[19129] = i[19129];
  assign o[19128] = i[19128];
  assign o[19127] = i[19127];
  assign o[19126] = i[19126];
  assign o[19125] = i[19125];
  assign o[19124] = i[19124];
  assign o[19123] = i[19123];
  assign o[19122] = i[19122];
  assign o[19121] = i[19121];
  assign o[19120] = i[19120];
  assign o[19119] = i[19119];
  assign o[19118] = i[19118];
  assign o[19117] = i[19117];
  assign o[19116] = i[19116];
  assign o[19115] = i[19115];
  assign o[19114] = i[19114];
  assign o[19113] = i[19113];
  assign o[19112] = i[19112];
  assign o[19111] = i[19111];
  assign o[19110] = i[19110];
  assign o[19109] = i[19109];
  assign o[19108] = i[19108];
  assign o[19107] = i[19107];
  assign o[19106] = i[19106];
  assign o[19105] = i[19105];
  assign o[19104] = i[19104];
  assign o[19103] = i[19103];
  assign o[19102] = i[19102];
  assign o[19101] = i[19101];
  assign o[19100] = i[19100];
  assign o[19099] = i[19099];
  assign o[19098] = i[19098];
  assign o[19097] = i[19097];
  assign o[19096] = i[19096];
  assign o[19095] = i[19095];
  assign o[19094] = i[19094];
  assign o[19093] = i[19093];
  assign o[19092] = i[19092];
  assign o[19091] = i[19091];
  assign o[19090] = i[19090];
  assign o[19089] = i[19089];
  assign o[19088] = i[19088];
  assign o[19087] = i[19087];
  assign o[19086] = i[19086];
  assign o[19085] = i[19085];
  assign o[19084] = i[19084];
  assign o[19083] = i[19083];
  assign o[19082] = i[19082];
  assign o[19081] = i[19081];
  assign o[19080] = i[19080];
  assign o[19079] = i[19079];
  assign o[19078] = i[19078];
  assign o[19077] = i[19077];
  assign o[19076] = i[19076];
  assign o[19075] = i[19075];
  assign o[19074] = i[19074];
  assign o[19073] = i[19073];
  assign o[19072] = i[19072];
  assign o[19071] = i[19071];
  assign o[19070] = i[19070];
  assign o[19069] = i[19069];
  assign o[19068] = i[19068];
  assign o[19067] = i[19067];
  assign o[19066] = i[19066];
  assign o[19065] = i[19065];
  assign o[19064] = i[19064];
  assign o[19063] = i[19063];
  assign o[19062] = i[19062];
  assign o[19061] = i[19061];
  assign o[19060] = i[19060];
  assign o[19059] = i[19059];
  assign o[19058] = i[19058];
  assign o[19057] = i[19057];
  assign o[19056] = i[19056];
  assign o[19055] = i[19055];
  assign o[19054] = i[19054];
  assign o[19053] = i[19053];
  assign o[19052] = i[19052];
  assign o[19051] = i[19051];
  assign o[19050] = i[19050];
  assign o[19049] = i[19049];
  assign o[19048] = i[19048];
  assign o[19047] = i[19047];
  assign o[19046] = i[19046];
  assign o[19045] = i[19045];
  assign o[19044] = i[19044];
  assign o[19043] = i[19043];
  assign o[19042] = i[19042];
  assign o[19041] = i[19041];
  assign o[19040] = i[19040];
  assign o[19039] = i[19039];
  assign o[19038] = i[19038];
  assign o[19037] = i[19037];
  assign o[19036] = i[19036];
  assign o[19035] = i[19035];
  assign o[19034] = i[19034];
  assign o[19033] = i[19033];
  assign o[19032] = i[19032];
  assign o[19031] = i[19031];
  assign o[19030] = i[19030];
  assign o[19029] = i[19029];
  assign o[19028] = i[19028];
  assign o[19027] = i[19027];
  assign o[19026] = i[19026];
  assign o[19025] = i[19025];
  assign o[19024] = i[19024];
  assign o[19023] = i[19023];
  assign o[19022] = i[19022];
  assign o[19021] = i[19021];
  assign o[19020] = i[19020];
  assign o[19019] = i[19019];
  assign o[19018] = i[19018];
  assign o[19017] = i[19017];
  assign o[19016] = i[19016];
  assign o[19015] = i[19015];
  assign o[19014] = i[19014];
  assign o[19013] = i[19013];
  assign o[19012] = i[19012];
  assign o[19011] = i[19011];
  assign o[19010] = i[19010];
  assign o[19009] = i[19009];
  assign o[19008] = i[19008];
  assign o[19007] = i[19007];
  assign o[19006] = i[19006];
  assign o[19005] = i[19005];
  assign o[19004] = i[19004];
  assign o[19003] = i[19003];
  assign o[19002] = i[19002];
  assign o[19001] = i[19001];
  assign o[19000] = i[19000];
  assign o[18999] = i[18999];
  assign o[18998] = i[18998];
  assign o[18997] = i[18997];
  assign o[18996] = i[18996];
  assign o[18995] = i[18995];
  assign o[18994] = i[18994];
  assign o[18993] = i[18993];
  assign o[18992] = i[18992];
  assign o[18991] = i[18991];
  assign o[18990] = i[18990];
  assign o[18989] = i[18989];
  assign o[18988] = i[18988];
  assign o[18987] = i[18987];
  assign o[18986] = i[18986];
  assign o[18985] = i[18985];
  assign o[18984] = i[18984];
  assign o[18983] = i[18983];
  assign o[18982] = i[18982];
  assign o[18981] = i[18981];
  assign o[18980] = i[18980];
  assign o[18979] = i[18979];
  assign o[18978] = i[18978];
  assign o[18977] = i[18977];
  assign o[18976] = i[18976];
  assign o[18975] = i[18975];
  assign o[18974] = i[18974];
  assign o[18973] = i[18973];
  assign o[18972] = i[18972];
  assign o[18971] = i[18971];
  assign o[18970] = i[18970];
  assign o[18969] = i[18969];
  assign o[18968] = i[18968];
  assign o[18967] = i[18967];
  assign o[18966] = i[18966];
  assign o[18965] = i[18965];
  assign o[18964] = i[18964];
  assign o[18963] = i[18963];
  assign o[18962] = i[18962];
  assign o[18961] = i[18961];
  assign o[18960] = i[18960];
  assign o[18959] = i[18959];
  assign o[18958] = i[18958];
  assign o[18957] = i[18957];
  assign o[18956] = i[18956];
  assign o[18955] = i[18955];
  assign o[18954] = i[18954];
  assign o[18953] = i[18953];
  assign o[18952] = i[18952];
  assign o[18951] = i[18951];
  assign o[18950] = i[18950];
  assign o[18949] = i[18949];
  assign o[18948] = i[18948];
  assign o[18947] = i[18947];
  assign o[18946] = i[18946];
  assign o[18945] = i[18945];
  assign o[18944] = i[18944];
  assign o[18943] = i[18943];
  assign o[18942] = i[18942];
  assign o[18941] = i[18941];
  assign o[18940] = i[18940];
  assign o[18939] = i[18939];
  assign o[18938] = i[18938];
  assign o[18937] = i[18937];
  assign o[18936] = i[18936];
  assign o[18935] = i[18935];
  assign o[18934] = i[18934];
  assign o[18933] = i[18933];
  assign o[18932] = i[18932];
  assign o[18931] = i[18931];
  assign o[18930] = i[18930];
  assign o[18929] = i[18929];
  assign o[18928] = i[18928];
  assign o[18927] = i[18927];
  assign o[18926] = i[18926];
  assign o[18925] = i[18925];
  assign o[18924] = i[18924];
  assign o[18923] = i[18923];
  assign o[18922] = i[18922];
  assign o[18921] = i[18921];
  assign o[18920] = i[18920];
  assign o[18919] = i[18919];
  assign o[18918] = i[18918];
  assign o[18917] = i[18917];
  assign o[18916] = i[18916];
  assign o[18915] = i[18915];
  assign o[18914] = i[18914];
  assign o[18913] = i[18913];
  assign o[18912] = i[18912];
  assign o[18911] = i[18911];
  assign o[18910] = i[18910];
  assign o[18909] = i[18909];
  assign o[18908] = i[18908];
  assign o[18907] = i[18907];
  assign o[18906] = i[18906];
  assign o[18905] = i[18905];
  assign o[18904] = i[18904];
  assign o[18903] = i[18903];
  assign o[18902] = i[18902];
  assign o[18901] = i[18901];
  assign o[18900] = i[18900];
  assign o[18899] = i[18899];
  assign o[18898] = i[18898];
  assign o[18897] = i[18897];
  assign o[18896] = i[18896];
  assign o[18895] = i[18895];
  assign o[18894] = i[18894];
  assign o[18893] = i[18893];
  assign o[18892] = i[18892];
  assign o[18891] = i[18891];
  assign o[18890] = i[18890];
  assign o[18889] = i[18889];
  assign o[18888] = i[18888];
  assign o[18887] = i[18887];
  assign o[18886] = i[18886];
  assign o[18885] = i[18885];
  assign o[18884] = i[18884];
  assign o[18883] = i[18883];
  assign o[18882] = i[18882];
  assign o[18881] = i[18881];
  assign o[18880] = i[18880];
  assign o[18879] = i[18879];
  assign o[18878] = i[18878];
  assign o[18877] = i[18877];
  assign o[18876] = i[18876];
  assign o[18875] = i[18875];
  assign o[18874] = i[18874];
  assign o[18873] = i[18873];
  assign o[18872] = i[18872];
  assign o[18871] = i[18871];
  assign o[18870] = i[18870];
  assign o[18869] = i[18869];
  assign o[18868] = i[18868];
  assign o[18867] = i[18867];
  assign o[18866] = i[18866];
  assign o[18865] = i[18865];
  assign o[18864] = i[18864];
  assign o[18863] = i[18863];
  assign o[18862] = i[18862];
  assign o[18861] = i[18861];
  assign o[18860] = i[18860];
  assign o[18859] = i[18859];
  assign o[18858] = i[18858];
  assign o[18857] = i[18857];
  assign o[18856] = i[18856];
  assign o[18855] = i[18855];
  assign o[18854] = i[18854];
  assign o[18853] = i[18853];
  assign o[18852] = i[18852];
  assign o[18851] = i[18851];
  assign o[18850] = i[18850];
  assign o[18849] = i[18849];
  assign o[18848] = i[18848];
  assign o[18847] = i[18847];
  assign o[18846] = i[18846];
  assign o[18845] = i[18845];
  assign o[18844] = i[18844];
  assign o[18843] = i[18843];
  assign o[18842] = i[18842];
  assign o[18841] = i[18841];
  assign o[18840] = i[18840];
  assign o[18839] = i[18839];
  assign o[18838] = i[18838];
  assign o[18837] = i[18837];
  assign o[18836] = i[18836];
  assign o[18835] = i[18835];
  assign o[18834] = i[18834];
  assign o[18833] = i[18833];
  assign o[18832] = i[18832];
  assign o[18831] = i[18831];
  assign o[18830] = i[18830];
  assign o[18829] = i[18829];
  assign o[18828] = i[18828];
  assign o[18827] = i[18827];
  assign o[18826] = i[18826];
  assign o[18825] = i[18825];
  assign o[18824] = i[18824];
  assign o[18823] = i[18823];
  assign o[18822] = i[18822];
  assign o[18821] = i[18821];
  assign o[18820] = i[18820];
  assign o[18819] = i[18819];
  assign o[18818] = i[18818];
  assign o[18817] = i[18817];
  assign o[18816] = i[18816];
  assign o[18815] = i[18815];
  assign o[18814] = i[18814];
  assign o[18813] = i[18813];
  assign o[18812] = i[18812];
  assign o[18811] = i[18811];
  assign o[18810] = i[18810];
  assign o[18809] = i[18809];
  assign o[18808] = i[18808];
  assign o[18807] = i[18807];
  assign o[18806] = i[18806];
  assign o[18805] = i[18805];
  assign o[18804] = i[18804];
  assign o[18803] = i[18803];
  assign o[18802] = i[18802];
  assign o[18801] = i[18801];
  assign o[18800] = i[18800];
  assign o[18799] = i[18799];
  assign o[18798] = i[18798];
  assign o[18797] = i[18797];
  assign o[18796] = i[18796];
  assign o[18795] = i[18795];
  assign o[18794] = i[18794];
  assign o[18793] = i[18793];
  assign o[18792] = i[18792];
  assign o[18791] = i[18791];
  assign o[18790] = i[18790];
  assign o[18789] = i[18789];
  assign o[18788] = i[18788];
  assign o[18787] = i[18787];
  assign o[18786] = i[18786];
  assign o[18785] = i[18785];
  assign o[18784] = i[18784];
  assign o[18783] = i[18783];
  assign o[18782] = i[18782];
  assign o[18781] = i[18781];
  assign o[18780] = i[18780];
  assign o[18779] = i[18779];
  assign o[18778] = i[18778];
  assign o[18777] = i[18777];
  assign o[18776] = i[18776];
  assign o[18775] = i[18775];
  assign o[18774] = i[18774];
  assign o[18773] = i[18773];
  assign o[18772] = i[18772];
  assign o[18771] = i[18771];
  assign o[18770] = i[18770];
  assign o[18769] = i[18769];
  assign o[18768] = i[18768];
  assign o[18767] = i[18767];
  assign o[18766] = i[18766];
  assign o[18765] = i[18765];
  assign o[18764] = i[18764];
  assign o[18763] = i[18763];
  assign o[18762] = i[18762];
  assign o[18761] = i[18761];
  assign o[18760] = i[18760];
  assign o[18759] = i[18759];
  assign o[18758] = i[18758];
  assign o[18757] = i[18757];
  assign o[18756] = i[18756];
  assign o[18755] = i[18755];
  assign o[18754] = i[18754];
  assign o[18753] = i[18753];
  assign o[18752] = i[18752];
  assign o[18751] = i[18751];
  assign o[18750] = i[18750];
  assign o[18749] = i[18749];
  assign o[18748] = i[18748];
  assign o[18747] = i[18747];
  assign o[18746] = i[18746];
  assign o[18745] = i[18745];
  assign o[18744] = i[18744];
  assign o[18743] = i[18743];
  assign o[18742] = i[18742];
  assign o[18741] = i[18741];
  assign o[18740] = i[18740];
  assign o[18739] = i[18739];
  assign o[18738] = i[18738];
  assign o[18737] = i[18737];
  assign o[18736] = i[18736];
  assign o[18735] = i[18735];
  assign o[18734] = i[18734];
  assign o[18733] = i[18733];
  assign o[18732] = i[18732];
  assign o[18731] = i[18731];
  assign o[18730] = i[18730];
  assign o[18729] = i[18729];
  assign o[18728] = i[18728];
  assign o[18727] = i[18727];
  assign o[18726] = i[18726];
  assign o[18725] = i[18725];
  assign o[18724] = i[18724];
  assign o[18723] = i[18723];
  assign o[18722] = i[18722];
  assign o[18721] = i[18721];
  assign o[18720] = i[18720];
  assign o[18719] = i[18719];
  assign o[18718] = i[18718];
  assign o[18717] = i[18717];
  assign o[18716] = i[18716];
  assign o[18715] = i[18715];
  assign o[18714] = i[18714];
  assign o[18713] = i[18713];
  assign o[18712] = i[18712];
  assign o[18711] = i[18711];
  assign o[18710] = i[18710];
  assign o[18709] = i[18709];
  assign o[18708] = i[18708];
  assign o[18707] = i[18707];
  assign o[18706] = i[18706];
  assign o[18705] = i[18705];
  assign o[18704] = i[18704];
  assign o[18703] = i[18703];
  assign o[18702] = i[18702];
  assign o[18701] = i[18701];
  assign o[18700] = i[18700];
  assign o[18699] = i[18699];
  assign o[18698] = i[18698];
  assign o[18697] = i[18697];
  assign o[18696] = i[18696];
  assign o[18695] = i[18695];
  assign o[18694] = i[18694];
  assign o[18693] = i[18693];
  assign o[18692] = i[18692];
  assign o[18691] = i[18691];
  assign o[18690] = i[18690];
  assign o[18689] = i[18689];
  assign o[18688] = i[18688];
  assign o[18687] = i[18687];
  assign o[18686] = i[18686];
  assign o[18685] = i[18685];
  assign o[18684] = i[18684];
  assign o[18683] = i[18683];
  assign o[18682] = i[18682];
  assign o[18681] = i[18681];
  assign o[18680] = i[18680];
  assign o[18679] = i[18679];
  assign o[18678] = i[18678];
  assign o[18677] = i[18677];
  assign o[18676] = i[18676];
  assign o[18675] = i[18675];
  assign o[18674] = i[18674];
  assign o[18673] = i[18673];
  assign o[18672] = i[18672];
  assign o[18671] = i[18671];
  assign o[18670] = i[18670];
  assign o[18669] = i[18669];
  assign o[18668] = i[18668];
  assign o[18667] = i[18667];
  assign o[18666] = i[18666];
  assign o[18665] = i[18665];
  assign o[18664] = i[18664];
  assign o[18663] = i[18663];
  assign o[18662] = i[18662];
  assign o[18661] = i[18661];
  assign o[18660] = i[18660];
  assign o[18659] = i[18659];
  assign o[18658] = i[18658];
  assign o[18657] = i[18657];
  assign o[18656] = i[18656];
  assign o[18655] = i[18655];
  assign o[18654] = i[18654];
  assign o[18653] = i[18653];
  assign o[18652] = i[18652];
  assign o[18651] = i[18651];
  assign o[18650] = i[18650];
  assign o[18649] = i[18649];
  assign o[18648] = i[18648];
  assign o[18647] = i[18647];
  assign o[18646] = i[18646];
  assign o[18645] = i[18645];
  assign o[18644] = i[18644];
  assign o[18643] = i[18643];
  assign o[18642] = i[18642];
  assign o[18641] = i[18641];
  assign o[18640] = i[18640];
  assign o[18639] = i[18639];
  assign o[18638] = i[18638];
  assign o[18637] = i[18637];
  assign o[18636] = i[18636];
  assign o[18635] = i[18635];
  assign o[18634] = i[18634];
  assign o[18633] = i[18633];
  assign o[18632] = i[18632];
  assign o[18631] = i[18631];
  assign o[18630] = i[18630];
  assign o[18629] = i[18629];
  assign o[18628] = i[18628];
  assign o[18627] = i[18627];
  assign o[18626] = i[18626];
  assign o[18625] = i[18625];
  assign o[18624] = i[18624];
  assign o[18623] = i[18623];
  assign o[18622] = i[18622];
  assign o[18621] = i[18621];
  assign o[18620] = i[18620];
  assign o[18619] = i[18619];
  assign o[18618] = i[18618];
  assign o[18617] = i[18617];
  assign o[18616] = i[18616];
  assign o[18615] = i[18615];
  assign o[18614] = i[18614];
  assign o[18613] = i[18613];
  assign o[18612] = i[18612];
  assign o[18611] = i[18611];
  assign o[18610] = i[18610];
  assign o[18609] = i[18609];
  assign o[18608] = i[18608];
  assign o[18607] = i[18607];
  assign o[18606] = i[18606];
  assign o[18605] = i[18605];
  assign o[18604] = i[18604];
  assign o[18603] = i[18603];
  assign o[18602] = i[18602];
  assign o[18601] = i[18601];
  assign o[18600] = i[18600];
  assign o[18599] = i[18599];
  assign o[18598] = i[18598];
  assign o[18597] = i[18597];
  assign o[18596] = i[18596];
  assign o[18595] = i[18595];
  assign o[18594] = i[18594];
  assign o[18593] = i[18593];
  assign o[18592] = i[18592];
  assign o[18591] = i[18591];
  assign o[18590] = i[18590];
  assign o[18589] = i[18589];
  assign o[18588] = i[18588];
  assign o[18587] = i[18587];
  assign o[18586] = i[18586];
  assign o[18585] = i[18585];
  assign o[18584] = i[18584];
  assign o[18583] = i[18583];
  assign o[18582] = i[18582];
  assign o[18581] = i[18581];
  assign o[18580] = i[18580];
  assign o[18579] = i[18579];
  assign o[18578] = i[18578];
  assign o[18577] = i[18577];
  assign o[18576] = i[18576];
  assign o[18575] = i[18575];
  assign o[18574] = i[18574];
  assign o[18573] = i[18573];
  assign o[18572] = i[18572];
  assign o[18571] = i[18571];
  assign o[18570] = i[18570];
  assign o[18569] = i[18569];
  assign o[18568] = i[18568];
  assign o[18567] = i[18567];
  assign o[18566] = i[18566];
  assign o[18565] = i[18565];
  assign o[18564] = i[18564];
  assign o[18563] = i[18563];
  assign o[18562] = i[18562];
  assign o[18561] = i[18561];
  assign o[18560] = i[18560];
  assign o[18559] = i[18559];
  assign o[18558] = i[18558];
  assign o[18557] = i[18557];
  assign o[18556] = i[18556];
  assign o[18555] = i[18555];
  assign o[18554] = i[18554];
  assign o[18553] = i[18553];
  assign o[18552] = i[18552];
  assign o[18551] = i[18551];
  assign o[18550] = i[18550];
  assign o[18549] = i[18549];
  assign o[18548] = i[18548];
  assign o[18547] = i[18547];
  assign o[18546] = i[18546];
  assign o[18545] = i[18545];
  assign o[18544] = i[18544];
  assign o[18543] = i[18543];
  assign o[18542] = i[18542];
  assign o[18541] = i[18541];
  assign o[18540] = i[18540];
  assign o[18539] = i[18539];
  assign o[18538] = i[18538];
  assign o[18537] = i[18537];
  assign o[18536] = i[18536];
  assign o[18535] = i[18535];
  assign o[18534] = i[18534];
  assign o[18533] = i[18533];
  assign o[18532] = i[18532];
  assign o[18531] = i[18531];
  assign o[18530] = i[18530];
  assign o[18529] = i[18529];
  assign o[18528] = i[18528];
  assign o[18527] = i[18527];
  assign o[18526] = i[18526];
  assign o[18525] = i[18525];
  assign o[18524] = i[18524];
  assign o[18523] = i[18523];
  assign o[18522] = i[18522];
  assign o[18521] = i[18521];
  assign o[18520] = i[18520];
  assign o[18519] = i[18519];
  assign o[18518] = i[18518];
  assign o[18517] = i[18517];
  assign o[18516] = i[18516];
  assign o[18515] = i[18515];
  assign o[18514] = i[18514];
  assign o[18513] = i[18513];
  assign o[18512] = i[18512];
  assign o[18511] = i[18511];
  assign o[18510] = i[18510];
  assign o[18509] = i[18509];
  assign o[18508] = i[18508];
  assign o[18507] = i[18507];
  assign o[18506] = i[18506];
  assign o[18505] = i[18505];
  assign o[18504] = i[18504];
  assign o[18503] = i[18503];
  assign o[18502] = i[18502];
  assign o[18501] = i[18501];
  assign o[18500] = i[18500];
  assign o[18499] = i[18499];
  assign o[18498] = i[18498];
  assign o[18497] = i[18497];
  assign o[18496] = i[18496];
  assign o[18495] = i[18495];
  assign o[18494] = i[18494];
  assign o[18493] = i[18493];
  assign o[18492] = i[18492];
  assign o[18491] = i[18491];
  assign o[18490] = i[18490];
  assign o[18489] = i[18489];
  assign o[18488] = i[18488];
  assign o[18487] = i[18487];
  assign o[18486] = i[18486];
  assign o[18485] = i[18485];
  assign o[18484] = i[18484];
  assign o[18483] = i[18483];
  assign o[18482] = i[18482];
  assign o[18481] = i[18481];
  assign o[18480] = i[18480];
  assign o[18479] = i[18479];
  assign o[18478] = i[18478];
  assign o[18477] = i[18477];
  assign o[18476] = i[18476];
  assign o[18475] = i[18475];
  assign o[18474] = i[18474];
  assign o[18473] = i[18473];
  assign o[18472] = i[18472];
  assign o[18471] = i[18471];
  assign o[18470] = i[18470];
  assign o[18469] = i[18469];
  assign o[18468] = i[18468];
  assign o[18467] = i[18467];
  assign o[18466] = i[18466];
  assign o[18465] = i[18465];
  assign o[18464] = i[18464];
  assign o[18463] = i[18463];
  assign o[18462] = i[18462];
  assign o[18461] = i[18461];
  assign o[18460] = i[18460];
  assign o[18459] = i[18459];
  assign o[18458] = i[18458];
  assign o[18457] = i[18457];
  assign o[18456] = i[18456];
  assign o[18455] = i[18455];
  assign o[18454] = i[18454];
  assign o[18453] = i[18453];
  assign o[18452] = i[18452];
  assign o[18451] = i[18451];
  assign o[18450] = i[18450];
  assign o[18449] = i[18449];
  assign o[18448] = i[18448];
  assign o[18447] = i[18447];
  assign o[18446] = i[18446];
  assign o[18445] = i[18445];
  assign o[18444] = i[18444];
  assign o[18443] = i[18443];
  assign o[18442] = i[18442];
  assign o[18441] = i[18441];
  assign o[18440] = i[18440];
  assign o[18439] = i[18439];
  assign o[18438] = i[18438];
  assign o[18437] = i[18437];
  assign o[18436] = i[18436];
  assign o[18435] = i[18435];
  assign o[18434] = i[18434];
  assign o[18433] = i[18433];
  assign o[18432] = i[18432];
  assign o[18431] = i[18431];
  assign o[18430] = i[18430];
  assign o[18429] = i[18429];
  assign o[18428] = i[18428];
  assign o[18427] = i[18427];
  assign o[18426] = i[18426];
  assign o[18425] = i[18425];
  assign o[18424] = i[18424];
  assign o[18423] = i[18423];
  assign o[18422] = i[18422];
  assign o[18421] = i[18421];
  assign o[18420] = i[18420];
  assign o[18419] = i[18419];
  assign o[18418] = i[18418];
  assign o[18417] = i[18417];
  assign o[18416] = i[18416];
  assign o[18415] = i[18415];
  assign o[18414] = i[18414];
  assign o[18413] = i[18413];
  assign o[18412] = i[18412];
  assign o[18411] = i[18411];
  assign o[18410] = i[18410];
  assign o[18409] = i[18409];
  assign o[18408] = i[18408];
  assign o[18407] = i[18407];
  assign o[18406] = i[18406];
  assign o[18405] = i[18405];
  assign o[18404] = i[18404];
  assign o[18403] = i[18403];
  assign o[18402] = i[18402];
  assign o[18401] = i[18401];
  assign o[18400] = i[18400];
  assign o[18399] = i[18399];
  assign o[18398] = i[18398];
  assign o[18397] = i[18397];
  assign o[18396] = i[18396];
  assign o[18395] = i[18395];
  assign o[18394] = i[18394];
  assign o[18393] = i[18393];
  assign o[18392] = i[18392];
  assign o[18391] = i[18391];
  assign o[18390] = i[18390];
  assign o[18389] = i[18389];
  assign o[18388] = i[18388];
  assign o[18387] = i[18387];
  assign o[18386] = i[18386];
  assign o[18385] = i[18385];
  assign o[18384] = i[18384];
  assign o[18383] = i[18383];
  assign o[18382] = i[18382];
  assign o[18381] = i[18381];
  assign o[18380] = i[18380];
  assign o[18379] = i[18379];
  assign o[18378] = i[18378];
  assign o[18377] = i[18377];
  assign o[18376] = i[18376];
  assign o[18375] = i[18375];
  assign o[18374] = i[18374];
  assign o[18373] = i[18373];
  assign o[18372] = i[18372];
  assign o[18371] = i[18371];
  assign o[18370] = i[18370];
  assign o[18369] = i[18369];
  assign o[18368] = i[18368];
  assign o[18367] = i[18367];
  assign o[18366] = i[18366];
  assign o[18365] = i[18365];
  assign o[18364] = i[18364];
  assign o[18363] = i[18363];
  assign o[18362] = i[18362];
  assign o[18361] = i[18361];
  assign o[18360] = i[18360];
  assign o[18359] = i[18359];
  assign o[18358] = i[18358];
  assign o[18357] = i[18357];
  assign o[18356] = i[18356];
  assign o[18355] = i[18355];
  assign o[18354] = i[18354];
  assign o[18353] = i[18353];
  assign o[18352] = i[18352];
  assign o[18351] = i[18351];
  assign o[18350] = i[18350];
  assign o[18349] = i[18349];
  assign o[18348] = i[18348];
  assign o[18347] = i[18347];
  assign o[18346] = i[18346];
  assign o[18345] = i[18345];
  assign o[18344] = i[18344];
  assign o[18343] = i[18343];
  assign o[18342] = i[18342];
  assign o[18341] = i[18341];
  assign o[18340] = i[18340];
  assign o[18339] = i[18339];
  assign o[18338] = i[18338];
  assign o[18337] = i[18337];
  assign o[18336] = i[18336];
  assign o[18335] = i[18335];
  assign o[18334] = i[18334];
  assign o[18333] = i[18333];
  assign o[18332] = i[18332];
  assign o[18331] = i[18331];
  assign o[18330] = i[18330];
  assign o[18329] = i[18329];
  assign o[18328] = i[18328];
  assign o[18327] = i[18327];
  assign o[18326] = i[18326];
  assign o[18325] = i[18325];
  assign o[18324] = i[18324];
  assign o[18323] = i[18323];
  assign o[18322] = i[18322];
  assign o[18321] = i[18321];
  assign o[18320] = i[18320];
  assign o[18319] = i[18319];
  assign o[18318] = i[18318];
  assign o[18317] = i[18317];
  assign o[18316] = i[18316];
  assign o[18315] = i[18315];
  assign o[18314] = i[18314];
  assign o[18313] = i[18313];
  assign o[18312] = i[18312];
  assign o[18311] = i[18311];
  assign o[18310] = i[18310];
  assign o[18309] = i[18309];
  assign o[18308] = i[18308];
  assign o[18307] = i[18307];
  assign o[18306] = i[18306];
  assign o[18305] = i[18305];
  assign o[18304] = i[18304];
  assign o[18303] = i[18303];
  assign o[18302] = i[18302];
  assign o[18301] = i[18301];
  assign o[18300] = i[18300];
  assign o[18299] = i[18299];
  assign o[18298] = i[18298];
  assign o[18297] = i[18297];
  assign o[18296] = i[18296];
  assign o[18295] = i[18295];
  assign o[18294] = i[18294];
  assign o[18293] = i[18293];
  assign o[18292] = i[18292];
  assign o[18291] = i[18291];
  assign o[18290] = i[18290];
  assign o[18289] = i[18289];
  assign o[18288] = i[18288];
  assign o[18287] = i[18287];
  assign o[18286] = i[18286];
  assign o[18285] = i[18285];
  assign o[18284] = i[18284];
  assign o[18283] = i[18283];
  assign o[18282] = i[18282];
  assign o[18281] = i[18281];
  assign o[18280] = i[18280];
  assign o[18279] = i[18279];
  assign o[18278] = i[18278];
  assign o[18277] = i[18277];
  assign o[18276] = i[18276];
  assign o[18275] = i[18275];
  assign o[18274] = i[18274];
  assign o[18273] = i[18273];
  assign o[18272] = i[18272];
  assign o[18271] = i[18271];
  assign o[18270] = i[18270];
  assign o[18269] = i[18269];
  assign o[18268] = i[18268];
  assign o[18267] = i[18267];
  assign o[18266] = i[18266];
  assign o[18265] = i[18265];
  assign o[18264] = i[18264];
  assign o[18263] = i[18263];
  assign o[18262] = i[18262];
  assign o[18261] = i[18261];
  assign o[18260] = i[18260];
  assign o[18259] = i[18259];
  assign o[18258] = i[18258];
  assign o[18257] = i[18257];
  assign o[18256] = i[18256];
  assign o[18255] = i[18255];
  assign o[18254] = i[18254];
  assign o[18253] = i[18253];
  assign o[18252] = i[18252];
  assign o[18251] = i[18251];
  assign o[18250] = i[18250];
  assign o[18249] = i[18249];
  assign o[18248] = i[18248];
  assign o[18247] = i[18247];
  assign o[18246] = i[18246];
  assign o[18245] = i[18245];
  assign o[18244] = i[18244];
  assign o[18243] = i[18243];
  assign o[18242] = i[18242];
  assign o[18241] = i[18241];
  assign o[18240] = i[18240];
  assign o[18239] = i[18239];
  assign o[18238] = i[18238];
  assign o[18237] = i[18237];
  assign o[18236] = i[18236];
  assign o[18235] = i[18235];
  assign o[18234] = i[18234];
  assign o[18233] = i[18233];
  assign o[18232] = i[18232];
  assign o[18231] = i[18231];
  assign o[18230] = i[18230];
  assign o[18229] = i[18229];
  assign o[18228] = i[18228];
  assign o[18227] = i[18227];
  assign o[18226] = i[18226];
  assign o[18225] = i[18225];
  assign o[18224] = i[18224];
  assign o[18223] = i[18223];
  assign o[18222] = i[18222];
  assign o[18221] = i[18221];
  assign o[18220] = i[18220];
  assign o[18219] = i[18219];
  assign o[18218] = i[18218];
  assign o[18217] = i[18217];
  assign o[18216] = i[18216];
  assign o[18215] = i[18215];
  assign o[18214] = i[18214];
  assign o[18213] = i[18213];
  assign o[18212] = i[18212];
  assign o[18211] = i[18211];
  assign o[18210] = i[18210];
  assign o[18209] = i[18209];
  assign o[18208] = i[18208];
  assign o[18207] = i[18207];
  assign o[18206] = i[18206];
  assign o[18205] = i[18205];
  assign o[18204] = i[18204];
  assign o[18203] = i[18203];
  assign o[18202] = i[18202];
  assign o[18201] = i[18201];
  assign o[18200] = i[18200];
  assign o[18199] = i[18199];
  assign o[18198] = i[18198];
  assign o[18197] = i[18197];
  assign o[18196] = i[18196];
  assign o[18195] = i[18195];
  assign o[18194] = i[18194];
  assign o[18193] = i[18193];
  assign o[18192] = i[18192];
  assign o[18191] = i[18191];
  assign o[18190] = i[18190];
  assign o[18189] = i[18189];
  assign o[18188] = i[18188];
  assign o[18187] = i[18187];
  assign o[18186] = i[18186];
  assign o[18185] = i[18185];
  assign o[18184] = i[18184];
  assign o[18183] = i[18183];
  assign o[18182] = i[18182];
  assign o[18181] = i[18181];
  assign o[18180] = i[18180];
  assign o[18179] = i[18179];
  assign o[18178] = i[18178];
  assign o[18177] = i[18177];
  assign o[18176] = i[18176];
  assign o[18175] = i[18175];
  assign o[18174] = i[18174];
  assign o[18173] = i[18173];
  assign o[18172] = i[18172];
  assign o[18171] = i[18171];
  assign o[18170] = i[18170];
  assign o[18169] = i[18169];
  assign o[18168] = i[18168];
  assign o[18167] = i[18167];
  assign o[18166] = i[18166];
  assign o[18165] = i[18165];
  assign o[18164] = i[18164];
  assign o[18163] = i[18163];
  assign o[18162] = i[18162];
  assign o[18161] = i[18161];
  assign o[18160] = i[18160];
  assign o[18159] = i[18159];
  assign o[18158] = i[18158];
  assign o[18157] = i[18157];
  assign o[18156] = i[18156];
  assign o[18155] = i[18155];
  assign o[18154] = i[18154];
  assign o[18153] = i[18153];
  assign o[18152] = i[18152];
  assign o[18151] = i[18151];
  assign o[18150] = i[18150];
  assign o[18149] = i[18149];
  assign o[18148] = i[18148];
  assign o[18147] = i[18147];
  assign o[18146] = i[18146];
  assign o[18145] = i[18145];
  assign o[18144] = i[18144];
  assign o[18143] = i[18143];
  assign o[18142] = i[18142];
  assign o[18141] = i[18141];
  assign o[18140] = i[18140];
  assign o[18139] = i[18139];
  assign o[18138] = i[18138];
  assign o[18137] = i[18137];
  assign o[18136] = i[18136];
  assign o[18135] = i[18135];
  assign o[18134] = i[18134];
  assign o[18133] = i[18133];
  assign o[18132] = i[18132];
  assign o[18131] = i[18131];
  assign o[18130] = i[18130];
  assign o[18129] = i[18129];
  assign o[18128] = i[18128];
  assign o[18127] = i[18127];
  assign o[18126] = i[18126];
  assign o[18125] = i[18125];
  assign o[18124] = i[18124];
  assign o[18123] = i[18123];
  assign o[18122] = i[18122];
  assign o[18121] = i[18121];
  assign o[18120] = i[18120];
  assign o[18119] = i[18119];
  assign o[18118] = i[18118];
  assign o[18117] = i[18117];
  assign o[18116] = i[18116];
  assign o[18115] = i[18115];
  assign o[18114] = i[18114];
  assign o[18113] = i[18113];
  assign o[18112] = i[18112];
  assign o[18111] = i[18111];
  assign o[18110] = i[18110];
  assign o[18109] = i[18109];
  assign o[18108] = i[18108];
  assign o[18107] = i[18107];
  assign o[18106] = i[18106];
  assign o[18105] = i[18105];
  assign o[18104] = i[18104];
  assign o[18103] = i[18103];
  assign o[18102] = i[18102];
  assign o[18101] = i[18101];
  assign o[18100] = i[18100];
  assign o[18099] = i[18099];
  assign o[18098] = i[18098];
  assign o[18097] = i[18097];
  assign o[18096] = i[18096];
  assign o[18095] = i[18095];
  assign o[18094] = i[18094];
  assign o[18093] = i[18093];
  assign o[18092] = i[18092];
  assign o[18091] = i[18091];
  assign o[18090] = i[18090];
  assign o[18089] = i[18089];
  assign o[18088] = i[18088];
  assign o[18087] = i[18087];
  assign o[18086] = i[18086];
  assign o[18085] = i[18085];
  assign o[18084] = i[18084];
  assign o[18083] = i[18083];
  assign o[18082] = i[18082];
  assign o[18081] = i[18081];
  assign o[18080] = i[18080];
  assign o[18079] = i[18079];
  assign o[18078] = i[18078];
  assign o[18077] = i[18077];
  assign o[18076] = i[18076];
  assign o[18075] = i[18075];
  assign o[18074] = i[18074];
  assign o[18073] = i[18073];
  assign o[18072] = i[18072];
  assign o[18071] = i[18071];
  assign o[18070] = i[18070];
  assign o[18069] = i[18069];
  assign o[18068] = i[18068];
  assign o[18067] = i[18067];
  assign o[18066] = i[18066];
  assign o[18065] = i[18065];
  assign o[18064] = i[18064];
  assign o[18063] = i[18063];
  assign o[18062] = i[18062];
  assign o[18061] = i[18061];
  assign o[18060] = i[18060];
  assign o[18059] = i[18059];
  assign o[18058] = i[18058];
  assign o[18057] = i[18057];
  assign o[18056] = i[18056];
  assign o[18055] = i[18055];
  assign o[18054] = i[18054];
  assign o[18053] = i[18053];
  assign o[18052] = i[18052];
  assign o[18051] = i[18051];
  assign o[18050] = i[18050];
  assign o[18049] = i[18049];
  assign o[18048] = i[18048];
  assign o[18047] = i[18047];
  assign o[18046] = i[18046];
  assign o[18045] = i[18045];
  assign o[18044] = i[18044];
  assign o[18043] = i[18043];
  assign o[18042] = i[18042];
  assign o[18041] = i[18041];
  assign o[18040] = i[18040];
  assign o[18039] = i[18039];
  assign o[18038] = i[18038];
  assign o[18037] = i[18037];
  assign o[18036] = i[18036];
  assign o[18035] = i[18035];
  assign o[18034] = i[18034];
  assign o[18033] = i[18033];
  assign o[18032] = i[18032];
  assign o[18031] = i[18031];
  assign o[18030] = i[18030];
  assign o[18029] = i[18029];
  assign o[18028] = i[18028];
  assign o[18027] = i[18027];
  assign o[18026] = i[18026];
  assign o[18025] = i[18025];
  assign o[18024] = i[18024];
  assign o[18023] = i[18023];
  assign o[18022] = i[18022];
  assign o[18021] = i[18021];
  assign o[18020] = i[18020];
  assign o[18019] = i[18019];
  assign o[18018] = i[18018];
  assign o[18017] = i[18017];
  assign o[18016] = i[18016];
  assign o[18015] = i[18015];
  assign o[18014] = i[18014];
  assign o[18013] = i[18013];
  assign o[18012] = i[18012];
  assign o[18011] = i[18011];
  assign o[18010] = i[18010];
  assign o[18009] = i[18009];
  assign o[18008] = i[18008];
  assign o[18007] = i[18007];
  assign o[18006] = i[18006];
  assign o[18005] = i[18005];
  assign o[18004] = i[18004];
  assign o[18003] = i[18003];
  assign o[18002] = i[18002];
  assign o[18001] = i[18001];
  assign o[18000] = i[18000];
  assign o[17999] = i[17999];
  assign o[17998] = i[17998];
  assign o[17997] = i[17997];
  assign o[17996] = i[17996];
  assign o[17995] = i[17995];
  assign o[17994] = i[17994];
  assign o[17993] = i[17993];
  assign o[17992] = i[17992];
  assign o[17991] = i[17991];
  assign o[17990] = i[17990];
  assign o[17989] = i[17989];
  assign o[17988] = i[17988];
  assign o[17987] = i[17987];
  assign o[17986] = i[17986];
  assign o[17985] = i[17985];
  assign o[17984] = i[17984];
  assign o[17983] = i[17983];
  assign o[17982] = i[17982];
  assign o[17981] = i[17981];
  assign o[17980] = i[17980];
  assign o[17979] = i[17979];
  assign o[17978] = i[17978];
  assign o[17977] = i[17977];
  assign o[17976] = i[17976];
  assign o[17975] = i[17975];
  assign o[17974] = i[17974];
  assign o[17973] = i[17973];
  assign o[17972] = i[17972];
  assign o[17971] = i[17971];
  assign o[17970] = i[17970];
  assign o[17969] = i[17969];
  assign o[17968] = i[17968];
  assign o[17967] = i[17967];
  assign o[17966] = i[17966];
  assign o[17965] = i[17965];
  assign o[17964] = i[17964];
  assign o[17963] = i[17963];
  assign o[17962] = i[17962];
  assign o[17961] = i[17961];
  assign o[17960] = i[17960];
  assign o[17959] = i[17959];
  assign o[17958] = i[17958];
  assign o[17957] = i[17957];
  assign o[17956] = i[17956];
  assign o[17955] = i[17955];
  assign o[17954] = i[17954];
  assign o[17953] = i[17953];
  assign o[17952] = i[17952];
  assign o[17951] = i[17951];
  assign o[17950] = i[17950];
  assign o[17949] = i[17949];
  assign o[17948] = i[17948];
  assign o[17947] = i[17947];
  assign o[17946] = i[17946];
  assign o[17945] = i[17945];
  assign o[17944] = i[17944];
  assign o[17943] = i[17943];
  assign o[17942] = i[17942];
  assign o[17941] = i[17941];
  assign o[17940] = i[17940];
  assign o[17939] = i[17939];
  assign o[17938] = i[17938];
  assign o[17937] = i[17937];
  assign o[17936] = i[17936];
  assign o[17935] = i[17935];
  assign o[17934] = i[17934];
  assign o[17933] = i[17933];
  assign o[17932] = i[17932];
  assign o[17931] = i[17931];
  assign o[17930] = i[17930];
  assign o[17929] = i[17929];
  assign o[17928] = i[17928];
  assign o[17927] = i[17927];
  assign o[17926] = i[17926];
  assign o[17925] = i[17925];
  assign o[17924] = i[17924];
  assign o[17923] = i[17923];
  assign o[17922] = i[17922];
  assign o[17921] = i[17921];
  assign o[17920] = i[17920];
  assign o[17919] = i[17919];
  assign o[17918] = i[17918];
  assign o[17917] = i[17917];
  assign o[17916] = i[17916];
  assign o[17915] = i[17915];
  assign o[17914] = i[17914];
  assign o[17913] = i[17913];
  assign o[17912] = i[17912];
  assign o[17911] = i[17911];
  assign o[17910] = i[17910];
  assign o[17909] = i[17909];
  assign o[17908] = i[17908];
  assign o[17907] = i[17907];
  assign o[17906] = i[17906];
  assign o[17905] = i[17905];
  assign o[17904] = i[17904];
  assign o[17903] = i[17903];
  assign o[17902] = i[17902];
  assign o[17901] = i[17901];
  assign o[17900] = i[17900];
  assign o[17899] = i[17899];
  assign o[17898] = i[17898];
  assign o[17897] = i[17897];
  assign o[17896] = i[17896];
  assign o[17895] = i[17895];
  assign o[17894] = i[17894];
  assign o[17893] = i[17893];
  assign o[17892] = i[17892];
  assign o[17891] = i[17891];
  assign o[17890] = i[17890];
  assign o[17889] = i[17889];
  assign o[17888] = i[17888];
  assign o[17887] = i[17887];
  assign o[17886] = i[17886];
  assign o[17885] = i[17885];
  assign o[17884] = i[17884];
  assign o[17883] = i[17883];
  assign o[17882] = i[17882];
  assign o[17881] = i[17881];
  assign o[17880] = i[17880];
  assign o[17879] = i[17879];
  assign o[17878] = i[17878];
  assign o[17877] = i[17877];
  assign o[17876] = i[17876];
  assign o[17875] = i[17875];
  assign o[17874] = i[17874];
  assign o[17873] = i[17873];
  assign o[17872] = i[17872];
  assign o[17871] = i[17871];
  assign o[17870] = i[17870];
  assign o[17869] = i[17869];
  assign o[17868] = i[17868];
  assign o[17867] = i[17867];
  assign o[17866] = i[17866];
  assign o[17865] = i[17865];
  assign o[17864] = i[17864];
  assign o[17863] = i[17863];
  assign o[17862] = i[17862];
  assign o[17861] = i[17861];
  assign o[17860] = i[17860];
  assign o[17859] = i[17859];
  assign o[17858] = i[17858];
  assign o[17857] = i[17857];
  assign o[17856] = i[17856];
  assign o[17855] = i[17855];
  assign o[17854] = i[17854];
  assign o[17853] = i[17853];
  assign o[17852] = i[17852];
  assign o[17851] = i[17851];
  assign o[17850] = i[17850];
  assign o[17849] = i[17849];
  assign o[17848] = i[17848];
  assign o[17847] = i[17847];
  assign o[17846] = i[17846];
  assign o[17845] = i[17845];
  assign o[17844] = i[17844];
  assign o[17843] = i[17843];
  assign o[17842] = i[17842];
  assign o[17841] = i[17841];
  assign o[17840] = i[17840];
  assign o[17839] = i[17839];
  assign o[17838] = i[17838];
  assign o[17837] = i[17837];
  assign o[17836] = i[17836];
  assign o[17835] = i[17835];
  assign o[17834] = i[17834];
  assign o[17833] = i[17833];
  assign o[17832] = i[17832];
  assign o[17831] = i[17831];
  assign o[17830] = i[17830];
  assign o[17829] = i[17829];
  assign o[17828] = i[17828];
  assign o[17827] = i[17827];
  assign o[17826] = i[17826];
  assign o[17825] = i[17825];
  assign o[17824] = i[17824];
  assign o[17823] = i[17823];
  assign o[17822] = i[17822];
  assign o[17821] = i[17821];
  assign o[17820] = i[17820];
  assign o[17819] = i[17819];
  assign o[17818] = i[17818];
  assign o[17817] = i[17817];
  assign o[17816] = i[17816];
  assign o[17815] = i[17815];
  assign o[17814] = i[17814];
  assign o[17813] = i[17813];
  assign o[17812] = i[17812];
  assign o[17811] = i[17811];
  assign o[17810] = i[17810];
  assign o[17809] = i[17809];
  assign o[17808] = i[17808];
  assign o[17807] = i[17807];
  assign o[17806] = i[17806];
  assign o[17805] = i[17805];
  assign o[17804] = i[17804];
  assign o[17803] = i[17803];
  assign o[17802] = i[17802];
  assign o[17801] = i[17801];
  assign o[17800] = i[17800];
  assign o[17799] = i[17799];
  assign o[17798] = i[17798];
  assign o[17797] = i[17797];
  assign o[17796] = i[17796];
  assign o[17795] = i[17795];
  assign o[17794] = i[17794];
  assign o[17793] = i[17793];
  assign o[17792] = i[17792];
  assign o[17791] = i[17791];
  assign o[17790] = i[17790];
  assign o[17789] = i[17789];
  assign o[17788] = i[17788];
  assign o[17787] = i[17787];
  assign o[17786] = i[17786];
  assign o[17785] = i[17785];
  assign o[17784] = i[17784];
  assign o[17783] = i[17783];
  assign o[17782] = i[17782];
  assign o[17781] = i[17781];
  assign o[17780] = i[17780];
  assign o[17779] = i[17779];
  assign o[17778] = i[17778];
  assign o[17777] = i[17777];
  assign o[17776] = i[17776];
  assign o[17775] = i[17775];
  assign o[17774] = i[17774];
  assign o[17773] = i[17773];
  assign o[17772] = i[17772];
  assign o[17771] = i[17771];
  assign o[17770] = i[17770];
  assign o[17769] = i[17769];
  assign o[17768] = i[17768];
  assign o[17767] = i[17767];
  assign o[17766] = i[17766];
  assign o[17765] = i[17765];
  assign o[17764] = i[17764];
  assign o[17763] = i[17763];
  assign o[17762] = i[17762];
  assign o[17761] = i[17761];
  assign o[17760] = i[17760];
  assign o[17759] = i[17759];
  assign o[17758] = i[17758];
  assign o[17757] = i[17757];
  assign o[17756] = i[17756];
  assign o[17755] = i[17755];
  assign o[17754] = i[17754];
  assign o[17753] = i[17753];
  assign o[17752] = i[17752];
  assign o[17751] = i[17751];
  assign o[17750] = i[17750];
  assign o[17749] = i[17749];
  assign o[17748] = i[17748];
  assign o[17747] = i[17747];
  assign o[17746] = i[17746];
  assign o[17745] = i[17745];
  assign o[17744] = i[17744];
  assign o[17743] = i[17743];
  assign o[17742] = i[17742];
  assign o[17741] = i[17741];
  assign o[17740] = i[17740];
  assign o[17739] = i[17739];
  assign o[17738] = i[17738];
  assign o[17737] = i[17737];
  assign o[17736] = i[17736];
  assign o[17735] = i[17735];
  assign o[17734] = i[17734];
  assign o[17733] = i[17733];
  assign o[17732] = i[17732];
  assign o[17731] = i[17731];
  assign o[17730] = i[17730];
  assign o[17729] = i[17729];
  assign o[17728] = i[17728];
  assign o[17727] = i[17727];
  assign o[17726] = i[17726];
  assign o[17725] = i[17725];
  assign o[17724] = i[17724];
  assign o[17723] = i[17723];
  assign o[17722] = i[17722];
  assign o[17721] = i[17721];
  assign o[17720] = i[17720];
  assign o[17719] = i[17719];
  assign o[17718] = i[17718];
  assign o[17717] = i[17717];
  assign o[17716] = i[17716];
  assign o[17715] = i[17715];
  assign o[17714] = i[17714];
  assign o[17713] = i[17713];
  assign o[17712] = i[17712];
  assign o[17711] = i[17711];
  assign o[17710] = i[17710];
  assign o[17709] = i[17709];
  assign o[17708] = i[17708];
  assign o[17707] = i[17707];
  assign o[17706] = i[17706];
  assign o[17705] = i[17705];
  assign o[17704] = i[17704];
  assign o[17703] = i[17703];
  assign o[17702] = i[17702];
  assign o[17701] = i[17701];
  assign o[17700] = i[17700];
  assign o[17699] = i[17699];
  assign o[17698] = i[17698];
  assign o[17697] = i[17697];
  assign o[17696] = i[17696];
  assign o[17695] = i[17695];
  assign o[17694] = i[17694];
  assign o[17693] = i[17693];
  assign o[17692] = i[17692];
  assign o[17691] = i[17691];
  assign o[17690] = i[17690];
  assign o[17689] = i[17689];
  assign o[17688] = i[17688];
  assign o[17687] = i[17687];
  assign o[17686] = i[17686];
  assign o[17685] = i[17685];
  assign o[17684] = i[17684];
  assign o[17683] = i[17683];
  assign o[17682] = i[17682];
  assign o[17681] = i[17681];
  assign o[17680] = i[17680];
  assign o[17679] = i[17679];
  assign o[17678] = i[17678];
  assign o[17677] = i[17677];
  assign o[17676] = i[17676];
  assign o[17675] = i[17675];
  assign o[17674] = i[17674];
  assign o[17673] = i[17673];
  assign o[17672] = i[17672];
  assign o[17671] = i[17671];
  assign o[17670] = i[17670];
  assign o[17669] = i[17669];
  assign o[17668] = i[17668];
  assign o[17667] = i[17667];
  assign o[17666] = i[17666];
  assign o[17665] = i[17665];
  assign o[17664] = i[17664];
  assign o[17663] = i[17663];
  assign o[17662] = i[17662];
  assign o[17661] = i[17661];
  assign o[17660] = i[17660];
  assign o[17659] = i[17659];
  assign o[17658] = i[17658];
  assign o[17657] = i[17657];
  assign o[17656] = i[17656];
  assign o[17655] = i[17655];
  assign o[17654] = i[17654];
  assign o[17653] = i[17653];
  assign o[17652] = i[17652];
  assign o[17651] = i[17651];
  assign o[17650] = i[17650];
  assign o[17649] = i[17649];
  assign o[17648] = i[17648];
  assign o[17647] = i[17647];
  assign o[17646] = i[17646];
  assign o[17645] = i[17645];
  assign o[17644] = i[17644];
  assign o[17643] = i[17643];
  assign o[17642] = i[17642];
  assign o[17641] = i[17641];
  assign o[17640] = i[17640];
  assign o[17639] = i[17639];
  assign o[17638] = i[17638];
  assign o[17637] = i[17637];
  assign o[17636] = i[17636];
  assign o[17635] = i[17635];
  assign o[17634] = i[17634];
  assign o[17633] = i[17633];
  assign o[17632] = i[17632];
  assign o[17631] = i[17631];
  assign o[17630] = i[17630];
  assign o[17629] = i[17629];
  assign o[17628] = i[17628];
  assign o[17627] = i[17627];
  assign o[17626] = i[17626];
  assign o[17625] = i[17625];
  assign o[17624] = i[17624];
  assign o[17623] = i[17623];
  assign o[17622] = i[17622];
  assign o[17621] = i[17621];
  assign o[17620] = i[17620];
  assign o[17619] = i[17619];
  assign o[17618] = i[17618];
  assign o[17617] = i[17617];
  assign o[17616] = i[17616];
  assign o[17615] = i[17615];
  assign o[17614] = i[17614];
  assign o[17613] = i[17613];
  assign o[17612] = i[17612];
  assign o[17611] = i[17611];
  assign o[17610] = i[17610];
  assign o[17609] = i[17609];
  assign o[17608] = i[17608];
  assign o[17607] = i[17607];
  assign o[17606] = i[17606];
  assign o[17605] = i[17605];
  assign o[17604] = i[17604];
  assign o[17603] = i[17603];
  assign o[17602] = i[17602];
  assign o[17601] = i[17601];
  assign o[17600] = i[17600];
  assign o[17599] = i[17599];
  assign o[17598] = i[17598];
  assign o[17597] = i[17597];
  assign o[17596] = i[17596];
  assign o[17595] = i[17595];
  assign o[17594] = i[17594];
  assign o[17593] = i[17593];
  assign o[17592] = i[17592];
  assign o[17591] = i[17591];
  assign o[17590] = i[17590];
  assign o[17589] = i[17589];
  assign o[17588] = i[17588];
  assign o[17587] = i[17587];
  assign o[17586] = i[17586];
  assign o[17585] = i[17585];
  assign o[17584] = i[17584];
  assign o[17583] = i[17583];
  assign o[17582] = i[17582];
  assign o[17581] = i[17581];
  assign o[17580] = i[17580];
  assign o[17579] = i[17579];
  assign o[17578] = i[17578];
  assign o[17577] = i[17577];
  assign o[17576] = i[17576];
  assign o[17575] = i[17575];
  assign o[17574] = i[17574];
  assign o[17573] = i[17573];
  assign o[17572] = i[17572];
  assign o[17571] = i[17571];
  assign o[17570] = i[17570];
  assign o[17569] = i[17569];
  assign o[17568] = i[17568];
  assign o[17567] = i[17567];
  assign o[17566] = i[17566];
  assign o[17565] = i[17565];
  assign o[17564] = i[17564];
  assign o[17563] = i[17563];
  assign o[17562] = i[17562];
  assign o[17561] = i[17561];
  assign o[17560] = i[17560];
  assign o[17559] = i[17559];
  assign o[17558] = i[17558];
  assign o[17557] = i[17557];
  assign o[17556] = i[17556];
  assign o[17555] = i[17555];
  assign o[17554] = i[17554];
  assign o[17553] = i[17553];
  assign o[17552] = i[17552];
  assign o[17551] = i[17551];
  assign o[17550] = i[17550];
  assign o[17549] = i[17549];
  assign o[17548] = i[17548];
  assign o[17547] = i[17547];
  assign o[17546] = i[17546];
  assign o[17545] = i[17545];
  assign o[17544] = i[17544];
  assign o[17543] = i[17543];
  assign o[17542] = i[17542];
  assign o[17541] = i[17541];
  assign o[17540] = i[17540];
  assign o[17539] = i[17539];
  assign o[17538] = i[17538];
  assign o[17537] = i[17537];
  assign o[17536] = i[17536];
  assign o[17535] = i[17535];
  assign o[17534] = i[17534];
  assign o[17533] = i[17533];
  assign o[17532] = i[17532];
  assign o[17531] = i[17531];
  assign o[17530] = i[17530];
  assign o[17529] = i[17529];
  assign o[17528] = i[17528];
  assign o[17527] = i[17527];
  assign o[17526] = i[17526];
  assign o[17525] = i[17525];
  assign o[17524] = i[17524];
  assign o[17523] = i[17523];
  assign o[17522] = i[17522];
  assign o[17521] = i[17521];
  assign o[17520] = i[17520];
  assign o[17519] = i[17519];
  assign o[17518] = i[17518];
  assign o[17517] = i[17517];
  assign o[17516] = i[17516];
  assign o[17515] = i[17515];
  assign o[17514] = i[17514];
  assign o[17513] = i[17513];
  assign o[17512] = i[17512];
  assign o[17511] = i[17511];
  assign o[17510] = i[17510];
  assign o[17509] = i[17509];
  assign o[17508] = i[17508];
  assign o[17507] = i[17507];
  assign o[17506] = i[17506];
  assign o[17505] = i[17505];
  assign o[17504] = i[17504];
  assign o[17503] = i[17503];
  assign o[17502] = i[17502];
  assign o[17501] = i[17501];
  assign o[17500] = i[17500];
  assign o[17499] = i[17499];
  assign o[17498] = i[17498];
  assign o[17497] = i[17497];
  assign o[17496] = i[17496];
  assign o[17495] = i[17495];
  assign o[17494] = i[17494];
  assign o[17493] = i[17493];
  assign o[17492] = i[17492];
  assign o[17491] = i[17491];
  assign o[17490] = i[17490];
  assign o[17489] = i[17489];
  assign o[17488] = i[17488];
  assign o[17487] = i[17487];
  assign o[17486] = i[17486];
  assign o[17485] = i[17485];
  assign o[17484] = i[17484];
  assign o[17483] = i[17483];
  assign o[17482] = i[17482];
  assign o[17481] = i[17481];
  assign o[17480] = i[17480];
  assign o[17479] = i[17479];
  assign o[17478] = i[17478];
  assign o[17477] = i[17477];
  assign o[17476] = i[17476];
  assign o[17475] = i[17475];
  assign o[17474] = i[17474];
  assign o[17473] = i[17473];
  assign o[17472] = i[17472];
  assign o[17471] = i[17471];
  assign o[17470] = i[17470];
  assign o[17469] = i[17469];
  assign o[17468] = i[17468];
  assign o[17467] = i[17467];
  assign o[17466] = i[17466];
  assign o[17465] = i[17465];
  assign o[17464] = i[17464];
  assign o[17463] = i[17463];
  assign o[17462] = i[17462];
  assign o[17461] = i[17461];
  assign o[17460] = i[17460];
  assign o[17459] = i[17459];
  assign o[17458] = i[17458];
  assign o[17457] = i[17457];
  assign o[17456] = i[17456];
  assign o[17455] = i[17455];
  assign o[17454] = i[17454];
  assign o[17453] = i[17453];
  assign o[17452] = i[17452];
  assign o[17451] = i[17451];
  assign o[17450] = i[17450];
  assign o[17449] = i[17449];
  assign o[17448] = i[17448];
  assign o[17447] = i[17447];
  assign o[17446] = i[17446];
  assign o[17445] = i[17445];
  assign o[17444] = i[17444];
  assign o[17443] = i[17443];
  assign o[17442] = i[17442];
  assign o[17441] = i[17441];
  assign o[17440] = i[17440];
  assign o[17439] = i[17439];
  assign o[17438] = i[17438];
  assign o[17437] = i[17437];
  assign o[17436] = i[17436];
  assign o[17435] = i[17435];
  assign o[17434] = i[17434];
  assign o[17433] = i[17433];
  assign o[17432] = i[17432];
  assign o[17431] = i[17431];
  assign o[17430] = i[17430];
  assign o[17429] = i[17429];
  assign o[17428] = i[17428];
  assign o[17427] = i[17427];
  assign o[17426] = i[17426];
  assign o[17425] = i[17425];
  assign o[17424] = i[17424];
  assign o[17423] = i[17423];
  assign o[17422] = i[17422];
  assign o[17421] = i[17421];
  assign o[17420] = i[17420];
  assign o[17419] = i[17419];
  assign o[17418] = i[17418];
  assign o[17417] = i[17417];
  assign o[17416] = i[17416];
  assign o[17415] = i[17415];
  assign o[17414] = i[17414];
  assign o[17413] = i[17413];
  assign o[17412] = i[17412];
  assign o[17411] = i[17411];
  assign o[17410] = i[17410];
  assign o[17409] = i[17409];
  assign o[17408] = i[17408];
  assign o[17407] = i[17407];
  assign o[17406] = i[17406];
  assign o[17405] = i[17405];
  assign o[17404] = i[17404];
  assign o[17403] = i[17403];
  assign o[17402] = i[17402];
  assign o[17401] = i[17401];
  assign o[17400] = i[17400];
  assign o[17399] = i[17399];
  assign o[17398] = i[17398];
  assign o[17397] = i[17397];
  assign o[17396] = i[17396];
  assign o[17395] = i[17395];
  assign o[17394] = i[17394];
  assign o[17393] = i[17393];
  assign o[17392] = i[17392];
  assign o[17391] = i[17391];
  assign o[17390] = i[17390];
  assign o[17389] = i[17389];
  assign o[17388] = i[17388];
  assign o[17387] = i[17387];
  assign o[17386] = i[17386];
  assign o[17385] = i[17385];
  assign o[17384] = i[17384];
  assign o[17383] = i[17383];
  assign o[17382] = i[17382];
  assign o[17381] = i[17381];
  assign o[17380] = i[17380];
  assign o[17379] = i[17379];
  assign o[17378] = i[17378];
  assign o[17377] = i[17377];
  assign o[17376] = i[17376];
  assign o[17375] = i[17375];
  assign o[17374] = i[17374];
  assign o[17373] = i[17373];
  assign o[17372] = i[17372];
  assign o[17371] = i[17371];
  assign o[17370] = i[17370];
  assign o[17369] = i[17369];
  assign o[17368] = i[17368];
  assign o[17367] = i[17367];
  assign o[17366] = i[17366];
  assign o[17365] = i[17365];
  assign o[17364] = i[17364];
  assign o[17363] = i[17363];
  assign o[17362] = i[17362];
  assign o[17361] = i[17361];
  assign o[17360] = i[17360];
  assign o[17359] = i[17359];
  assign o[17358] = i[17358];
  assign o[17357] = i[17357];
  assign o[17356] = i[17356];
  assign o[17355] = i[17355];
  assign o[17354] = i[17354];
  assign o[17353] = i[17353];
  assign o[17352] = i[17352];
  assign o[17351] = i[17351];
  assign o[17350] = i[17350];
  assign o[17349] = i[17349];
  assign o[17348] = i[17348];
  assign o[17347] = i[17347];
  assign o[17346] = i[17346];
  assign o[17345] = i[17345];
  assign o[17344] = i[17344];
  assign o[17343] = i[17343];
  assign o[17342] = i[17342];
  assign o[17341] = i[17341];
  assign o[17340] = i[17340];
  assign o[17339] = i[17339];
  assign o[17338] = i[17338];
  assign o[17337] = i[17337];
  assign o[17336] = i[17336];
  assign o[17335] = i[17335];
  assign o[17334] = i[17334];
  assign o[17333] = i[17333];
  assign o[17332] = i[17332];
  assign o[17331] = i[17331];
  assign o[17330] = i[17330];
  assign o[17329] = i[17329];
  assign o[17328] = i[17328];
  assign o[17327] = i[17327];
  assign o[17326] = i[17326];
  assign o[17325] = i[17325];
  assign o[17324] = i[17324];
  assign o[17323] = i[17323];
  assign o[17322] = i[17322];
  assign o[17321] = i[17321];
  assign o[17320] = i[17320];
  assign o[17319] = i[17319];
  assign o[17318] = i[17318];
  assign o[17317] = i[17317];
  assign o[17316] = i[17316];
  assign o[17315] = i[17315];
  assign o[17314] = i[17314];
  assign o[17313] = i[17313];
  assign o[17312] = i[17312];
  assign o[17311] = i[17311];
  assign o[17310] = i[17310];
  assign o[17309] = i[17309];
  assign o[17308] = i[17308];
  assign o[17307] = i[17307];
  assign o[17306] = i[17306];
  assign o[17305] = i[17305];
  assign o[17304] = i[17304];
  assign o[17303] = i[17303];
  assign o[17302] = i[17302];
  assign o[17301] = i[17301];
  assign o[17300] = i[17300];
  assign o[17299] = i[17299];
  assign o[17298] = i[17298];
  assign o[17297] = i[17297];
  assign o[17296] = i[17296];
  assign o[17295] = i[17295];
  assign o[17294] = i[17294];
  assign o[17293] = i[17293];
  assign o[17292] = i[17292];
  assign o[17291] = i[17291];
  assign o[17290] = i[17290];
  assign o[17289] = i[17289];
  assign o[17288] = i[17288];
  assign o[17287] = i[17287];
  assign o[17286] = i[17286];
  assign o[17285] = i[17285];
  assign o[17284] = i[17284];
  assign o[17283] = i[17283];
  assign o[17282] = i[17282];
  assign o[17281] = i[17281];
  assign o[17280] = i[17280];
  assign o[17279] = i[17279];
  assign o[17278] = i[17278];
  assign o[17277] = i[17277];
  assign o[17276] = i[17276];
  assign o[17275] = i[17275];
  assign o[17274] = i[17274];
  assign o[17273] = i[17273];
  assign o[17272] = i[17272];
  assign o[17271] = i[17271];
  assign o[17270] = i[17270];
  assign o[17269] = i[17269];
  assign o[17268] = i[17268];
  assign o[17267] = i[17267];
  assign o[17266] = i[17266];
  assign o[17265] = i[17265];
  assign o[17264] = i[17264];
  assign o[17263] = i[17263];
  assign o[17262] = i[17262];
  assign o[17261] = i[17261];
  assign o[17260] = i[17260];
  assign o[17259] = i[17259];
  assign o[17258] = i[17258];
  assign o[17257] = i[17257];
  assign o[17256] = i[17256];
  assign o[17255] = i[17255];
  assign o[17254] = i[17254];
  assign o[17253] = i[17253];
  assign o[17252] = i[17252];
  assign o[17251] = i[17251];
  assign o[17250] = i[17250];
  assign o[17249] = i[17249];
  assign o[17248] = i[17248];
  assign o[17247] = i[17247];
  assign o[17246] = i[17246];
  assign o[17245] = i[17245];
  assign o[17244] = i[17244];
  assign o[17243] = i[17243];
  assign o[17242] = i[17242];
  assign o[17241] = i[17241];
  assign o[17240] = i[17240];
  assign o[17239] = i[17239];
  assign o[17238] = i[17238];
  assign o[17237] = i[17237];
  assign o[17236] = i[17236];
  assign o[17235] = i[17235];
  assign o[17234] = i[17234];
  assign o[17233] = i[17233];
  assign o[17232] = i[17232];
  assign o[17231] = i[17231];
  assign o[17230] = i[17230];
  assign o[17229] = i[17229];
  assign o[17228] = i[17228];
  assign o[17227] = i[17227];
  assign o[17226] = i[17226];
  assign o[17225] = i[17225];
  assign o[17224] = i[17224];
  assign o[17223] = i[17223];
  assign o[17222] = i[17222];
  assign o[17221] = i[17221];
  assign o[17220] = i[17220];
  assign o[17219] = i[17219];
  assign o[17218] = i[17218];
  assign o[17217] = i[17217];
  assign o[17216] = i[17216];
  assign o[17215] = i[17215];
  assign o[17214] = i[17214];
  assign o[17213] = i[17213];
  assign o[17212] = i[17212];
  assign o[17211] = i[17211];
  assign o[17210] = i[17210];
  assign o[17209] = i[17209];
  assign o[17208] = i[17208];
  assign o[17207] = i[17207];
  assign o[17206] = i[17206];
  assign o[17205] = i[17205];
  assign o[17204] = i[17204];
  assign o[17203] = i[17203];
  assign o[17202] = i[17202];
  assign o[17201] = i[17201];
  assign o[17200] = i[17200];
  assign o[17199] = i[17199];
  assign o[17198] = i[17198];
  assign o[17197] = i[17197];
  assign o[17196] = i[17196];
  assign o[17195] = i[17195];
  assign o[17194] = i[17194];
  assign o[17193] = i[17193];
  assign o[17192] = i[17192];
  assign o[17191] = i[17191];
  assign o[17190] = i[17190];
  assign o[17189] = i[17189];
  assign o[17188] = i[17188];
  assign o[17187] = i[17187];
  assign o[17186] = i[17186];
  assign o[17185] = i[17185];
  assign o[17184] = i[17184];
  assign o[17183] = i[17183];
  assign o[17182] = i[17182];
  assign o[17181] = i[17181];
  assign o[17180] = i[17180];
  assign o[17179] = i[17179];
  assign o[17178] = i[17178];
  assign o[17177] = i[17177];
  assign o[17176] = i[17176];
  assign o[17175] = i[17175];
  assign o[17174] = i[17174];
  assign o[17173] = i[17173];
  assign o[17172] = i[17172];
  assign o[17171] = i[17171];
  assign o[17170] = i[17170];
  assign o[17169] = i[17169];
  assign o[17168] = i[17168];
  assign o[17167] = i[17167];
  assign o[17166] = i[17166];
  assign o[17165] = i[17165];
  assign o[17164] = i[17164];
  assign o[17163] = i[17163];
  assign o[17162] = i[17162];
  assign o[17161] = i[17161];
  assign o[17160] = i[17160];
  assign o[17159] = i[17159];
  assign o[17158] = i[17158];
  assign o[17157] = i[17157];
  assign o[17156] = i[17156];
  assign o[17155] = i[17155];
  assign o[17154] = i[17154];
  assign o[17153] = i[17153];
  assign o[17152] = i[17152];
  assign o[17151] = i[17151];
  assign o[17150] = i[17150];
  assign o[17149] = i[17149];
  assign o[17148] = i[17148];
  assign o[17147] = i[17147];
  assign o[17146] = i[17146];
  assign o[17145] = i[17145];
  assign o[17144] = i[17144];
  assign o[17143] = i[17143];
  assign o[17142] = i[17142];
  assign o[17141] = i[17141];
  assign o[17140] = i[17140];
  assign o[17139] = i[17139];
  assign o[17138] = i[17138];
  assign o[17137] = i[17137];
  assign o[17136] = i[17136];
  assign o[17135] = i[17135];
  assign o[17134] = i[17134];
  assign o[17133] = i[17133];
  assign o[17132] = i[17132];
  assign o[17131] = i[17131];
  assign o[17130] = i[17130];
  assign o[17129] = i[17129];
  assign o[17128] = i[17128];
  assign o[17127] = i[17127];
  assign o[17126] = i[17126];
  assign o[17125] = i[17125];
  assign o[17124] = i[17124];
  assign o[17123] = i[17123];
  assign o[17122] = i[17122];
  assign o[17121] = i[17121];
  assign o[17120] = i[17120];
  assign o[17119] = i[17119];
  assign o[17118] = i[17118];
  assign o[17117] = i[17117];
  assign o[17116] = i[17116];
  assign o[17115] = i[17115];
  assign o[17114] = i[17114];
  assign o[17113] = i[17113];
  assign o[17112] = i[17112];
  assign o[17111] = i[17111];
  assign o[17110] = i[17110];
  assign o[17109] = i[17109];
  assign o[17108] = i[17108];
  assign o[17107] = i[17107];
  assign o[17106] = i[17106];
  assign o[17105] = i[17105];
  assign o[17104] = i[17104];
  assign o[17103] = i[17103];
  assign o[17102] = i[17102];
  assign o[17101] = i[17101];
  assign o[17100] = i[17100];
  assign o[17099] = i[17099];
  assign o[17098] = i[17098];
  assign o[17097] = i[17097];
  assign o[17096] = i[17096];
  assign o[17095] = i[17095];
  assign o[17094] = i[17094];
  assign o[17093] = i[17093];
  assign o[17092] = i[17092];
  assign o[17091] = i[17091];
  assign o[17090] = i[17090];
  assign o[17089] = i[17089];
  assign o[17088] = i[17088];
  assign o[17087] = i[17087];
  assign o[17086] = i[17086];
  assign o[17085] = i[17085];
  assign o[17084] = i[17084];
  assign o[17083] = i[17083];
  assign o[17082] = i[17082];
  assign o[17081] = i[17081];
  assign o[17080] = i[17080];
  assign o[17079] = i[17079];
  assign o[17078] = i[17078];
  assign o[17077] = i[17077];
  assign o[17076] = i[17076];
  assign o[17075] = i[17075];
  assign o[17074] = i[17074];
  assign o[17073] = i[17073];
  assign o[17072] = i[17072];
  assign o[17071] = i[17071];
  assign o[17070] = i[17070];
  assign o[17069] = i[17069];
  assign o[17068] = i[17068];
  assign o[17067] = i[17067];
  assign o[17066] = i[17066];
  assign o[17065] = i[17065];
  assign o[17064] = i[17064];
  assign o[17063] = i[17063];
  assign o[17062] = i[17062];
  assign o[17061] = i[17061];
  assign o[17060] = i[17060];
  assign o[17059] = i[17059];
  assign o[17058] = i[17058];
  assign o[17057] = i[17057];
  assign o[17056] = i[17056];
  assign o[17055] = i[17055];
  assign o[17054] = i[17054];
  assign o[17053] = i[17053];
  assign o[17052] = i[17052];
  assign o[17051] = i[17051];
  assign o[17050] = i[17050];
  assign o[17049] = i[17049];
  assign o[17048] = i[17048];
  assign o[17047] = i[17047];
  assign o[17046] = i[17046];
  assign o[17045] = i[17045];
  assign o[17044] = i[17044];
  assign o[17043] = i[17043];
  assign o[17042] = i[17042];
  assign o[17041] = i[17041];
  assign o[17040] = i[17040];
  assign o[17039] = i[17039];
  assign o[17038] = i[17038];
  assign o[17037] = i[17037];
  assign o[17036] = i[17036];
  assign o[17035] = i[17035];
  assign o[17034] = i[17034];
  assign o[17033] = i[17033];
  assign o[17032] = i[17032];
  assign o[17031] = i[17031];
  assign o[17030] = i[17030];
  assign o[17029] = i[17029];
  assign o[17028] = i[17028];
  assign o[17027] = i[17027];
  assign o[17026] = i[17026];
  assign o[17025] = i[17025];
  assign o[17024] = i[17024];
  assign o[17023] = i[17023];
  assign o[17022] = i[17022];
  assign o[17021] = i[17021];
  assign o[17020] = i[17020];
  assign o[17019] = i[17019];
  assign o[17018] = i[17018];
  assign o[17017] = i[17017];
  assign o[17016] = i[17016];
  assign o[17015] = i[17015];
  assign o[17014] = i[17014];
  assign o[17013] = i[17013];
  assign o[17012] = i[17012];
  assign o[17011] = i[17011];
  assign o[17010] = i[17010];
  assign o[17009] = i[17009];
  assign o[17008] = i[17008];
  assign o[17007] = i[17007];
  assign o[17006] = i[17006];
  assign o[17005] = i[17005];
  assign o[17004] = i[17004];
  assign o[17003] = i[17003];
  assign o[17002] = i[17002];
  assign o[17001] = i[17001];
  assign o[17000] = i[17000];
  assign o[16999] = i[16999];
  assign o[16998] = i[16998];
  assign o[16997] = i[16997];
  assign o[16996] = i[16996];
  assign o[16995] = i[16995];
  assign o[16994] = i[16994];
  assign o[16993] = i[16993];
  assign o[16992] = i[16992];
  assign o[16991] = i[16991];
  assign o[16990] = i[16990];
  assign o[16989] = i[16989];
  assign o[16988] = i[16988];
  assign o[16987] = i[16987];
  assign o[16986] = i[16986];
  assign o[16985] = i[16985];
  assign o[16984] = i[16984];
  assign o[16983] = i[16983];
  assign o[16982] = i[16982];
  assign o[16981] = i[16981];
  assign o[16980] = i[16980];
  assign o[16979] = i[16979];
  assign o[16978] = i[16978];
  assign o[16977] = i[16977];
  assign o[16976] = i[16976];
  assign o[16975] = i[16975];
  assign o[16974] = i[16974];
  assign o[16973] = i[16973];
  assign o[16972] = i[16972];
  assign o[16971] = i[16971];
  assign o[16970] = i[16970];
  assign o[16969] = i[16969];
  assign o[16968] = i[16968];
  assign o[16967] = i[16967];
  assign o[16966] = i[16966];
  assign o[16965] = i[16965];
  assign o[16964] = i[16964];
  assign o[16963] = i[16963];
  assign o[16962] = i[16962];
  assign o[16961] = i[16961];
  assign o[16960] = i[16960];
  assign o[16959] = i[16959];
  assign o[16958] = i[16958];
  assign o[16957] = i[16957];
  assign o[16956] = i[16956];
  assign o[16955] = i[16955];
  assign o[16954] = i[16954];
  assign o[16953] = i[16953];
  assign o[16952] = i[16952];
  assign o[16951] = i[16951];
  assign o[16950] = i[16950];
  assign o[16949] = i[16949];
  assign o[16948] = i[16948];
  assign o[16947] = i[16947];
  assign o[16946] = i[16946];
  assign o[16945] = i[16945];
  assign o[16944] = i[16944];
  assign o[16943] = i[16943];
  assign o[16942] = i[16942];
  assign o[16941] = i[16941];
  assign o[16940] = i[16940];
  assign o[16939] = i[16939];
  assign o[16938] = i[16938];
  assign o[16937] = i[16937];
  assign o[16936] = i[16936];
  assign o[16935] = i[16935];
  assign o[16934] = i[16934];
  assign o[16933] = i[16933];
  assign o[16932] = i[16932];
  assign o[16931] = i[16931];
  assign o[16930] = i[16930];
  assign o[16929] = i[16929];
  assign o[16928] = i[16928];
  assign o[16927] = i[16927];
  assign o[16926] = i[16926];
  assign o[16925] = i[16925];
  assign o[16924] = i[16924];
  assign o[16923] = i[16923];
  assign o[16922] = i[16922];
  assign o[16921] = i[16921];
  assign o[16920] = i[16920];
  assign o[16919] = i[16919];
  assign o[16918] = i[16918];
  assign o[16917] = i[16917];
  assign o[16916] = i[16916];
  assign o[16915] = i[16915];
  assign o[16914] = i[16914];
  assign o[16913] = i[16913];
  assign o[16912] = i[16912];
  assign o[16911] = i[16911];
  assign o[16910] = i[16910];
  assign o[16909] = i[16909];
  assign o[16908] = i[16908];
  assign o[16907] = i[16907];
  assign o[16906] = i[16906];
  assign o[16905] = i[16905];
  assign o[16904] = i[16904];
  assign o[16903] = i[16903];
  assign o[16902] = i[16902];
  assign o[16901] = i[16901];
  assign o[16900] = i[16900];
  assign o[16899] = i[16899];
  assign o[16898] = i[16898];
  assign o[16897] = i[16897];
  assign o[16896] = i[16896];
  assign o[16895] = i[16895];
  assign o[16894] = i[16894];
  assign o[16893] = i[16893];
  assign o[16892] = i[16892];
  assign o[16891] = i[16891];
  assign o[16890] = i[16890];
  assign o[16889] = i[16889];
  assign o[16888] = i[16888];
  assign o[16887] = i[16887];
  assign o[16886] = i[16886];
  assign o[16885] = i[16885];
  assign o[16884] = i[16884];
  assign o[16883] = i[16883];
  assign o[16882] = i[16882];
  assign o[16881] = i[16881];
  assign o[16880] = i[16880];
  assign o[16879] = i[16879];
  assign o[16878] = i[16878];
  assign o[16877] = i[16877];
  assign o[16876] = i[16876];
  assign o[16875] = i[16875];
  assign o[16874] = i[16874];
  assign o[16873] = i[16873];
  assign o[16872] = i[16872];
  assign o[16871] = i[16871];
  assign o[16870] = i[16870];
  assign o[16869] = i[16869];
  assign o[16868] = i[16868];
  assign o[16867] = i[16867];
  assign o[16866] = i[16866];
  assign o[16865] = i[16865];
  assign o[16864] = i[16864];
  assign o[16863] = i[16863];
  assign o[16862] = i[16862];
  assign o[16861] = i[16861];
  assign o[16860] = i[16860];
  assign o[16859] = i[16859];
  assign o[16858] = i[16858];
  assign o[16857] = i[16857];
  assign o[16856] = i[16856];
  assign o[16855] = i[16855];
  assign o[16854] = i[16854];
  assign o[16853] = i[16853];
  assign o[16852] = i[16852];
  assign o[16851] = i[16851];
  assign o[16850] = i[16850];
  assign o[16849] = i[16849];
  assign o[16848] = i[16848];
  assign o[16847] = i[16847];
  assign o[16846] = i[16846];
  assign o[16845] = i[16845];
  assign o[16844] = i[16844];
  assign o[16843] = i[16843];
  assign o[16842] = i[16842];
  assign o[16841] = i[16841];
  assign o[16840] = i[16840];
  assign o[16839] = i[16839];
  assign o[16838] = i[16838];
  assign o[16837] = i[16837];
  assign o[16836] = i[16836];
  assign o[16835] = i[16835];
  assign o[16834] = i[16834];
  assign o[16833] = i[16833];
  assign o[16832] = i[16832];
  assign o[16831] = i[16831];
  assign o[16830] = i[16830];
  assign o[16829] = i[16829];
  assign o[16828] = i[16828];
  assign o[16827] = i[16827];
  assign o[16826] = i[16826];
  assign o[16825] = i[16825];
  assign o[16824] = i[16824];
  assign o[16823] = i[16823];
  assign o[16822] = i[16822];
  assign o[16821] = i[16821];
  assign o[16820] = i[16820];
  assign o[16819] = i[16819];
  assign o[16818] = i[16818];
  assign o[16817] = i[16817];
  assign o[16816] = i[16816];
  assign o[16815] = i[16815];
  assign o[16814] = i[16814];
  assign o[16813] = i[16813];
  assign o[16812] = i[16812];
  assign o[16811] = i[16811];
  assign o[16810] = i[16810];
  assign o[16809] = i[16809];
  assign o[16808] = i[16808];
  assign o[16807] = i[16807];
  assign o[16806] = i[16806];
  assign o[16805] = i[16805];
  assign o[16804] = i[16804];
  assign o[16803] = i[16803];
  assign o[16802] = i[16802];
  assign o[16801] = i[16801];
  assign o[16800] = i[16800];
  assign o[16799] = i[16799];
  assign o[16798] = i[16798];
  assign o[16797] = i[16797];
  assign o[16796] = i[16796];
  assign o[16795] = i[16795];
  assign o[16794] = i[16794];
  assign o[16793] = i[16793];
  assign o[16792] = i[16792];
  assign o[16791] = i[16791];
  assign o[16790] = i[16790];
  assign o[16789] = i[16789];
  assign o[16788] = i[16788];
  assign o[16787] = i[16787];
  assign o[16786] = i[16786];
  assign o[16785] = i[16785];
  assign o[16784] = i[16784];
  assign o[16783] = i[16783];
  assign o[16782] = i[16782];
  assign o[16781] = i[16781];
  assign o[16780] = i[16780];
  assign o[16779] = i[16779];
  assign o[16778] = i[16778];
  assign o[16777] = i[16777];
  assign o[16776] = i[16776];
  assign o[16775] = i[16775];
  assign o[16774] = i[16774];
  assign o[16773] = i[16773];
  assign o[16772] = i[16772];
  assign o[16771] = i[16771];
  assign o[16770] = i[16770];
  assign o[16769] = i[16769];
  assign o[16768] = i[16768];
  assign o[16767] = i[16767];
  assign o[16766] = i[16766];
  assign o[16765] = i[16765];
  assign o[16764] = i[16764];
  assign o[16763] = i[16763];
  assign o[16762] = i[16762];
  assign o[16761] = i[16761];
  assign o[16760] = i[16760];
  assign o[16759] = i[16759];
  assign o[16758] = i[16758];
  assign o[16757] = i[16757];
  assign o[16756] = i[16756];
  assign o[16755] = i[16755];
  assign o[16754] = i[16754];
  assign o[16753] = i[16753];
  assign o[16752] = i[16752];
  assign o[16751] = i[16751];
  assign o[16750] = i[16750];
  assign o[16749] = i[16749];
  assign o[16748] = i[16748];
  assign o[16747] = i[16747];
  assign o[16746] = i[16746];
  assign o[16745] = i[16745];
  assign o[16744] = i[16744];
  assign o[16743] = i[16743];
  assign o[16742] = i[16742];
  assign o[16741] = i[16741];
  assign o[16740] = i[16740];
  assign o[16739] = i[16739];
  assign o[16738] = i[16738];
  assign o[16737] = i[16737];
  assign o[16736] = i[16736];
  assign o[16735] = i[16735];
  assign o[16734] = i[16734];
  assign o[16733] = i[16733];
  assign o[16732] = i[16732];
  assign o[16731] = i[16731];
  assign o[16730] = i[16730];
  assign o[16729] = i[16729];
  assign o[16728] = i[16728];
  assign o[16727] = i[16727];
  assign o[16726] = i[16726];
  assign o[16725] = i[16725];
  assign o[16724] = i[16724];
  assign o[16723] = i[16723];
  assign o[16722] = i[16722];
  assign o[16721] = i[16721];
  assign o[16720] = i[16720];
  assign o[16719] = i[16719];
  assign o[16718] = i[16718];
  assign o[16717] = i[16717];
  assign o[16716] = i[16716];
  assign o[16715] = i[16715];
  assign o[16714] = i[16714];
  assign o[16713] = i[16713];
  assign o[16712] = i[16712];
  assign o[16711] = i[16711];
  assign o[16710] = i[16710];
  assign o[16709] = i[16709];
  assign o[16708] = i[16708];
  assign o[16707] = i[16707];
  assign o[16706] = i[16706];
  assign o[16705] = i[16705];
  assign o[16704] = i[16704];
  assign o[16703] = i[16703];
  assign o[16702] = i[16702];
  assign o[16701] = i[16701];
  assign o[16700] = i[16700];
  assign o[16699] = i[16699];
  assign o[16698] = i[16698];
  assign o[16697] = i[16697];
  assign o[16696] = i[16696];
  assign o[16695] = i[16695];
  assign o[16694] = i[16694];
  assign o[16693] = i[16693];
  assign o[16692] = i[16692];
  assign o[16691] = i[16691];
  assign o[16690] = i[16690];
  assign o[16689] = i[16689];
  assign o[16688] = i[16688];
  assign o[16687] = i[16687];
  assign o[16686] = i[16686];
  assign o[16685] = i[16685];
  assign o[16684] = i[16684];
  assign o[16683] = i[16683];
  assign o[16682] = i[16682];
  assign o[16681] = i[16681];
  assign o[16680] = i[16680];
  assign o[16679] = i[16679];
  assign o[16678] = i[16678];
  assign o[16677] = i[16677];
  assign o[16676] = i[16676];
  assign o[16675] = i[16675];
  assign o[16674] = i[16674];
  assign o[16673] = i[16673];
  assign o[16672] = i[16672];
  assign o[16671] = i[16671];
  assign o[16670] = i[16670];
  assign o[16669] = i[16669];
  assign o[16668] = i[16668];
  assign o[16667] = i[16667];
  assign o[16666] = i[16666];
  assign o[16665] = i[16665];
  assign o[16664] = i[16664];
  assign o[16663] = i[16663];
  assign o[16662] = i[16662];
  assign o[16661] = i[16661];
  assign o[16660] = i[16660];
  assign o[16659] = i[16659];
  assign o[16658] = i[16658];
  assign o[16657] = i[16657];
  assign o[16656] = i[16656];
  assign o[16655] = i[16655];
  assign o[16654] = i[16654];
  assign o[16653] = i[16653];
  assign o[16652] = i[16652];
  assign o[16651] = i[16651];
  assign o[16650] = i[16650];
  assign o[16649] = i[16649];
  assign o[16648] = i[16648];
  assign o[16647] = i[16647];
  assign o[16646] = i[16646];
  assign o[16645] = i[16645];
  assign o[16644] = i[16644];
  assign o[16643] = i[16643];
  assign o[16642] = i[16642];
  assign o[16641] = i[16641];
  assign o[16640] = i[16640];
  assign o[16639] = i[16639];
  assign o[16638] = i[16638];
  assign o[16637] = i[16637];
  assign o[16636] = i[16636];
  assign o[16635] = i[16635];
  assign o[16634] = i[16634];
  assign o[16633] = i[16633];
  assign o[16632] = i[16632];
  assign o[16631] = i[16631];
  assign o[16630] = i[16630];
  assign o[16629] = i[16629];
  assign o[16628] = i[16628];
  assign o[16627] = i[16627];
  assign o[16626] = i[16626];
  assign o[16625] = i[16625];
  assign o[16624] = i[16624];
  assign o[16623] = i[16623];
  assign o[16622] = i[16622];
  assign o[16621] = i[16621];
  assign o[16620] = i[16620];
  assign o[16619] = i[16619];
  assign o[16618] = i[16618];
  assign o[16617] = i[16617];
  assign o[16616] = i[16616];
  assign o[16615] = i[16615];
  assign o[16614] = i[16614];
  assign o[16613] = i[16613];
  assign o[16612] = i[16612];
  assign o[16611] = i[16611];
  assign o[16610] = i[16610];
  assign o[16609] = i[16609];
  assign o[16608] = i[16608];
  assign o[16607] = i[16607];
  assign o[16606] = i[16606];
  assign o[16605] = i[16605];
  assign o[16604] = i[16604];
  assign o[16603] = i[16603];
  assign o[16602] = i[16602];
  assign o[16601] = i[16601];
  assign o[16600] = i[16600];
  assign o[16599] = i[16599];
  assign o[16598] = i[16598];
  assign o[16597] = i[16597];
  assign o[16596] = i[16596];
  assign o[16595] = i[16595];
  assign o[16594] = i[16594];
  assign o[16593] = i[16593];
  assign o[16592] = i[16592];
  assign o[16591] = i[16591];
  assign o[16590] = i[16590];
  assign o[16589] = i[16589];
  assign o[16588] = i[16588];
  assign o[16587] = i[16587];
  assign o[16586] = i[16586];
  assign o[16585] = i[16585];
  assign o[16584] = i[16584];
  assign o[16583] = i[16583];
  assign o[16582] = i[16582];
  assign o[16581] = i[16581];
  assign o[16580] = i[16580];
  assign o[16579] = i[16579];
  assign o[16578] = i[16578];
  assign o[16577] = i[16577];
  assign o[16576] = i[16576];
  assign o[16575] = i[16575];
  assign o[16574] = i[16574];
  assign o[16573] = i[16573];
  assign o[16572] = i[16572];
  assign o[16571] = i[16571];
  assign o[16570] = i[16570];
  assign o[16569] = i[16569];
  assign o[16568] = i[16568];
  assign o[16567] = i[16567];
  assign o[16566] = i[16566];
  assign o[16565] = i[16565];
  assign o[16564] = i[16564];
  assign o[16563] = i[16563];
  assign o[16562] = i[16562];
  assign o[16561] = i[16561];
  assign o[16560] = i[16560];
  assign o[16559] = i[16559];
  assign o[16558] = i[16558];
  assign o[16557] = i[16557];
  assign o[16556] = i[16556];
  assign o[16555] = i[16555];
  assign o[16554] = i[16554];
  assign o[16553] = i[16553];
  assign o[16552] = i[16552];
  assign o[16551] = i[16551];
  assign o[16550] = i[16550];
  assign o[16549] = i[16549];
  assign o[16548] = i[16548];
  assign o[16547] = i[16547];
  assign o[16546] = i[16546];
  assign o[16545] = i[16545];
  assign o[16544] = i[16544];
  assign o[16543] = i[16543];
  assign o[16542] = i[16542];
  assign o[16541] = i[16541];
  assign o[16540] = i[16540];
  assign o[16539] = i[16539];
  assign o[16538] = i[16538];
  assign o[16537] = i[16537];
  assign o[16536] = i[16536];
  assign o[16535] = i[16535];
  assign o[16534] = i[16534];
  assign o[16533] = i[16533];
  assign o[16532] = i[16532];
  assign o[16531] = i[16531];
  assign o[16530] = i[16530];
  assign o[16529] = i[16529];
  assign o[16528] = i[16528];
  assign o[16527] = i[16527];
  assign o[16526] = i[16526];
  assign o[16525] = i[16525];
  assign o[16524] = i[16524];
  assign o[16523] = i[16523];
  assign o[16522] = i[16522];
  assign o[16521] = i[16521];
  assign o[16520] = i[16520];
  assign o[16519] = i[16519];
  assign o[16518] = i[16518];
  assign o[16517] = i[16517];
  assign o[16516] = i[16516];
  assign o[16515] = i[16515];
  assign o[16514] = i[16514];
  assign o[16513] = i[16513];
  assign o[16512] = i[16512];
  assign o[16511] = i[16511];
  assign o[16510] = i[16510];
  assign o[16509] = i[16509];
  assign o[16508] = i[16508];
  assign o[16507] = i[16507];
  assign o[16506] = i[16506];
  assign o[16505] = i[16505];
  assign o[16504] = i[16504];
  assign o[16503] = i[16503];
  assign o[16502] = i[16502];
  assign o[16501] = i[16501];
  assign o[16500] = i[16500];
  assign o[16499] = i[16499];
  assign o[16498] = i[16498];
  assign o[16497] = i[16497];
  assign o[16496] = i[16496];
  assign o[16495] = i[16495];
  assign o[16494] = i[16494];
  assign o[16493] = i[16493];
  assign o[16492] = i[16492];
  assign o[16491] = i[16491];
  assign o[16490] = i[16490];
  assign o[16489] = i[16489];
  assign o[16488] = i[16488];
  assign o[16487] = i[16487];
  assign o[16486] = i[16486];
  assign o[16485] = i[16485];
  assign o[16484] = i[16484];
  assign o[16483] = i[16483];
  assign o[16482] = i[16482];
  assign o[16481] = i[16481];
  assign o[16480] = i[16480];
  assign o[16479] = i[16479];
  assign o[16478] = i[16478];
  assign o[16477] = i[16477];
  assign o[16476] = i[16476];
  assign o[16475] = i[16475];
  assign o[16474] = i[16474];
  assign o[16473] = i[16473];
  assign o[16472] = i[16472];
  assign o[16471] = i[16471];
  assign o[16470] = i[16470];
  assign o[16469] = i[16469];
  assign o[16468] = i[16468];
  assign o[16467] = i[16467];
  assign o[16466] = i[16466];
  assign o[16465] = i[16465];
  assign o[16464] = i[16464];
  assign o[16463] = i[16463];
  assign o[16462] = i[16462];
  assign o[16461] = i[16461];
  assign o[16460] = i[16460];
  assign o[16459] = i[16459];
  assign o[16458] = i[16458];
  assign o[16457] = i[16457];
  assign o[16456] = i[16456];
  assign o[16455] = i[16455];
  assign o[16454] = i[16454];
  assign o[16453] = i[16453];
  assign o[16452] = i[16452];
  assign o[16451] = i[16451];
  assign o[16450] = i[16450];
  assign o[16449] = i[16449];
  assign o[16448] = i[16448];
  assign o[16447] = i[16447];
  assign o[16446] = i[16446];
  assign o[16445] = i[16445];
  assign o[16444] = i[16444];
  assign o[16443] = i[16443];
  assign o[16442] = i[16442];
  assign o[16441] = i[16441];
  assign o[16440] = i[16440];
  assign o[16439] = i[16439];
  assign o[16438] = i[16438];
  assign o[16437] = i[16437];
  assign o[16436] = i[16436];
  assign o[16435] = i[16435];
  assign o[16434] = i[16434];
  assign o[16433] = i[16433];
  assign o[16432] = i[16432];
  assign o[16431] = i[16431];
  assign o[16430] = i[16430];
  assign o[16429] = i[16429];
  assign o[16428] = i[16428];
  assign o[16427] = i[16427];
  assign o[16426] = i[16426];
  assign o[16425] = i[16425];
  assign o[16424] = i[16424];
  assign o[16423] = i[16423];
  assign o[16422] = i[16422];
  assign o[16421] = i[16421];
  assign o[16420] = i[16420];
  assign o[16419] = i[16419];
  assign o[16418] = i[16418];
  assign o[16417] = i[16417];
  assign o[16416] = i[16416];
  assign o[16415] = i[16415];
  assign o[16414] = i[16414];
  assign o[16413] = i[16413];
  assign o[16412] = i[16412];
  assign o[16411] = i[16411];
  assign o[16410] = i[16410];
  assign o[16409] = i[16409];
  assign o[16408] = i[16408];
  assign o[16407] = i[16407];
  assign o[16406] = i[16406];
  assign o[16405] = i[16405];
  assign o[16404] = i[16404];
  assign o[16403] = i[16403];
  assign o[16402] = i[16402];
  assign o[16401] = i[16401];
  assign o[16400] = i[16400];
  assign o[16399] = i[16399];
  assign o[16398] = i[16398];
  assign o[16397] = i[16397];
  assign o[16396] = i[16396];
  assign o[16395] = i[16395];
  assign o[16394] = i[16394];
  assign o[16393] = i[16393];
  assign o[16392] = i[16392];
  assign o[16391] = i[16391];
  assign o[16390] = i[16390];
  assign o[16389] = i[16389];
  assign o[16388] = i[16388];
  assign o[16387] = i[16387];
  assign o[16386] = i[16386];
  assign o[16385] = i[16385];
  assign o[16384] = i[16384];
  assign o[16383] = i[16383];
  assign o[16382] = i[16382];
  assign o[16381] = i[16381];
  assign o[16380] = i[16380];
  assign o[16379] = i[16379];
  assign o[16378] = i[16378];
  assign o[16377] = i[16377];
  assign o[16376] = i[16376];
  assign o[16375] = i[16375];
  assign o[16374] = i[16374];
  assign o[16373] = i[16373];
  assign o[16372] = i[16372];
  assign o[16371] = i[16371];
  assign o[16370] = i[16370];
  assign o[16369] = i[16369];
  assign o[16368] = i[16368];
  assign o[16367] = i[16367];
  assign o[16366] = i[16366];
  assign o[16365] = i[16365];
  assign o[16364] = i[16364];
  assign o[16363] = i[16363];
  assign o[16362] = i[16362];
  assign o[16361] = i[16361];
  assign o[16360] = i[16360];
  assign o[16359] = i[16359];
  assign o[16358] = i[16358];
  assign o[16357] = i[16357];
  assign o[16356] = i[16356];
  assign o[16355] = i[16355];
  assign o[16354] = i[16354];
  assign o[16353] = i[16353];
  assign o[16352] = i[16352];
  assign o[16351] = i[16351];
  assign o[16350] = i[16350];
  assign o[16349] = i[16349];
  assign o[16348] = i[16348];
  assign o[16347] = i[16347];
  assign o[16346] = i[16346];
  assign o[16345] = i[16345];
  assign o[16344] = i[16344];
  assign o[16343] = i[16343];
  assign o[16342] = i[16342];
  assign o[16341] = i[16341];
  assign o[16340] = i[16340];
  assign o[16339] = i[16339];
  assign o[16338] = i[16338];
  assign o[16337] = i[16337];
  assign o[16336] = i[16336];
  assign o[16335] = i[16335];
  assign o[16334] = i[16334];
  assign o[16333] = i[16333];
  assign o[16332] = i[16332];
  assign o[16331] = i[16331];
  assign o[16330] = i[16330];
  assign o[16329] = i[16329];
  assign o[16328] = i[16328];
  assign o[16327] = i[16327];
  assign o[16326] = i[16326];
  assign o[16325] = i[16325];
  assign o[16324] = i[16324];
  assign o[16323] = i[16323];
  assign o[16322] = i[16322];
  assign o[16321] = i[16321];
  assign o[16320] = i[16320];
  assign o[16319] = i[16319];
  assign o[16318] = i[16318];
  assign o[16317] = i[16317];
  assign o[16316] = i[16316];
  assign o[16315] = i[16315];
  assign o[16314] = i[16314];
  assign o[16313] = i[16313];
  assign o[16312] = i[16312];
  assign o[16311] = i[16311];
  assign o[16310] = i[16310];
  assign o[16309] = i[16309];
  assign o[16308] = i[16308];
  assign o[16307] = i[16307];
  assign o[16306] = i[16306];
  assign o[16305] = i[16305];
  assign o[16304] = i[16304];
  assign o[16303] = i[16303];
  assign o[16302] = i[16302];
  assign o[16301] = i[16301];
  assign o[16300] = i[16300];
  assign o[16299] = i[16299];
  assign o[16298] = i[16298];
  assign o[16297] = i[16297];
  assign o[16296] = i[16296];
  assign o[16295] = i[16295];
  assign o[16294] = i[16294];
  assign o[16293] = i[16293];
  assign o[16292] = i[16292];
  assign o[16291] = i[16291];
  assign o[16290] = i[16290];
  assign o[16289] = i[16289];
  assign o[16288] = i[16288];
  assign o[16287] = i[16287];
  assign o[16286] = i[16286];
  assign o[16285] = i[16285];
  assign o[16284] = i[16284];
  assign o[16283] = i[16283];
  assign o[16282] = i[16282];
  assign o[16281] = i[16281];
  assign o[16280] = i[16280];
  assign o[16279] = i[16279];
  assign o[16278] = i[16278];
  assign o[16277] = i[16277];
  assign o[16276] = i[16276];
  assign o[16275] = i[16275];
  assign o[16274] = i[16274];
  assign o[16273] = i[16273];
  assign o[16272] = i[16272];
  assign o[16271] = i[16271];
  assign o[16270] = i[16270];
  assign o[16269] = i[16269];
  assign o[16268] = i[16268];
  assign o[16267] = i[16267];
  assign o[16266] = i[16266];
  assign o[16265] = i[16265];
  assign o[16264] = i[16264];
  assign o[16263] = i[16263];
  assign o[16262] = i[16262];
  assign o[16261] = i[16261];
  assign o[16260] = i[16260];
  assign o[16259] = i[16259];
  assign o[16258] = i[16258];
  assign o[16257] = i[16257];
  assign o[16256] = i[16256];
  assign o[16255] = i[16255];
  assign o[16254] = i[16254];
  assign o[16253] = i[16253];
  assign o[16252] = i[16252];
  assign o[16251] = i[16251];
  assign o[16250] = i[16250];
  assign o[16249] = i[16249];
  assign o[16248] = i[16248];
  assign o[16247] = i[16247];
  assign o[16246] = i[16246];
  assign o[16245] = i[16245];
  assign o[16244] = i[16244];
  assign o[16243] = i[16243];
  assign o[16242] = i[16242];
  assign o[16241] = i[16241];
  assign o[16240] = i[16240];
  assign o[16239] = i[16239];
  assign o[16238] = i[16238];
  assign o[16237] = i[16237];
  assign o[16236] = i[16236];
  assign o[16235] = i[16235];
  assign o[16234] = i[16234];
  assign o[16233] = i[16233];
  assign o[16232] = i[16232];
  assign o[16231] = i[16231];
  assign o[16230] = i[16230];
  assign o[16229] = i[16229];
  assign o[16228] = i[16228];
  assign o[16227] = i[16227];
  assign o[16226] = i[16226];
  assign o[16225] = i[16225];
  assign o[16224] = i[16224];
  assign o[16223] = i[16223];
  assign o[16222] = i[16222];
  assign o[16221] = i[16221];
  assign o[16220] = i[16220];
  assign o[16219] = i[16219];
  assign o[16218] = i[16218];
  assign o[16217] = i[16217];
  assign o[16216] = i[16216];
  assign o[16215] = i[16215];
  assign o[16214] = i[16214];
  assign o[16213] = i[16213];
  assign o[16212] = i[16212];
  assign o[16211] = i[16211];
  assign o[16210] = i[16210];
  assign o[16209] = i[16209];
  assign o[16208] = i[16208];
  assign o[16207] = i[16207];
  assign o[16206] = i[16206];
  assign o[16205] = i[16205];
  assign o[16204] = i[16204];
  assign o[16203] = i[16203];
  assign o[16202] = i[16202];
  assign o[16201] = i[16201];
  assign o[16200] = i[16200];
  assign o[16199] = i[16199];
  assign o[16198] = i[16198];
  assign o[16197] = i[16197];
  assign o[16196] = i[16196];
  assign o[16195] = i[16195];
  assign o[16194] = i[16194];
  assign o[16193] = i[16193];
  assign o[16192] = i[16192];
  assign o[16191] = i[16191];
  assign o[16190] = i[16190];
  assign o[16189] = i[16189];
  assign o[16188] = i[16188];
  assign o[16187] = i[16187];
  assign o[16186] = i[16186];
  assign o[16185] = i[16185];
  assign o[16184] = i[16184];
  assign o[16183] = i[16183];
  assign o[16182] = i[16182];
  assign o[16181] = i[16181];
  assign o[16180] = i[16180];
  assign o[16179] = i[16179];
  assign o[16178] = i[16178];
  assign o[16177] = i[16177];
  assign o[16176] = i[16176];
  assign o[16175] = i[16175];
  assign o[16174] = i[16174];
  assign o[16173] = i[16173];
  assign o[16172] = i[16172];
  assign o[16171] = i[16171];
  assign o[16170] = i[16170];
  assign o[16169] = i[16169];
  assign o[16168] = i[16168];
  assign o[16167] = i[16167];
  assign o[16166] = i[16166];
  assign o[16165] = i[16165];
  assign o[16164] = i[16164];
  assign o[16163] = i[16163];
  assign o[16162] = i[16162];
  assign o[16161] = i[16161];
  assign o[16160] = i[16160];
  assign o[16159] = i[16159];
  assign o[16158] = i[16158];
  assign o[16157] = i[16157];
  assign o[16156] = i[16156];
  assign o[16155] = i[16155];
  assign o[16154] = i[16154];
  assign o[16153] = i[16153];
  assign o[16152] = i[16152];
  assign o[16151] = i[16151];
  assign o[16150] = i[16150];
  assign o[16149] = i[16149];
  assign o[16148] = i[16148];
  assign o[16147] = i[16147];
  assign o[16146] = i[16146];
  assign o[16145] = i[16145];
  assign o[16144] = i[16144];
  assign o[16143] = i[16143];
  assign o[16142] = i[16142];
  assign o[16141] = i[16141];
  assign o[16140] = i[16140];
  assign o[16139] = i[16139];
  assign o[16138] = i[16138];
  assign o[16137] = i[16137];
  assign o[16136] = i[16136];
  assign o[16135] = i[16135];
  assign o[16134] = i[16134];
  assign o[16133] = i[16133];
  assign o[16132] = i[16132];
  assign o[16131] = i[16131];
  assign o[16130] = i[16130];
  assign o[16129] = i[16129];
  assign o[16128] = i[16128];
  assign o[16127] = i[16127];
  assign o[16126] = i[16126];
  assign o[16125] = i[16125];
  assign o[16124] = i[16124];
  assign o[16123] = i[16123];
  assign o[16122] = i[16122];
  assign o[16121] = i[16121];
  assign o[16120] = i[16120];
  assign o[16119] = i[16119];
  assign o[16118] = i[16118];
  assign o[16117] = i[16117];
  assign o[16116] = i[16116];
  assign o[16115] = i[16115];
  assign o[16114] = i[16114];
  assign o[16113] = i[16113];
  assign o[16112] = i[16112];
  assign o[16111] = i[16111];
  assign o[16110] = i[16110];
  assign o[16109] = i[16109];
  assign o[16108] = i[16108];
  assign o[16107] = i[16107];
  assign o[16106] = i[16106];
  assign o[16105] = i[16105];
  assign o[16104] = i[16104];
  assign o[16103] = i[16103];
  assign o[16102] = i[16102];
  assign o[16101] = i[16101];
  assign o[16100] = i[16100];
  assign o[16099] = i[16099];
  assign o[16098] = i[16098];
  assign o[16097] = i[16097];
  assign o[16096] = i[16096];
  assign o[16095] = i[16095];
  assign o[16094] = i[16094];
  assign o[16093] = i[16093];
  assign o[16092] = i[16092];
  assign o[16091] = i[16091];
  assign o[16090] = i[16090];
  assign o[16089] = i[16089];
  assign o[16088] = i[16088];
  assign o[16087] = i[16087];
  assign o[16086] = i[16086];
  assign o[16085] = i[16085];
  assign o[16084] = i[16084];
  assign o[16083] = i[16083];
  assign o[16082] = i[16082];
  assign o[16081] = i[16081];
  assign o[16080] = i[16080];
  assign o[16079] = i[16079];
  assign o[16078] = i[16078];
  assign o[16077] = i[16077];
  assign o[16076] = i[16076];
  assign o[16075] = i[16075];
  assign o[16074] = i[16074];
  assign o[16073] = i[16073];
  assign o[16072] = i[16072];
  assign o[16071] = i[16071];
  assign o[16070] = i[16070];
  assign o[16069] = i[16069];
  assign o[16068] = i[16068];
  assign o[16067] = i[16067];
  assign o[16066] = i[16066];
  assign o[16065] = i[16065];
  assign o[16064] = i[16064];
  assign o[16063] = i[16063];
  assign o[16062] = i[16062];
  assign o[16061] = i[16061];
  assign o[16060] = i[16060];
  assign o[16059] = i[16059];
  assign o[16058] = i[16058];
  assign o[16057] = i[16057];
  assign o[16056] = i[16056];
  assign o[16055] = i[16055];
  assign o[16054] = i[16054];
  assign o[16053] = i[16053];
  assign o[16052] = i[16052];
  assign o[16051] = i[16051];
  assign o[16050] = i[16050];
  assign o[16049] = i[16049];
  assign o[16048] = i[16048];
  assign o[16047] = i[16047];
  assign o[16046] = i[16046];
  assign o[16045] = i[16045];
  assign o[16044] = i[16044];
  assign o[16043] = i[16043];
  assign o[16042] = i[16042];
  assign o[16041] = i[16041];
  assign o[16040] = i[16040];
  assign o[16039] = i[16039];
  assign o[16038] = i[16038];
  assign o[16037] = i[16037];
  assign o[16036] = i[16036];
  assign o[16035] = i[16035];
  assign o[16034] = i[16034];
  assign o[16033] = i[16033];
  assign o[16032] = i[16032];
  assign o[16031] = i[16031];
  assign o[16030] = i[16030];
  assign o[16029] = i[16029];
  assign o[16028] = i[16028];
  assign o[16027] = i[16027];
  assign o[16026] = i[16026];
  assign o[16025] = i[16025];
  assign o[16024] = i[16024];
  assign o[16023] = i[16023];
  assign o[16022] = i[16022];
  assign o[16021] = i[16021];
  assign o[16020] = i[16020];
  assign o[16019] = i[16019];
  assign o[16018] = i[16018];
  assign o[16017] = i[16017];
  assign o[16016] = i[16016];
  assign o[16015] = i[16015];
  assign o[16014] = i[16014];
  assign o[16013] = i[16013];
  assign o[16012] = i[16012];
  assign o[16011] = i[16011];
  assign o[16010] = i[16010];
  assign o[16009] = i[16009];
  assign o[16008] = i[16008];
  assign o[16007] = i[16007];
  assign o[16006] = i[16006];
  assign o[16005] = i[16005];
  assign o[16004] = i[16004];
  assign o[16003] = i[16003];
  assign o[16002] = i[16002];
  assign o[16001] = i[16001];
  assign o[16000] = i[16000];
  assign o[15999] = i[15999];
  assign o[15998] = i[15998];
  assign o[15997] = i[15997];
  assign o[15996] = i[15996];
  assign o[15995] = i[15995];
  assign o[15994] = i[15994];
  assign o[15993] = i[15993];
  assign o[15992] = i[15992];
  assign o[15991] = i[15991];
  assign o[15990] = i[15990];
  assign o[15989] = i[15989];
  assign o[15988] = i[15988];
  assign o[15987] = i[15987];
  assign o[15986] = i[15986];
  assign o[15985] = i[15985];
  assign o[15984] = i[15984];
  assign o[15983] = i[15983];
  assign o[15982] = i[15982];
  assign o[15981] = i[15981];
  assign o[15980] = i[15980];
  assign o[15979] = i[15979];
  assign o[15978] = i[15978];
  assign o[15977] = i[15977];
  assign o[15976] = i[15976];
  assign o[15975] = i[15975];
  assign o[15974] = i[15974];
  assign o[15973] = i[15973];
  assign o[15972] = i[15972];
  assign o[15971] = i[15971];
  assign o[15970] = i[15970];
  assign o[15969] = i[15969];
  assign o[15968] = i[15968];
  assign o[15967] = i[15967];
  assign o[15966] = i[15966];
  assign o[15965] = i[15965];
  assign o[15964] = i[15964];
  assign o[15963] = i[15963];
  assign o[15962] = i[15962];
  assign o[15961] = i[15961];
  assign o[15960] = i[15960];
  assign o[15959] = i[15959];
  assign o[15958] = i[15958];
  assign o[15957] = i[15957];
  assign o[15956] = i[15956];
  assign o[15955] = i[15955];
  assign o[15954] = i[15954];
  assign o[15953] = i[15953];
  assign o[15952] = i[15952];
  assign o[15951] = i[15951];
  assign o[15950] = i[15950];
  assign o[15949] = i[15949];
  assign o[15948] = i[15948];
  assign o[15947] = i[15947];
  assign o[15946] = i[15946];
  assign o[15945] = i[15945];
  assign o[15944] = i[15944];
  assign o[15943] = i[15943];
  assign o[15942] = i[15942];
  assign o[15941] = i[15941];
  assign o[15940] = i[15940];
  assign o[15939] = i[15939];
  assign o[15938] = i[15938];
  assign o[15937] = i[15937];
  assign o[15936] = i[15936];
  assign o[15935] = i[15935];
  assign o[15934] = i[15934];
  assign o[15933] = i[15933];
  assign o[15932] = i[15932];
  assign o[15931] = i[15931];
  assign o[15930] = i[15930];
  assign o[15929] = i[15929];
  assign o[15928] = i[15928];
  assign o[15927] = i[15927];
  assign o[15926] = i[15926];
  assign o[15925] = i[15925];
  assign o[15924] = i[15924];
  assign o[15923] = i[15923];
  assign o[15922] = i[15922];
  assign o[15921] = i[15921];
  assign o[15920] = i[15920];
  assign o[15919] = i[15919];
  assign o[15918] = i[15918];
  assign o[15917] = i[15917];
  assign o[15916] = i[15916];
  assign o[15915] = i[15915];
  assign o[15914] = i[15914];
  assign o[15913] = i[15913];
  assign o[15912] = i[15912];
  assign o[15911] = i[15911];
  assign o[15910] = i[15910];
  assign o[15909] = i[15909];
  assign o[15908] = i[15908];
  assign o[15907] = i[15907];
  assign o[15906] = i[15906];
  assign o[15905] = i[15905];
  assign o[15904] = i[15904];
  assign o[15903] = i[15903];
  assign o[15902] = i[15902];
  assign o[15901] = i[15901];
  assign o[15900] = i[15900];
  assign o[15899] = i[15899];
  assign o[15898] = i[15898];
  assign o[15897] = i[15897];
  assign o[15896] = i[15896];
  assign o[15895] = i[15895];
  assign o[15894] = i[15894];
  assign o[15893] = i[15893];
  assign o[15892] = i[15892];
  assign o[15891] = i[15891];
  assign o[15890] = i[15890];
  assign o[15889] = i[15889];
  assign o[15888] = i[15888];
  assign o[15887] = i[15887];
  assign o[15886] = i[15886];
  assign o[15885] = i[15885];
  assign o[15884] = i[15884];
  assign o[15883] = i[15883];
  assign o[15882] = i[15882];
  assign o[15881] = i[15881];
  assign o[15880] = i[15880];
  assign o[15879] = i[15879];
  assign o[15878] = i[15878];
  assign o[15877] = i[15877];
  assign o[15876] = i[15876];
  assign o[15875] = i[15875];
  assign o[15874] = i[15874];
  assign o[15873] = i[15873];
  assign o[15872] = i[15872];
  assign o[15871] = i[15871];
  assign o[15870] = i[15870];
  assign o[15869] = i[15869];
  assign o[15868] = i[15868];
  assign o[15867] = i[15867];
  assign o[15866] = i[15866];
  assign o[15865] = i[15865];
  assign o[15864] = i[15864];
  assign o[15863] = i[15863];
  assign o[15862] = i[15862];
  assign o[15861] = i[15861];
  assign o[15860] = i[15860];
  assign o[15859] = i[15859];
  assign o[15858] = i[15858];
  assign o[15857] = i[15857];
  assign o[15856] = i[15856];
  assign o[15855] = i[15855];
  assign o[15854] = i[15854];
  assign o[15853] = i[15853];
  assign o[15852] = i[15852];
  assign o[15851] = i[15851];
  assign o[15850] = i[15850];
  assign o[15849] = i[15849];
  assign o[15848] = i[15848];
  assign o[15847] = i[15847];
  assign o[15846] = i[15846];
  assign o[15845] = i[15845];
  assign o[15844] = i[15844];
  assign o[15843] = i[15843];
  assign o[15842] = i[15842];
  assign o[15841] = i[15841];
  assign o[15840] = i[15840];
  assign o[15839] = i[15839];
  assign o[15838] = i[15838];
  assign o[15837] = i[15837];
  assign o[15836] = i[15836];
  assign o[15835] = i[15835];
  assign o[15834] = i[15834];
  assign o[15833] = i[15833];
  assign o[15832] = i[15832];
  assign o[15831] = i[15831];
  assign o[15830] = i[15830];
  assign o[15829] = i[15829];
  assign o[15828] = i[15828];
  assign o[15827] = i[15827];
  assign o[15826] = i[15826];
  assign o[15825] = i[15825];
  assign o[15824] = i[15824];
  assign o[15823] = i[15823];
  assign o[15822] = i[15822];
  assign o[15821] = i[15821];
  assign o[15820] = i[15820];
  assign o[15819] = i[15819];
  assign o[15818] = i[15818];
  assign o[15817] = i[15817];
  assign o[15816] = i[15816];
  assign o[15815] = i[15815];
  assign o[15814] = i[15814];
  assign o[15813] = i[15813];
  assign o[15812] = i[15812];
  assign o[15811] = i[15811];
  assign o[15810] = i[15810];
  assign o[15809] = i[15809];
  assign o[15808] = i[15808];
  assign o[15807] = i[15807];
  assign o[15806] = i[15806];
  assign o[15805] = i[15805];
  assign o[15804] = i[15804];
  assign o[15803] = i[15803];
  assign o[15802] = i[15802];
  assign o[15801] = i[15801];
  assign o[15800] = i[15800];
  assign o[15799] = i[15799];
  assign o[15798] = i[15798];
  assign o[15797] = i[15797];
  assign o[15796] = i[15796];
  assign o[15795] = i[15795];
  assign o[15794] = i[15794];
  assign o[15793] = i[15793];
  assign o[15792] = i[15792];
  assign o[15791] = i[15791];
  assign o[15790] = i[15790];
  assign o[15789] = i[15789];
  assign o[15788] = i[15788];
  assign o[15787] = i[15787];
  assign o[15786] = i[15786];
  assign o[15785] = i[15785];
  assign o[15784] = i[15784];
  assign o[15783] = i[15783];
  assign o[15782] = i[15782];
  assign o[15781] = i[15781];
  assign o[15780] = i[15780];
  assign o[15779] = i[15779];
  assign o[15778] = i[15778];
  assign o[15777] = i[15777];
  assign o[15776] = i[15776];
  assign o[15775] = i[15775];
  assign o[15774] = i[15774];
  assign o[15773] = i[15773];
  assign o[15772] = i[15772];
  assign o[15771] = i[15771];
  assign o[15770] = i[15770];
  assign o[15769] = i[15769];
  assign o[15768] = i[15768];
  assign o[15767] = i[15767];
  assign o[15766] = i[15766];
  assign o[15765] = i[15765];
  assign o[15764] = i[15764];
  assign o[15763] = i[15763];
  assign o[15762] = i[15762];
  assign o[15761] = i[15761];
  assign o[15760] = i[15760];
  assign o[15759] = i[15759];
  assign o[15758] = i[15758];
  assign o[15757] = i[15757];
  assign o[15756] = i[15756];
  assign o[15755] = i[15755];
  assign o[15754] = i[15754];
  assign o[15753] = i[15753];
  assign o[15752] = i[15752];
  assign o[15751] = i[15751];
  assign o[15750] = i[15750];
  assign o[15749] = i[15749];
  assign o[15748] = i[15748];
  assign o[15747] = i[15747];
  assign o[15746] = i[15746];
  assign o[15745] = i[15745];
  assign o[15744] = i[15744];
  assign o[15743] = i[15743];
  assign o[15742] = i[15742];
  assign o[15741] = i[15741];
  assign o[15740] = i[15740];
  assign o[15739] = i[15739];
  assign o[15738] = i[15738];
  assign o[15737] = i[15737];
  assign o[15736] = i[15736];
  assign o[15735] = i[15735];
  assign o[15734] = i[15734];
  assign o[15733] = i[15733];
  assign o[15732] = i[15732];
  assign o[15731] = i[15731];
  assign o[15730] = i[15730];
  assign o[15729] = i[15729];
  assign o[15728] = i[15728];
  assign o[15727] = i[15727];
  assign o[15726] = i[15726];
  assign o[15725] = i[15725];
  assign o[15724] = i[15724];
  assign o[15723] = i[15723];
  assign o[15722] = i[15722];
  assign o[15721] = i[15721];
  assign o[15720] = i[15720];
  assign o[15719] = i[15719];
  assign o[15718] = i[15718];
  assign o[15717] = i[15717];
  assign o[15716] = i[15716];
  assign o[15715] = i[15715];
  assign o[15714] = i[15714];
  assign o[15713] = i[15713];
  assign o[15712] = i[15712];
  assign o[15711] = i[15711];
  assign o[15710] = i[15710];
  assign o[15709] = i[15709];
  assign o[15708] = i[15708];
  assign o[15707] = i[15707];
  assign o[15706] = i[15706];
  assign o[15705] = i[15705];
  assign o[15704] = i[15704];
  assign o[15703] = i[15703];
  assign o[15702] = i[15702];
  assign o[15701] = i[15701];
  assign o[15700] = i[15700];
  assign o[15699] = i[15699];
  assign o[15698] = i[15698];
  assign o[15697] = i[15697];
  assign o[15696] = i[15696];
  assign o[15695] = i[15695];
  assign o[15694] = i[15694];
  assign o[15693] = i[15693];
  assign o[15692] = i[15692];
  assign o[15691] = i[15691];
  assign o[15690] = i[15690];
  assign o[15689] = i[15689];
  assign o[15688] = i[15688];
  assign o[15687] = i[15687];
  assign o[15686] = i[15686];
  assign o[15685] = i[15685];
  assign o[15684] = i[15684];
  assign o[15683] = i[15683];
  assign o[15682] = i[15682];
  assign o[15681] = i[15681];
  assign o[15680] = i[15680];
  assign o[15679] = i[15679];
  assign o[15678] = i[15678];
  assign o[15677] = i[15677];
  assign o[15676] = i[15676];
  assign o[15675] = i[15675];
  assign o[15674] = i[15674];
  assign o[15673] = i[15673];
  assign o[15672] = i[15672];
  assign o[15671] = i[15671];
  assign o[15670] = i[15670];
  assign o[15669] = i[15669];
  assign o[15668] = i[15668];
  assign o[15667] = i[15667];
  assign o[15666] = i[15666];
  assign o[15665] = i[15665];
  assign o[15664] = i[15664];
  assign o[15663] = i[15663];
  assign o[15662] = i[15662];
  assign o[15661] = i[15661];
  assign o[15660] = i[15660];
  assign o[15659] = i[15659];
  assign o[15658] = i[15658];
  assign o[15657] = i[15657];
  assign o[15656] = i[15656];
  assign o[15655] = i[15655];
  assign o[15654] = i[15654];
  assign o[15653] = i[15653];
  assign o[15652] = i[15652];
  assign o[15651] = i[15651];
  assign o[15650] = i[15650];
  assign o[15649] = i[15649];
  assign o[15648] = i[15648];
  assign o[15647] = i[15647];
  assign o[15646] = i[15646];
  assign o[15645] = i[15645];
  assign o[15644] = i[15644];
  assign o[15643] = i[15643];
  assign o[15642] = i[15642];
  assign o[15641] = i[15641];
  assign o[15640] = i[15640];
  assign o[15639] = i[15639];
  assign o[15638] = i[15638];
  assign o[15637] = i[15637];
  assign o[15636] = i[15636];
  assign o[15635] = i[15635];
  assign o[15634] = i[15634];
  assign o[15633] = i[15633];
  assign o[15632] = i[15632];
  assign o[15631] = i[15631];
  assign o[15630] = i[15630];
  assign o[15629] = i[15629];
  assign o[15628] = i[15628];
  assign o[15627] = i[15627];
  assign o[15626] = i[15626];
  assign o[15625] = i[15625];
  assign o[15624] = i[15624];
  assign o[15623] = i[15623];
  assign o[15622] = i[15622];
  assign o[15621] = i[15621];
  assign o[15620] = i[15620];
  assign o[15619] = i[15619];
  assign o[15618] = i[15618];
  assign o[15617] = i[15617];
  assign o[15616] = i[15616];
  assign o[15615] = i[15615];
  assign o[15614] = i[15614];
  assign o[15613] = i[15613];
  assign o[15612] = i[15612];
  assign o[15611] = i[15611];
  assign o[15610] = i[15610];
  assign o[15609] = i[15609];
  assign o[15608] = i[15608];
  assign o[15607] = i[15607];
  assign o[15606] = i[15606];
  assign o[15605] = i[15605];
  assign o[15604] = i[15604];
  assign o[15603] = i[15603];
  assign o[15602] = i[15602];
  assign o[15601] = i[15601];
  assign o[15600] = i[15600];
  assign o[15599] = i[15599];
  assign o[15598] = i[15598];
  assign o[15597] = i[15597];
  assign o[15596] = i[15596];
  assign o[15595] = i[15595];
  assign o[15594] = i[15594];
  assign o[15593] = i[15593];
  assign o[15592] = i[15592];
  assign o[15591] = i[15591];
  assign o[15590] = i[15590];
  assign o[15589] = i[15589];
  assign o[15588] = i[15588];
  assign o[15587] = i[15587];
  assign o[15586] = i[15586];
  assign o[15585] = i[15585];
  assign o[15584] = i[15584];
  assign o[15583] = i[15583];
  assign o[15582] = i[15582];
  assign o[15581] = i[15581];
  assign o[15580] = i[15580];
  assign o[15579] = i[15579];
  assign o[15578] = i[15578];
  assign o[15577] = i[15577];
  assign o[15576] = i[15576];
  assign o[15575] = i[15575];
  assign o[15574] = i[15574];
  assign o[15573] = i[15573];
  assign o[15572] = i[15572];
  assign o[15571] = i[15571];
  assign o[15570] = i[15570];
  assign o[15569] = i[15569];
  assign o[15568] = i[15568];
  assign o[15567] = i[15567];
  assign o[15566] = i[15566];
  assign o[15565] = i[15565];
  assign o[15564] = i[15564];
  assign o[15563] = i[15563];
  assign o[15562] = i[15562];
  assign o[15561] = i[15561];
  assign o[15560] = i[15560];
  assign o[15559] = i[15559];
  assign o[15558] = i[15558];
  assign o[15557] = i[15557];
  assign o[15556] = i[15556];
  assign o[15555] = i[15555];
  assign o[15554] = i[15554];
  assign o[15553] = i[15553];
  assign o[15552] = i[15552];
  assign o[15551] = i[15551];
  assign o[15550] = i[15550];
  assign o[15549] = i[15549];
  assign o[15548] = i[15548];
  assign o[15547] = i[15547];
  assign o[15546] = i[15546];
  assign o[15545] = i[15545];
  assign o[15544] = i[15544];
  assign o[15543] = i[15543];
  assign o[15542] = i[15542];
  assign o[15541] = i[15541];
  assign o[15540] = i[15540];
  assign o[15539] = i[15539];
  assign o[15538] = i[15538];
  assign o[15537] = i[15537];
  assign o[15536] = i[15536];
  assign o[15535] = i[15535];
  assign o[15534] = i[15534];
  assign o[15533] = i[15533];
  assign o[15532] = i[15532];
  assign o[15531] = i[15531];
  assign o[15530] = i[15530];
  assign o[15529] = i[15529];
  assign o[15528] = i[15528];
  assign o[15527] = i[15527];
  assign o[15526] = i[15526];
  assign o[15525] = i[15525];
  assign o[15524] = i[15524];
  assign o[15523] = i[15523];
  assign o[15522] = i[15522];
  assign o[15521] = i[15521];
  assign o[15520] = i[15520];
  assign o[15519] = i[15519];
  assign o[15518] = i[15518];
  assign o[15517] = i[15517];
  assign o[15516] = i[15516];
  assign o[15515] = i[15515];
  assign o[15514] = i[15514];
  assign o[15513] = i[15513];
  assign o[15512] = i[15512];
  assign o[15511] = i[15511];
  assign o[15510] = i[15510];
  assign o[15509] = i[15509];
  assign o[15508] = i[15508];
  assign o[15507] = i[15507];
  assign o[15506] = i[15506];
  assign o[15505] = i[15505];
  assign o[15504] = i[15504];
  assign o[15503] = i[15503];
  assign o[15502] = i[15502];
  assign o[15501] = i[15501];
  assign o[15500] = i[15500];
  assign o[15499] = i[15499];
  assign o[15498] = i[15498];
  assign o[15497] = i[15497];
  assign o[15496] = i[15496];
  assign o[15495] = i[15495];
  assign o[15494] = i[15494];
  assign o[15493] = i[15493];
  assign o[15492] = i[15492];
  assign o[15491] = i[15491];
  assign o[15490] = i[15490];
  assign o[15489] = i[15489];
  assign o[15488] = i[15488];
  assign o[15487] = i[15487];
  assign o[15486] = i[15486];
  assign o[15485] = i[15485];
  assign o[15484] = i[15484];
  assign o[15483] = i[15483];
  assign o[15482] = i[15482];
  assign o[15481] = i[15481];
  assign o[15480] = i[15480];
  assign o[15479] = i[15479];
  assign o[15478] = i[15478];
  assign o[15477] = i[15477];
  assign o[15476] = i[15476];
  assign o[15475] = i[15475];
  assign o[15474] = i[15474];
  assign o[15473] = i[15473];
  assign o[15472] = i[15472];
  assign o[15471] = i[15471];
  assign o[15470] = i[15470];
  assign o[15469] = i[15469];
  assign o[15468] = i[15468];
  assign o[15467] = i[15467];
  assign o[15466] = i[15466];
  assign o[15465] = i[15465];
  assign o[15464] = i[15464];
  assign o[15463] = i[15463];
  assign o[15462] = i[15462];
  assign o[15461] = i[15461];
  assign o[15460] = i[15460];
  assign o[15459] = i[15459];
  assign o[15458] = i[15458];
  assign o[15457] = i[15457];
  assign o[15456] = i[15456];
  assign o[15455] = i[15455];
  assign o[15454] = i[15454];
  assign o[15453] = i[15453];
  assign o[15452] = i[15452];
  assign o[15451] = i[15451];
  assign o[15450] = i[15450];
  assign o[15449] = i[15449];
  assign o[15448] = i[15448];
  assign o[15447] = i[15447];
  assign o[15446] = i[15446];
  assign o[15445] = i[15445];
  assign o[15444] = i[15444];
  assign o[15443] = i[15443];
  assign o[15442] = i[15442];
  assign o[15441] = i[15441];
  assign o[15440] = i[15440];
  assign o[15439] = i[15439];
  assign o[15438] = i[15438];
  assign o[15437] = i[15437];
  assign o[15436] = i[15436];
  assign o[15435] = i[15435];
  assign o[15434] = i[15434];
  assign o[15433] = i[15433];
  assign o[15432] = i[15432];
  assign o[15431] = i[15431];
  assign o[15430] = i[15430];
  assign o[15429] = i[15429];
  assign o[15428] = i[15428];
  assign o[15427] = i[15427];
  assign o[15426] = i[15426];
  assign o[15425] = i[15425];
  assign o[15424] = i[15424];
  assign o[15423] = i[15423];
  assign o[15422] = i[15422];
  assign o[15421] = i[15421];
  assign o[15420] = i[15420];
  assign o[15419] = i[15419];
  assign o[15418] = i[15418];
  assign o[15417] = i[15417];
  assign o[15416] = i[15416];
  assign o[15415] = i[15415];
  assign o[15414] = i[15414];
  assign o[15413] = i[15413];
  assign o[15412] = i[15412];
  assign o[15411] = i[15411];
  assign o[15410] = i[15410];
  assign o[15409] = i[15409];
  assign o[15408] = i[15408];
  assign o[15407] = i[15407];
  assign o[15406] = i[15406];
  assign o[15405] = i[15405];
  assign o[15404] = i[15404];
  assign o[15403] = i[15403];
  assign o[15402] = i[15402];
  assign o[15401] = i[15401];
  assign o[15400] = i[15400];
  assign o[15399] = i[15399];
  assign o[15398] = i[15398];
  assign o[15397] = i[15397];
  assign o[15396] = i[15396];
  assign o[15395] = i[15395];
  assign o[15394] = i[15394];
  assign o[15393] = i[15393];
  assign o[15392] = i[15392];
  assign o[15391] = i[15391];
  assign o[15390] = i[15390];
  assign o[15389] = i[15389];
  assign o[15388] = i[15388];
  assign o[15387] = i[15387];
  assign o[15386] = i[15386];
  assign o[15385] = i[15385];
  assign o[15384] = i[15384];
  assign o[15383] = i[15383];
  assign o[15382] = i[15382];
  assign o[15381] = i[15381];
  assign o[15380] = i[15380];
  assign o[15379] = i[15379];
  assign o[15378] = i[15378];
  assign o[15377] = i[15377];
  assign o[15376] = i[15376];
  assign o[15375] = i[15375];
  assign o[15374] = i[15374];
  assign o[15373] = i[15373];
  assign o[15372] = i[15372];
  assign o[15371] = i[15371];
  assign o[15370] = i[15370];
  assign o[15369] = i[15369];
  assign o[15368] = i[15368];
  assign o[15367] = i[15367];
  assign o[15366] = i[15366];
  assign o[15365] = i[15365];
  assign o[15364] = i[15364];
  assign o[15363] = i[15363];
  assign o[15362] = i[15362];
  assign o[15361] = i[15361];
  assign o[15360] = i[15360];
  assign o[15359] = i[15359];
  assign o[15358] = i[15358];
  assign o[15357] = i[15357];
  assign o[15356] = i[15356];
  assign o[15355] = i[15355];
  assign o[15354] = i[15354];
  assign o[15353] = i[15353];
  assign o[15352] = i[15352];
  assign o[15351] = i[15351];
  assign o[15350] = i[15350];
  assign o[15349] = i[15349];
  assign o[15348] = i[15348];
  assign o[15347] = i[15347];
  assign o[15346] = i[15346];
  assign o[15345] = i[15345];
  assign o[15344] = i[15344];
  assign o[15343] = i[15343];
  assign o[15342] = i[15342];
  assign o[15341] = i[15341];
  assign o[15340] = i[15340];
  assign o[15339] = i[15339];
  assign o[15338] = i[15338];
  assign o[15337] = i[15337];
  assign o[15336] = i[15336];
  assign o[15335] = i[15335];
  assign o[15334] = i[15334];
  assign o[15333] = i[15333];
  assign o[15332] = i[15332];
  assign o[15331] = i[15331];
  assign o[15330] = i[15330];
  assign o[15329] = i[15329];
  assign o[15328] = i[15328];
  assign o[15327] = i[15327];
  assign o[15326] = i[15326];
  assign o[15325] = i[15325];
  assign o[15324] = i[15324];
  assign o[15323] = i[15323];
  assign o[15322] = i[15322];
  assign o[15321] = i[15321];
  assign o[15320] = i[15320];
  assign o[15319] = i[15319];
  assign o[15318] = i[15318];
  assign o[15317] = i[15317];
  assign o[15316] = i[15316];
  assign o[15315] = i[15315];
  assign o[15314] = i[15314];
  assign o[15313] = i[15313];
  assign o[15312] = i[15312];
  assign o[15311] = i[15311];
  assign o[15310] = i[15310];
  assign o[15309] = i[15309];
  assign o[15308] = i[15308];
  assign o[15307] = i[15307];
  assign o[15306] = i[15306];
  assign o[15305] = i[15305];
  assign o[15304] = i[15304];
  assign o[15303] = i[15303];
  assign o[15302] = i[15302];
  assign o[15301] = i[15301];
  assign o[15300] = i[15300];
  assign o[15299] = i[15299];
  assign o[15298] = i[15298];
  assign o[15297] = i[15297];
  assign o[15296] = i[15296];
  assign o[15295] = i[15295];
  assign o[15294] = i[15294];
  assign o[15293] = i[15293];
  assign o[15292] = i[15292];
  assign o[15291] = i[15291];
  assign o[15290] = i[15290];
  assign o[15289] = i[15289];
  assign o[15288] = i[15288];
  assign o[15287] = i[15287];
  assign o[15286] = i[15286];
  assign o[15285] = i[15285];
  assign o[15284] = i[15284];
  assign o[15283] = i[15283];
  assign o[15282] = i[15282];
  assign o[15281] = i[15281];
  assign o[15280] = i[15280];
  assign o[15279] = i[15279];
  assign o[15278] = i[15278];
  assign o[15277] = i[15277];
  assign o[15276] = i[15276];
  assign o[15275] = i[15275];
  assign o[15274] = i[15274];
  assign o[15273] = i[15273];
  assign o[15272] = i[15272];
  assign o[15271] = i[15271];
  assign o[15270] = i[15270];
  assign o[15269] = i[15269];
  assign o[15268] = i[15268];
  assign o[15267] = i[15267];
  assign o[15266] = i[15266];
  assign o[15265] = i[15265];
  assign o[15264] = i[15264];
  assign o[15263] = i[15263];
  assign o[15262] = i[15262];
  assign o[15261] = i[15261];
  assign o[15260] = i[15260];
  assign o[15259] = i[15259];
  assign o[15258] = i[15258];
  assign o[15257] = i[15257];
  assign o[15256] = i[15256];
  assign o[15255] = i[15255];
  assign o[15254] = i[15254];
  assign o[15253] = i[15253];
  assign o[15252] = i[15252];
  assign o[15251] = i[15251];
  assign o[15250] = i[15250];
  assign o[15249] = i[15249];
  assign o[15248] = i[15248];
  assign o[15247] = i[15247];
  assign o[15246] = i[15246];
  assign o[15245] = i[15245];
  assign o[15244] = i[15244];
  assign o[15243] = i[15243];
  assign o[15242] = i[15242];
  assign o[15241] = i[15241];
  assign o[15240] = i[15240];
  assign o[15239] = i[15239];
  assign o[15238] = i[15238];
  assign o[15237] = i[15237];
  assign o[15236] = i[15236];
  assign o[15235] = i[15235];
  assign o[15234] = i[15234];
  assign o[15233] = i[15233];
  assign o[15232] = i[15232];
  assign o[15231] = i[15231];
  assign o[15230] = i[15230];
  assign o[15229] = i[15229];
  assign o[15228] = i[15228];
  assign o[15227] = i[15227];
  assign o[15226] = i[15226];
  assign o[15225] = i[15225];
  assign o[15224] = i[15224];
  assign o[15223] = i[15223];
  assign o[15222] = i[15222];
  assign o[15221] = i[15221];
  assign o[15220] = i[15220];
  assign o[15219] = i[15219];
  assign o[15218] = i[15218];
  assign o[15217] = i[15217];
  assign o[15216] = i[15216];
  assign o[15215] = i[15215];
  assign o[15214] = i[15214];
  assign o[15213] = i[15213];
  assign o[15212] = i[15212];
  assign o[15211] = i[15211];
  assign o[15210] = i[15210];
  assign o[15209] = i[15209];
  assign o[15208] = i[15208];
  assign o[15207] = i[15207];
  assign o[15206] = i[15206];
  assign o[15205] = i[15205];
  assign o[15204] = i[15204];
  assign o[15203] = i[15203];
  assign o[15202] = i[15202];
  assign o[15201] = i[15201];
  assign o[15200] = i[15200];
  assign o[15199] = i[15199];
  assign o[15198] = i[15198];
  assign o[15197] = i[15197];
  assign o[15196] = i[15196];
  assign o[15195] = i[15195];
  assign o[15194] = i[15194];
  assign o[15193] = i[15193];
  assign o[15192] = i[15192];
  assign o[15191] = i[15191];
  assign o[15190] = i[15190];
  assign o[15189] = i[15189];
  assign o[15188] = i[15188];
  assign o[15187] = i[15187];
  assign o[15186] = i[15186];
  assign o[15185] = i[15185];
  assign o[15184] = i[15184];
  assign o[15183] = i[15183];
  assign o[15182] = i[15182];
  assign o[15181] = i[15181];
  assign o[15180] = i[15180];
  assign o[15179] = i[15179];
  assign o[15178] = i[15178];
  assign o[15177] = i[15177];
  assign o[15176] = i[15176];
  assign o[15175] = i[15175];
  assign o[15174] = i[15174];
  assign o[15173] = i[15173];
  assign o[15172] = i[15172];
  assign o[15171] = i[15171];
  assign o[15170] = i[15170];
  assign o[15169] = i[15169];
  assign o[15168] = i[15168];
  assign o[15167] = i[15167];
  assign o[15166] = i[15166];
  assign o[15165] = i[15165];
  assign o[15164] = i[15164];
  assign o[15163] = i[15163];
  assign o[15162] = i[15162];
  assign o[15161] = i[15161];
  assign o[15160] = i[15160];
  assign o[15159] = i[15159];
  assign o[15158] = i[15158];
  assign o[15157] = i[15157];
  assign o[15156] = i[15156];
  assign o[15155] = i[15155];
  assign o[15154] = i[15154];
  assign o[15153] = i[15153];
  assign o[15152] = i[15152];
  assign o[15151] = i[15151];
  assign o[15150] = i[15150];
  assign o[15149] = i[15149];
  assign o[15148] = i[15148];
  assign o[15147] = i[15147];
  assign o[15146] = i[15146];
  assign o[15145] = i[15145];
  assign o[15144] = i[15144];
  assign o[15143] = i[15143];
  assign o[15142] = i[15142];
  assign o[15141] = i[15141];
  assign o[15140] = i[15140];
  assign o[15139] = i[15139];
  assign o[15138] = i[15138];
  assign o[15137] = i[15137];
  assign o[15136] = i[15136];
  assign o[15135] = i[15135];
  assign o[15134] = i[15134];
  assign o[15133] = i[15133];
  assign o[15132] = i[15132];
  assign o[15131] = i[15131];
  assign o[15130] = i[15130];
  assign o[15129] = i[15129];
  assign o[15128] = i[15128];
  assign o[15127] = i[15127];
  assign o[15126] = i[15126];
  assign o[15125] = i[15125];
  assign o[15124] = i[15124];
  assign o[15123] = i[15123];
  assign o[15122] = i[15122];
  assign o[15121] = i[15121];
  assign o[15120] = i[15120];
  assign o[15119] = i[15119];
  assign o[15118] = i[15118];
  assign o[15117] = i[15117];
  assign o[15116] = i[15116];
  assign o[15115] = i[15115];
  assign o[15114] = i[15114];
  assign o[15113] = i[15113];
  assign o[15112] = i[15112];
  assign o[15111] = i[15111];
  assign o[15110] = i[15110];
  assign o[15109] = i[15109];
  assign o[15108] = i[15108];
  assign o[15107] = i[15107];
  assign o[15106] = i[15106];
  assign o[15105] = i[15105];
  assign o[15104] = i[15104];
  assign o[15103] = i[15103];
  assign o[15102] = i[15102];
  assign o[15101] = i[15101];
  assign o[15100] = i[15100];
  assign o[15099] = i[15099];
  assign o[15098] = i[15098];
  assign o[15097] = i[15097];
  assign o[15096] = i[15096];
  assign o[15095] = i[15095];
  assign o[15094] = i[15094];
  assign o[15093] = i[15093];
  assign o[15092] = i[15092];
  assign o[15091] = i[15091];
  assign o[15090] = i[15090];
  assign o[15089] = i[15089];
  assign o[15088] = i[15088];
  assign o[15087] = i[15087];
  assign o[15086] = i[15086];
  assign o[15085] = i[15085];
  assign o[15084] = i[15084];
  assign o[15083] = i[15083];
  assign o[15082] = i[15082];
  assign o[15081] = i[15081];
  assign o[15080] = i[15080];
  assign o[15079] = i[15079];
  assign o[15078] = i[15078];
  assign o[15077] = i[15077];
  assign o[15076] = i[15076];
  assign o[15075] = i[15075];
  assign o[15074] = i[15074];
  assign o[15073] = i[15073];
  assign o[15072] = i[15072];
  assign o[15071] = i[15071];
  assign o[15070] = i[15070];
  assign o[15069] = i[15069];
  assign o[15068] = i[15068];
  assign o[15067] = i[15067];
  assign o[15066] = i[15066];
  assign o[15065] = i[15065];
  assign o[15064] = i[15064];
  assign o[15063] = i[15063];
  assign o[15062] = i[15062];
  assign o[15061] = i[15061];
  assign o[15060] = i[15060];
  assign o[15059] = i[15059];
  assign o[15058] = i[15058];
  assign o[15057] = i[15057];
  assign o[15056] = i[15056];
  assign o[15055] = i[15055];
  assign o[15054] = i[15054];
  assign o[15053] = i[15053];
  assign o[15052] = i[15052];
  assign o[15051] = i[15051];
  assign o[15050] = i[15050];
  assign o[15049] = i[15049];
  assign o[15048] = i[15048];
  assign o[15047] = i[15047];
  assign o[15046] = i[15046];
  assign o[15045] = i[15045];
  assign o[15044] = i[15044];
  assign o[15043] = i[15043];
  assign o[15042] = i[15042];
  assign o[15041] = i[15041];
  assign o[15040] = i[15040];
  assign o[15039] = i[15039];
  assign o[15038] = i[15038];
  assign o[15037] = i[15037];
  assign o[15036] = i[15036];
  assign o[15035] = i[15035];
  assign o[15034] = i[15034];
  assign o[15033] = i[15033];
  assign o[15032] = i[15032];
  assign o[15031] = i[15031];
  assign o[15030] = i[15030];
  assign o[15029] = i[15029];
  assign o[15028] = i[15028];
  assign o[15027] = i[15027];
  assign o[15026] = i[15026];
  assign o[15025] = i[15025];
  assign o[15024] = i[15024];
  assign o[15023] = i[15023];
  assign o[15022] = i[15022];
  assign o[15021] = i[15021];
  assign o[15020] = i[15020];
  assign o[15019] = i[15019];
  assign o[15018] = i[15018];
  assign o[15017] = i[15017];
  assign o[15016] = i[15016];
  assign o[15015] = i[15015];
  assign o[15014] = i[15014];
  assign o[15013] = i[15013];
  assign o[15012] = i[15012];
  assign o[15011] = i[15011];
  assign o[15010] = i[15010];
  assign o[15009] = i[15009];
  assign o[15008] = i[15008];
  assign o[15007] = i[15007];
  assign o[15006] = i[15006];
  assign o[15005] = i[15005];
  assign o[15004] = i[15004];
  assign o[15003] = i[15003];
  assign o[15002] = i[15002];
  assign o[15001] = i[15001];
  assign o[15000] = i[15000];
  assign o[14999] = i[14999];
  assign o[14998] = i[14998];
  assign o[14997] = i[14997];
  assign o[14996] = i[14996];
  assign o[14995] = i[14995];
  assign o[14994] = i[14994];
  assign o[14993] = i[14993];
  assign o[14992] = i[14992];
  assign o[14991] = i[14991];
  assign o[14990] = i[14990];
  assign o[14989] = i[14989];
  assign o[14988] = i[14988];
  assign o[14987] = i[14987];
  assign o[14986] = i[14986];
  assign o[14985] = i[14985];
  assign o[14984] = i[14984];
  assign o[14983] = i[14983];
  assign o[14982] = i[14982];
  assign o[14981] = i[14981];
  assign o[14980] = i[14980];
  assign o[14979] = i[14979];
  assign o[14978] = i[14978];
  assign o[14977] = i[14977];
  assign o[14976] = i[14976];
  assign o[14975] = i[14975];
  assign o[14974] = i[14974];
  assign o[14973] = i[14973];
  assign o[14972] = i[14972];
  assign o[14971] = i[14971];
  assign o[14970] = i[14970];
  assign o[14969] = i[14969];
  assign o[14968] = i[14968];
  assign o[14967] = i[14967];
  assign o[14966] = i[14966];
  assign o[14965] = i[14965];
  assign o[14964] = i[14964];
  assign o[14963] = i[14963];
  assign o[14962] = i[14962];
  assign o[14961] = i[14961];
  assign o[14960] = i[14960];
  assign o[14959] = i[14959];
  assign o[14958] = i[14958];
  assign o[14957] = i[14957];
  assign o[14956] = i[14956];
  assign o[14955] = i[14955];
  assign o[14954] = i[14954];
  assign o[14953] = i[14953];
  assign o[14952] = i[14952];
  assign o[14951] = i[14951];
  assign o[14950] = i[14950];
  assign o[14949] = i[14949];
  assign o[14948] = i[14948];
  assign o[14947] = i[14947];
  assign o[14946] = i[14946];
  assign o[14945] = i[14945];
  assign o[14944] = i[14944];
  assign o[14943] = i[14943];
  assign o[14942] = i[14942];
  assign o[14941] = i[14941];
  assign o[14940] = i[14940];
  assign o[14939] = i[14939];
  assign o[14938] = i[14938];
  assign o[14937] = i[14937];
  assign o[14936] = i[14936];
  assign o[14935] = i[14935];
  assign o[14934] = i[14934];
  assign o[14933] = i[14933];
  assign o[14932] = i[14932];
  assign o[14931] = i[14931];
  assign o[14930] = i[14930];
  assign o[14929] = i[14929];
  assign o[14928] = i[14928];
  assign o[14927] = i[14927];
  assign o[14926] = i[14926];
  assign o[14925] = i[14925];
  assign o[14924] = i[14924];
  assign o[14923] = i[14923];
  assign o[14922] = i[14922];
  assign o[14921] = i[14921];
  assign o[14920] = i[14920];
  assign o[14919] = i[14919];
  assign o[14918] = i[14918];
  assign o[14917] = i[14917];
  assign o[14916] = i[14916];
  assign o[14915] = i[14915];
  assign o[14914] = i[14914];
  assign o[14913] = i[14913];
  assign o[14912] = i[14912];
  assign o[14911] = i[14911];
  assign o[14910] = i[14910];
  assign o[14909] = i[14909];
  assign o[14908] = i[14908];
  assign o[14907] = i[14907];
  assign o[14906] = i[14906];
  assign o[14905] = i[14905];
  assign o[14904] = i[14904];
  assign o[14903] = i[14903];
  assign o[14902] = i[14902];
  assign o[14901] = i[14901];
  assign o[14900] = i[14900];
  assign o[14899] = i[14899];
  assign o[14898] = i[14898];
  assign o[14897] = i[14897];
  assign o[14896] = i[14896];
  assign o[14895] = i[14895];
  assign o[14894] = i[14894];
  assign o[14893] = i[14893];
  assign o[14892] = i[14892];
  assign o[14891] = i[14891];
  assign o[14890] = i[14890];
  assign o[14889] = i[14889];
  assign o[14888] = i[14888];
  assign o[14887] = i[14887];
  assign o[14886] = i[14886];
  assign o[14885] = i[14885];
  assign o[14884] = i[14884];
  assign o[14883] = i[14883];
  assign o[14882] = i[14882];
  assign o[14881] = i[14881];
  assign o[14880] = i[14880];
  assign o[14879] = i[14879];
  assign o[14878] = i[14878];
  assign o[14877] = i[14877];
  assign o[14876] = i[14876];
  assign o[14875] = i[14875];
  assign o[14874] = i[14874];
  assign o[14873] = i[14873];
  assign o[14872] = i[14872];
  assign o[14871] = i[14871];
  assign o[14870] = i[14870];
  assign o[14869] = i[14869];
  assign o[14868] = i[14868];
  assign o[14867] = i[14867];
  assign o[14866] = i[14866];
  assign o[14865] = i[14865];
  assign o[14864] = i[14864];
  assign o[14863] = i[14863];
  assign o[14862] = i[14862];
  assign o[14861] = i[14861];
  assign o[14860] = i[14860];
  assign o[14859] = i[14859];
  assign o[14858] = i[14858];
  assign o[14857] = i[14857];
  assign o[14856] = i[14856];
  assign o[14855] = i[14855];
  assign o[14854] = i[14854];
  assign o[14853] = i[14853];
  assign o[14852] = i[14852];
  assign o[14851] = i[14851];
  assign o[14850] = i[14850];
  assign o[14849] = i[14849];
  assign o[14848] = i[14848];
  assign o[14847] = i[14847];
  assign o[14846] = i[14846];
  assign o[14845] = i[14845];
  assign o[14844] = i[14844];
  assign o[14843] = i[14843];
  assign o[14842] = i[14842];
  assign o[14841] = i[14841];
  assign o[14840] = i[14840];
  assign o[14839] = i[14839];
  assign o[14838] = i[14838];
  assign o[14837] = i[14837];
  assign o[14836] = i[14836];
  assign o[14835] = i[14835];
  assign o[14834] = i[14834];
  assign o[14833] = i[14833];
  assign o[14832] = i[14832];
  assign o[14831] = i[14831];
  assign o[14830] = i[14830];
  assign o[14829] = i[14829];
  assign o[14828] = i[14828];
  assign o[14827] = i[14827];
  assign o[14826] = i[14826];
  assign o[14825] = i[14825];
  assign o[14824] = i[14824];
  assign o[14823] = i[14823];
  assign o[14822] = i[14822];
  assign o[14821] = i[14821];
  assign o[14820] = i[14820];
  assign o[14819] = i[14819];
  assign o[14818] = i[14818];
  assign o[14817] = i[14817];
  assign o[14816] = i[14816];
  assign o[14815] = i[14815];
  assign o[14814] = i[14814];
  assign o[14813] = i[14813];
  assign o[14812] = i[14812];
  assign o[14811] = i[14811];
  assign o[14810] = i[14810];
  assign o[14809] = i[14809];
  assign o[14808] = i[14808];
  assign o[14807] = i[14807];
  assign o[14806] = i[14806];
  assign o[14805] = i[14805];
  assign o[14804] = i[14804];
  assign o[14803] = i[14803];
  assign o[14802] = i[14802];
  assign o[14801] = i[14801];
  assign o[14800] = i[14800];
  assign o[14799] = i[14799];
  assign o[14798] = i[14798];
  assign o[14797] = i[14797];
  assign o[14796] = i[14796];
  assign o[14795] = i[14795];
  assign o[14794] = i[14794];
  assign o[14793] = i[14793];
  assign o[14792] = i[14792];
  assign o[14791] = i[14791];
  assign o[14790] = i[14790];
  assign o[14789] = i[14789];
  assign o[14788] = i[14788];
  assign o[14787] = i[14787];
  assign o[14786] = i[14786];
  assign o[14785] = i[14785];
  assign o[14784] = i[14784];
  assign o[14783] = i[14783];
  assign o[14782] = i[14782];
  assign o[14781] = i[14781];
  assign o[14780] = i[14780];
  assign o[14779] = i[14779];
  assign o[14778] = i[14778];
  assign o[14777] = i[14777];
  assign o[14776] = i[14776];
  assign o[14775] = i[14775];
  assign o[14774] = i[14774];
  assign o[14773] = i[14773];
  assign o[14772] = i[14772];
  assign o[14771] = i[14771];
  assign o[14770] = i[14770];
  assign o[14769] = i[14769];
  assign o[14768] = i[14768];
  assign o[14767] = i[14767];
  assign o[14766] = i[14766];
  assign o[14765] = i[14765];
  assign o[14764] = i[14764];
  assign o[14763] = i[14763];
  assign o[14762] = i[14762];
  assign o[14761] = i[14761];
  assign o[14760] = i[14760];
  assign o[14759] = i[14759];
  assign o[14758] = i[14758];
  assign o[14757] = i[14757];
  assign o[14756] = i[14756];
  assign o[14755] = i[14755];
  assign o[14754] = i[14754];
  assign o[14753] = i[14753];
  assign o[14752] = i[14752];
  assign o[14751] = i[14751];
  assign o[14750] = i[14750];
  assign o[14749] = i[14749];
  assign o[14748] = i[14748];
  assign o[14747] = i[14747];
  assign o[14746] = i[14746];
  assign o[14745] = i[14745];
  assign o[14744] = i[14744];
  assign o[14743] = i[14743];
  assign o[14742] = i[14742];
  assign o[14741] = i[14741];
  assign o[14740] = i[14740];
  assign o[14739] = i[14739];
  assign o[14738] = i[14738];
  assign o[14737] = i[14737];
  assign o[14736] = i[14736];
  assign o[14735] = i[14735];
  assign o[14734] = i[14734];
  assign o[14733] = i[14733];
  assign o[14732] = i[14732];
  assign o[14731] = i[14731];
  assign o[14730] = i[14730];
  assign o[14729] = i[14729];
  assign o[14728] = i[14728];
  assign o[14727] = i[14727];
  assign o[14726] = i[14726];
  assign o[14725] = i[14725];
  assign o[14724] = i[14724];
  assign o[14723] = i[14723];
  assign o[14722] = i[14722];
  assign o[14721] = i[14721];
  assign o[14720] = i[14720];
  assign o[14719] = i[14719];
  assign o[14718] = i[14718];
  assign o[14717] = i[14717];
  assign o[14716] = i[14716];
  assign o[14715] = i[14715];
  assign o[14714] = i[14714];
  assign o[14713] = i[14713];
  assign o[14712] = i[14712];
  assign o[14711] = i[14711];
  assign o[14710] = i[14710];
  assign o[14709] = i[14709];
  assign o[14708] = i[14708];
  assign o[14707] = i[14707];
  assign o[14706] = i[14706];
  assign o[14705] = i[14705];
  assign o[14704] = i[14704];
  assign o[14703] = i[14703];
  assign o[14702] = i[14702];
  assign o[14701] = i[14701];
  assign o[14700] = i[14700];
  assign o[14699] = i[14699];
  assign o[14698] = i[14698];
  assign o[14697] = i[14697];
  assign o[14696] = i[14696];
  assign o[14695] = i[14695];
  assign o[14694] = i[14694];
  assign o[14693] = i[14693];
  assign o[14692] = i[14692];
  assign o[14691] = i[14691];
  assign o[14690] = i[14690];
  assign o[14689] = i[14689];
  assign o[14688] = i[14688];
  assign o[14687] = i[14687];
  assign o[14686] = i[14686];
  assign o[14685] = i[14685];
  assign o[14684] = i[14684];
  assign o[14683] = i[14683];
  assign o[14682] = i[14682];
  assign o[14681] = i[14681];
  assign o[14680] = i[14680];
  assign o[14679] = i[14679];
  assign o[14678] = i[14678];
  assign o[14677] = i[14677];
  assign o[14676] = i[14676];
  assign o[14675] = i[14675];
  assign o[14674] = i[14674];
  assign o[14673] = i[14673];
  assign o[14672] = i[14672];
  assign o[14671] = i[14671];
  assign o[14670] = i[14670];
  assign o[14669] = i[14669];
  assign o[14668] = i[14668];
  assign o[14667] = i[14667];
  assign o[14666] = i[14666];
  assign o[14665] = i[14665];
  assign o[14664] = i[14664];
  assign o[14663] = i[14663];
  assign o[14662] = i[14662];
  assign o[14661] = i[14661];
  assign o[14660] = i[14660];
  assign o[14659] = i[14659];
  assign o[14658] = i[14658];
  assign o[14657] = i[14657];
  assign o[14656] = i[14656];
  assign o[14655] = i[14655];
  assign o[14654] = i[14654];
  assign o[14653] = i[14653];
  assign o[14652] = i[14652];
  assign o[14651] = i[14651];
  assign o[14650] = i[14650];
  assign o[14649] = i[14649];
  assign o[14648] = i[14648];
  assign o[14647] = i[14647];
  assign o[14646] = i[14646];
  assign o[14645] = i[14645];
  assign o[14644] = i[14644];
  assign o[14643] = i[14643];
  assign o[14642] = i[14642];
  assign o[14641] = i[14641];
  assign o[14640] = i[14640];
  assign o[14639] = i[14639];
  assign o[14638] = i[14638];
  assign o[14637] = i[14637];
  assign o[14636] = i[14636];
  assign o[14635] = i[14635];
  assign o[14634] = i[14634];
  assign o[14633] = i[14633];
  assign o[14632] = i[14632];
  assign o[14631] = i[14631];
  assign o[14630] = i[14630];
  assign o[14629] = i[14629];
  assign o[14628] = i[14628];
  assign o[14627] = i[14627];
  assign o[14626] = i[14626];
  assign o[14625] = i[14625];
  assign o[14624] = i[14624];
  assign o[14623] = i[14623];
  assign o[14622] = i[14622];
  assign o[14621] = i[14621];
  assign o[14620] = i[14620];
  assign o[14619] = i[14619];
  assign o[14618] = i[14618];
  assign o[14617] = i[14617];
  assign o[14616] = i[14616];
  assign o[14615] = i[14615];
  assign o[14614] = i[14614];
  assign o[14613] = i[14613];
  assign o[14612] = i[14612];
  assign o[14611] = i[14611];
  assign o[14610] = i[14610];
  assign o[14609] = i[14609];
  assign o[14608] = i[14608];
  assign o[14607] = i[14607];
  assign o[14606] = i[14606];
  assign o[14605] = i[14605];
  assign o[14604] = i[14604];
  assign o[14603] = i[14603];
  assign o[14602] = i[14602];
  assign o[14601] = i[14601];
  assign o[14600] = i[14600];
  assign o[14599] = i[14599];
  assign o[14598] = i[14598];
  assign o[14597] = i[14597];
  assign o[14596] = i[14596];
  assign o[14595] = i[14595];
  assign o[14594] = i[14594];
  assign o[14593] = i[14593];
  assign o[14592] = i[14592];
  assign o[14591] = i[14591];
  assign o[14590] = i[14590];
  assign o[14589] = i[14589];
  assign o[14588] = i[14588];
  assign o[14587] = i[14587];
  assign o[14586] = i[14586];
  assign o[14585] = i[14585];
  assign o[14584] = i[14584];
  assign o[14583] = i[14583];
  assign o[14582] = i[14582];
  assign o[14581] = i[14581];
  assign o[14580] = i[14580];
  assign o[14579] = i[14579];
  assign o[14578] = i[14578];
  assign o[14577] = i[14577];
  assign o[14576] = i[14576];
  assign o[14575] = i[14575];
  assign o[14574] = i[14574];
  assign o[14573] = i[14573];
  assign o[14572] = i[14572];
  assign o[14571] = i[14571];
  assign o[14570] = i[14570];
  assign o[14569] = i[14569];
  assign o[14568] = i[14568];
  assign o[14567] = i[14567];
  assign o[14566] = i[14566];
  assign o[14565] = i[14565];
  assign o[14564] = i[14564];
  assign o[14563] = i[14563];
  assign o[14562] = i[14562];
  assign o[14561] = i[14561];
  assign o[14560] = i[14560];
  assign o[14559] = i[14559];
  assign o[14558] = i[14558];
  assign o[14557] = i[14557];
  assign o[14556] = i[14556];
  assign o[14555] = i[14555];
  assign o[14554] = i[14554];
  assign o[14553] = i[14553];
  assign o[14552] = i[14552];
  assign o[14551] = i[14551];
  assign o[14550] = i[14550];
  assign o[14549] = i[14549];
  assign o[14548] = i[14548];
  assign o[14547] = i[14547];
  assign o[14546] = i[14546];
  assign o[14545] = i[14545];
  assign o[14544] = i[14544];
  assign o[14543] = i[14543];
  assign o[14542] = i[14542];
  assign o[14541] = i[14541];
  assign o[14540] = i[14540];
  assign o[14539] = i[14539];
  assign o[14538] = i[14538];
  assign o[14537] = i[14537];
  assign o[14536] = i[14536];
  assign o[14535] = i[14535];
  assign o[14534] = i[14534];
  assign o[14533] = i[14533];
  assign o[14532] = i[14532];
  assign o[14531] = i[14531];
  assign o[14530] = i[14530];
  assign o[14529] = i[14529];
  assign o[14528] = i[14528];
  assign o[14527] = i[14527];
  assign o[14526] = i[14526];
  assign o[14525] = i[14525];
  assign o[14524] = i[14524];
  assign o[14523] = i[14523];
  assign o[14522] = i[14522];
  assign o[14521] = i[14521];
  assign o[14520] = i[14520];
  assign o[14519] = i[14519];
  assign o[14518] = i[14518];
  assign o[14517] = i[14517];
  assign o[14516] = i[14516];
  assign o[14515] = i[14515];
  assign o[14514] = i[14514];
  assign o[14513] = i[14513];
  assign o[14512] = i[14512];
  assign o[14511] = i[14511];
  assign o[14510] = i[14510];
  assign o[14509] = i[14509];
  assign o[14508] = i[14508];
  assign o[14507] = i[14507];
  assign o[14506] = i[14506];
  assign o[14505] = i[14505];
  assign o[14504] = i[14504];
  assign o[14503] = i[14503];
  assign o[14502] = i[14502];
  assign o[14501] = i[14501];
  assign o[14500] = i[14500];
  assign o[14499] = i[14499];
  assign o[14498] = i[14498];
  assign o[14497] = i[14497];
  assign o[14496] = i[14496];
  assign o[14495] = i[14495];
  assign o[14494] = i[14494];
  assign o[14493] = i[14493];
  assign o[14492] = i[14492];
  assign o[14491] = i[14491];
  assign o[14490] = i[14490];
  assign o[14489] = i[14489];
  assign o[14488] = i[14488];
  assign o[14487] = i[14487];
  assign o[14486] = i[14486];
  assign o[14485] = i[14485];
  assign o[14484] = i[14484];
  assign o[14483] = i[14483];
  assign o[14482] = i[14482];
  assign o[14481] = i[14481];
  assign o[14480] = i[14480];
  assign o[14479] = i[14479];
  assign o[14478] = i[14478];
  assign o[14477] = i[14477];
  assign o[14476] = i[14476];
  assign o[14475] = i[14475];
  assign o[14474] = i[14474];
  assign o[14473] = i[14473];
  assign o[14472] = i[14472];
  assign o[14471] = i[14471];
  assign o[14470] = i[14470];
  assign o[14469] = i[14469];
  assign o[14468] = i[14468];
  assign o[14467] = i[14467];
  assign o[14466] = i[14466];
  assign o[14465] = i[14465];
  assign o[14464] = i[14464];
  assign o[14463] = i[14463];
  assign o[14462] = i[14462];
  assign o[14461] = i[14461];
  assign o[14460] = i[14460];
  assign o[14459] = i[14459];
  assign o[14458] = i[14458];
  assign o[14457] = i[14457];
  assign o[14456] = i[14456];
  assign o[14455] = i[14455];
  assign o[14454] = i[14454];
  assign o[14453] = i[14453];
  assign o[14452] = i[14452];
  assign o[14451] = i[14451];
  assign o[14450] = i[14450];
  assign o[14449] = i[14449];
  assign o[14448] = i[14448];
  assign o[14447] = i[14447];
  assign o[14446] = i[14446];
  assign o[14445] = i[14445];
  assign o[14444] = i[14444];
  assign o[14443] = i[14443];
  assign o[14442] = i[14442];
  assign o[14441] = i[14441];
  assign o[14440] = i[14440];
  assign o[14439] = i[14439];
  assign o[14438] = i[14438];
  assign o[14437] = i[14437];
  assign o[14436] = i[14436];
  assign o[14435] = i[14435];
  assign o[14434] = i[14434];
  assign o[14433] = i[14433];
  assign o[14432] = i[14432];
  assign o[14431] = i[14431];
  assign o[14430] = i[14430];
  assign o[14429] = i[14429];
  assign o[14428] = i[14428];
  assign o[14427] = i[14427];
  assign o[14426] = i[14426];
  assign o[14425] = i[14425];
  assign o[14424] = i[14424];
  assign o[14423] = i[14423];
  assign o[14422] = i[14422];
  assign o[14421] = i[14421];
  assign o[14420] = i[14420];
  assign o[14419] = i[14419];
  assign o[14418] = i[14418];
  assign o[14417] = i[14417];
  assign o[14416] = i[14416];
  assign o[14415] = i[14415];
  assign o[14414] = i[14414];
  assign o[14413] = i[14413];
  assign o[14412] = i[14412];
  assign o[14411] = i[14411];
  assign o[14410] = i[14410];
  assign o[14409] = i[14409];
  assign o[14408] = i[14408];
  assign o[14407] = i[14407];
  assign o[14406] = i[14406];
  assign o[14405] = i[14405];
  assign o[14404] = i[14404];
  assign o[14403] = i[14403];
  assign o[14402] = i[14402];
  assign o[14401] = i[14401];
  assign o[14400] = i[14400];
  assign o[14399] = i[14399];
  assign o[14398] = i[14398];
  assign o[14397] = i[14397];
  assign o[14396] = i[14396];
  assign o[14395] = i[14395];
  assign o[14394] = i[14394];
  assign o[14393] = i[14393];
  assign o[14392] = i[14392];
  assign o[14391] = i[14391];
  assign o[14390] = i[14390];
  assign o[14389] = i[14389];
  assign o[14388] = i[14388];
  assign o[14387] = i[14387];
  assign o[14386] = i[14386];
  assign o[14385] = i[14385];
  assign o[14384] = i[14384];
  assign o[14383] = i[14383];
  assign o[14382] = i[14382];
  assign o[14381] = i[14381];
  assign o[14380] = i[14380];
  assign o[14379] = i[14379];
  assign o[14378] = i[14378];
  assign o[14377] = i[14377];
  assign o[14376] = i[14376];
  assign o[14375] = i[14375];
  assign o[14374] = i[14374];
  assign o[14373] = i[14373];
  assign o[14372] = i[14372];
  assign o[14371] = i[14371];
  assign o[14370] = i[14370];
  assign o[14369] = i[14369];
  assign o[14368] = i[14368];
  assign o[14367] = i[14367];
  assign o[14366] = i[14366];
  assign o[14365] = i[14365];
  assign o[14364] = i[14364];
  assign o[14363] = i[14363];
  assign o[14362] = i[14362];
  assign o[14361] = i[14361];
  assign o[14360] = i[14360];
  assign o[14359] = i[14359];
  assign o[14358] = i[14358];
  assign o[14357] = i[14357];
  assign o[14356] = i[14356];
  assign o[14355] = i[14355];
  assign o[14354] = i[14354];
  assign o[14353] = i[14353];
  assign o[14352] = i[14352];
  assign o[14351] = i[14351];
  assign o[14350] = i[14350];
  assign o[14349] = i[14349];
  assign o[14348] = i[14348];
  assign o[14347] = i[14347];
  assign o[14346] = i[14346];
  assign o[14345] = i[14345];
  assign o[14344] = i[14344];
  assign o[14343] = i[14343];
  assign o[14342] = i[14342];
  assign o[14341] = i[14341];
  assign o[14340] = i[14340];
  assign o[14339] = i[14339];
  assign o[14338] = i[14338];
  assign o[14337] = i[14337];
  assign o[14336] = i[14336];
  assign o[14335] = i[14335];
  assign o[14334] = i[14334];
  assign o[14333] = i[14333];
  assign o[14332] = i[14332];
  assign o[14331] = i[14331];
  assign o[14330] = i[14330];
  assign o[14329] = i[14329];
  assign o[14328] = i[14328];
  assign o[14327] = i[14327];
  assign o[14326] = i[14326];
  assign o[14325] = i[14325];
  assign o[14324] = i[14324];
  assign o[14323] = i[14323];
  assign o[14322] = i[14322];
  assign o[14321] = i[14321];
  assign o[14320] = i[14320];
  assign o[14319] = i[14319];
  assign o[14318] = i[14318];
  assign o[14317] = i[14317];
  assign o[14316] = i[14316];
  assign o[14315] = i[14315];
  assign o[14314] = i[14314];
  assign o[14313] = i[14313];
  assign o[14312] = i[14312];
  assign o[14311] = i[14311];
  assign o[14310] = i[14310];
  assign o[14309] = i[14309];
  assign o[14308] = i[14308];
  assign o[14307] = i[14307];
  assign o[14306] = i[14306];
  assign o[14305] = i[14305];
  assign o[14304] = i[14304];
  assign o[14303] = i[14303];
  assign o[14302] = i[14302];
  assign o[14301] = i[14301];
  assign o[14300] = i[14300];
  assign o[14299] = i[14299];
  assign o[14298] = i[14298];
  assign o[14297] = i[14297];
  assign o[14296] = i[14296];
  assign o[14295] = i[14295];
  assign o[14294] = i[14294];
  assign o[14293] = i[14293];
  assign o[14292] = i[14292];
  assign o[14291] = i[14291];
  assign o[14290] = i[14290];
  assign o[14289] = i[14289];
  assign o[14288] = i[14288];
  assign o[14287] = i[14287];
  assign o[14286] = i[14286];
  assign o[14285] = i[14285];
  assign o[14284] = i[14284];
  assign o[14283] = i[14283];
  assign o[14282] = i[14282];
  assign o[14281] = i[14281];
  assign o[14280] = i[14280];
  assign o[14279] = i[14279];
  assign o[14278] = i[14278];
  assign o[14277] = i[14277];
  assign o[14276] = i[14276];
  assign o[14275] = i[14275];
  assign o[14274] = i[14274];
  assign o[14273] = i[14273];
  assign o[14272] = i[14272];
  assign o[14271] = i[14271];
  assign o[14270] = i[14270];
  assign o[14269] = i[14269];
  assign o[14268] = i[14268];
  assign o[14267] = i[14267];
  assign o[14266] = i[14266];
  assign o[14265] = i[14265];
  assign o[14264] = i[14264];
  assign o[14263] = i[14263];
  assign o[14262] = i[14262];
  assign o[14261] = i[14261];
  assign o[14260] = i[14260];
  assign o[14259] = i[14259];
  assign o[14258] = i[14258];
  assign o[14257] = i[14257];
  assign o[14256] = i[14256];
  assign o[14255] = i[14255];
  assign o[14254] = i[14254];
  assign o[14253] = i[14253];
  assign o[14252] = i[14252];
  assign o[14251] = i[14251];
  assign o[14250] = i[14250];
  assign o[14249] = i[14249];
  assign o[14248] = i[14248];
  assign o[14247] = i[14247];
  assign o[14246] = i[14246];
  assign o[14245] = i[14245];
  assign o[14244] = i[14244];
  assign o[14243] = i[14243];
  assign o[14242] = i[14242];
  assign o[14241] = i[14241];
  assign o[14240] = i[14240];
  assign o[14239] = i[14239];
  assign o[14238] = i[14238];
  assign o[14237] = i[14237];
  assign o[14236] = i[14236];
  assign o[14235] = i[14235];
  assign o[14234] = i[14234];
  assign o[14233] = i[14233];
  assign o[14232] = i[14232];
  assign o[14231] = i[14231];
  assign o[14230] = i[14230];
  assign o[14229] = i[14229];
  assign o[14228] = i[14228];
  assign o[14227] = i[14227];
  assign o[14226] = i[14226];
  assign o[14225] = i[14225];
  assign o[14224] = i[14224];
  assign o[14223] = i[14223];
  assign o[14222] = i[14222];
  assign o[14221] = i[14221];
  assign o[14220] = i[14220];
  assign o[14219] = i[14219];
  assign o[14218] = i[14218];
  assign o[14217] = i[14217];
  assign o[14216] = i[14216];
  assign o[14215] = i[14215];
  assign o[14214] = i[14214];
  assign o[14213] = i[14213];
  assign o[14212] = i[14212];
  assign o[14211] = i[14211];
  assign o[14210] = i[14210];
  assign o[14209] = i[14209];
  assign o[14208] = i[14208];
  assign o[14207] = i[14207];
  assign o[14206] = i[14206];
  assign o[14205] = i[14205];
  assign o[14204] = i[14204];
  assign o[14203] = i[14203];
  assign o[14202] = i[14202];
  assign o[14201] = i[14201];
  assign o[14200] = i[14200];
  assign o[14199] = i[14199];
  assign o[14198] = i[14198];
  assign o[14197] = i[14197];
  assign o[14196] = i[14196];
  assign o[14195] = i[14195];
  assign o[14194] = i[14194];
  assign o[14193] = i[14193];
  assign o[14192] = i[14192];
  assign o[14191] = i[14191];
  assign o[14190] = i[14190];
  assign o[14189] = i[14189];
  assign o[14188] = i[14188];
  assign o[14187] = i[14187];
  assign o[14186] = i[14186];
  assign o[14185] = i[14185];
  assign o[14184] = i[14184];
  assign o[14183] = i[14183];
  assign o[14182] = i[14182];
  assign o[14181] = i[14181];
  assign o[14180] = i[14180];
  assign o[14179] = i[14179];
  assign o[14178] = i[14178];
  assign o[14177] = i[14177];
  assign o[14176] = i[14176];
  assign o[14175] = i[14175];
  assign o[14174] = i[14174];
  assign o[14173] = i[14173];
  assign o[14172] = i[14172];
  assign o[14171] = i[14171];
  assign o[14170] = i[14170];
  assign o[14169] = i[14169];
  assign o[14168] = i[14168];
  assign o[14167] = i[14167];
  assign o[14166] = i[14166];
  assign o[14165] = i[14165];
  assign o[14164] = i[14164];
  assign o[14163] = i[14163];
  assign o[14162] = i[14162];
  assign o[14161] = i[14161];
  assign o[14160] = i[14160];
  assign o[14159] = i[14159];
  assign o[14158] = i[14158];
  assign o[14157] = i[14157];
  assign o[14156] = i[14156];
  assign o[14155] = i[14155];
  assign o[14154] = i[14154];
  assign o[14153] = i[14153];
  assign o[14152] = i[14152];
  assign o[14151] = i[14151];
  assign o[14150] = i[14150];
  assign o[14149] = i[14149];
  assign o[14148] = i[14148];
  assign o[14147] = i[14147];
  assign o[14146] = i[14146];
  assign o[14145] = i[14145];
  assign o[14144] = i[14144];
  assign o[14143] = i[14143];
  assign o[14142] = i[14142];
  assign o[14141] = i[14141];
  assign o[14140] = i[14140];
  assign o[14139] = i[14139];
  assign o[14138] = i[14138];
  assign o[14137] = i[14137];
  assign o[14136] = i[14136];
  assign o[14135] = i[14135];
  assign o[14134] = i[14134];
  assign o[14133] = i[14133];
  assign o[14132] = i[14132];
  assign o[14131] = i[14131];
  assign o[14130] = i[14130];
  assign o[14129] = i[14129];
  assign o[14128] = i[14128];
  assign o[14127] = i[14127];
  assign o[14126] = i[14126];
  assign o[14125] = i[14125];
  assign o[14124] = i[14124];
  assign o[14123] = i[14123];
  assign o[14122] = i[14122];
  assign o[14121] = i[14121];
  assign o[14120] = i[14120];
  assign o[14119] = i[14119];
  assign o[14118] = i[14118];
  assign o[14117] = i[14117];
  assign o[14116] = i[14116];
  assign o[14115] = i[14115];
  assign o[14114] = i[14114];
  assign o[14113] = i[14113];
  assign o[14112] = i[14112];
  assign o[14111] = i[14111];
  assign o[14110] = i[14110];
  assign o[14109] = i[14109];
  assign o[14108] = i[14108];
  assign o[14107] = i[14107];
  assign o[14106] = i[14106];
  assign o[14105] = i[14105];
  assign o[14104] = i[14104];
  assign o[14103] = i[14103];
  assign o[14102] = i[14102];
  assign o[14101] = i[14101];
  assign o[14100] = i[14100];
  assign o[14099] = i[14099];
  assign o[14098] = i[14098];
  assign o[14097] = i[14097];
  assign o[14096] = i[14096];
  assign o[14095] = i[14095];
  assign o[14094] = i[14094];
  assign o[14093] = i[14093];
  assign o[14092] = i[14092];
  assign o[14091] = i[14091];
  assign o[14090] = i[14090];
  assign o[14089] = i[14089];
  assign o[14088] = i[14088];
  assign o[14087] = i[14087];
  assign o[14086] = i[14086];
  assign o[14085] = i[14085];
  assign o[14084] = i[14084];
  assign o[14083] = i[14083];
  assign o[14082] = i[14082];
  assign o[14081] = i[14081];
  assign o[14080] = i[14080];
  assign o[14079] = i[14079];
  assign o[14078] = i[14078];
  assign o[14077] = i[14077];
  assign o[14076] = i[14076];
  assign o[14075] = i[14075];
  assign o[14074] = i[14074];
  assign o[14073] = i[14073];
  assign o[14072] = i[14072];
  assign o[14071] = i[14071];
  assign o[14070] = i[14070];
  assign o[14069] = i[14069];
  assign o[14068] = i[14068];
  assign o[14067] = i[14067];
  assign o[14066] = i[14066];
  assign o[14065] = i[14065];
  assign o[14064] = i[14064];
  assign o[14063] = i[14063];
  assign o[14062] = i[14062];
  assign o[14061] = i[14061];
  assign o[14060] = i[14060];
  assign o[14059] = i[14059];
  assign o[14058] = i[14058];
  assign o[14057] = i[14057];
  assign o[14056] = i[14056];
  assign o[14055] = i[14055];
  assign o[14054] = i[14054];
  assign o[14053] = i[14053];
  assign o[14052] = i[14052];
  assign o[14051] = i[14051];
  assign o[14050] = i[14050];
  assign o[14049] = i[14049];
  assign o[14048] = i[14048];
  assign o[14047] = i[14047];
  assign o[14046] = i[14046];
  assign o[14045] = i[14045];
  assign o[14044] = i[14044];
  assign o[14043] = i[14043];
  assign o[14042] = i[14042];
  assign o[14041] = i[14041];
  assign o[14040] = i[14040];
  assign o[14039] = i[14039];
  assign o[14038] = i[14038];
  assign o[14037] = i[14037];
  assign o[14036] = i[14036];
  assign o[14035] = i[14035];
  assign o[14034] = i[14034];
  assign o[14033] = i[14033];
  assign o[14032] = i[14032];
  assign o[14031] = i[14031];
  assign o[14030] = i[14030];
  assign o[14029] = i[14029];
  assign o[14028] = i[14028];
  assign o[14027] = i[14027];
  assign o[14026] = i[14026];
  assign o[14025] = i[14025];
  assign o[14024] = i[14024];
  assign o[14023] = i[14023];
  assign o[14022] = i[14022];
  assign o[14021] = i[14021];
  assign o[14020] = i[14020];
  assign o[14019] = i[14019];
  assign o[14018] = i[14018];
  assign o[14017] = i[14017];
  assign o[14016] = i[14016];
  assign o[14015] = i[14015];
  assign o[14014] = i[14014];
  assign o[14013] = i[14013];
  assign o[14012] = i[14012];
  assign o[14011] = i[14011];
  assign o[14010] = i[14010];
  assign o[14009] = i[14009];
  assign o[14008] = i[14008];
  assign o[14007] = i[14007];
  assign o[14006] = i[14006];
  assign o[14005] = i[14005];
  assign o[14004] = i[14004];
  assign o[14003] = i[14003];
  assign o[14002] = i[14002];
  assign o[14001] = i[14001];
  assign o[14000] = i[14000];
  assign o[13999] = i[13999];
  assign o[13998] = i[13998];
  assign o[13997] = i[13997];
  assign o[13996] = i[13996];
  assign o[13995] = i[13995];
  assign o[13994] = i[13994];
  assign o[13993] = i[13993];
  assign o[13992] = i[13992];
  assign o[13991] = i[13991];
  assign o[13990] = i[13990];
  assign o[13989] = i[13989];
  assign o[13988] = i[13988];
  assign o[13987] = i[13987];
  assign o[13986] = i[13986];
  assign o[13985] = i[13985];
  assign o[13984] = i[13984];
  assign o[13983] = i[13983];
  assign o[13982] = i[13982];
  assign o[13981] = i[13981];
  assign o[13980] = i[13980];
  assign o[13979] = i[13979];
  assign o[13978] = i[13978];
  assign o[13977] = i[13977];
  assign o[13976] = i[13976];
  assign o[13975] = i[13975];
  assign o[13974] = i[13974];
  assign o[13973] = i[13973];
  assign o[13972] = i[13972];
  assign o[13971] = i[13971];
  assign o[13970] = i[13970];
  assign o[13969] = i[13969];
  assign o[13968] = i[13968];
  assign o[13967] = i[13967];
  assign o[13966] = i[13966];
  assign o[13965] = i[13965];
  assign o[13964] = i[13964];
  assign o[13963] = i[13963];
  assign o[13962] = i[13962];
  assign o[13961] = i[13961];
  assign o[13960] = i[13960];
  assign o[13959] = i[13959];
  assign o[13958] = i[13958];
  assign o[13957] = i[13957];
  assign o[13956] = i[13956];
  assign o[13955] = i[13955];
  assign o[13954] = i[13954];
  assign o[13953] = i[13953];
  assign o[13952] = i[13952];
  assign o[13951] = i[13951];
  assign o[13950] = i[13950];
  assign o[13949] = i[13949];
  assign o[13948] = i[13948];
  assign o[13947] = i[13947];
  assign o[13946] = i[13946];
  assign o[13945] = i[13945];
  assign o[13944] = i[13944];
  assign o[13943] = i[13943];
  assign o[13942] = i[13942];
  assign o[13941] = i[13941];
  assign o[13940] = i[13940];
  assign o[13939] = i[13939];
  assign o[13938] = i[13938];
  assign o[13937] = i[13937];
  assign o[13936] = i[13936];
  assign o[13935] = i[13935];
  assign o[13934] = i[13934];
  assign o[13933] = i[13933];
  assign o[13932] = i[13932];
  assign o[13931] = i[13931];
  assign o[13930] = i[13930];
  assign o[13929] = i[13929];
  assign o[13928] = i[13928];
  assign o[13927] = i[13927];
  assign o[13926] = i[13926];
  assign o[13925] = i[13925];
  assign o[13924] = i[13924];
  assign o[13923] = i[13923];
  assign o[13922] = i[13922];
  assign o[13921] = i[13921];
  assign o[13920] = i[13920];
  assign o[13919] = i[13919];
  assign o[13918] = i[13918];
  assign o[13917] = i[13917];
  assign o[13916] = i[13916];
  assign o[13915] = i[13915];
  assign o[13914] = i[13914];
  assign o[13913] = i[13913];
  assign o[13912] = i[13912];
  assign o[13911] = i[13911];
  assign o[13910] = i[13910];
  assign o[13909] = i[13909];
  assign o[13908] = i[13908];
  assign o[13907] = i[13907];
  assign o[13906] = i[13906];
  assign o[13905] = i[13905];
  assign o[13904] = i[13904];
  assign o[13903] = i[13903];
  assign o[13902] = i[13902];
  assign o[13901] = i[13901];
  assign o[13900] = i[13900];
  assign o[13899] = i[13899];
  assign o[13898] = i[13898];
  assign o[13897] = i[13897];
  assign o[13896] = i[13896];
  assign o[13895] = i[13895];
  assign o[13894] = i[13894];
  assign o[13893] = i[13893];
  assign o[13892] = i[13892];
  assign o[13891] = i[13891];
  assign o[13890] = i[13890];
  assign o[13889] = i[13889];
  assign o[13888] = i[13888];
  assign o[13887] = i[13887];
  assign o[13886] = i[13886];
  assign o[13885] = i[13885];
  assign o[13884] = i[13884];
  assign o[13883] = i[13883];
  assign o[13882] = i[13882];
  assign o[13881] = i[13881];
  assign o[13880] = i[13880];
  assign o[13879] = i[13879];
  assign o[13878] = i[13878];
  assign o[13877] = i[13877];
  assign o[13876] = i[13876];
  assign o[13875] = i[13875];
  assign o[13874] = i[13874];
  assign o[13873] = i[13873];
  assign o[13872] = i[13872];
  assign o[13871] = i[13871];
  assign o[13870] = i[13870];
  assign o[13869] = i[13869];
  assign o[13868] = i[13868];
  assign o[13867] = i[13867];
  assign o[13866] = i[13866];
  assign o[13865] = i[13865];
  assign o[13864] = i[13864];
  assign o[13863] = i[13863];
  assign o[13862] = i[13862];
  assign o[13861] = i[13861];
  assign o[13860] = i[13860];
  assign o[13859] = i[13859];
  assign o[13858] = i[13858];
  assign o[13857] = i[13857];
  assign o[13856] = i[13856];
  assign o[13855] = i[13855];
  assign o[13854] = i[13854];
  assign o[13853] = i[13853];
  assign o[13852] = i[13852];
  assign o[13851] = i[13851];
  assign o[13850] = i[13850];
  assign o[13849] = i[13849];
  assign o[13848] = i[13848];
  assign o[13847] = i[13847];
  assign o[13846] = i[13846];
  assign o[13845] = i[13845];
  assign o[13844] = i[13844];
  assign o[13843] = i[13843];
  assign o[13842] = i[13842];
  assign o[13841] = i[13841];
  assign o[13840] = i[13840];
  assign o[13839] = i[13839];
  assign o[13838] = i[13838];
  assign o[13837] = i[13837];
  assign o[13836] = i[13836];
  assign o[13835] = i[13835];
  assign o[13834] = i[13834];
  assign o[13833] = i[13833];
  assign o[13832] = i[13832];
  assign o[13831] = i[13831];
  assign o[13830] = i[13830];
  assign o[13829] = i[13829];
  assign o[13828] = i[13828];
  assign o[13827] = i[13827];
  assign o[13826] = i[13826];
  assign o[13825] = i[13825];
  assign o[13824] = i[13824];
  assign o[13823] = i[13823];
  assign o[13822] = i[13822];
  assign o[13821] = i[13821];
  assign o[13820] = i[13820];
  assign o[13819] = i[13819];
  assign o[13818] = i[13818];
  assign o[13817] = i[13817];
  assign o[13816] = i[13816];
  assign o[13815] = i[13815];
  assign o[13814] = i[13814];
  assign o[13813] = i[13813];
  assign o[13812] = i[13812];
  assign o[13811] = i[13811];
  assign o[13810] = i[13810];
  assign o[13809] = i[13809];
  assign o[13808] = i[13808];
  assign o[13807] = i[13807];
  assign o[13806] = i[13806];
  assign o[13805] = i[13805];
  assign o[13804] = i[13804];
  assign o[13803] = i[13803];
  assign o[13802] = i[13802];
  assign o[13801] = i[13801];
  assign o[13800] = i[13800];
  assign o[13799] = i[13799];
  assign o[13798] = i[13798];
  assign o[13797] = i[13797];
  assign o[13796] = i[13796];
  assign o[13795] = i[13795];
  assign o[13794] = i[13794];
  assign o[13793] = i[13793];
  assign o[13792] = i[13792];
  assign o[13791] = i[13791];
  assign o[13790] = i[13790];
  assign o[13789] = i[13789];
  assign o[13788] = i[13788];
  assign o[13787] = i[13787];
  assign o[13786] = i[13786];
  assign o[13785] = i[13785];
  assign o[13784] = i[13784];
  assign o[13783] = i[13783];
  assign o[13782] = i[13782];
  assign o[13781] = i[13781];
  assign o[13780] = i[13780];
  assign o[13779] = i[13779];
  assign o[13778] = i[13778];
  assign o[13777] = i[13777];
  assign o[13776] = i[13776];
  assign o[13775] = i[13775];
  assign o[13774] = i[13774];
  assign o[13773] = i[13773];
  assign o[13772] = i[13772];
  assign o[13771] = i[13771];
  assign o[13770] = i[13770];
  assign o[13769] = i[13769];
  assign o[13768] = i[13768];
  assign o[13767] = i[13767];
  assign o[13766] = i[13766];
  assign o[13765] = i[13765];
  assign o[13764] = i[13764];
  assign o[13763] = i[13763];
  assign o[13762] = i[13762];
  assign o[13761] = i[13761];
  assign o[13760] = i[13760];
  assign o[13759] = i[13759];
  assign o[13758] = i[13758];
  assign o[13757] = i[13757];
  assign o[13756] = i[13756];
  assign o[13755] = i[13755];
  assign o[13754] = i[13754];
  assign o[13753] = i[13753];
  assign o[13752] = i[13752];
  assign o[13751] = i[13751];
  assign o[13750] = i[13750];
  assign o[13749] = i[13749];
  assign o[13748] = i[13748];
  assign o[13747] = i[13747];
  assign o[13746] = i[13746];
  assign o[13745] = i[13745];
  assign o[13744] = i[13744];
  assign o[13743] = i[13743];
  assign o[13742] = i[13742];
  assign o[13741] = i[13741];
  assign o[13740] = i[13740];
  assign o[13739] = i[13739];
  assign o[13738] = i[13738];
  assign o[13737] = i[13737];
  assign o[13736] = i[13736];
  assign o[13735] = i[13735];
  assign o[13734] = i[13734];
  assign o[13733] = i[13733];
  assign o[13732] = i[13732];
  assign o[13731] = i[13731];
  assign o[13730] = i[13730];
  assign o[13729] = i[13729];
  assign o[13728] = i[13728];
  assign o[13727] = i[13727];
  assign o[13726] = i[13726];
  assign o[13725] = i[13725];
  assign o[13724] = i[13724];
  assign o[13723] = i[13723];
  assign o[13722] = i[13722];
  assign o[13721] = i[13721];
  assign o[13720] = i[13720];
  assign o[13719] = i[13719];
  assign o[13718] = i[13718];
  assign o[13717] = i[13717];
  assign o[13716] = i[13716];
  assign o[13715] = i[13715];
  assign o[13714] = i[13714];
  assign o[13713] = i[13713];
  assign o[13712] = i[13712];
  assign o[13711] = i[13711];
  assign o[13710] = i[13710];
  assign o[13709] = i[13709];
  assign o[13708] = i[13708];
  assign o[13707] = i[13707];
  assign o[13706] = i[13706];
  assign o[13705] = i[13705];
  assign o[13704] = i[13704];
  assign o[13703] = i[13703];
  assign o[13702] = i[13702];
  assign o[13701] = i[13701];
  assign o[13700] = i[13700];
  assign o[13699] = i[13699];
  assign o[13698] = i[13698];
  assign o[13697] = i[13697];
  assign o[13696] = i[13696];
  assign o[13695] = i[13695];
  assign o[13694] = i[13694];
  assign o[13693] = i[13693];
  assign o[13692] = i[13692];
  assign o[13691] = i[13691];
  assign o[13690] = i[13690];
  assign o[13689] = i[13689];
  assign o[13688] = i[13688];
  assign o[13687] = i[13687];
  assign o[13686] = i[13686];
  assign o[13685] = i[13685];
  assign o[13684] = i[13684];
  assign o[13683] = i[13683];
  assign o[13682] = i[13682];
  assign o[13681] = i[13681];
  assign o[13680] = i[13680];
  assign o[13679] = i[13679];
  assign o[13678] = i[13678];
  assign o[13677] = i[13677];
  assign o[13676] = i[13676];
  assign o[13675] = i[13675];
  assign o[13674] = i[13674];
  assign o[13673] = i[13673];
  assign o[13672] = i[13672];
  assign o[13671] = i[13671];
  assign o[13670] = i[13670];
  assign o[13669] = i[13669];
  assign o[13668] = i[13668];
  assign o[13667] = i[13667];
  assign o[13666] = i[13666];
  assign o[13665] = i[13665];
  assign o[13664] = i[13664];
  assign o[13663] = i[13663];
  assign o[13662] = i[13662];
  assign o[13661] = i[13661];
  assign o[13660] = i[13660];
  assign o[13659] = i[13659];
  assign o[13658] = i[13658];
  assign o[13657] = i[13657];
  assign o[13656] = i[13656];
  assign o[13655] = i[13655];
  assign o[13654] = i[13654];
  assign o[13653] = i[13653];
  assign o[13652] = i[13652];
  assign o[13651] = i[13651];
  assign o[13650] = i[13650];
  assign o[13649] = i[13649];
  assign o[13648] = i[13648];
  assign o[13647] = i[13647];
  assign o[13646] = i[13646];
  assign o[13645] = i[13645];
  assign o[13644] = i[13644];
  assign o[13643] = i[13643];
  assign o[13642] = i[13642];
  assign o[13641] = i[13641];
  assign o[13640] = i[13640];
  assign o[13639] = i[13639];
  assign o[13638] = i[13638];
  assign o[13637] = i[13637];
  assign o[13636] = i[13636];
  assign o[13635] = i[13635];
  assign o[13634] = i[13634];
  assign o[13633] = i[13633];
  assign o[13632] = i[13632];
  assign o[13631] = i[13631];
  assign o[13630] = i[13630];
  assign o[13629] = i[13629];
  assign o[13628] = i[13628];
  assign o[13627] = i[13627];
  assign o[13626] = i[13626];
  assign o[13625] = i[13625];
  assign o[13624] = i[13624];
  assign o[13623] = i[13623];
  assign o[13622] = i[13622];
  assign o[13621] = i[13621];
  assign o[13620] = i[13620];
  assign o[13619] = i[13619];
  assign o[13618] = i[13618];
  assign o[13617] = i[13617];
  assign o[13616] = i[13616];
  assign o[13615] = i[13615];
  assign o[13614] = i[13614];
  assign o[13613] = i[13613];
  assign o[13612] = i[13612];
  assign o[13611] = i[13611];
  assign o[13610] = i[13610];
  assign o[13609] = i[13609];
  assign o[13608] = i[13608];
  assign o[13607] = i[13607];
  assign o[13606] = i[13606];
  assign o[13605] = i[13605];
  assign o[13604] = i[13604];
  assign o[13603] = i[13603];
  assign o[13602] = i[13602];
  assign o[13601] = i[13601];
  assign o[13600] = i[13600];
  assign o[13599] = i[13599];
  assign o[13598] = i[13598];
  assign o[13597] = i[13597];
  assign o[13596] = i[13596];
  assign o[13595] = i[13595];
  assign o[13594] = i[13594];
  assign o[13593] = i[13593];
  assign o[13592] = i[13592];
  assign o[13591] = i[13591];
  assign o[13590] = i[13590];
  assign o[13589] = i[13589];
  assign o[13588] = i[13588];
  assign o[13587] = i[13587];
  assign o[13586] = i[13586];
  assign o[13585] = i[13585];
  assign o[13584] = i[13584];
  assign o[13583] = i[13583];
  assign o[13582] = i[13582];
  assign o[13581] = i[13581];
  assign o[13580] = i[13580];
  assign o[13579] = i[13579];
  assign o[13578] = i[13578];
  assign o[13577] = i[13577];
  assign o[13576] = i[13576];
  assign o[13575] = i[13575];
  assign o[13574] = i[13574];
  assign o[13573] = i[13573];
  assign o[13572] = i[13572];
  assign o[13571] = i[13571];
  assign o[13570] = i[13570];
  assign o[13569] = i[13569];
  assign o[13568] = i[13568];
  assign o[13567] = i[13567];
  assign o[13566] = i[13566];
  assign o[13565] = i[13565];
  assign o[13564] = i[13564];
  assign o[13563] = i[13563];
  assign o[13562] = i[13562];
  assign o[13561] = i[13561];
  assign o[13560] = i[13560];
  assign o[13559] = i[13559];
  assign o[13558] = i[13558];
  assign o[13557] = i[13557];
  assign o[13556] = i[13556];
  assign o[13555] = i[13555];
  assign o[13554] = i[13554];
  assign o[13553] = i[13553];
  assign o[13552] = i[13552];
  assign o[13551] = i[13551];
  assign o[13550] = i[13550];
  assign o[13549] = i[13549];
  assign o[13548] = i[13548];
  assign o[13547] = i[13547];
  assign o[13546] = i[13546];
  assign o[13545] = i[13545];
  assign o[13544] = i[13544];
  assign o[13543] = i[13543];
  assign o[13542] = i[13542];
  assign o[13541] = i[13541];
  assign o[13540] = i[13540];
  assign o[13539] = i[13539];
  assign o[13538] = i[13538];
  assign o[13537] = i[13537];
  assign o[13536] = i[13536];
  assign o[13535] = i[13535];
  assign o[13534] = i[13534];
  assign o[13533] = i[13533];
  assign o[13532] = i[13532];
  assign o[13531] = i[13531];
  assign o[13530] = i[13530];
  assign o[13529] = i[13529];
  assign o[13528] = i[13528];
  assign o[13527] = i[13527];
  assign o[13526] = i[13526];
  assign o[13525] = i[13525];
  assign o[13524] = i[13524];
  assign o[13523] = i[13523];
  assign o[13522] = i[13522];
  assign o[13521] = i[13521];
  assign o[13520] = i[13520];
  assign o[13519] = i[13519];
  assign o[13518] = i[13518];
  assign o[13517] = i[13517];
  assign o[13516] = i[13516];
  assign o[13515] = i[13515];
  assign o[13514] = i[13514];
  assign o[13513] = i[13513];
  assign o[13512] = i[13512];
  assign o[13511] = i[13511];
  assign o[13510] = i[13510];
  assign o[13509] = i[13509];
  assign o[13508] = i[13508];
  assign o[13507] = i[13507];
  assign o[13506] = i[13506];
  assign o[13505] = i[13505];
  assign o[13504] = i[13504];
  assign o[13503] = i[13503];
  assign o[13502] = i[13502];
  assign o[13501] = i[13501];
  assign o[13500] = i[13500];
  assign o[13499] = i[13499];
  assign o[13498] = i[13498];
  assign o[13497] = i[13497];
  assign o[13496] = i[13496];
  assign o[13495] = i[13495];
  assign o[13494] = i[13494];
  assign o[13493] = i[13493];
  assign o[13492] = i[13492];
  assign o[13491] = i[13491];
  assign o[13490] = i[13490];
  assign o[13489] = i[13489];
  assign o[13488] = i[13488];
  assign o[13487] = i[13487];
  assign o[13486] = i[13486];
  assign o[13485] = i[13485];
  assign o[13484] = i[13484];
  assign o[13483] = i[13483];
  assign o[13482] = i[13482];
  assign o[13481] = i[13481];
  assign o[13480] = i[13480];
  assign o[13479] = i[13479];
  assign o[13478] = i[13478];
  assign o[13477] = i[13477];
  assign o[13476] = i[13476];
  assign o[13475] = i[13475];
  assign o[13474] = i[13474];
  assign o[13473] = i[13473];
  assign o[13472] = i[13472];
  assign o[13471] = i[13471];
  assign o[13470] = i[13470];
  assign o[13469] = i[13469];
  assign o[13468] = i[13468];
  assign o[13467] = i[13467];
  assign o[13466] = i[13466];
  assign o[13465] = i[13465];
  assign o[13464] = i[13464];
  assign o[13463] = i[13463];
  assign o[13462] = i[13462];
  assign o[13461] = i[13461];
  assign o[13460] = i[13460];
  assign o[13459] = i[13459];
  assign o[13458] = i[13458];
  assign o[13457] = i[13457];
  assign o[13456] = i[13456];
  assign o[13455] = i[13455];
  assign o[13454] = i[13454];
  assign o[13453] = i[13453];
  assign o[13452] = i[13452];
  assign o[13451] = i[13451];
  assign o[13450] = i[13450];
  assign o[13449] = i[13449];
  assign o[13448] = i[13448];
  assign o[13447] = i[13447];
  assign o[13446] = i[13446];
  assign o[13445] = i[13445];
  assign o[13444] = i[13444];
  assign o[13443] = i[13443];
  assign o[13442] = i[13442];
  assign o[13441] = i[13441];
  assign o[13440] = i[13440];
  assign o[13439] = i[13439];
  assign o[13438] = i[13438];
  assign o[13437] = i[13437];
  assign o[13436] = i[13436];
  assign o[13435] = i[13435];
  assign o[13434] = i[13434];
  assign o[13433] = i[13433];
  assign o[13432] = i[13432];
  assign o[13431] = i[13431];
  assign o[13430] = i[13430];
  assign o[13429] = i[13429];
  assign o[13428] = i[13428];
  assign o[13427] = i[13427];
  assign o[13426] = i[13426];
  assign o[13425] = i[13425];
  assign o[13424] = i[13424];
  assign o[13423] = i[13423];
  assign o[13422] = i[13422];
  assign o[13421] = i[13421];
  assign o[13420] = i[13420];
  assign o[13419] = i[13419];
  assign o[13418] = i[13418];
  assign o[13417] = i[13417];
  assign o[13416] = i[13416];
  assign o[13415] = i[13415];
  assign o[13414] = i[13414];
  assign o[13413] = i[13413];
  assign o[13412] = i[13412];
  assign o[13411] = i[13411];
  assign o[13410] = i[13410];
  assign o[13409] = i[13409];
  assign o[13408] = i[13408];
  assign o[13407] = i[13407];
  assign o[13406] = i[13406];
  assign o[13405] = i[13405];
  assign o[13404] = i[13404];
  assign o[13403] = i[13403];
  assign o[13402] = i[13402];
  assign o[13401] = i[13401];
  assign o[13400] = i[13400];
  assign o[13399] = i[13399];
  assign o[13398] = i[13398];
  assign o[13397] = i[13397];
  assign o[13396] = i[13396];
  assign o[13395] = i[13395];
  assign o[13394] = i[13394];
  assign o[13393] = i[13393];
  assign o[13392] = i[13392];
  assign o[13391] = i[13391];
  assign o[13390] = i[13390];
  assign o[13389] = i[13389];
  assign o[13388] = i[13388];
  assign o[13387] = i[13387];
  assign o[13386] = i[13386];
  assign o[13385] = i[13385];
  assign o[13384] = i[13384];
  assign o[13383] = i[13383];
  assign o[13382] = i[13382];
  assign o[13381] = i[13381];
  assign o[13380] = i[13380];
  assign o[13379] = i[13379];
  assign o[13378] = i[13378];
  assign o[13377] = i[13377];
  assign o[13376] = i[13376];
  assign o[13375] = i[13375];
  assign o[13374] = i[13374];
  assign o[13373] = i[13373];
  assign o[13372] = i[13372];
  assign o[13371] = i[13371];
  assign o[13370] = i[13370];
  assign o[13369] = i[13369];
  assign o[13368] = i[13368];
  assign o[13367] = i[13367];
  assign o[13366] = i[13366];
  assign o[13365] = i[13365];
  assign o[13364] = i[13364];
  assign o[13363] = i[13363];
  assign o[13362] = i[13362];
  assign o[13361] = i[13361];
  assign o[13360] = i[13360];
  assign o[13359] = i[13359];
  assign o[13358] = i[13358];
  assign o[13357] = i[13357];
  assign o[13356] = i[13356];
  assign o[13355] = i[13355];
  assign o[13354] = i[13354];
  assign o[13353] = i[13353];
  assign o[13352] = i[13352];
  assign o[13351] = i[13351];
  assign o[13350] = i[13350];
  assign o[13349] = i[13349];
  assign o[13348] = i[13348];
  assign o[13347] = i[13347];
  assign o[13346] = i[13346];
  assign o[13345] = i[13345];
  assign o[13344] = i[13344];
  assign o[13343] = i[13343];
  assign o[13342] = i[13342];
  assign o[13341] = i[13341];
  assign o[13340] = i[13340];
  assign o[13339] = i[13339];
  assign o[13338] = i[13338];
  assign o[13337] = i[13337];
  assign o[13336] = i[13336];
  assign o[13335] = i[13335];
  assign o[13334] = i[13334];
  assign o[13333] = i[13333];
  assign o[13332] = i[13332];
  assign o[13331] = i[13331];
  assign o[13330] = i[13330];
  assign o[13329] = i[13329];
  assign o[13328] = i[13328];
  assign o[13327] = i[13327];
  assign o[13326] = i[13326];
  assign o[13325] = i[13325];
  assign o[13324] = i[13324];
  assign o[13323] = i[13323];
  assign o[13322] = i[13322];
  assign o[13321] = i[13321];
  assign o[13320] = i[13320];
  assign o[13319] = i[13319];
  assign o[13318] = i[13318];
  assign o[13317] = i[13317];
  assign o[13316] = i[13316];
  assign o[13315] = i[13315];
  assign o[13314] = i[13314];
  assign o[13313] = i[13313];
  assign o[13312] = i[13312];
  assign o[13311] = i[13311];
  assign o[13310] = i[13310];
  assign o[13309] = i[13309];
  assign o[13308] = i[13308];
  assign o[13307] = i[13307];
  assign o[13306] = i[13306];
  assign o[13305] = i[13305];
  assign o[13304] = i[13304];
  assign o[13303] = i[13303];
  assign o[13302] = i[13302];
  assign o[13301] = i[13301];
  assign o[13300] = i[13300];
  assign o[13299] = i[13299];
  assign o[13298] = i[13298];
  assign o[13297] = i[13297];
  assign o[13296] = i[13296];
  assign o[13295] = i[13295];
  assign o[13294] = i[13294];
  assign o[13293] = i[13293];
  assign o[13292] = i[13292];
  assign o[13291] = i[13291];
  assign o[13290] = i[13290];
  assign o[13289] = i[13289];
  assign o[13288] = i[13288];
  assign o[13287] = i[13287];
  assign o[13286] = i[13286];
  assign o[13285] = i[13285];
  assign o[13284] = i[13284];
  assign o[13283] = i[13283];
  assign o[13282] = i[13282];
  assign o[13281] = i[13281];
  assign o[13280] = i[13280];
  assign o[13279] = i[13279];
  assign o[13278] = i[13278];
  assign o[13277] = i[13277];
  assign o[13276] = i[13276];
  assign o[13275] = i[13275];
  assign o[13274] = i[13274];
  assign o[13273] = i[13273];
  assign o[13272] = i[13272];
  assign o[13271] = i[13271];
  assign o[13270] = i[13270];
  assign o[13269] = i[13269];
  assign o[13268] = i[13268];
  assign o[13267] = i[13267];
  assign o[13266] = i[13266];
  assign o[13265] = i[13265];
  assign o[13264] = i[13264];
  assign o[13263] = i[13263];
  assign o[13262] = i[13262];
  assign o[13261] = i[13261];
  assign o[13260] = i[13260];
  assign o[13259] = i[13259];
  assign o[13258] = i[13258];
  assign o[13257] = i[13257];
  assign o[13256] = i[13256];
  assign o[13255] = i[13255];
  assign o[13254] = i[13254];
  assign o[13253] = i[13253];
  assign o[13252] = i[13252];
  assign o[13251] = i[13251];
  assign o[13250] = i[13250];
  assign o[13249] = i[13249];
  assign o[13248] = i[13248];
  assign o[13247] = i[13247];
  assign o[13246] = i[13246];
  assign o[13245] = i[13245];
  assign o[13244] = i[13244];
  assign o[13243] = i[13243];
  assign o[13242] = i[13242];
  assign o[13241] = i[13241];
  assign o[13240] = i[13240];
  assign o[13239] = i[13239];
  assign o[13238] = i[13238];
  assign o[13237] = i[13237];
  assign o[13236] = i[13236];
  assign o[13235] = i[13235];
  assign o[13234] = i[13234];
  assign o[13233] = i[13233];
  assign o[13232] = i[13232];
  assign o[13231] = i[13231];
  assign o[13230] = i[13230];
  assign o[13229] = i[13229];
  assign o[13228] = i[13228];
  assign o[13227] = i[13227];
  assign o[13226] = i[13226];
  assign o[13225] = i[13225];
  assign o[13224] = i[13224];
  assign o[13223] = i[13223];
  assign o[13222] = i[13222];
  assign o[13221] = i[13221];
  assign o[13220] = i[13220];
  assign o[13219] = i[13219];
  assign o[13218] = i[13218];
  assign o[13217] = i[13217];
  assign o[13216] = i[13216];
  assign o[13215] = i[13215];
  assign o[13214] = i[13214];
  assign o[13213] = i[13213];
  assign o[13212] = i[13212];
  assign o[13211] = i[13211];
  assign o[13210] = i[13210];
  assign o[13209] = i[13209];
  assign o[13208] = i[13208];
  assign o[13207] = i[13207];
  assign o[13206] = i[13206];
  assign o[13205] = i[13205];
  assign o[13204] = i[13204];
  assign o[13203] = i[13203];
  assign o[13202] = i[13202];
  assign o[13201] = i[13201];
  assign o[13200] = i[13200];
  assign o[13199] = i[13199];
  assign o[13198] = i[13198];
  assign o[13197] = i[13197];
  assign o[13196] = i[13196];
  assign o[13195] = i[13195];
  assign o[13194] = i[13194];
  assign o[13193] = i[13193];
  assign o[13192] = i[13192];
  assign o[13191] = i[13191];
  assign o[13190] = i[13190];
  assign o[13189] = i[13189];
  assign o[13188] = i[13188];
  assign o[13187] = i[13187];
  assign o[13186] = i[13186];
  assign o[13185] = i[13185];
  assign o[13184] = i[13184];
  assign o[13183] = i[13183];
  assign o[13182] = i[13182];
  assign o[13181] = i[13181];
  assign o[13180] = i[13180];
  assign o[13179] = i[13179];
  assign o[13178] = i[13178];
  assign o[13177] = i[13177];
  assign o[13176] = i[13176];
  assign o[13175] = i[13175];
  assign o[13174] = i[13174];
  assign o[13173] = i[13173];
  assign o[13172] = i[13172];
  assign o[13171] = i[13171];
  assign o[13170] = i[13170];
  assign o[13169] = i[13169];
  assign o[13168] = i[13168];
  assign o[13167] = i[13167];
  assign o[13166] = i[13166];
  assign o[13165] = i[13165];
  assign o[13164] = i[13164];
  assign o[13163] = i[13163];
  assign o[13162] = i[13162];
  assign o[13161] = i[13161];
  assign o[13160] = i[13160];
  assign o[13159] = i[13159];
  assign o[13158] = i[13158];
  assign o[13157] = i[13157];
  assign o[13156] = i[13156];
  assign o[13155] = i[13155];
  assign o[13154] = i[13154];
  assign o[13153] = i[13153];
  assign o[13152] = i[13152];
  assign o[13151] = i[13151];
  assign o[13150] = i[13150];
  assign o[13149] = i[13149];
  assign o[13148] = i[13148];
  assign o[13147] = i[13147];
  assign o[13146] = i[13146];
  assign o[13145] = i[13145];
  assign o[13144] = i[13144];
  assign o[13143] = i[13143];
  assign o[13142] = i[13142];
  assign o[13141] = i[13141];
  assign o[13140] = i[13140];
  assign o[13139] = i[13139];
  assign o[13138] = i[13138];
  assign o[13137] = i[13137];
  assign o[13136] = i[13136];
  assign o[13135] = i[13135];
  assign o[13134] = i[13134];
  assign o[13133] = i[13133];
  assign o[13132] = i[13132];
  assign o[13131] = i[13131];
  assign o[13130] = i[13130];
  assign o[13129] = i[13129];
  assign o[13128] = i[13128];
  assign o[13127] = i[13127];
  assign o[13126] = i[13126];
  assign o[13125] = i[13125];
  assign o[13124] = i[13124];
  assign o[13123] = i[13123];
  assign o[13122] = i[13122];
  assign o[13121] = i[13121];
  assign o[13120] = i[13120];
  assign o[13119] = i[13119];
  assign o[13118] = i[13118];
  assign o[13117] = i[13117];
  assign o[13116] = i[13116];
  assign o[13115] = i[13115];
  assign o[13114] = i[13114];
  assign o[13113] = i[13113];
  assign o[13112] = i[13112];
  assign o[13111] = i[13111];
  assign o[13110] = i[13110];
  assign o[13109] = i[13109];
  assign o[13108] = i[13108];
  assign o[13107] = i[13107];
  assign o[13106] = i[13106];
  assign o[13105] = i[13105];
  assign o[13104] = i[13104];
  assign o[13103] = i[13103];
  assign o[13102] = i[13102];
  assign o[13101] = i[13101];
  assign o[13100] = i[13100];
  assign o[13099] = i[13099];
  assign o[13098] = i[13098];
  assign o[13097] = i[13097];
  assign o[13096] = i[13096];
  assign o[13095] = i[13095];
  assign o[13094] = i[13094];
  assign o[13093] = i[13093];
  assign o[13092] = i[13092];
  assign o[13091] = i[13091];
  assign o[13090] = i[13090];
  assign o[13089] = i[13089];
  assign o[13088] = i[13088];
  assign o[13087] = i[13087];
  assign o[13086] = i[13086];
  assign o[13085] = i[13085];
  assign o[13084] = i[13084];
  assign o[13083] = i[13083];
  assign o[13082] = i[13082];
  assign o[13081] = i[13081];
  assign o[13080] = i[13080];
  assign o[13079] = i[13079];
  assign o[13078] = i[13078];
  assign o[13077] = i[13077];
  assign o[13076] = i[13076];
  assign o[13075] = i[13075];
  assign o[13074] = i[13074];
  assign o[13073] = i[13073];
  assign o[13072] = i[13072];
  assign o[13071] = i[13071];
  assign o[13070] = i[13070];
  assign o[13069] = i[13069];
  assign o[13068] = i[13068];
  assign o[13067] = i[13067];
  assign o[13066] = i[13066];
  assign o[13065] = i[13065];
  assign o[13064] = i[13064];
  assign o[13063] = i[13063];
  assign o[13062] = i[13062];
  assign o[13061] = i[13061];
  assign o[13060] = i[13060];
  assign o[13059] = i[13059];
  assign o[13058] = i[13058];
  assign o[13057] = i[13057];
  assign o[13056] = i[13056];
  assign o[13055] = i[13055];
  assign o[13054] = i[13054];
  assign o[13053] = i[13053];
  assign o[13052] = i[13052];
  assign o[13051] = i[13051];
  assign o[13050] = i[13050];
  assign o[13049] = i[13049];
  assign o[13048] = i[13048];
  assign o[13047] = i[13047];
  assign o[13046] = i[13046];
  assign o[13045] = i[13045];
  assign o[13044] = i[13044];
  assign o[13043] = i[13043];
  assign o[13042] = i[13042];
  assign o[13041] = i[13041];
  assign o[13040] = i[13040];
  assign o[13039] = i[13039];
  assign o[13038] = i[13038];
  assign o[13037] = i[13037];
  assign o[13036] = i[13036];
  assign o[13035] = i[13035];
  assign o[13034] = i[13034];
  assign o[13033] = i[13033];
  assign o[13032] = i[13032];
  assign o[13031] = i[13031];
  assign o[13030] = i[13030];
  assign o[13029] = i[13029];
  assign o[13028] = i[13028];
  assign o[13027] = i[13027];
  assign o[13026] = i[13026];
  assign o[13025] = i[13025];
  assign o[13024] = i[13024];
  assign o[13023] = i[13023];
  assign o[13022] = i[13022];
  assign o[13021] = i[13021];
  assign o[13020] = i[13020];
  assign o[13019] = i[13019];
  assign o[13018] = i[13018];
  assign o[13017] = i[13017];
  assign o[13016] = i[13016];
  assign o[13015] = i[13015];
  assign o[13014] = i[13014];
  assign o[13013] = i[13013];
  assign o[13012] = i[13012];
  assign o[13011] = i[13011];
  assign o[13010] = i[13010];
  assign o[13009] = i[13009];
  assign o[13008] = i[13008];
  assign o[13007] = i[13007];
  assign o[13006] = i[13006];
  assign o[13005] = i[13005];
  assign o[13004] = i[13004];
  assign o[13003] = i[13003];
  assign o[13002] = i[13002];
  assign o[13001] = i[13001];
  assign o[13000] = i[13000];
  assign o[12999] = i[12999];
  assign o[12998] = i[12998];
  assign o[12997] = i[12997];
  assign o[12996] = i[12996];
  assign o[12995] = i[12995];
  assign o[12994] = i[12994];
  assign o[12993] = i[12993];
  assign o[12992] = i[12992];
  assign o[12991] = i[12991];
  assign o[12990] = i[12990];
  assign o[12989] = i[12989];
  assign o[12988] = i[12988];
  assign o[12987] = i[12987];
  assign o[12986] = i[12986];
  assign o[12985] = i[12985];
  assign o[12984] = i[12984];
  assign o[12983] = i[12983];
  assign o[12982] = i[12982];
  assign o[12981] = i[12981];
  assign o[12980] = i[12980];
  assign o[12979] = i[12979];
  assign o[12978] = i[12978];
  assign o[12977] = i[12977];
  assign o[12976] = i[12976];
  assign o[12975] = i[12975];
  assign o[12974] = i[12974];
  assign o[12973] = i[12973];
  assign o[12972] = i[12972];
  assign o[12971] = i[12971];
  assign o[12970] = i[12970];
  assign o[12969] = i[12969];
  assign o[12968] = i[12968];
  assign o[12967] = i[12967];
  assign o[12966] = i[12966];
  assign o[12965] = i[12965];
  assign o[12964] = i[12964];
  assign o[12963] = i[12963];
  assign o[12962] = i[12962];
  assign o[12961] = i[12961];
  assign o[12960] = i[12960];
  assign o[12959] = i[12959];
  assign o[12958] = i[12958];
  assign o[12957] = i[12957];
  assign o[12956] = i[12956];
  assign o[12955] = i[12955];
  assign o[12954] = i[12954];
  assign o[12953] = i[12953];
  assign o[12952] = i[12952];
  assign o[12951] = i[12951];
  assign o[12950] = i[12950];
  assign o[12949] = i[12949];
  assign o[12948] = i[12948];
  assign o[12947] = i[12947];
  assign o[12946] = i[12946];
  assign o[12945] = i[12945];
  assign o[12944] = i[12944];
  assign o[12943] = i[12943];
  assign o[12942] = i[12942];
  assign o[12941] = i[12941];
  assign o[12940] = i[12940];
  assign o[12939] = i[12939];
  assign o[12938] = i[12938];
  assign o[12937] = i[12937];
  assign o[12936] = i[12936];
  assign o[12935] = i[12935];
  assign o[12934] = i[12934];
  assign o[12933] = i[12933];
  assign o[12932] = i[12932];
  assign o[12931] = i[12931];
  assign o[12930] = i[12930];
  assign o[12929] = i[12929];
  assign o[12928] = i[12928];
  assign o[12927] = i[12927];
  assign o[12926] = i[12926];
  assign o[12925] = i[12925];
  assign o[12924] = i[12924];
  assign o[12923] = i[12923];
  assign o[12922] = i[12922];
  assign o[12921] = i[12921];
  assign o[12920] = i[12920];
  assign o[12919] = i[12919];
  assign o[12918] = i[12918];
  assign o[12917] = i[12917];
  assign o[12916] = i[12916];
  assign o[12915] = i[12915];
  assign o[12914] = i[12914];
  assign o[12913] = i[12913];
  assign o[12912] = i[12912];
  assign o[12911] = i[12911];
  assign o[12910] = i[12910];
  assign o[12909] = i[12909];
  assign o[12908] = i[12908];
  assign o[12907] = i[12907];
  assign o[12906] = i[12906];
  assign o[12905] = i[12905];
  assign o[12904] = i[12904];
  assign o[12903] = i[12903];
  assign o[12902] = i[12902];
  assign o[12901] = i[12901];
  assign o[12900] = i[12900];
  assign o[12899] = i[12899];
  assign o[12898] = i[12898];
  assign o[12897] = i[12897];
  assign o[12896] = i[12896];
  assign o[12895] = i[12895];
  assign o[12894] = i[12894];
  assign o[12893] = i[12893];
  assign o[12892] = i[12892];
  assign o[12891] = i[12891];
  assign o[12890] = i[12890];
  assign o[12889] = i[12889];
  assign o[12888] = i[12888];
  assign o[12887] = i[12887];
  assign o[12886] = i[12886];
  assign o[12885] = i[12885];
  assign o[12884] = i[12884];
  assign o[12883] = i[12883];
  assign o[12882] = i[12882];
  assign o[12881] = i[12881];
  assign o[12880] = i[12880];
  assign o[12879] = i[12879];
  assign o[12878] = i[12878];
  assign o[12877] = i[12877];
  assign o[12876] = i[12876];
  assign o[12875] = i[12875];
  assign o[12874] = i[12874];
  assign o[12873] = i[12873];
  assign o[12872] = i[12872];
  assign o[12871] = i[12871];
  assign o[12870] = i[12870];
  assign o[12869] = i[12869];
  assign o[12868] = i[12868];
  assign o[12867] = i[12867];
  assign o[12866] = i[12866];
  assign o[12865] = i[12865];
  assign o[12864] = i[12864];
  assign o[12863] = i[12863];
  assign o[12862] = i[12862];
  assign o[12861] = i[12861];
  assign o[12860] = i[12860];
  assign o[12859] = i[12859];
  assign o[12858] = i[12858];
  assign o[12857] = i[12857];
  assign o[12856] = i[12856];
  assign o[12855] = i[12855];
  assign o[12854] = i[12854];
  assign o[12853] = i[12853];
  assign o[12852] = i[12852];
  assign o[12851] = i[12851];
  assign o[12850] = i[12850];
  assign o[12849] = i[12849];
  assign o[12848] = i[12848];
  assign o[12847] = i[12847];
  assign o[12846] = i[12846];
  assign o[12845] = i[12845];
  assign o[12844] = i[12844];
  assign o[12843] = i[12843];
  assign o[12842] = i[12842];
  assign o[12841] = i[12841];
  assign o[12840] = i[12840];
  assign o[12839] = i[12839];
  assign o[12838] = i[12838];
  assign o[12837] = i[12837];
  assign o[12836] = i[12836];
  assign o[12835] = i[12835];
  assign o[12834] = i[12834];
  assign o[12833] = i[12833];
  assign o[12832] = i[12832];
  assign o[12831] = i[12831];
  assign o[12830] = i[12830];
  assign o[12829] = i[12829];
  assign o[12828] = i[12828];
  assign o[12827] = i[12827];
  assign o[12826] = i[12826];
  assign o[12825] = i[12825];
  assign o[12824] = i[12824];
  assign o[12823] = i[12823];
  assign o[12822] = i[12822];
  assign o[12821] = i[12821];
  assign o[12820] = i[12820];
  assign o[12819] = i[12819];
  assign o[12818] = i[12818];
  assign o[12817] = i[12817];
  assign o[12816] = i[12816];
  assign o[12815] = i[12815];
  assign o[12814] = i[12814];
  assign o[12813] = i[12813];
  assign o[12812] = i[12812];
  assign o[12811] = i[12811];
  assign o[12810] = i[12810];
  assign o[12809] = i[12809];
  assign o[12808] = i[12808];
  assign o[12807] = i[12807];
  assign o[12806] = i[12806];
  assign o[12805] = i[12805];
  assign o[12804] = i[12804];
  assign o[12803] = i[12803];
  assign o[12802] = i[12802];
  assign o[12801] = i[12801];
  assign o[12800] = i[12800];
  assign o[12799] = i[12799];
  assign o[12798] = i[12798];
  assign o[12797] = i[12797];
  assign o[12796] = i[12796];
  assign o[12795] = i[12795];
  assign o[12794] = i[12794];
  assign o[12793] = i[12793];
  assign o[12792] = i[12792];
  assign o[12791] = i[12791];
  assign o[12790] = i[12790];
  assign o[12789] = i[12789];
  assign o[12788] = i[12788];
  assign o[12787] = i[12787];
  assign o[12786] = i[12786];
  assign o[12785] = i[12785];
  assign o[12784] = i[12784];
  assign o[12783] = i[12783];
  assign o[12782] = i[12782];
  assign o[12781] = i[12781];
  assign o[12780] = i[12780];
  assign o[12779] = i[12779];
  assign o[12778] = i[12778];
  assign o[12777] = i[12777];
  assign o[12776] = i[12776];
  assign o[12775] = i[12775];
  assign o[12774] = i[12774];
  assign o[12773] = i[12773];
  assign o[12772] = i[12772];
  assign o[12771] = i[12771];
  assign o[12770] = i[12770];
  assign o[12769] = i[12769];
  assign o[12768] = i[12768];
  assign o[12767] = i[12767];
  assign o[12766] = i[12766];
  assign o[12765] = i[12765];
  assign o[12764] = i[12764];
  assign o[12763] = i[12763];
  assign o[12762] = i[12762];
  assign o[12761] = i[12761];
  assign o[12760] = i[12760];
  assign o[12759] = i[12759];
  assign o[12758] = i[12758];
  assign o[12757] = i[12757];
  assign o[12756] = i[12756];
  assign o[12755] = i[12755];
  assign o[12754] = i[12754];
  assign o[12753] = i[12753];
  assign o[12752] = i[12752];
  assign o[12751] = i[12751];
  assign o[12750] = i[12750];
  assign o[12749] = i[12749];
  assign o[12748] = i[12748];
  assign o[12747] = i[12747];
  assign o[12746] = i[12746];
  assign o[12745] = i[12745];
  assign o[12744] = i[12744];
  assign o[12743] = i[12743];
  assign o[12742] = i[12742];
  assign o[12741] = i[12741];
  assign o[12740] = i[12740];
  assign o[12739] = i[12739];
  assign o[12738] = i[12738];
  assign o[12737] = i[12737];
  assign o[12736] = i[12736];
  assign o[12735] = i[12735];
  assign o[12734] = i[12734];
  assign o[12733] = i[12733];
  assign o[12732] = i[12732];
  assign o[12731] = i[12731];
  assign o[12730] = i[12730];
  assign o[12729] = i[12729];
  assign o[12728] = i[12728];
  assign o[12727] = i[12727];
  assign o[12726] = i[12726];
  assign o[12725] = i[12725];
  assign o[12724] = i[12724];
  assign o[12723] = i[12723];
  assign o[12722] = i[12722];
  assign o[12721] = i[12721];
  assign o[12720] = i[12720];
  assign o[12719] = i[12719];
  assign o[12718] = i[12718];
  assign o[12717] = i[12717];
  assign o[12716] = i[12716];
  assign o[12715] = i[12715];
  assign o[12714] = i[12714];
  assign o[12713] = i[12713];
  assign o[12712] = i[12712];
  assign o[12711] = i[12711];
  assign o[12710] = i[12710];
  assign o[12709] = i[12709];
  assign o[12708] = i[12708];
  assign o[12707] = i[12707];
  assign o[12706] = i[12706];
  assign o[12705] = i[12705];
  assign o[12704] = i[12704];
  assign o[12703] = i[12703];
  assign o[12702] = i[12702];
  assign o[12701] = i[12701];
  assign o[12700] = i[12700];
  assign o[12699] = i[12699];
  assign o[12698] = i[12698];
  assign o[12697] = i[12697];
  assign o[12696] = i[12696];
  assign o[12695] = i[12695];
  assign o[12694] = i[12694];
  assign o[12693] = i[12693];
  assign o[12692] = i[12692];
  assign o[12691] = i[12691];
  assign o[12690] = i[12690];
  assign o[12689] = i[12689];
  assign o[12688] = i[12688];
  assign o[12687] = i[12687];
  assign o[12686] = i[12686];
  assign o[12685] = i[12685];
  assign o[12684] = i[12684];
  assign o[12683] = i[12683];
  assign o[12682] = i[12682];
  assign o[12681] = i[12681];
  assign o[12680] = i[12680];
  assign o[12679] = i[12679];
  assign o[12678] = i[12678];
  assign o[12677] = i[12677];
  assign o[12676] = i[12676];
  assign o[12675] = i[12675];
  assign o[12674] = i[12674];
  assign o[12673] = i[12673];
  assign o[12672] = i[12672];
  assign o[12671] = i[12671];
  assign o[12670] = i[12670];
  assign o[12669] = i[12669];
  assign o[12668] = i[12668];
  assign o[12667] = i[12667];
  assign o[12666] = i[12666];
  assign o[12665] = i[12665];
  assign o[12664] = i[12664];
  assign o[12663] = i[12663];
  assign o[12662] = i[12662];
  assign o[12661] = i[12661];
  assign o[12660] = i[12660];
  assign o[12659] = i[12659];
  assign o[12658] = i[12658];
  assign o[12657] = i[12657];
  assign o[12656] = i[12656];
  assign o[12655] = i[12655];
  assign o[12654] = i[12654];
  assign o[12653] = i[12653];
  assign o[12652] = i[12652];
  assign o[12651] = i[12651];
  assign o[12650] = i[12650];
  assign o[12649] = i[12649];
  assign o[12648] = i[12648];
  assign o[12647] = i[12647];
  assign o[12646] = i[12646];
  assign o[12645] = i[12645];
  assign o[12644] = i[12644];
  assign o[12643] = i[12643];
  assign o[12642] = i[12642];
  assign o[12641] = i[12641];
  assign o[12640] = i[12640];
  assign o[12639] = i[12639];
  assign o[12638] = i[12638];
  assign o[12637] = i[12637];
  assign o[12636] = i[12636];
  assign o[12635] = i[12635];
  assign o[12634] = i[12634];
  assign o[12633] = i[12633];
  assign o[12632] = i[12632];
  assign o[12631] = i[12631];
  assign o[12630] = i[12630];
  assign o[12629] = i[12629];
  assign o[12628] = i[12628];
  assign o[12627] = i[12627];
  assign o[12626] = i[12626];
  assign o[12625] = i[12625];
  assign o[12624] = i[12624];
  assign o[12623] = i[12623];
  assign o[12622] = i[12622];
  assign o[12621] = i[12621];
  assign o[12620] = i[12620];
  assign o[12619] = i[12619];
  assign o[12618] = i[12618];
  assign o[12617] = i[12617];
  assign o[12616] = i[12616];
  assign o[12615] = i[12615];
  assign o[12614] = i[12614];
  assign o[12613] = i[12613];
  assign o[12612] = i[12612];
  assign o[12611] = i[12611];
  assign o[12610] = i[12610];
  assign o[12609] = i[12609];
  assign o[12608] = i[12608];
  assign o[12607] = i[12607];
  assign o[12606] = i[12606];
  assign o[12605] = i[12605];
  assign o[12604] = i[12604];
  assign o[12603] = i[12603];
  assign o[12602] = i[12602];
  assign o[12601] = i[12601];
  assign o[12600] = i[12600];
  assign o[12599] = i[12599];
  assign o[12598] = i[12598];
  assign o[12597] = i[12597];
  assign o[12596] = i[12596];
  assign o[12595] = i[12595];
  assign o[12594] = i[12594];
  assign o[12593] = i[12593];
  assign o[12592] = i[12592];
  assign o[12591] = i[12591];
  assign o[12590] = i[12590];
  assign o[12589] = i[12589];
  assign o[12588] = i[12588];
  assign o[12587] = i[12587];
  assign o[12586] = i[12586];
  assign o[12585] = i[12585];
  assign o[12584] = i[12584];
  assign o[12583] = i[12583];
  assign o[12582] = i[12582];
  assign o[12581] = i[12581];
  assign o[12580] = i[12580];
  assign o[12579] = i[12579];
  assign o[12578] = i[12578];
  assign o[12577] = i[12577];
  assign o[12576] = i[12576];
  assign o[12575] = i[12575];
  assign o[12574] = i[12574];
  assign o[12573] = i[12573];
  assign o[12572] = i[12572];
  assign o[12571] = i[12571];
  assign o[12570] = i[12570];
  assign o[12569] = i[12569];
  assign o[12568] = i[12568];
  assign o[12567] = i[12567];
  assign o[12566] = i[12566];
  assign o[12565] = i[12565];
  assign o[12564] = i[12564];
  assign o[12563] = i[12563];
  assign o[12562] = i[12562];
  assign o[12561] = i[12561];
  assign o[12560] = i[12560];
  assign o[12559] = i[12559];
  assign o[12558] = i[12558];
  assign o[12557] = i[12557];
  assign o[12556] = i[12556];
  assign o[12555] = i[12555];
  assign o[12554] = i[12554];
  assign o[12553] = i[12553];
  assign o[12552] = i[12552];
  assign o[12551] = i[12551];
  assign o[12550] = i[12550];
  assign o[12549] = i[12549];
  assign o[12548] = i[12548];
  assign o[12547] = i[12547];
  assign o[12546] = i[12546];
  assign o[12545] = i[12545];
  assign o[12544] = i[12544];
  assign o[12543] = i[12543];
  assign o[12542] = i[12542];
  assign o[12541] = i[12541];
  assign o[12540] = i[12540];
  assign o[12539] = i[12539];
  assign o[12538] = i[12538];
  assign o[12537] = i[12537];
  assign o[12536] = i[12536];
  assign o[12535] = i[12535];
  assign o[12534] = i[12534];
  assign o[12533] = i[12533];
  assign o[12532] = i[12532];
  assign o[12531] = i[12531];
  assign o[12530] = i[12530];
  assign o[12529] = i[12529];
  assign o[12528] = i[12528];
  assign o[12527] = i[12527];
  assign o[12526] = i[12526];
  assign o[12525] = i[12525];
  assign o[12524] = i[12524];
  assign o[12523] = i[12523];
  assign o[12522] = i[12522];
  assign o[12521] = i[12521];
  assign o[12520] = i[12520];
  assign o[12519] = i[12519];
  assign o[12518] = i[12518];
  assign o[12517] = i[12517];
  assign o[12516] = i[12516];
  assign o[12515] = i[12515];
  assign o[12514] = i[12514];
  assign o[12513] = i[12513];
  assign o[12512] = i[12512];
  assign o[12511] = i[12511];
  assign o[12510] = i[12510];
  assign o[12509] = i[12509];
  assign o[12508] = i[12508];
  assign o[12507] = i[12507];
  assign o[12506] = i[12506];
  assign o[12505] = i[12505];
  assign o[12504] = i[12504];
  assign o[12503] = i[12503];
  assign o[12502] = i[12502];
  assign o[12501] = i[12501];
  assign o[12500] = i[12500];
  assign o[12499] = i[12499];
  assign o[12498] = i[12498];
  assign o[12497] = i[12497];
  assign o[12496] = i[12496];
  assign o[12495] = i[12495];
  assign o[12494] = i[12494];
  assign o[12493] = i[12493];
  assign o[12492] = i[12492];
  assign o[12491] = i[12491];
  assign o[12490] = i[12490];
  assign o[12489] = i[12489];
  assign o[12488] = i[12488];
  assign o[12487] = i[12487];
  assign o[12486] = i[12486];
  assign o[12485] = i[12485];
  assign o[12484] = i[12484];
  assign o[12483] = i[12483];
  assign o[12482] = i[12482];
  assign o[12481] = i[12481];
  assign o[12480] = i[12480];
  assign o[12479] = i[12479];
  assign o[12478] = i[12478];
  assign o[12477] = i[12477];
  assign o[12476] = i[12476];
  assign o[12475] = i[12475];
  assign o[12474] = i[12474];
  assign o[12473] = i[12473];
  assign o[12472] = i[12472];
  assign o[12471] = i[12471];
  assign o[12470] = i[12470];
  assign o[12469] = i[12469];
  assign o[12468] = i[12468];
  assign o[12467] = i[12467];
  assign o[12466] = i[12466];
  assign o[12465] = i[12465];
  assign o[12464] = i[12464];
  assign o[12463] = i[12463];
  assign o[12462] = i[12462];
  assign o[12461] = i[12461];
  assign o[12460] = i[12460];
  assign o[12459] = i[12459];
  assign o[12458] = i[12458];
  assign o[12457] = i[12457];
  assign o[12456] = i[12456];
  assign o[12455] = i[12455];
  assign o[12454] = i[12454];
  assign o[12453] = i[12453];
  assign o[12452] = i[12452];
  assign o[12451] = i[12451];
  assign o[12450] = i[12450];
  assign o[12449] = i[12449];
  assign o[12448] = i[12448];
  assign o[12447] = i[12447];
  assign o[12446] = i[12446];
  assign o[12445] = i[12445];
  assign o[12444] = i[12444];
  assign o[12443] = i[12443];
  assign o[12442] = i[12442];
  assign o[12441] = i[12441];
  assign o[12440] = i[12440];
  assign o[12439] = i[12439];
  assign o[12438] = i[12438];
  assign o[12437] = i[12437];
  assign o[12436] = i[12436];
  assign o[12435] = i[12435];
  assign o[12434] = i[12434];
  assign o[12433] = i[12433];
  assign o[12432] = i[12432];
  assign o[12431] = i[12431];
  assign o[12430] = i[12430];
  assign o[12429] = i[12429];
  assign o[12428] = i[12428];
  assign o[12427] = i[12427];
  assign o[12426] = i[12426];
  assign o[12425] = i[12425];
  assign o[12424] = i[12424];
  assign o[12423] = i[12423];
  assign o[12422] = i[12422];
  assign o[12421] = i[12421];
  assign o[12420] = i[12420];
  assign o[12419] = i[12419];
  assign o[12418] = i[12418];
  assign o[12417] = i[12417];
  assign o[12416] = i[12416];
  assign o[12415] = i[12415];
  assign o[12414] = i[12414];
  assign o[12413] = i[12413];
  assign o[12412] = i[12412];
  assign o[12411] = i[12411];
  assign o[12410] = i[12410];
  assign o[12409] = i[12409];
  assign o[12408] = i[12408];
  assign o[12407] = i[12407];
  assign o[12406] = i[12406];
  assign o[12405] = i[12405];
  assign o[12404] = i[12404];
  assign o[12403] = i[12403];
  assign o[12402] = i[12402];
  assign o[12401] = i[12401];
  assign o[12400] = i[12400];
  assign o[12399] = i[12399];
  assign o[12398] = i[12398];
  assign o[12397] = i[12397];
  assign o[12396] = i[12396];
  assign o[12395] = i[12395];
  assign o[12394] = i[12394];
  assign o[12393] = i[12393];
  assign o[12392] = i[12392];
  assign o[12391] = i[12391];
  assign o[12390] = i[12390];
  assign o[12389] = i[12389];
  assign o[12388] = i[12388];
  assign o[12387] = i[12387];
  assign o[12386] = i[12386];
  assign o[12385] = i[12385];
  assign o[12384] = i[12384];
  assign o[12383] = i[12383];
  assign o[12382] = i[12382];
  assign o[12381] = i[12381];
  assign o[12380] = i[12380];
  assign o[12379] = i[12379];
  assign o[12378] = i[12378];
  assign o[12377] = i[12377];
  assign o[12376] = i[12376];
  assign o[12375] = i[12375];
  assign o[12374] = i[12374];
  assign o[12373] = i[12373];
  assign o[12372] = i[12372];
  assign o[12371] = i[12371];
  assign o[12370] = i[12370];
  assign o[12369] = i[12369];
  assign o[12368] = i[12368];
  assign o[12367] = i[12367];
  assign o[12366] = i[12366];
  assign o[12365] = i[12365];
  assign o[12364] = i[12364];
  assign o[12363] = i[12363];
  assign o[12362] = i[12362];
  assign o[12361] = i[12361];
  assign o[12360] = i[12360];
  assign o[12359] = i[12359];
  assign o[12358] = i[12358];
  assign o[12357] = i[12357];
  assign o[12356] = i[12356];
  assign o[12355] = i[12355];
  assign o[12354] = i[12354];
  assign o[12353] = i[12353];
  assign o[12352] = i[12352];
  assign o[12351] = i[12351];
  assign o[12350] = i[12350];
  assign o[12349] = i[12349];
  assign o[12348] = i[12348];
  assign o[12347] = i[12347];
  assign o[12346] = i[12346];
  assign o[12345] = i[12345];
  assign o[12344] = i[12344];
  assign o[12343] = i[12343];
  assign o[12342] = i[12342];
  assign o[12341] = i[12341];
  assign o[12340] = i[12340];
  assign o[12339] = i[12339];
  assign o[12338] = i[12338];
  assign o[12337] = i[12337];
  assign o[12336] = i[12336];
  assign o[12335] = i[12335];
  assign o[12334] = i[12334];
  assign o[12333] = i[12333];
  assign o[12332] = i[12332];
  assign o[12331] = i[12331];
  assign o[12330] = i[12330];
  assign o[12329] = i[12329];
  assign o[12328] = i[12328];
  assign o[12327] = i[12327];
  assign o[12326] = i[12326];
  assign o[12325] = i[12325];
  assign o[12324] = i[12324];
  assign o[12323] = i[12323];
  assign o[12322] = i[12322];
  assign o[12321] = i[12321];
  assign o[12320] = i[12320];
  assign o[12319] = i[12319];
  assign o[12318] = i[12318];
  assign o[12317] = i[12317];
  assign o[12316] = i[12316];
  assign o[12315] = i[12315];
  assign o[12314] = i[12314];
  assign o[12313] = i[12313];
  assign o[12312] = i[12312];
  assign o[12311] = i[12311];
  assign o[12310] = i[12310];
  assign o[12309] = i[12309];
  assign o[12308] = i[12308];
  assign o[12307] = i[12307];
  assign o[12306] = i[12306];
  assign o[12305] = i[12305];
  assign o[12304] = i[12304];
  assign o[12303] = i[12303];
  assign o[12302] = i[12302];
  assign o[12301] = i[12301];
  assign o[12300] = i[12300];
  assign o[12299] = i[12299];
  assign o[12298] = i[12298];
  assign o[12297] = i[12297];
  assign o[12296] = i[12296];
  assign o[12295] = i[12295];
  assign o[12294] = i[12294];
  assign o[12293] = i[12293];
  assign o[12292] = i[12292];
  assign o[12291] = i[12291];
  assign o[12290] = i[12290];
  assign o[12289] = i[12289];
  assign o[12288] = i[12288];
  assign o[12287] = i[12287];
  assign o[12286] = i[12286];
  assign o[12285] = i[12285];
  assign o[12284] = i[12284];
  assign o[12283] = i[12283];
  assign o[12282] = i[12282];
  assign o[12281] = i[12281];
  assign o[12280] = i[12280];
  assign o[12279] = i[12279];
  assign o[12278] = i[12278];
  assign o[12277] = i[12277];
  assign o[12276] = i[12276];
  assign o[12275] = i[12275];
  assign o[12274] = i[12274];
  assign o[12273] = i[12273];
  assign o[12272] = i[12272];
  assign o[12271] = i[12271];
  assign o[12270] = i[12270];
  assign o[12269] = i[12269];
  assign o[12268] = i[12268];
  assign o[12267] = i[12267];
  assign o[12266] = i[12266];
  assign o[12265] = i[12265];
  assign o[12264] = i[12264];
  assign o[12263] = i[12263];
  assign o[12262] = i[12262];
  assign o[12261] = i[12261];
  assign o[12260] = i[12260];
  assign o[12259] = i[12259];
  assign o[12258] = i[12258];
  assign o[12257] = i[12257];
  assign o[12256] = i[12256];
  assign o[12255] = i[12255];
  assign o[12254] = i[12254];
  assign o[12253] = i[12253];
  assign o[12252] = i[12252];
  assign o[12251] = i[12251];
  assign o[12250] = i[12250];
  assign o[12249] = i[12249];
  assign o[12248] = i[12248];
  assign o[12247] = i[12247];
  assign o[12246] = i[12246];
  assign o[12245] = i[12245];
  assign o[12244] = i[12244];
  assign o[12243] = i[12243];
  assign o[12242] = i[12242];
  assign o[12241] = i[12241];
  assign o[12240] = i[12240];
  assign o[12239] = i[12239];
  assign o[12238] = i[12238];
  assign o[12237] = i[12237];
  assign o[12236] = i[12236];
  assign o[12235] = i[12235];
  assign o[12234] = i[12234];
  assign o[12233] = i[12233];
  assign o[12232] = i[12232];
  assign o[12231] = i[12231];
  assign o[12230] = i[12230];
  assign o[12229] = i[12229];
  assign o[12228] = i[12228];
  assign o[12227] = i[12227];
  assign o[12226] = i[12226];
  assign o[12225] = i[12225];
  assign o[12224] = i[12224];
  assign o[12223] = i[12223];
  assign o[12222] = i[12222];
  assign o[12221] = i[12221];
  assign o[12220] = i[12220];
  assign o[12219] = i[12219];
  assign o[12218] = i[12218];
  assign o[12217] = i[12217];
  assign o[12216] = i[12216];
  assign o[12215] = i[12215];
  assign o[12214] = i[12214];
  assign o[12213] = i[12213];
  assign o[12212] = i[12212];
  assign o[12211] = i[12211];
  assign o[12210] = i[12210];
  assign o[12209] = i[12209];
  assign o[12208] = i[12208];
  assign o[12207] = i[12207];
  assign o[12206] = i[12206];
  assign o[12205] = i[12205];
  assign o[12204] = i[12204];
  assign o[12203] = i[12203];
  assign o[12202] = i[12202];
  assign o[12201] = i[12201];
  assign o[12200] = i[12200];
  assign o[12199] = i[12199];
  assign o[12198] = i[12198];
  assign o[12197] = i[12197];
  assign o[12196] = i[12196];
  assign o[12195] = i[12195];
  assign o[12194] = i[12194];
  assign o[12193] = i[12193];
  assign o[12192] = i[12192];
  assign o[12191] = i[12191];
  assign o[12190] = i[12190];
  assign o[12189] = i[12189];
  assign o[12188] = i[12188];
  assign o[12187] = i[12187];
  assign o[12186] = i[12186];
  assign o[12185] = i[12185];
  assign o[12184] = i[12184];
  assign o[12183] = i[12183];
  assign o[12182] = i[12182];
  assign o[12181] = i[12181];
  assign o[12180] = i[12180];
  assign o[12179] = i[12179];
  assign o[12178] = i[12178];
  assign o[12177] = i[12177];
  assign o[12176] = i[12176];
  assign o[12175] = i[12175];
  assign o[12174] = i[12174];
  assign o[12173] = i[12173];
  assign o[12172] = i[12172];
  assign o[12171] = i[12171];
  assign o[12170] = i[12170];
  assign o[12169] = i[12169];
  assign o[12168] = i[12168];
  assign o[12167] = i[12167];
  assign o[12166] = i[12166];
  assign o[12165] = i[12165];
  assign o[12164] = i[12164];
  assign o[12163] = i[12163];
  assign o[12162] = i[12162];
  assign o[12161] = i[12161];
  assign o[12160] = i[12160];
  assign o[12159] = i[12159];
  assign o[12158] = i[12158];
  assign o[12157] = i[12157];
  assign o[12156] = i[12156];
  assign o[12155] = i[12155];
  assign o[12154] = i[12154];
  assign o[12153] = i[12153];
  assign o[12152] = i[12152];
  assign o[12151] = i[12151];
  assign o[12150] = i[12150];
  assign o[12149] = i[12149];
  assign o[12148] = i[12148];
  assign o[12147] = i[12147];
  assign o[12146] = i[12146];
  assign o[12145] = i[12145];
  assign o[12144] = i[12144];
  assign o[12143] = i[12143];
  assign o[12142] = i[12142];
  assign o[12141] = i[12141];
  assign o[12140] = i[12140];
  assign o[12139] = i[12139];
  assign o[12138] = i[12138];
  assign o[12137] = i[12137];
  assign o[12136] = i[12136];
  assign o[12135] = i[12135];
  assign o[12134] = i[12134];
  assign o[12133] = i[12133];
  assign o[12132] = i[12132];
  assign o[12131] = i[12131];
  assign o[12130] = i[12130];
  assign o[12129] = i[12129];
  assign o[12128] = i[12128];
  assign o[12127] = i[12127];
  assign o[12126] = i[12126];
  assign o[12125] = i[12125];
  assign o[12124] = i[12124];
  assign o[12123] = i[12123];
  assign o[12122] = i[12122];
  assign o[12121] = i[12121];
  assign o[12120] = i[12120];
  assign o[12119] = i[12119];
  assign o[12118] = i[12118];
  assign o[12117] = i[12117];
  assign o[12116] = i[12116];
  assign o[12115] = i[12115];
  assign o[12114] = i[12114];
  assign o[12113] = i[12113];
  assign o[12112] = i[12112];
  assign o[12111] = i[12111];
  assign o[12110] = i[12110];
  assign o[12109] = i[12109];
  assign o[12108] = i[12108];
  assign o[12107] = i[12107];
  assign o[12106] = i[12106];
  assign o[12105] = i[12105];
  assign o[12104] = i[12104];
  assign o[12103] = i[12103];
  assign o[12102] = i[12102];
  assign o[12101] = i[12101];
  assign o[12100] = i[12100];
  assign o[12099] = i[12099];
  assign o[12098] = i[12098];
  assign o[12097] = i[12097];
  assign o[12096] = i[12096];
  assign o[12095] = i[12095];
  assign o[12094] = i[12094];
  assign o[12093] = i[12093];
  assign o[12092] = i[12092];
  assign o[12091] = i[12091];
  assign o[12090] = i[12090];
  assign o[12089] = i[12089];
  assign o[12088] = i[12088];
  assign o[12087] = i[12087];
  assign o[12086] = i[12086];
  assign o[12085] = i[12085];
  assign o[12084] = i[12084];
  assign o[12083] = i[12083];
  assign o[12082] = i[12082];
  assign o[12081] = i[12081];
  assign o[12080] = i[12080];
  assign o[12079] = i[12079];
  assign o[12078] = i[12078];
  assign o[12077] = i[12077];
  assign o[12076] = i[12076];
  assign o[12075] = i[12075];
  assign o[12074] = i[12074];
  assign o[12073] = i[12073];
  assign o[12072] = i[12072];
  assign o[12071] = i[12071];
  assign o[12070] = i[12070];
  assign o[12069] = i[12069];
  assign o[12068] = i[12068];
  assign o[12067] = i[12067];
  assign o[12066] = i[12066];
  assign o[12065] = i[12065];
  assign o[12064] = i[12064];
  assign o[12063] = i[12063];
  assign o[12062] = i[12062];
  assign o[12061] = i[12061];
  assign o[12060] = i[12060];
  assign o[12059] = i[12059];
  assign o[12058] = i[12058];
  assign o[12057] = i[12057];
  assign o[12056] = i[12056];
  assign o[12055] = i[12055];
  assign o[12054] = i[12054];
  assign o[12053] = i[12053];
  assign o[12052] = i[12052];
  assign o[12051] = i[12051];
  assign o[12050] = i[12050];
  assign o[12049] = i[12049];
  assign o[12048] = i[12048];
  assign o[12047] = i[12047];
  assign o[12046] = i[12046];
  assign o[12045] = i[12045];
  assign o[12044] = i[12044];
  assign o[12043] = i[12043];
  assign o[12042] = i[12042];
  assign o[12041] = i[12041];
  assign o[12040] = i[12040];
  assign o[12039] = i[12039];
  assign o[12038] = i[12038];
  assign o[12037] = i[12037];
  assign o[12036] = i[12036];
  assign o[12035] = i[12035];
  assign o[12034] = i[12034];
  assign o[12033] = i[12033];
  assign o[12032] = i[12032];
  assign o[12031] = i[12031];
  assign o[12030] = i[12030];
  assign o[12029] = i[12029];
  assign o[12028] = i[12028];
  assign o[12027] = i[12027];
  assign o[12026] = i[12026];
  assign o[12025] = i[12025];
  assign o[12024] = i[12024];
  assign o[12023] = i[12023];
  assign o[12022] = i[12022];
  assign o[12021] = i[12021];
  assign o[12020] = i[12020];
  assign o[12019] = i[12019];
  assign o[12018] = i[12018];
  assign o[12017] = i[12017];
  assign o[12016] = i[12016];
  assign o[12015] = i[12015];
  assign o[12014] = i[12014];
  assign o[12013] = i[12013];
  assign o[12012] = i[12012];
  assign o[12011] = i[12011];
  assign o[12010] = i[12010];
  assign o[12009] = i[12009];
  assign o[12008] = i[12008];
  assign o[12007] = i[12007];
  assign o[12006] = i[12006];
  assign o[12005] = i[12005];
  assign o[12004] = i[12004];
  assign o[12003] = i[12003];
  assign o[12002] = i[12002];
  assign o[12001] = i[12001];
  assign o[12000] = i[12000];
  assign o[11999] = i[11999];
  assign o[11998] = i[11998];
  assign o[11997] = i[11997];
  assign o[11996] = i[11996];
  assign o[11995] = i[11995];
  assign o[11994] = i[11994];
  assign o[11993] = i[11993];
  assign o[11992] = i[11992];
  assign o[11991] = i[11991];
  assign o[11990] = i[11990];
  assign o[11989] = i[11989];
  assign o[11988] = i[11988];
  assign o[11987] = i[11987];
  assign o[11986] = i[11986];
  assign o[11985] = i[11985];
  assign o[11984] = i[11984];
  assign o[11983] = i[11983];
  assign o[11982] = i[11982];
  assign o[11981] = i[11981];
  assign o[11980] = i[11980];
  assign o[11979] = i[11979];
  assign o[11978] = i[11978];
  assign o[11977] = i[11977];
  assign o[11976] = i[11976];
  assign o[11975] = i[11975];
  assign o[11974] = i[11974];
  assign o[11973] = i[11973];
  assign o[11972] = i[11972];
  assign o[11971] = i[11971];
  assign o[11970] = i[11970];
  assign o[11969] = i[11969];
  assign o[11968] = i[11968];
  assign o[11967] = i[11967];
  assign o[11966] = i[11966];
  assign o[11965] = i[11965];
  assign o[11964] = i[11964];
  assign o[11963] = i[11963];
  assign o[11962] = i[11962];
  assign o[11961] = i[11961];
  assign o[11960] = i[11960];
  assign o[11959] = i[11959];
  assign o[11958] = i[11958];
  assign o[11957] = i[11957];
  assign o[11956] = i[11956];
  assign o[11955] = i[11955];
  assign o[11954] = i[11954];
  assign o[11953] = i[11953];
  assign o[11952] = i[11952];
  assign o[11951] = i[11951];
  assign o[11950] = i[11950];
  assign o[11949] = i[11949];
  assign o[11948] = i[11948];
  assign o[11947] = i[11947];
  assign o[11946] = i[11946];
  assign o[11945] = i[11945];
  assign o[11944] = i[11944];
  assign o[11943] = i[11943];
  assign o[11942] = i[11942];
  assign o[11941] = i[11941];
  assign o[11940] = i[11940];
  assign o[11939] = i[11939];
  assign o[11938] = i[11938];
  assign o[11937] = i[11937];
  assign o[11936] = i[11936];
  assign o[11935] = i[11935];
  assign o[11934] = i[11934];
  assign o[11933] = i[11933];
  assign o[11932] = i[11932];
  assign o[11931] = i[11931];
  assign o[11930] = i[11930];
  assign o[11929] = i[11929];
  assign o[11928] = i[11928];
  assign o[11927] = i[11927];
  assign o[11926] = i[11926];
  assign o[11925] = i[11925];
  assign o[11924] = i[11924];
  assign o[11923] = i[11923];
  assign o[11922] = i[11922];
  assign o[11921] = i[11921];
  assign o[11920] = i[11920];
  assign o[11919] = i[11919];
  assign o[11918] = i[11918];
  assign o[11917] = i[11917];
  assign o[11916] = i[11916];
  assign o[11915] = i[11915];
  assign o[11914] = i[11914];
  assign o[11913] = i[11913];
  assign o[11912] = i[11912];
  assign o[11911] = i[11911];
  assign o[11910] = i[11910];
  assign o[11909] = i[11909];
  assign o[11908] = i[11908];
  assign o[11907] = i[11907];
  assign o[11906] = i[11906];
  assign o[11905] = i[11905];
  assign o[11904] = i[11904];
  assign o[11903] = i[11903];
  assign o[11902] = i[11902];
  assign o[11901] = i[11901];
  assign o[11900] = i[11900];
  assign o[11899] = i[11899];
  assign o[11898] = i[11898];
  assign o[11897] = i[11897];
  assign o[11896] = i[11896];
  assign o[11895] = i[11895];
  assign o[11894] = i[11894];
  assign o[11893] = i[11893];
  assign o[11892] = i[11892];
  assign o[11891] = i[11891];
  assign o[11890] = i[11890];
  assign o[11889] = i[11889];
  assign o[11888] = i[11888];
  assign o[11887] = i[11887];
  assign o[11886] = i[11886];
  assign o[11885] = i[11885];
  assign o[11884] = i[11884];
  assign o[11883] = i[11883];
  assign o[11882] = i[11882];
  assign o[11881] = i[11881];
  assign o[11880] = i[11880];
  assign o[11879] = i[11879];
  assign o[11878] = i[11878];
  assign o[11877] = i[11877];
  assign o[11876] = i[11876];
  assign o[11875] = i[11875];
  assign o[11874] = i[11874];
  assign o[11873] = i[11873];
  assign o[11872] = i[11872];
  assign o[11871] = i[11871];
  assign o[11870] = i[11870];
  assign o[11869] = i[11869];
  assign o[11868] = i[11868];
  assign o[11867] = i[11867];
  assign o[11866] = i[11866];
  assign o[11865] = i[11865];
  assign o[11864] = i[11864];
  assign o[11863] = i[11863];
  assign o[11862] = i[11862];
  assign o[11861] = i[11861];
  assign o[11860] = i[11860];
  assign o[11859] = i[11859];
  assign o[11858] = i[11858];
  assign o[11857] = i[11857];
  assign o[11856] = i[11856];
  assign o[11855] = i[11855];
  assign o[11854] = i[11854];
  assign o[11853] = i[11853];
  assign o[11852] = i[11852];
  assign o[11851] = i[11851];
  assign o[11850] = i[11850];
  assign o[11849] = i[11849];
  assign o[11848] = i[11848];
  assign o[11847] = i[11847];
  assign o[11846] = i[11846];
  assign o[11845] = i[11845];
  assign o[11844] = i[11844];
  assign o[11843] = i[11843];
  assign o[11842] = i[11842];
  assign o[11841] = i[11841];
  assign o[11840] = i[11840];
  assign o[11839] = i[11839];
  assign o[11838] = i[11838];
  assign o[11837] = i[11837];
  assign o[11836] = i[11836];
  assign o[11835] = i[11835];
  assign o[11834] = i[11834];
  assign o[11833] = i[11833];
  assign o[11832] = i[11832];
  assign o[11831] = i[11831];
  assign o[11830] = i[11830];
  assign o[11829] = i[11829];
  assign o[11828] = i[11828];
  assign o[11827] = i[11827];
  assign o[11826] = i[11826];
  assign o[11825] = i[11825];
  assign o[11824] = i[11824];
  assign o[11823] = i[11823];
  assign o[11822] = i[11822];
  assign o[11821] = i[11821];
  assign o[11820] = i[11820];
  assign o[11819] = i[11819];
  assign o[11818] = i[11818];
  assign o[11817] = i[11817];
  assign o[11816] = i[11816];
  assign o[11815] = i[11815];
  assign o[11814] = i[11814];
  assign o[11813] = i[11813];
  assign o[11812] = i[11812];
  assign o[11811] = i[11811];
  assign o[11810] = i[11810];
  assign o[11809] = i[11809];
  assign o[11808] = i[11808];
  assign o[11807] = i[11807];
  assign o[11806] = i[11806];
  assign o[11805] = i[11805];
  assign o[11804] = i[11804];
  assign o[11803] = i[11803];
  assign o[11802] = i[11802];
  assign o[11801] = i[11801];
  assign o[11800] = i[11800];
  assign o[11799] = i[11799];
  assign o[11798] = i[11798];
  assign o[11797] = i[11797];
  assign o[11796] = i[11796];
  assign o[11795] = i[11795];
  assign o[11794] = i[11794];
  assign o[11793] = i[11793];
  assign o[11792] = i[11792];
  assign o[11791] = i[11791];
  assign o[11790] = i[11790];
  assign o[11789] = i[11789];
  assign o[11788] = i[11788];
  assign o[11787] = i[11787];
  assign o[11786] = i[11786];
  assign o[11785] = i[11785];
  assign o[11784] = i[11784];
  assign o[11783] = i[11783];
  assign o[11782] = i[11782];
  assign o[11781] = i[11781];
  assign o[11780] = i[11780];
  assign o[11779] = i[11779];
  assign o[11778] = i[11778];
  assign o[11777] = i[11777];
  assign o[11776] = i[11776];
  assign o[11775] = i[11775];
  assign o[11774] = i[11774];
  assign o[11773] = i[11773];
  assign o[11772] = i[11772];
  assign o[11771] = i[11771];
  assign o[11770] = i[11770];
  assign o[11769] = i[11769];
  assign o[11768] = i[11768];
  assign o[11767] = i[11767];
  assign o[11766] = i[11766];
  assign o[11765] = i[11765];
  assign o[11764] = i[11764];
  assign o[11763] = i[11763];
  assign o[11762] = i[11762];
  assign o[11761] = i[11761];
  assign o[11760] = i[11760];
  assign o[11759] = i[11759];
  assign o[11758] = i[11758];
  assign o[11757] = i[11757];
  assign o[11756] = i[11756];
  assign o[11755] = i[11755];
  assign o[11754] = i[11754];
  assign o[11753] = i[11753];
  assign o[11752] = i[11752];
  assign o[11751] = i[11751];
  assign o[11750] = i[11750];
  assign o[11749] = i[11749];
  assign o[11748] = i[11748];
  assign o[11747] = i[11747];
  assign o[11746] = i[11746];
  assign o[11745] = i[11745];
  assign o[11744] = i[11744];
  assign o[11743] = i[11743];
  assign o[11742] = i[11742];
  assign o[11741] = i[11741];
  assign o[11740] = i[11740];
  assign o[11739] = i[11739];
  assign o[11738] = i[11738];
  assign o[11737] = i[11737];
  assign o[11736] = i[11736];
  assign o[11735] = i[11735];
  assign o[11734] = i[11734];
  assign o[11733] = i[11733];
  assign o[11732] = i[11732];
  assign o[11731] = i[11731];
  assign o[11730] = i[11730];
  assign o[11729] = i[11729];
  assign o[11728] = i[11728];
  assign o[11727] = i[11727];
  assign o[11726] = i[11726];
  assign o[11725] = i[11725];
  assign o[11724] = i[11724];
  assign o[11723] = i[11723];
  assign o[11722] = i[11722];
  assign o[11721] = i[11721];
  assign o[11720] = i[11720];
  assign o[11719] = i[11719];
  assign o[11718] = i[11718];
  assign o[11717] = i[11717];
  assign o[11716] = i[11716];
  assign o[11715] = i[11715];
  assign o[11714] = i[11714];
  assign o[11713] = i[11713];
  assign o[11712] = i[11712];
  assign o[11711] = i[11711];
  assign o[11710] = i[11710];
  assign o[11709] = i[11709];
  assign o[11708] = i[11708];
  assign o[11707] = i[11707];
  assign o[11706] = i[11706];
  assign o[11705] = i[11705];
  assign o[11704] = i[11704];
  assign o[11703] = i[11703];
  assign o[11702] = i[11702];
  assign o[11701] = i[11701];
  assign o[11700] = i[11700];
  assign o[11699] = i[11699];
  assign o[11698] = i[11698];
  assign o[11697] = i[11697];
  assign o[11696] = i[11696];
  assign o[11695] = i[11695];
  assign o[11694] = i[11694];
  assign o[11693] = i[11693];
  assign o[11692] = i[11692];
  assign o[11691] = i[11691];
  assign o[11690] = i[11690];
  assign o[11689] = i[11689];
  assign o[11688] = i[11688];
  assign o[11687] = i[11687];
  assign o[11686] = i[11686];
  assign o[11685] = i[11685];
  assign o[11684] = i[11684];
  assign o[11683] = i[11683];
  assign o[11682] = i[11682];
  assign o[11681] = i[11681];
  assign o[11680] = i[11680];
  assign o[11679] = i[11679];
  assign o[11678] = i[11678];
  assign o[11677] = i[11677];
  assign o[11676] = i[11676];
  assign o[11675] = i[11675];
  assign o[11674] = i[11674];
  assign o[11673] = i[11673];
  assign o[11672] = i[11672];
  assign o[11671] = i[11671];
  assign o[11670] = i[11670];
  assign o[11669] = i[11669];
  assign o[11668] = i[11668];
  assign o[11667] = i[11667];
  assign o[11666] = i[11666];
  assign o[11665] = i[11665];
  assign o[11664] = i[11664];
  assign o[11663] = i[11663];
  assign o[11662] = i[11662];
  assign o[11661] = i[11661];
  assign o[11660] = i[11660];
  assign o[11659] = i[11659];
  assign o[11658] = i[11658];
  assign o[11657] = i[11657];
  assign o[11656] = i[11656];
  assign o[11655] = i[11655];
  assign o[11654] = i[11654];
  assign o[11653] = i[11653];
  assign o[11652] = i[11652];
  assign o[11651] = i[11651];
  assign o[11650] = i[11650];
  assign o[11649] = i[11649];
  assign o[11648] = i[11648];
  assign o[11647] = i[11647];
  assign o[11646] = i[11646];
  assign o[11645] = i[11645];
  assign o[11644] = i[11644];
  assign o[11643] = i[11643];
  assign o[11642] = i[11642];
  assign o[11641] = i[11641];
  assign o[11640] = i[11640];
  assign o[11639] = i[11639];
  assign o[11638] = i[11638];
  assign o[11637] = i[11637];
  assign o[11636] = i[11636];
  assign o[11635] = i[11635];
  assign o[11634] = i[11634];
  assign o[11633] = i[11633];
  assign o[11632] = i[11632];
  assign o[11631] = i[11631];
  assign o[11630] = i[11630];
  assign o[11629] = i[11629];
  assign o[11628] = i[11628];
  assign o[11627] = i[11627];
  assign o[11626] = i[11626];
  assign o[11625] = i[11625];
  assign o[11624] = i[11624];
  assign o[11623] = i[11623];
  assign o[11622] = i[11622];
  assign o[11621] = i[11621];
  assign o[11620] = i[11620];
  assign o[11619] = i[11619];
  assign o[11618] = i[11618];
  assign o[11617] = i[11617];
  assign o[11616] = i[11616];
  assign o[11615] = i[11615];
  assign o[11614] = i[11614];
  assign o[11613] = i[11613];
  assign o[11612] = i[11612];
  assign o[11611] = i[11611];
  assign o[11610] = i[11610];
  assign o[11609] = i[11609];
  assign o[11608] = i[11608];
  assign o[11607] = i[11607];
  assign o[11606] = i[11606];
  assign o[11605] = i[11605];
  assign o[11604] = i[11604];
  assign o[11603] = i[11603];
  assign o[11602] = i[11602];
  assign o[11601] = i[11601];
  assign o[11600] = i[11600];
  assign o[11599] = i[11599];
  assign o[11598] = i[11598];
  assign o[11597] = i[11597];
  assign o[11596] = i[11596];
  assign o[11595] = i[11595];
  assign o[11594] = i[11594];
  assign o[11593] = i[11593];
  assign o[11592] = i[11592];
  assign o[11591] = i[11591];
  assign o[11590] = i[11590];
  assign o[11589] = i[11589];
  assign o[11588] = i[11588];
  assign o[11587] = i[11587];
  assign o[11586] = i[11586];
  assign o[11585] = i[11585];
  assign o[11584] = i[11584];
  assign o[11583] = i[11583];
  assign o[11582] = i[11582];
  assign o[11581] = i[11581];
  assign o[11580] = i[11580];
  assign o[11579] = i[11579];
  assign o[11578] = i[11578];
  assign o[11577] = i[11577];
  assign o[11576] = i[11576];
  assign o[11575] = i[11575];
  assign o[11574] = i[11574];
  assign o[11573] = i[11573];
  assign o[11572] = i[11572];
  assign o[11571] = i[11571];
  assign o[11570] = i[11570];
  assign o[11569] = i[11569];
  assign o[11568] = i[11568];
  assign o[11567] = i[11567];
  assign o[11566] = i[11566];
  assign o[11565] = i[11565];
  assign o[11564] = i[11564];
  assign o[11563] = i[11563];
  assign o[11562] = i[11562];
  assign o[11561] = i[11561];
  assign o[11560] = i[11560];
  assign o[11559] = i[11559];
  assign o[11558] = i[11558];
  assign o[11557] = i[11557];
  assign o[11556] = i[11556];
  assign o[11555] = i[11555];
  assign o[11554] = i[11554];
  assign o[11553] = i[11553];
  assign o[11552] = i[11552];
  assign o[11551] = i[11551];
  assign o[11550] = i[11550];
  assign o[11549] = i[11549];
  assign o[11548] = i[11548];
  assign o[11547] = i[11547];
  assign o[11546] = i[11546];
  assign o[11545] = i[11545];
  assign o[11544] = i[11544];
  assign o[11543] = i[11543];
  assign o[11542] = i[11542];
  assign o[11541] = i[11541];
  assign o[11540] = i[11540];
  assign o[11539] = i[11539];
  assign o[11538] = i[11538];
  assign o[11537] = i[11537];
  assign o[11536] = i[11536];
  assign o[11535] = i[11535];
  assign o[11534] = i[11534];
  assign o[11533] = i[11533];
  assign o[11532] = i[11532];
  assign o[11531] = i[11531];
  assign o[11530] = i[11530];
  assign o[11529] = i[11529];
  assign o[11528] = i[11528];
  assign o[11527] = i[11527];
  assign o[11526] = i[11526];
  assign o[11525] = i[11525];
  assign o[11524] = i[11524];
  assign o[11523] = i[11523];
  assign o[11522] = i[11522];
  assign o[11521] = i[11521];
  assign o[11520] = i[11520];
  assign o[11519] = i[11519];
  assign o[11518] = i[11518];
  assign o[11517] = i[11517];
  assign o[11516] = i[11516];
  assign o[11515] = i[11515];
  assign o[11514] = i[11514];
  assign o[11513] = i[11513];
  assign o[11512] = i[11512];
  assign o[11511] = i[11511];
  assign o[11510] = i[11510];
  assign o[11509] = i[11509];
  assign o[11508] = i[11508];
  assign o[11507] = i[11507];
  assign o[11506] = i[11506];
  assign o[11505] = i[11505];
  assign o[11504] = i[11504];
  assign o[11503] = i[11503];
  assign o[11502] = i[11502];
  assign o[11501] = i[11501];
  assign o[11500] = i[11500];
  assign o[11499] = i[11499];
  assign o[11498] = i[11498];
  assign o[11497] = i[11497];
  assign o[11496] = i[11496];
  assign o[11495] = i[11495];
  assign o[11494] = i[11494];
  assign o[11493] = i[11493];
  assign o[11492] = i[11492];
  assign o[11491] = i[11491];
  assign o[11490] = i[11490];
  assign o[11489] = i[11489];
  assign o[11488] = i[11488];
  assign o[11487] = i[11487];
  assign o[11486] = i[11486];
  assign o[11485] = i[11485];
  assign o[11484] = i[11484];
  assign o[11483] = i[11483];
  assign o[11482] = i[11482];
  assign o[11481] = i[11481];
  assign o[11480] = i[11480];
  assign o[11479] = i[11479];
  assign o[11478] = i[11478];
  assign o[11477] = i[11477];
  assign o[11476] = i[11476];
  assign o[11475] = i[11475];
  assign o[11474] = i[11474];
  assign o[11473] = i[11473];
  assign o[11472] = i[11472];
  assign o[11471] = i[11471];
  assign o[11470] = i[11470];
  assign o[11469] = i[11469];
  assign o[11468] = i[11468];
  assign o[11467] = i[11467];
  assign o[11466] = i[11466];
  assign o[11465] = i[11465];
  assign o[11464] = i[11464];
  assign o[11463] = i[11463];
  assign o[11462] = i[11462];
  assign o[11461] = i[11461];
  assign o[11460] = i[11460];
  assign o[11459] = i[11459];
  assign o[11458] = i[11458];
  assign o[11457] = i[11457];
  assign o[11456] = i[11456];
  assign o[11455] = i[11455];
  assign o[11454] = i[11454];
  assign o[11453] = i[11453];
  assign o[11452] = i[11452];
  assign o[11451] = i[11451];
  assign o[11450] = i[11450];
  assign o[11449] = i[11449];
  assign o[11448] = i[11448];
  assign o[11447] = i[11447];
  assign o[11446] = i[11446];
  assign o[11445] = i[11445];
  assign o[11444] = i[11444];
  assign o[11443] = i[11443];
  assign o[11442] = i[11442];
  assign o[11441] = i[11441];
  assign o[11440] = i[11440];
  assign o[11439] = i[11439];
  assign o[11438] = i[11438];
  assign o[11437] = i[11437];
  assign o[11436] = i[11436];
  assign o[11435] = i[11435];
  assign o[11434] = i[11434];
  assign o[11433] = i[11433];
  assign o[11432] = i[11432];
  assign o[11431] = i[11431];
  assign o[11430] = i[11430];
  assign o[11429] = i[11429];
  assign o[11428] = i[11428];
  assign o[11427] = i[11427];
  assign o[11426] = i[11426];
  assign o[11425] = i[11425];
  assign o[11424] = i[11424];
  assign o[11423] = i[11423];
  assign o[11422] = i[11422];
  assign o[11421] = i[11421];
  assign o[11420] = i[11420];
  assign o[11419] = i[11419];
  assign o[11418] = i[11418];
  assign o[11417] = i[11417];
  assign o[11416] = i[11416];
  assign o[11415] = i[11415];
  assign o[11414] = i[11414];
  assign o[11413] = i[11413];
  assign o[11412] = i[11412];
  assign o[11411] = i[11411];
  assign o[11410] = i[11410];
  assign o[11409] = i[11409];
  assign o[11408] = i[11408];
  assign o[11407] = i[11407];
  assign o[11406] = i[11406];
  assign o[11405] = i[11405];
  assign o[11404] = i[11404];
  assign o[11403] = i[11403];
  assign o[11402] = i[11402];
  assign o[11401] = i[11401];
  assign o[11400] = i[11400];
  assign o[11399] = i[11399];
  assign o[11398] = i[11398];
  assign o[11397] = i[11397];
  assign o[11396] = i[11396];
  assign o[11395] = i[11395];
  assign o[11394] = i[11394];
  assign o[11393] = i[11393];
  assign o[11392] = i[11392];
  assign o[11391] = i[11391];
  assign o[11390] = i[11390];
  assign o[11389] = i[11389];
  assign o[11388] = i[11388];
  assign o[11387] = i[11387];
  assign o[11386] = i[11386];
  assign o[11385] = i[11385];
  assign o[11384] = i[11384];
  assign o[11383] = i[11383];
  assign o[11382] = i[11382];
  assign o[11381] = i[11381];
  assign o[11380] = i[11380];
  assign o[11379] = i[11379];
  assign o[11378] = i[11378];
  assign o[11377] = i[11377];
  assign o[11376] = i[11376];
  assign o[11375] = i[11375];
  assign o[11374] = i[11374];
  assign o[11373] = i[11373];
  assign o[11372] = i[11372];
  assign o[11371] = i[11371];
  assign o[11370] = i[11370];
  assign o[11369] = i[11369];
  assign o[11368] = i[11368];
  assign o[11367] = i[11367];
  assign o[11366] = i[11366];
  assign o[11365] = i[11365];
  assign o[11364] = i[11364];
  assign o[11363] = i[11363];
  assign o[11362] = i[11362];
  assign o[11361] = i[11361];
  assign o[11360] = i[11360];
  assign o[11359] = i[11359];
  assign o[11358] = i[11358];
  assign o[11357] = i[11357];
  assign o[11356] = i[11356];
  assign o[11355] = i[11355];
  assign o[11354] = i[11354];
  assign o[11353] = i[11353];
  assign o[11352] = i[11352];
  assign o[11351] = i[11351];
  assign o[11350] = i[11350];
  assign o[11349] = i[11349];
  assign o[11348] = i[11348];
  assign o[11347] = i[11347];
  assign o[11346] = i[11346];
  assign o[11345] = i[11345];
  assign o[11344] = i[11344];
  assign o[11343] = i[11343];
  assign o[11342] = i[11342];
  assign o[11341] = i[11341];
  assign o[11340] = i[11340];
  assign o[11339] = i[11339];
  assign o[11338] = i[11338];
  assign o[11337] = i[11337];
  assign o[11336] = i[11336];
  assign o[11335] = i[11335];
  assign o[11334] = i[11334];
  assign o[11333] = i[11333];
  assign o[11332] = i[11332];
  assign o[11331] = i[11331];
  assign o[11330] = i[11330];
  assign o[11329] = i[11329];
  assign o[11328] = i[11328];
  assign o[11327] = i[11327];
  assign o[11326] = i[11326];
  assign o[11325] = i[11325];
  assign o[11324] = i[11324];
  assign o[11323] = i[11323];
  assign o[11322] = i[11322];
  assign o[11321] = i[11321];
  assign o[11320] = i[11320];
  assign o[11319] = i[11319];
  assign o[11318] = i[11318];
  assign o[11317] = i[11317];
  assign o[11316] = i[11316];
  assign o[11315] = i[11315];
  assign o[11314] = i[11314];
  assign o[11313] = i[11313];
  assign o[11312] = i[11312];
  assign o[11311] = i[11311];
  assign o[11310] = i[11310];
  assign o[11309] = i[11309];
  assign o[11308] = i[11308];
  assign o[11307] = i[11307];
  assign o[11306] = i[11306];
  assign o[11305] = i[11305];
  assign o[11304] = i[11304];
  assign o[11303] = i[11303];
  assign o[11302] = i[11302];
  assign o[11301] = i[11301];
  assign o[11300] = i[11300];
  assign o[11299] = i[11299];
  assign o[11298] = i[11298];
  assign o[11297] = i[11297];
  assign o[11296] = i[11296];
  assign o[11295] = i[11295];
  assign o[11294] = i[11294];
  assign o[11293] = i[11293];
  assign o[11292] = i[11292];
  assign o[11291] = i[11291];
  assign o[11290] = i[11290];
  assign o[11289] = i[11289];
  assign o[11288] = i[11288];
  assign o[11287] = i[11287];
  assign o[11286] = i[11286];
  assign o[11285] = i[11285];
  assign o[11284] = i[11284];
  assign o[11283] = i[11283];
  assign o[11282] = i[11282];
  assign o[11281] = i[11281];
  assign o[11280] = i[11280];
  assign o[11279] = i[11279];
  assign o[11278] = i[11278];
  assign o[11277] = i[11277];
  assign o[11276] = i[11276];
  assign o[11275] = i[11275];
  assign o[11274] = i[11274];
  assign o[11273] = i[11273];
  assign o[11272] = i[11272];
  assign o[11271] = i[11271];
  assign o[11270] = i[11270];
  assign o[11269] = i[11269];
  assign o[11268] = i[11268];
  assign o[11267] = i[11267];
  assign o[11266] = i[11266];
  assign o[11265] = i[11265];
  assign o[11264] = i[11264];
  assign o[11263] = i[11263];
  assign o[11262] = i[11262];
  assign o[11261] = i[11261];
  assign o[11260] = i[11260];
  assign o[11259] = i[11259];
  assign o[11258] = i[11258];
  assign o[11257] = i[11257];
  assign o[11256] = i[11256];
  assign o[11255] = i[11255];
  assign o[11254] = i[11254];
  assign o[11253] = i[11253];
  assign o[11252] = i[11252];
  assign o[11251] = i[11251];
  assign o[11250] = i[11250];
  assign o[11249] = i[11249];
  assign o[11248] = i[11248];
  assign o[11247] = i[11247];
  assign o[11246] = i[11246];
  assign o[11245] = i[11245];
  assign o[11244] = i[11244];
  assign o[11243] = i[11243];
  assign o[11242] = i[11242];
  assign o[11241] = i[11241];
  assign o[11240] = i[11240];
  assign o[11239] = i[11239];
  assign o[11238] = i[11238];
  assign o[11237] = i[11237];
  assign o[11236] = i[11236];
  assign o[11235] = i[11235];
  assign o[11234] = i[11234];
  assign o[11233] = i[11233];
  assign o[11232] = i[11232];
  assign o[11231] = i[11231];
  assign o[11230] = i[11230];
  assign o[11229] = i[11229];
  assign o[11228] = i[11228];
  assign o[11227] = i[11227];
  assign o[11226] = i[11226];
  assign o[11225] = i[11225];
  assign o[11224] = i[11224];
  assign o[11223] = i[11223];
  assign o[11222] = i[11222];
  assign o[11221] = i[11221];
  assign o[11220] = i[11220];
  assign o[11219] = i[11219];
  assign o[11218] = i[11218];
  assign o[11217] = i[11217];
  assign o[11216] = i[11216];
  assign o[11215] = i[11215];
  assign o[11214] = i[11214];
  assign o[11213] = i[11213];
  assign o[11212] = i[11212];
  assign o[11211] = i[11211];
  assign o[11210] = i[11210];
  assign o[11209] = i[11209];
  assign o[11208] = i[11208];
  assign o[11207] = i[11207];
  assign o[11206] = i[11206];
  assign o[11205] = i[11205];
  assign o[11204] = i[11204];
  assign o[11203] = i[11203];
  assign o[11202] = i[11202];
  assign o[11201] = i[11201];
  assign o[11200] = i[11200];
  assign o[11199] = i[11199];
  assign o[11198] = i[11198];
  assign o[11197] = i[11197];
  assign o[11196] = i[11196];
  assign o[11195] = i[11195];
  assign o[11194] = i[11194];
  assign o[11193] = i[11193];
  assign o[11192] = i[11192];
  assign o[11191] = i[11191];
  assign o[11190] = i[11190];
  assign o[11189] = i[11189];
  assign o[11188] = i[11188];
  assign o[11187] = i[11187];
  assign o[11186] = i[11186];
  assign o[11185] = i[11185];
  assign o[11184] = i[11184];
  assign o[11183] = i[11183];
  assign o[11182] = i[11182];
  assign o[11181] = i[11181];
  assign o[11180] = i[11180];
  assign o[11179] = i[11179];
  assign o[11178] = i[11178];
  assign o[11177] = i[11177];
  assign o[11176] = i[11176];
  assign o[11175] = i[11175];
  assign o[11174] = i[11174];
  assign o[11173] = i[11173];
  assign o[11172] = i[11172];
  assign o[11171] = i[11171];
  assign o[11170] = i[11170];
  assign o[11169] = i[11169];
  assign o[11168] = i[11168];
  assign o[11167] = i[11167];
  assign o[11166] = i[11166];
  assign o[11165] = i[11165];
  assign o[11164] = i[11164];
  assign o[11163] = i[11163];
  assign o[11162] = i[11162];
  assign o[11161] = i[11161];
  assign o[11160] = i[11160];
  assign o[11159] = i[11159];
  assign o[11158] = i[11158];
  assign o[11157] = i[11157];
  assign o[11156] = i[11156];
  assign o[11155] = i[11155];
  assign o[11154] = i[11154];
  assign o[11153] = i[11153];
  assign o[11152] = i[11152];
  assign o[11151] = i[11151];
  assign o[11150] = i[11150];
  assign o[11149] = i[11149];
  assign o[11148] = i[11148];
  assign o[11147] = i[11147];
  assign o[11146] = i[11146];
  assign o[11145] = i[11145];
  assign o[11144] = i[11144];
  assign o[11143] = i[11143];
  assign o[11142] = i[11142];
  assign o[11141] = i[11141];
  assign o[11140] = i[11140];
  assign o[11139] = i[11139];
  assign o[11138] = i[11138];
  assign o[11137] = i[11137];
  assign o[11136] = i[11136];
  assign o[11135] = i[11135];
  assign o[11134] = i[11134];
  assign o[11133] = i[11133];
  assign o[11132] = i[11132];
  assign o[11131] = i[11131];
  assign o[11130] = i[11130];
  assign o[11129] = i[11129];
  assign o[11128] = i[11128];
  assign o[11127] = i[11127];
  assign o[11126] = i[11126];
  assign o[11125] = i[11125];
  assign o[11124] = i[11124];
  assign o[11123] = i[11123];
  assign o[11122] = i[11122];
  assign o[11121] = i[11121];
  assign o[11120] = i[11120];
  assign o[11119] = i[11119];
  assign o[11118] = i[11118];
  assign o[11117] = i[11117];
  assign o[11116] = i[11116];
  assign o[11115] = i[11115];
  assign o[11114] = i[11114];
  assign o[11113] = i[11113];
  assign o[11112] = i[11112];
  assign o[11111] = i[11111];
  assign o[11110] = i[11110];
  assign o[11109] = i[11109];
  assign o[11108] = i[11108];
  assign o[11107] = i[11107];
  assign o[11106] = i[11106];
  assign o[11105] = i[11105];
  assign o[11104] = i[11104];
  assign o[11103] = i[11103];
  assign o[11102] = i[11102];
  assign o[11101] = i[11101];
  assign o[11100] = i[11100];
  assign o[11099] = i[11099];
  assign o[11098] = i[11098];
  assign o[11097] = i[11097];
  assign o[11096] = i[11096];
  assign o[11095] = i[11095];
  assign o[11094] = i[11094];
  assign o[11093] = i[11093];
  assign o[11092] = i[11092];
  assign o[11091] = i[11091];
  assign o[11090] = i[11090];
  assign o[11089] = i[11089];
  assign o[11088] = i[11088];
  assign o[11087] = i[11087];
  assign o[11086] = i[11086];
  assign o[11085] = i[11085];
  assign o[11084] = i[11084];
  assign o[11083] = i[11083];
  assign o[11082] = i[11082];
  assign o[11081] = i[11081];
  assign o[11080] = i[11080];
  assign o[11079] = i[11079];
  assign o[11078] = i[11078];
  assign o[11077] = i[11077];
  assign o[11076] = i[11076];
  assign o[11075] = i[11075];
  assign o[11074] = i[11074];
  assign o[11073] = i[11073];
  assign o[11072] = i[11072];
  assign o[11071] = i[11071];
  assign o[11070] = i[11070];
  assign o[11069] = i[11069];
  assign o[11068] = i[11068];
  assign o[11067] = i[11067];
  assign o[11066] = i[11066];
  assign o[11065] = i[11065];
  assign o[11064] = i[11064];
  assign o[11063] = i[11063];
  assign o[11062] = i[11062];
  assign o[11061] = i[11061];
  assign o[11060] = i[11060];
  assign o[11059] = i[11059];
  assign o[11058] = i[11058];
  assign o[11057] = i[11057];
  assign o[11056] = i[11056];
  assign o[11055] = i[11055];
  assign o[11054] = i[11054];
  assign o[11053] = i[11053];
  assign o[11052] = i[11052];
  assign o[11051] = i[11051];
  assign o[11050] = i[11050];
  assign o[11049] = i[11049];
  assign o[11048] = i[11048];
  assign o[11047] = i[11047];
  assign o[11046] = i[11046];
  assign o[11045] = i[11045];
  assign o[11044] = i[11044];
  assign o[11043] = i[11043];
  assign o[11042] = i[11042];
  assign o[11041] = i[11041];
  assign o[11040] = i[11040];
  assign o[11039] = i[11039];
  assign o[11038] = i[11038];
  assign o[11037] = i[11037];
  assign o[11036] = i[11036];
  assign o[11035] = i[11035];
  assign o[11034] = i[11034];
  assign o[11033] = i[11033];
  assign o[11032] = i[11032];
  assign o[11031] = i[11031];
  assign o[11030] = i[11030];
  assign o[11029] = i[11029];
  assign o[11028] = i[11028];
  assign o[11027] = i[11027];
  assign o[11026] = i[11026];
  assign o[11025] = i[11025];
  assign o[11024] = i[11024];
  assign o[11023] = i[11023];
  assign o[11022] = i[11022];
  assign o[11021] = i[11021];
  assign o[11020] = i[11020];
  assign o[11019] = i[11019];
  assign o[11018] = i[11018];
  assign o[11017] = i[11017];
  assign o[11016] = i[11016];
  assign o[11015] = i[11015];
  assign o[11014] = i[11014];
  assign o[11013] = i[11013];
  assign o[11012] = i[11012];
  assign o[11011] = i[11011];
  assign o[11010] = i[11010];
  assign o[11009] = i[11009];
  assign o[11008] = i[11008];
  assign o[11007] = i[11007];
  assign o[11006] = i[11006];
  assign o[11005] = i[11005];
  assign o[11004] = i[11004];
  assign o[11003] = i[11003];
  assign o[11002] = i[11002];
  assign o[11001] = i[11001];
  assign o[11000] = i[11000];
  assign o[10999] = i[10999];
  assign o[10998] = i[10998];
  assign o[10997] = i[10997];
  assign o[10996] = i[10996];
  assign o[10995] = i[10995];
  assign o[10994] = i[10994];
  assign o[10993] = i[10993];
  assign o[10992] = i[10992];
  assign o[10991] = i[10991];
  assign o[10990] = i[10990];
  assign o[10989] = i[10989];
  assign o[10988] = i[10988];
  assign o[10987] = i[10987];
  assign o[10986] = i[10986];
  assign o[10985] = i[10985];
  assign o[10984] = i[10984];
  assign o[10983] = i[10983];
  assign o[10982] = i[10982];
  assign o[10981] = i[10981];
  assign o[10980] = i[10980];
  assign o[10979] = i[10979];
  assign o[10978] = i[10978];
  assign o[10977] = i[10977];
  assign o[10976] = i[10976];
  assign o[10975] = i[10975];
  assign o[10974] = i[10974];
  assign o[10973] = i[10973];
  assign o[10972] = i[10972];
  assign o[10971] = i[10971];
  assign o[10970] = i[10970];
  assign o[10969] = i[10969];
  assign o[10968] = i[10968];
  assign o[10967] = i[10967];
  assign o[10966] = i[10966];
  assign o[10965] = i[10965];
  assign o[10964] = i[10964];
  assign o[10963] = i[10963];
  assign o[10962] = i[10962];
  assign o[10961] = i[10961];
  assign o[10960] = i[10960];
  assign o[10959] = i[10959];
  assign o[10958] = i[10958];
  assign o[10957] = i[10957];
  assign o[10956] = i[10956];
  assign o[10955] = i[10955];
  assign o[10954] = i[10954];
  assign o[10953] = i[10953];
  assign o[10952] = i[10952];
  assign o[10951] = i[10951];
  assign o[10950] = i[10950];
  assign o[10949] = i[10949];
  assign o[10948] = i[10948];
  assign o[10947] = i[10947];
  assign o[10946] = i[10946];
  assign o[10945] = i[10945];
  assign o[10944] = i[10944];
  assign o[10943] = i[10943];
  assign o[10942] = i[10942];
  assign o[10941] = i[10941];
  assign o[10940] = i[10940];
  assign o[10939] = i[10939];
  assign o[10938] = i[10938];
  assign o[10937] = i[10937];
  assign o[10936] = i[10936];
  assign o[10935] = i[10935];
  assign o[10934] = i[10934];
  assign o[10933] = i[10933];
  assign o[10932] = i[10932];
  assign o[10931] = i[10931];
  assign o[10930] = i[10930];
  assign o[10929] = i[10929];
  assign o[10928] = i[10928];
  assign o[10927] = i[10927];
  assign o[10926] = i[10926];
  assign o[10925] = i[10925];
  assign o[10924] = i[10924];
  assign o[10923] = i[10923];
  assign o[10922] = i[10922];
  assign o[10921] = i[10921];
  assign o[10920] = i[10920];
  assign o[10919] = i[10919];
  assign o[10918] = i[10918];
  assign o[10917] = i[10917];
  assign o[10916] = i[10916];
  assign o[10915] = i[10915];
  assign o[10914] = i[10914];
  assign o[10913] = i[10913];
  assign o[10912] = i[10912];
  assign o[10911] = i[10911];
  assign o[10910] = i[10910];
  assign o[10909] = i[10909];
  assign o[10908] = i[10908];
  assign o[10907] = i[10907];
  assign o[10906] = i[10906];
  assign o[10905] = i[10905];
  assign o[10904] = i[10904];
  assign o[10903] = i[10903];
  assign o[10902] = i[10902];
  assign o[10901] = i[10901];
  assign o[10900] = i[10900];
  assign o[10899] = i[10899];
  assign o[10898] = i[10898];
  assign o[10897] = i[10897];
  assign o[10896] = i[10896];
  assign o[10895] = i[10895];
  assign o[10894] = i[10894];
  assign o[10893] = i[10893];
  assign o[10892] = i[10892];
  assign o[10891] = i[10891];
  assign o[10890] = i[10890];
  assign o[10889] = i[10889];
  assign o[10888] = i[10888];
  assign o[10887] = i[10887];
  assign o[10886] = i[10886];
  assign o[10885] = i[10885];
  assign o[10884] = i[10884];
  assign o[10883] = i[10883];
  assign o[10882] = i[10882];
  assign o[10881] = i[10881];
  assign o[10880] = i[10880];
  assign o[10879] = i[10879];
  assign o[10878] = i[10878];
  assign o[10877] = i[10877];
  assign o[10876] = i[10876];
  assign o[10875] = i[10875];
  assign o[10874] = i[10874];
  assign o[10873] = i[10873];
  assign o[10872] = i[10872];
  assign o[10871] = i[10871];
  assign o[10870] = i[10870];
  assign o[10869] = i[10869];
  assign o[10868] = i[10868];
  assign o[10867] = i[10867];
  assign o[10866] = i[10866];
  assign o[10865] = i[10865];
  assign o[10864] = i[10864];
  assign o[10863] = i[10863];
  assign o[10862] = i[10862];
  assign o[10861] = i[10861];
  assign o[10860] = i[10860];
  assign o[10859] = i[10859];
  assign o[10858] = i[10858];
  assign o[10857] = i[10857];
  assign o[10856] = i[10856];
  assign o[10855] = i[10855];
  assign o[10854] = i[10854];
  assign o[10853] = i[10853];
  assign o[10852] = i[10852];
  assign o[10851] = i[10851];
  assign o[10850] = i[10850];
  assign o[10849] = i[10849];
  assign o[10848] = i[10848];
  assign o[10847] = i[10847];
  assign o[10846] = i[10846];
  assign o[10845] = i[10845];
  assign o[10844] = i[10844];
  assign o[10843] = i[10843];
  assign o[10842] = i[10842];
  assign o[10841] = i[10841];
  assign o[10840] = i[10840];
  assign o[10839] = i[10839];
  assign o[10838] = i[10838];
  assign o[10837] = i[10837];
  assign o[10836] = i[10836];
  assign o[10835] = i[10835];
  assign o[10834] = i[10834];
  assign o[10833] = i[10833];
  assign o[10832] = i[10832];
  assign o[10831] = i[10831];
  assign o[10830] = i[10830];
  assign o[10829] = i[10829];
  assign o[10828] = i[10828];
  assign o[10827] = i[10827];
  assign o[10826] = i[10826];
  assign o[10825] = i[10825];
  assign o[10824] = i[10824];
  assign o[10823] = i[10823];
  assign o[10822] = i[10822];
  assign o[10821] = i[10821];
  assign o[10820] = i[10820];
  assign o[10819] = i[10819];
  assign o[10818] = i[10818];
  assign o[10817] = i[10817];
  assign o[10816] = i[10816];
  assign o[10815] = i[10815];
  assign o[10814] = i[10814];
  assign o[10813] = i[10813];
  assign o[10812] = i[10812];
  assign o[10811] = i[10811];
  assign o[10810] = i[10810];
  assign o[10809] = i[10809];
  assign o[10808] = i[10808];
  assign o[10807] = i[10807];
  assign o[10806] = i[10806];
  assign o[10805] = i[10805];
  assign o[10804] = i[10804];
  assign o[10803] = i[10803];
  assign o[10802] = i[10802];
  assign o[10801] = i[10801];
  assign o[10800] = i[10800];
  assign o[10799] = i[10799];
  assign o[10798] = i[10798];
  assign o[10797] = i[10797];
  assign o[10796] = i[10796];
  assign o[10795] = i[10795];
  assign o[10794] = i[10794];
  assign o[10793] = i[10793];
  assign o[10792] = i[10792];
  assign o[10791] = i[10791];
  assign o[10790] = i[10790];
  assign o[10789] = i[10789];
  assign o[10788] = i[10788];
  assign o[10787] = i[10787];
  assign o[10786] = i[10786];
  assign o[10785] = i[10785];
  assign o[10784] = i[10784];
  assign o[10783] = i[10783];
  assign o[10782] = i[10782];
  assign o[10781] = i[10781];
  assign o[10780] = i[10780];
  assign o[10779] = i[10779];
  assign o[10778] = i[10778];
  assign o[10777] = i[10777];
  assign o[10776] = i[10776];
  assign o[10775] = i[10775];
  assign o[10774] = i[10774];
  assign o[10773] = i[10773];
  assign o[10772] = i[10772];
  assign o[10771] = i[10771];
  assign o[10770] = i[10770];
  assign o[10769] = i[10769];
  assign o[10768] = i[10768];
  assign o[10767] = i[10767];
  assign o[10766] = i[10766];
  assign o[10765] = i[10765];
  assign o[10764] = i[10764];
  assign o[10763] = i[10763];
  assign o[10762] = i[10762];
  assign o[10761] = i[10761];
  assign o[10760] = i[10760];
  assign o[10759] = i[10759];
  assign o[10758] = i[10758];
  assign o[10757] = i[10757];
  assign o[10756] = i[10756];
  assign o[10755] = i[10755];
  assign o[10754] = i[10754];
  assign o[10753] = i[10753];
  assign o[10752] = i[10752];
  assign o[10751] = i[10751];
  assign o[10750] = i[10750];
  assign o[10749] = i[10749];
  assign o[10748] = i[10748];
  assign o[10747] = i[10747];
  assign o[10746] = i[10746];
  assign o[10745] = i[10745];
  assign o[10744] = i[10744];
  assign o[10743] = i[10743];
  assign o[10742] = i[10742];
  assign o[10741] = i[10741];
  assign o[10740] = i[10740];
  assign o[10739] = i[10739];
  assign o[10738] = i[10738];
  assign o[10737] = i[10737];
  assign o[10736] = i[10736];
  assign o[10735] = i[10735];
  assign o[10734] = i[10734];
  assign o[10733] = i[10733];
  assign o[10732] = i[10732];
  assign o[10731] = i[10731];
  assign o[10730] = i[10730];
  assign o[10729] = i[10729];
  assign o[10728] = i[10728];
  assign o[10727] = i[10727];
  assign o[10726] = i[10726];
  assign o[10725] = i[10725];
  assign o[10724] = i[10724];
  assign o[10723] = i[10723];
  assign o[10722] = i[10722];
  assign o[10721] = i[10721];
  assign o[10720] = i[10720];
  assign o[10719] = i[10719];
  assign o[10718] = i[10718];
  assign o[10717] = i[10717];
  assign o[10716] = i[10716];
  assign o[10715] = i[10715];
  assign o[10714] = i[10714];
  assign o[10713] = i[10713];
  assign o[10712] = i[10712];
  assign o[10711] = i[10711];
  assign o[10710] = i[10710];
  assign o[10709] = i[10709];
  assign o[10708] = i[10708];
  assign o[10707] = i[10707];
  assign o[10706] = i[10706];
  assign o[10705] = i[10705];
  assign o[10704] = i[10704];
  assign o[10703] = i[10703];
  assign o[10702] = i[10702];
  assign o[10701] = i[10701];
  assign o[10700] = i[10700];
  assign o[10699] = i[10699];
  assign o[10698] = i[10698];
  assign o[10697] = i[10697];
  assign o[10696] = i[10696];
  assign o[10695] = i[10695];
  assign o[10694] = i[10694];
  assign o[10693] = i[10693];
  assign o[10692] = i[10692];
  assign o[10691] = i[10691];
  assign o[10690] = i[10690];
  assign o[10689] = i[10689];
  assign o[10688] = i[10688];
  assign o[10687] = i[10687];
  assign o[10686] = i[10686];
  assign o[10685] = i[10685];
  assign o[10684] = i[10684];
  assign o[10683] = i[10683];
  assign o[10682] = i[10682];
  assign o[10681] = i[10681];
  assign o[10680] = i[10680];
  assign o[10679] = i[10679];
  assign o[10678] = i[10678];
  assign o[10677] = i[10677];
  assign o[10676] = i[10676];
  assign o[10675] = i[10675];
  assign o[10674] = i[10674];
  assign o[10673] = i[10673];
  assign o[10672] = i[10672];
  assign o[10671] = i[10671];
  assign o[10670] = i[10670];
  assign o[10669] = i[10669];
  assign o[10668] = i[10668];
  assign o[10667] = i[10667];
  assign o[10666] = i[10666];
  assign o[10665] = i[10665];
  assign o[10664] = i[10664];
  assign o[10663] = i[10663];
  assign o[10662] = i[10662];
  assign o[10661] = i[10661];
  assign o[10660] = i[10660];
  assign o[10659] = i[10659];
  assign o[10658] = i[10658];
  assign o[10657] = i[10657];
  assign o[10656] = i[10656];
  assign o[10655] = i[10655];
  assign o[10654] = i[10654];
  assign o[10653] = i[10653];
  assign o[10652] = i[10652];
  assign o[10651] = i[10651];
  assign o[10650] = i[10650];
  assign o[10649] = i[10649];
  assign o[10648] = i[10648];
  assign o[10647] = i[10647];
  assign o[10646] = i[10646];
  assign o[10645] = i[10645];
  assign o[10644] = i[10644];
  assign o[10643] = i[10643];
  assign o[10642] = i[10642];
  assign o[10641] = i[10641];
  assign o[10640] = i[10640];
  assign o[10639] = i[10639];
  assign o[10638] = i[10638];
  assign o[10637] = i[10637];
  assign o[10636] = i[10636];
  assign o[10635] = i[10635];
  assign o[10634] = i[10634];
  assign o[10633] = i[10633];
  assign o[10632] = i[10632];
  assign o[10631] = i[10631];
  assign o[10630] = i[10630];
  assign o[10629] = i[10629];
  assign o[10628] = i[10628];
  assign o[10627] = i[10627];
  assign o[10626] = i[10626];
  assign o[10625] = i[10625];
  assign o[10624] = i[10624];
  assign o[10623] = i[10623];
  assign o[10622] = i[10622];
  assign o[10621] = i[10621];
  assign o[10620] = i[10620];
  assign o[10619] = i[10619];
  assign o[10618] = i[10618];
  assign o[10617] = i[10617];
  assign o[10616] = i[10616];
  assign o[10615] = i[10615];
  assign o[10614] = i[10614];
  assign o[10613] = i[10613];
  assign o[10612] = i[10612];
  assign o[10611] = i[10611];
  assign o[10610] = i[10610];
  assign o[10609] = i[10609];
  assign o[10608] = i[10608];
  assign o[10607] = i[10607];
  assign o[10606] = i[10606];
  assign o[10605] = i[10605];
  assign o[10604] = i[10604];
  assign o[10603] = i[10603];
  assign o[10602] = i[10602];
  assign o[10601] = i[10601];
  assign o[10600] = i[10600];
  assign o[10599] = i[10599];
  assign o[10598] = i[10598];
  assign o[10597] = i[10597];
  assign o[10596] = i[10596];
  assign o[10595] = i[10595];
  assign o[10594] = i[10594];
  assign o[10593] = i[10593];
  assign o[10592] = i[10592];
  assign o[10591] = i[10591];
  assign o[10590] = i[10590];
  assign o[10589] = i[10589];
  assign o[10588] = i[10588];
  assign o[10587] = i[10587];
  assign o[10586] = i[10586];
  assign o[10585] = i[10585];
  assign o[10584] = i[10584];
  assign o[10583] = i[10583];
  assign o[10582] = i[10582];
  assign o[10581] = i[10581];
  assign o[10580] = i[10580];
  assign o[10579] = i[10579];
  assign o[10578] = i[10578];
  assign o[10577] = i[10577];
  assign o[10576] = i[10576];
  assign o[10575] = i[10575];
  assign o[10574] = i[10574];
  assign o[10573] = i[10573];
  assign o[10572] = i[10572];
  assign o[10571] = i[10571];
  assign o[10570] = i[10570];
  assign o[10569] = i[10569];
  assign o[10568] = i[10568];
  assign o[10567] = i[10567];
  assign o[10566] = i[10566];
  assign o[10565] = i[10565];
  assign o[10564] = i[10564];
  assign o[10563] = i[10563];
  assign o[10562] = i[10562];
  assign o[10561] = i[10561];
  assign o[10560] = i[10560];
  assign o[10559] = i[10559];
  assign o[10558] = i[10558];
  assign o[10557] = i[10557];
  assign o[10556] = i[10556];
  assign o[10555] = i[10555];
  assign o[10554] = i[10554];
  assign o[10553] = i[10553];
  assign o[10552] = i[10552];
  assign o[10551] = i[10551];
  assign o[10550] = i[10550];
  assign o[10549] = i[10549];
  assign o[10548] = i[10548];
  assign o[10547] = i[10547];
  assign o[10546] = i[10546];
  assign o[10545] = i[10545];
  assign o[10544] = i[10544];
  assign o[10543] = i[10543];
  assign o[10542] = i[10542];
  assign o[10541] = i[10541];
  assign o[10540] = i[10540];
  assign o[10539] = i[10539];
  assign o[10538] = i[10538];
  assign o[10537] = i[10537];
  assign o[10536] = i[10536];
  assign o[10535] = i[10535];
  assign o[10534] = i[10534];
  assign o[10533] = i[10533];
  assign o[10532] = i[10532];
  assign o[10531] = i[10531];
  assign o[10530] = i[10530];
  assign o[10529] = i[10529];
  assign o[10528] = i[10528];
  assign o[10527] = i[10527];
  assign o[10526] = i[10526];
  assign o[10525] = i[10525];
  assign o[10524] = i[10524];
  assign o[10523] = i[10523];
  assign o[10522] = i[10522];
  assign o[10521] = i[10521];
  assign o[10520] = i[10520];
  assign o[10519] = i[10519];
  assign o[10518] = i[10518];
  assign o[10517] = i[10517];
  assign o[10516] = i[10516];
  assign o[10515] = i[10515];
  assign o[10514] = i[10514];
  assign o[10513] = i[10513];
  assign o[10512] = i[10512];
  assign o[10511] = i[10511];
  assign o[10510] = i[10510];
  assign o[10509] = i[10509];
  assign o[10508] = i[10508];
  assign o[10507] = i[10507];
  assign o[10506] = i[10506];
  assign o[10505] = i[10505];
  assign o[10504] = i[10504];
  assign o[10503] = i[10503];
  assign o[10502] = i[10502];
  assign o[10501] = i[10501];
  assign o[10500] = i[10500];
  assign o[10499] = i[10499];
  assign o[10498] = i[10498];
  assign o[10497] = i[10497];
  assign o[10496] = i[10496];
  assign o[10495] = i[10495];
  assign o[10494] = i[10494];
  assign o[10493] = i[10493];
  assign o[10492] = i[10492];
  assign o[10491] = i[10491];
  assign o[10490] = i[10490];
  assign o[10489] = i[10489];
  assign o[10488] = i[10488];
  assign o[10487] = i[10487];
  assign o[10486] = i[10486];
  assign o[10485] = i[10485];
  assign o[10484] = i[10484];
  assign o[10483] = i[10483];
  assign o[10482] = i[10482];
  assign o[10481] = i[10481];
  assign o[10480] = i[10480];
  assign o[10479] = i[10479];
  assign o[10478] = i[10478];
  assign o[10477] = i[10477];
  assign o[10476] = i[10476];
  assign o[10475] = i[10475];
  assign o[10474] = i[10474];
  assign o[10473] = i[10473];
  assign o[10472] = i[10472];
  assign o[10471] = i[10471];
  assign o[10470] = i[10470];
  assign o[10469] = i[10469];
  assign o[10468] = i[10468];
  assign o[10467] = i[10467];
  assign o[10466] = i[10466];
  assign o[10465] = i[10465];
  assign o[10464] = i[10464];
  assign o[10463] = i[10463];
  assign o[10462] = i[10462];
  assign o[10461] = i[10461];
  assign o[10460] = i[10460];
  assign o[10459] = i[10459];
  assign o[10458] = i[10458];
  assign o[10457] = i[10457];
  assign o[10456] = i[10456];
  assign o[10455] = i[10455];
  assign o[10454] = i[10454];
  assign o[10453] = i[10453];
  assign o[10452] = i[10452];
  assign o[10451] = i[10451];
  assign o[10450] = i[10450];
  assign o[10449] = i[10449];
  assign o[10448] = i[10448];
  assign o[10447] = i[10447];
  assign o[10446] = i[10446];
  assign o[10445] = i[10445];
  assign o[10444] = i[10444];
  assign o[10443] = i[10443];
  assign o[10442] = i[10442];
  assign o[10441] = i[10441];
  assign o[10440] = i[10440];
  assign o[10439] = i[10439];
  assign o[10438] = i[10438];
  assign o[10437] = i[10437];
  assign o[10436] = i[10436];
  assign o[10435] = i[10435];
  assign o[10434] = i[10434];
  assign o[10433] = i[10433];
  assign o[10432] = i[10432];
  assign o[10431] = i[10431];
  assign o[10430] = i[10430];
  assign o[10429] = i[10429];
  assign o[10428] = i[10428];
  assign o[10427] = i[10427];
  assign o[10426] = i[10426];
  assign o[10425] = i[10425];
  assign o[10424] = i[10424];
  assign o[10423] = i[10423];
  assign o[10422] = i[10422];
  assign o[10421] = i[10421];
  assign o[10420] = i[10420];
  assign o[10419] = i[10419];
  assign o[10418] = i[10418];
  assign o[10417] = i[10417];
  assign o[10416] = i[10416];
  assign o[10415] = i[10415];
  assign o[10414] = i[10414];
  assign o[10413] = i[10413];
  assign o[10412] = i[10412];
  assign o[10411] = i[10411];
  assign o[10410] = i[10410];
  assign o[10409] = i[10409];
  assign o[10408] = i[10408];
  assign o[10407] = i[10407];
  assign o[10406] = i[10406];
  assign o[10405] = i[10405];
  assign o[10404] = i[10404];
  assign o[10403] = i[10403];
  assign o[10402] = i[10402];
  assign o[10401] = i[10401];
  assign o[10400] = i[10400];
  assign o[10399] = i[10399];
  assign o[10398] = i[10398];
  assign o[10397] = i[10397];
  assign o[10396] = i[10396];
  assign o[10395] = i[10395];
  assign o[10394] = i[10394];
  assign o[10393] = i[10393];
  assign o[10392] = i[10392];
  assign o[10391] = i[10391];
  assign o[10390] = i[10390];
  assign o[10389] = i[10389];
  assign o[10388] = i[10388];
  assign o[10387] = i[10387];
  assign o[10386] = i[10386];
  assign o[10385] = i[10385];
  assign o[10384] = i[10384];
  assign o[10383] = i[10383];
  assign o[10382] = i[10382];
  assign o[10381] = i[10381];
  assign o[10380] = i[10380];
  assign o[10379] = i[10379];
  assign o[10378] = i[10378];
  assign o[10377] = i[10377];
  assign o[10376] = i[10376];
  assign o[10375] = i[10375];
  assign o[10374] = i[10374];
  assign o[10373] = i[10373];
  assign o[10372] = i[10372];
  assign o[10371] = i[10371];
  assign o[10370] = i[10370];
  assign o[10369] = i[10369];
  assign o[10368] = i[10368];
  assign o[10367] = i[10367];
  assign o[10366] = i[10366];
  assign o[10365] = i[10365];
  assign o[10364] = i[10364];
  assign o[10363] = i[10363];
  assign o[10362] = i[10362];
  assign o[10361] = i[10361];
  assign o[10360] = i[10360];
  assign o[10359] = i[10359];
  assign o[10358] = i[10358];
  assign o[10357] = i[10357];
  assign o[10356] = i[10356];
  assign o[10355] = i[10355];
  assign o[10354] = i[10354];
  assign o[10353] = i[10353];
  assign o[10352] = i[10352];
  assign o[10351] = i[10351];
  assign o[10350] = i[10350];
  assign o[10349] = i[10349];
  assign o[10348] = i[10348];
  assign o[10347] = i[10347];
  assign o[10346] = i[10346];
  assign o[10345] = i[10345];
  assign o[10344] = i[10344];
  assign o[10343] = i[10343];
  assign o[10342] = i[10342];
  assign o[10341] = i[10341];
  assign o[10340] = i[10340];
  assign o[10339] = i[10339];
  assign o[10338] = i[10338];
  assign o[10337] = i[10337];
  assign o[10336] = i[10336];
  assign o[10335] = i[10335];
  assign o[10334] = i[10334];
  assign o[10333] = i[10333];
  assign o[10332] = i[10332];
  assign o[10331] = i[10331];
  assign o[10330] = i[10330];
  assign o[10329] = i[10329];
  assign o[10328] = i[10328];
  assign o[10327] = i[10327];
  assign o[10326] = i[10326];
  assign o[10325] = i[10325];
  assign o[10324] = i[10324];
  assign o[10323] = i[10323];
  assign o[10322] = i[10322];
  assign o[10321] = i[10321];
  assign o[10320] = i[10320];
  assign o[10319] = i[10319];
  assign o[10318] = i[10318];
  assign o[10317] = i[10317];
  assign o[10316] = i[10316];
  assign o[10315] = i[10315];
  assign o[10314] = i[10314];
  assign o[10313] = i[10313];
  assign o[10312] = i[10312];
  assign o[10311] = i[10311];
  assign o[10310] = i[10310];
  assign o[10309] = i[10309];
  assign o[10308] = i[10308];
  assign o[10307] = i[10307];
  assign o[10306] = i[10306];
  assign o[10305] = i[10305];
  assign o[10304] = i[10304];
  assign o[10303] = i[10303];
  assign o[10302] = i[10302];
  assign o[10301] = i[10301];
  assign o[10300] = i[10300];
  assign o[10299] = i[10299];
  assign o[10298] = i[10298];
  assign o[10297] = i[10297];
  assign o[10296] = i[10296];
  assign o[10295] = i[10295];
  assign o[10294] = i[10294];
  assign o[10293] = i[10293];
  assign o[10292] = i[10292];
  assign o[10291] = i[10291];
  assign o[10290] = i[10290];
  assign o[10289] = i[10289];
  assign o[10288] = i[10288];
  assign o[10287] = i[10287];
  assign o[10286] = i[10286];
  assign o[10285] = i[10285];
  assign o[10284] = i[10284];
  assign o[10283] = i[10283];
  assign o[10282] = i[10282];
  assign o[10281] = i[10281];
  assign o[10280] = i[10280];
  assign o[10279] = i[10279];
  assign o[10278] = i[10278];
  assign o[10277] = i[10277];
  assign o[10276] = i[10276];
  assign o[10275] = i[10275];
  assign o[10274] = i[10274];
  assign o[10273] = i[10273];
  assign o[10272] = i[10272];
  assign o[10271] = i[10271];
  assign o[10270] = i[10270];
  assign o[10269] = i[10269];
  assign o[10268] = i[10268];
  assign o[10267] = i[10267];
  assign o[10266] = i[10266];
  assign o[10265] = i[10265];
  assign o[10264] = i[10264];
  assign o[10263] = i[10263];
  assign o[10262] = i[10262];
  assign o[10261] = i[10261];
  assign o[10260] = i[10260];
  assign o[10259] = i[10259];
  assign o[10258] = i[10258];
  assign o[10257] = i[10257];
  assign o[10256] = i[10256];
  assign o[10255] = i[10255];
  assign o[10254] = i[10254];
  assign o[10253] = i[10253];
  assign o[10252] = i[10252];
  assign o[10251] = i[10251];
  assign o[10250] = i[10250];
  assign o[10249] = i[10249];
  assign o[10248] = i[10248];
  assign o[10247] = i[10247];
  assign o[10246] = i[10246];
  assign o[10245] = i[10245];
  assign o[10244] = i[10244];
  assign o[10243] = i[10243];
  assign o[10242] = i[10242];
  assign o[10241] = i[10241];
  assign o[10240] = i[10240];
  assign o[10239] = i[10239];
  assign o[10238] = i[10238];
  assign o[10237] = i[10237];
  assign o[10236] = i[10236];
  assign o[10235] = i[10235];
  assign o[10234] = i[10234];
  assign o[10233] = i[10233];
  assign o[10232] = i[10232];
  assign o[10231] = i[10231];
  assign o[10230] = i[10230];
  assign o[10229] = i[10229];
  assign o[10228] = i[10228];
  assign o[10227] = i[10227];
  assign o[10226] = i[10226];
  assign o[10225] = i[10225];
  assign o[10224] = i[10224];
  assign o[10223] = i[10223];
  assign o[10222] = i[10222];
  assign o[10221] = i[10221];
  assign o[10220] = i[10220];
  assign o[10219] = i[10219];
  assign o[10218] = i[10218];
  assign o[10217] = i[10217];
  assign o[10216] = i[10216];
  assign o[10215] = i[10215];
  assign o[10214] = i[10214];
  assign o[10213] = i[10213];
  assign o[10212] = i[10212];
  assign o[10211] = i[10211];
  assign o[10210] = i[10210];
  assign o[10209] = i[10209];
  assign o[10208] = i[10208];
  assign o[10207] = i[10207];
  assign o[10206] = i[10206];
  assign o[10205] = i[10205];
  assign o[10204] = i[10204];
  assign o[10203] = i[10203];
  assign o[10202] = i[10202];
  assign o[10201] = i[10201];
  assign o[10200] = i[10200];
  assign o[10199] = i[10199];
  assign o[10198] = i[10198];
  assign o[10197] = i[10197];
  assign o[10196] = i[10196];
  assign o[10195] = i[10195];
  assign o[10194] = i[10194];
  assign o[10193] = i[10193];
  assign o[10192] = i[10192];
  assign o[10191] = i[10191];
  assign o[10190] = i[10190];
  assign o[10189] = i[10189];
  assign o[10188] = i[10188];
  assign o[10187] = i[10187];
  assign o[10186] = i[10186];
  assign o[10185] = i[10185];
  assign o[10184] = i[10184];
  assign o[10183] = i[10183];
  assign o[10182] = i[10182];
  assign o[10181] = i[10181];
  assign o[10180] = i[10180];
  assign o[10179] = i[10179];
  assign o[10178] = i[10178];
  assign o[10177] = i[10177];
  assign o[10176] = i[10176];
  assign o[10175] = i[10175];
  assign o[10174] = i[10174];
  assign o[10173] = i[10173];
  assign o[10172] = i[10172];
  assign o[10171] = i[10171];
  assign o[10170] = i[10170];
  assign o[10169] = i[10169];
  assign o[10168] = i[10168];
  assign o[10167] = i[10167];
  assign o[10166] = i[10166];
  assign o[10165] = i[10165];
  assign o[10164] = i[10164];
  assign o[10163] = i[10163];
  assign o[10162] = i[10162];
  assign o[10161] = i[10161];
  assign o[10160] = i[10160];
  assign o[10159] = i[10159];
  assign o[10158] = i[10158];
  assign o[10157] = i[10157];
  assign o[10156] = i[10156];
  assign o[10155] = i[10155];
  assign o[10154] = i[10154];
  assign o[10153] = i[10153];
  assign o[10152] = i[10152];
  assign o[10151] = i[10151];
  assign o[10150] = i[10150];
  assign o[10149] = i[10149];
  assign o[10148] = i[10148];
  assign o[10147] = i[10147];
  assign o[10146] = i[10146];
  assign o[10145] = i[10145];
  assign o[10144] = i[10144];
  assign o[10143] = i[10143];
  assign o[10142] = i[10142];
  assign o[10141] = i[10141];
  assign o[10140] = i[10140];
  assign o[10139] = i[10139];
  assign o[10138] = i[10138];
  assign o[10137] = i[10137];
  assign o[10136] = i[10136];
  assign o[10135] = i[10135];
  assign o[10134] = i[10134];
  assign o[10133] = i[10133];
  assign o[10132] = i[10132];
  assign o[10131] = i[10131];
  assign o[10130] = i[10130];
  assign o[10129] = i[10129];
  assign o[10128] = i[10128];
  assign o[10127] = i[10127];
  assign o[10126] = i[10126];
  assign o[10125] = i[10125];
  assign o[10124] = i[10124];
  assign o[10123] = i[10123];
  assign o[10122] = i[10122];
  assign o[10121] = i[10121];
  assign o[10120] = i[10120];
  assign o[10119] = i[10119];
  assign o[10118] = i[10118];
  assign o[10117] = i[10117];
  assign o[10116] = i[10116];
  assign o[10115] = i[10115];
  assign o[10114] = i[10114];
  assign o[10113] = i[10113];
  assign o[10112] = i[10112];
  assign o[10111] = i[10111];
  assign o[10110] = i[10110];
  assign o[10109] = i[10109];
  assign o[10108] = i[10108];
  assign o[10107] = i[10107];
  assign o[10106] = i[10106];
  assign o[10105] = i[10105];
  assign o[10104] = i[10104];
  assign o[10103] = i[10103];
  assign o[10102] = i[10102];
  assign o[10101] = i[10101];
  assign o[10100] = i[10100];
  assign o[10099] = i[10099];
  assign o[10098] = i[10098];
  assign o[10097] = i[10097];
  assign o[10096] = i[10096];
  assign o[10095] = i[10095];
  assign o[10094] = i[10094];
  assign o[10093] = i[10093];
  assign o[10092] = i[10092];
  assign o[10091] = i[10091];
  assign o[10090] = i[10090];
  assign o[10089] = i[10089];
  assign o[10088] = i[10088];
  assign o[10087] = i[10087];
  assign o[10086] = i[10086];
  assign o[10085] = i[10085];
  assign o[10084] = i[10084];
  assign o[10083] = i[10083];
  assign o[10082] = i[10082];
  assign o[10081] = i[10081];
  assign o[10080] = i[10080];
  assign o[10079] = i[10079];
  assign o[10078] = i[10078];
  assign o[10077] = i[10077];
  assign o[10076] = i[10076];
  assign o[10075] = i[10075];
  assign o[10074] = i[10074];
  assign o[10073] = i[10073];
  assign o[10072] = i[10072];
  assign o[10071] = i[10071];
  assign o[10070] = i[10070];
  assign o[10069] = i[10069];
  assign o[10068] = i[10068];
  assign o[10067] = i[10067];
  assign o[10066] = i[10066];
  assign o[10065] = i[10065];
  assign o[10064] = i[10064];
  assign o[10063] = i[10063];
  assign o[10062] = i[10062];
  assign o[10061] = i[10061];
  assign o[10060] = i[10060];
  assign o[10059] = i[10059];
  assign o[10058] = i[10058];
  assign o[10057] = i[10057];
  assign o[10056] = i[10056];
  assign o[10055] = i[10055];
  assign o[10054] = i[10054];
  assign o[10053] = i[10053];
  assign o[10052] = i[10052];
  assign o[10051] = i[10051];
  assign o[10050] = i[10050];
  assign o[10049] = i[10049];
  assign o[10048] = i[10048];
  assign o[10047] = i[10047];
  assign o[10046] = i[10046];
  assign o[10045] = i[10045];
  assign o[10044] = i[10044];
  assign o[10043] = i[10043];
  assign o[10042] = i[10042];
  assign o[10041] = i[10041];
  assign o[10040] = i[10040];
  assign o[10039] = i[10039];
  assign o[10038] = i[10038];
  assign o[10037] = i[10037];
  assign o[10036] = i[10036];
  assign o[10035] = i[10035];
  assign o[10034] = i[10034];
  assign o[10033] = i[10033];
  assign o[10032] = i[10032];
  assign o[10031] = i[10031];
  assign o[10030] = i[10030];
  assign o[10029] = i[10029];
  assign o[10028] = i[10028];
  assign o[10027] = i[10027];
  assign o[10026] = i[10026];
  assign o[10025] = i[10025];
  assign o[10024] = i[10024];
  assign o[10023] = i[10023];
  assign o[10022] = i[10022];
  assign o[10021] = i[10021];
  assign o[10020] = i[10020];
  assign o[10019] = i[10019];
  assign o[10018] = i[10018];
  assign o[10017] = i[10017];
  assign o[10016] = i[10016];
  assign o[10015] = i[10015];
  assign o[10014] = i[10014];
  assign o[10013] = i[10013];
  assign o[10012] = i[10012];
  assign o[10011] = i[10011];
  assign o[10010] = i[10010];
  assign o[10009] = i[10009];
  assign o[10008] = i[10008];
  assign o[10007] = i[10007];
  assign o[10006] = i[10006];
  assign o[10005] = i[10005];
  assign o[10004] = i[10004];
  assign o[10003] = i[10003];
  assign o[10002] = i[10002];
  assign o[10001] = i[10001];
  assign o[10000] = i[10000];
  assign o[9999] = i[9999];
  assign o[9998] = i[9998];
  assign o[9997] = i[9997];
  assign o[9996] = i[9996];
  assign o[9995] = i[9995];
  assign o[9994] = i[9994];
  assign o[9993] = i[9993];
  assign o[9992] = i[9992];
  assign o[9991] = i[9991];
  assign o[9990] = i[9990];
  assign o[9989] = i[9989];
  assign o[9988] = i[9988];
  assign o[9987] = i[9987];
  assign o[9986] = i[9986];
  assign o[9985] = i[9985];
  assign o[9984] = i[9984];
  assign o[9983] = i[9983];
  assign o[9982] = i[9982];
  assign o[9981] = i[9981];
  assign o[9980] = i[9980];
  assign o[9979] = i[9979];
  assign o[9978] = i[9978];
  assign o[9977] = i[9977];
  assign o[9976] = i[9976];
  assign o[9975] = i[9975];
  assign o[9974] = i[9974];
  assign o[9973] = i[9973];
  assign o[9972] = i[9972];
  assign o[9971] = i[9971];
  assign o[9970] = i[9970];
  assign o[9969] = i[9969];
  assign o[9968] = i[9968];
  assign o[9967] = i[9967];
  assign o[9966] = i[9966];
  assign o[9965] = i[9965];
  assign o[9964] = i[9964];
  assign o[9963] = i[9963];
  assign o[9962] = i[9962];
  assign o[9961] = i[9961];
  assign o[9960] = i[9960];
  assign o[9959] = i[9959];
  assign o[9958] = i[9958];
  assign o[9957] = i[9957];
  assign o[9956] = i[9956];
  assign o[9955] = i[9955];
  assign o[9954] = i[9954];
  assign o[9953] = i[9953];
  assign o[9952] = i[9952];
  assign o[9951] = i[9951];
  assign o[9950] = i[9950];
  assign o[9949] = i[9949];
  assign o[9948] = i[9948];
  assign o[9947] = i[9947];
  assign o[9946] = i[9946];
  assign o[9945] = i[9945];
  assign o[9944] = i[9944];
  assign o[9943] = i[9943];
  assign o[9942] = i[9942];
  assign o[9941] = i[9941];
  assign o[9940] = i[9940];
  assign o[9939] = i[9939];
  assign o[9938] = i[9938];
  assign o[9937] = i[9937];
  assign o[9936] = i[9936];
  assign o[9935] = i[9935];
  assign o[9934] = i[9934];
  assign o[9933] = i[9933];
  assign o[9932] = i[9932];
  assign o[9931] = i[9931];
  assign o[9930] = i[9930];
  assign o[9929] = i[9929];
  assign o[9928] = i[9928];
  assign o[9927] = i[9927];
  assign o[9926] = i[9926];
  assign o[9925] = i[9925];
  assign o[9924] = i[9924];
  assign o[9923] = i[9923];
  assign o[9922] = i[9922];
  assign o[9921] = i[9921];
  assign o[9920] = i[9920];
  assign o[9919] = i[9919];
  assign o[9918] = i[9918];
  assign o[9917] = i[9917];
  assign o[9916] = i[9916];
  assign o[9915] = i[9915];
  assign o[9914] = i[9914];
  assign o[9913] = i[9913];
  assign o[9912] = i[9912];
  assign o[9911] = i[9911];
  assign o[9910] = i[9910];
  assign o[9909] = i[9909];
  assign o[9908] = i[9908];
  assign o[9907] = i[9907];
  assign o[9906] = i[9906];
  assign o[9905] = i[9905];
  assign o[9904] = i[9904];
  assign o[9903] = i[9903];
  assign o[9902] = i[9902];
  assign o[9901] = i[9901];
  assign o[9900] = i[9900];
  assign o[9899] = i[9899];
  assign o[9898] = i[9898];
  assign o[9897] = i[9897];
  assign o[9896] = i[9896];
  assign o[9895] = i[9895];
  assign o[9894] = i[9894];
  assign o[9893] = i[9893];
  assign o[9892] = i[9892];
  assign o[9891] = i[9891];
  assign o[9890] = i[9890];
  assign o[9889] = i[9889];
  assign o[9888] = i[9888];
  assign o[9887] = i[9887];
  assign o[9886] = i[9886];
  assign o[9885] = i[9885];
  assign o[9884] = i[9884];
  assign o[9883] = i[9883];
  assign o[9882] = i[9882];
  assign o[9881] = i[9881];
  assign o[9880] = i[9880];
  assign o[9879] = i[9879];
  assign o[9878] = i[9878];
  assign o[9877] = i[9877];
  assign o[9876] = i[9876];
  assign o[9875] = i[9875];
  assign o[9874] = i[9874];
  assign o[9873] = i[9873];
  assign o[9872] = i[9872];
  assign o[9871] = i[9871];
  assign o[9870] = i[9870];
  assign o[9869] = i[9869];
  assign o[9868] = i[9868];
  assign o[9867] = i[9867];
  assign o[9866] = i[9866];
  assign o[9865] = i[9865];
  assign o[9864] = i[9864];
  assign o[9863] = i[9863];
  assign o[9862] = i[9862];
  assign o[9861] = i[9861];
  assign o[9860] = i[9860];
  assign o[9859] = i[9859];
  assign o[9858] = i[9858];
  assign o[9857] = i[9857];
  assign o[9856] = i[9856];
  assign o[9855] = i[9855];
  assign o[9854] = i[9854];
  assign o[9853] = i[9853];
  assign o[9852] = i[9852];
  assign o[9851] = i[9851];
  assign o[9850] = i[9850];
  assign o[9849] = i[9849];
  assign o[9848] = i[9848];
  assign o[9847] = i[9847];
  assign o[9846] = i[9846];
  assign o[9845] = i[9845];
  assign o[9844] = i[9844];
  assign o[9843] = i[9843];
  assign o[9842] = i[9842];
  assign o[9841] = i[9841];
  assign o[9840] = i[9840];
  assign o[9839] = i[9839];
  assign o[9838] = i[9838];
  assign o[9837] = i[9837];
  assign o[9836] = i[9836];
  assign o[9835] = i[9835];
  assign o[9834] = i[9834];
  assign o[9833] = i[9833];
  assign o[9832] = i[9832];
  assign o[9831] = i[9831];
  assign o[9830] = i[9830];
  assign o[9829] = i[9829];
  assign o[9828] = i[9828];
  assign o[9827] = i[9827];
  assign o[9826] = i[9826];
  assign o[9825] = i[9825];
  assign o[9824] = i[9824];
  assign o[9823] = i[9823];
  assign o[9822] = i[9822];
  assign o[9821] = i[9821];
  assign o[9820] = i[9820];
  assign o[9819] = i[9819];
  assign o[9818] = i[9818];
  assign o[9817] = i[9817];
  assign o[9816] = i[9816];
  assign o[9815] = i[9815];
  assign o[9814] = i[9814];
  assign o[9813] = i[9813];
  assign o[9812] = i[9812];
  assign o[9811] = i[9811];
  assign o[9810] = i[9810];
  assign o[9809] = i[9809];
  assign o[9808] = i[9808];
  assign o[9807] = i[9807];
  assign o[9806] = i[9806];
  assign o[9805] = i[9805];
  assign o[9804] = i[9804];
  assign o[9803] = i[9803];
  assign o[9802] = i[9802];
  assign o[9801] = i[9801];
  assign o[9800] = i[9800];
  assign o[9799] = i[9799];
  assign o[9798] = i[9798];
  assign o[9797] = i[9797];
  assign o[9796] = i[9796];
  assign o[9795] = i[9795];
  assign o[9794] = i[9794];
  assign o[9793] = i[9793];
  assign o[9792] = i[9792];
  assign o[9791] = i[9791];
  assign o[9790] = i[9790];
  assign o[9789] = i[9789];
  assign o[9788] = i[9788];
  assign o[9787] = i[9787];
  assign o[9786] = i[9786];
  assign o[9785] = i[9785];
  assign o[9784] = i[9784];
  assign o[9783] = i[9783];
  assign o[9782] = i[9782];
  assign o[9781] = i[9781];
  assign o[9780] = i[9780];
  assign o[9779] = i[9779];
  assign o[9778] = i[9778];
  assign o[9777] = i[9777];
  assign o[9776] = i[9776];
  assign o[9775] = i[9775];
  assign o[9774] = i[9774];
  assign o[9773] = i[9773];
  assign o[9772] = i[9772];
  assign o[9771] = i[9771];
  assign o[9770] = i[9770];
  assign o[9769] = i[9769];
  assign o[9768] = i[9768];
  assign o[9767] = i[9767];
  assign o[9766] = i[9766];
  assign o[9765] = i[9765];
  assign o[9764] = i[9764];
  assign o[9763] = i[9763];
  assign o[9762] = i[9762];
  assign o[9761] = i[9761];
  assign o[9760] = i[9760];
  assign o[9759] = i[9759];
  assign o[9758] = i[9758];
  assign o[9757] = i[9757];
  assign o[9756] = i[9756];
  assign o[9755] = i[9755];
  assign o[9754] = i[9754];
  assign o[9753] = i[9753];
  assign o[9752] = i[9752];
  assign o[9751] = i[9751];
  assign o[9750] = i[9750];
  assign o[9749] = i[9749];
  assign o[9748] = i[9748];
  assign o[9747] = i[9747];
  assign o[9746] = i[9746];
  assign o[9745] = i[9745];
  assign o[9744] = i[9744];
  assign o[9743] = i[9743];
  assign o[9742] = i[9742];
  assign o[9741] = i[9741];
  assign o[9740] = i[9740];
  assign o[9739] = i[9739];
  assign o[9738] = i[9738];
  assign o[9737] = i[9737];
  assign o[9736] = i[9736];
  assign o[9735] = i[9735];
  assign o[9734] = i[9734];
  assign o[9733] = i[9733];
  assign o[9732] = i[9732];
  assign o[9731] = i[9731];
  assign o[9730] = i[9730];
  assign o[9729] = i[9729];
  assign o[9728] = i[9728];
  assign o[9727] = i[9727];
  assign o[9726] = i[9726];
  assign o[9725] = i[9725];
  assign o[9724] = i[9724];
  assign o[9723] = i[9723];
  assign o[9722] = i[9722];
  assign o[9721] = i[9721];
  assign o[9720] = i[9720];
  assign o[9719] = i[9719];
  assign o[9718] = i[9718];
  assign o[9717] = i[9717];
  assign o[9716] = i[9716];
  assign o[9715] = i[9715];
  assign o[9714] = i[9714];
  assign o[9713] = i[9713];
  assign o[9712] = i[9712];
  assign o[9711] = i[9711];
  assign o[9710] = i[9710];
  assign o[9709] = i[9709];
  assign o[9708] = i[9708];
  assign o[9707] = i[9707];
  assign o[9706] = i[9706];
  assign o[9705] = i[9705];
  assign o[9704] = i[9704];
  assign o[9703] = i[9703];
  assign o[9702] = i[9702];
  assign o[9701] = i[9701];
  assign o[9700] = i[9700];
  assign o[9699] = i[9699];
  assign o[9698] = i[9698];
  assign o[9697] = i[9697];
  assign o[9696] = i[9696];
  assign o[9695] = i[9695];
  assign o[9694] = i[9694];
  assign o[9693] = i[9693];
  assign o[9692] = i[9692];
  assign o[9691] = i[9691];
  assign o[9690] = i[9690];
  assign o[9689] = i[9689];
  assign o[9688] = i[9688];
  assign o[9687] = i[9687];
  assign o[9686] = i[9686];
  assign o[9685] = i[9685];
  assign o[9684] = i[9684];
  assign o[9683] = i[9683];
  assign o[9682] = i[9682];
  assign o[9681] = i[9681];
  assign o[9680] = i[9680];
  assign o[9679] = i[9679];
  assign o[9678] = i[9678];
  assign o[9677] = i[9677];
  assign o[9676] = i[9676];
  assign o[9675] = i[9675];
  assign o[9674] = i[9674];
  assign o[9673] = i[9673];
  assign o[9672] = i[9672];
  assign o[9671] = i[9671];
  assign o[9670] = i[9670];
  assign o[9669] = i[9669];
  assign o[9668] = i[9668];
  assign o[9667] = i[9667];
  assign o[9666] = i[9666];
  assign o[9665] = i[9665];
  assign o[9664] = i[9664];
  assign o[9663] = i[9663];
  assign o[9662] = i[9662];
  assign o[9661] = i[9661];
  assign o[9660] = i[9660];
  assign o[9659] = i[9659];
  assign o[9658] = i[9658];
  assign o[9657] = i[9657];
  assign o[9656] = i[9656];
  assign o[9655] = i[9655];
  assign o[9654] = i[9654];
  assign o[9653] = i[9653];
  assign o[9652] = i[9652];
  assign o[9651] = i[9651];
  assign o[9650] = i[9650];
  assign o[9649] = i[9649];
  assign o[9648] = i[9648];
  assign o[9647] = i[9647];
  assign o[9646] = i[9646];
  assign o[9645] = i[9645];
  assign o[9644] = i[9644];
  assign o[9643] = i[9643];
  assign o[9642] = i[9642];
  assign o[9641] = i[9641];
  assign o[9640] = i[9640];
  assign o[9639] = i[9639];
  assign o[9638] = i[9638];
  assign o[9637] = i[9637];
  assign o[9636] = i[9636];
  assign o[9635] = i[9635];
  assign o[9634] = i[9634];
  assign o[9633] = i[9633];
  assign o[9632] = i[9632];
  assign o[9631] = i[9631];
  assign o[9630] = i[9630];
  assign o[9629] = i[9629];
  assign o[9628] = i[9628];
  assign o[9627] = i[9627];
  assign o[9626] = i[9626];
  assign o[9625] = i[9625];
  assign o[9624] = i[9624];
  assign o[9623] = i[9623];
  assign o[9622] = i[9622];
  assign o[9621] = i[9621];
  assign o[9620] = i[9620];
  assign o[9619] = i[9619];
  assign o[9618] = i[9618];
  assign o[9617] = i[9617];
  assign o[9616] = i[9616];
  assign o[9615] = i[9615];
  assign o[9614] = i[9614];
  assign o[9613] = i[9613];
  assign o[9612] = i[9612];
  assign o[9611] = i[9611];
  assign o[9610] = i[9610];
  assign o[9609] = i[9609];
  assign o[9608] = i[9608];
  assign o[9607] = i[9607];
  assign o[9606] = i[9606];
  assign o[9605] = i[9605];
  assign o[9604] = i[9604];
  assign o[9603] = i[9603];
  assign o[9602] = i[9602];
  assign o[9601] = i[9601];
  assign o[9600] = i[9600];
  assign o[9599] = i[9599];
  assign o[9598] = i[9598];
  assign o[9597] = i[9597];
  assign o[9596] = i[9596];
  assign o[9595] = i[9595];
  assign o[9594] = i[9594];
  assign o[9593] = i[9593];
  assign o[9592] = i[9592];
  assign o[9591] = i[9591];
  assign o[9590] = i[9590];
  assign o[9589] = i[9589];
  assign o[9588] = i[9588];
  assign o[9587] = i[9587];
  assign o[9586] = i[9586];
  assign o[9585] = i[9585];
  assign o[9584] = i[9584];
  assign o[9583] = i[9583];
  assign o[9582] = i[9582];
  assign o[9581] = i[9581];
  assign o[9580] = i[9580];
  assign o[9579] = i[9579];
  assign o[9578] = i[9578];
  assign o[9577] = i[9577];
  assign o[9576] = i[9576];
  assign o[9575] = i[9575];
  assign o[9574] = i[9574];
  assign o[9573] = i[9573];
  assign o[9572] = i[9572];
  assign o[9571] = i[9571];
  assign o[9570] = i[9570];
  assign o[9569] = i[9569];
  assign o[9568] = i[9568];
  assign o[9567] = i[9567];
  assign o[9566] = i[9566];
  assign o[9565] = i[9565];
  assign o[9564] = i[9564];
  assign o[9563] = i[9563];
  assign o[9562] = i[9562];
  assign o[9561] = i[9561];
  assign o[9560] = i[9560];
  assign o[9559] = i[9559];
  assign o[9558] = i[9558];
  assign o[9557] = i[9557];
  assign o[9556] = i[9556];
  assign o[9555] = i[9555];
  assign o[9554] = i[9554];
  assign o[9553] = i[9553];
  assign o[9552] = i[9552];
  assign o[9551] = i[9551];
  assign o[9550] = i[9550];
  assign o[9549] = i[9549];
  assign o[9548] = i[9548];
  assign o[9547] = i[9547];
  assign o[9546] = i[9546];
  assign o[9545] = i[9545];
  assign o[9544] = i[9544];
  assign o[9543] = i[9543];
  assign o[9542] = i[9542];
  assign o[9541] = i[9541];
  assign o[9540] = i[9540];
  assign o[9539] = i[9539];
  assign o[9538] = i[9538];
  assign o[9537] = i[9537];
  assign o[9536] = i[9536];
  assign o[9535] = i[9535];
  assign o[9534] = i[9534];
  assign o[9533] = i[9533];
  assign o[9532] = i[9532];
  assign o[9531] = i[9531];
  assign o[9530] = i[9530];
  assign o[9529] = i[9529];
  assign o[9528] = i[9528];
  assign o[9527] = i[9527];
  assign o[9526] = i[9526];
  assign o[9525] = i[9525];
  assign o[9524] = i[9524];
  assign o[9523] = i[9523];
  assign o[9522] = i[9522];
  assign o[9521] = i[9521];
  assign o[9520] = i[9520];
  assign o[9519] = i[9519];
  assign o[9518] = i[9518];
  assign o[9517] = i[9517];
  assign o[9516] = i[9516];
  assign o[9515] = i[9515];
  assign o[9514] = i[9514];
  assign o[9513] = i[9513];
  assign o[9512] = i[9512];
  assign o[9511] = i[9511];
  assign o[9510] = i[9510];
  assign o[9509] = i[9509];
  assign o[9508] = i[9508];
  assign o[9507] = i[9507];
  assign o[9506] = i[9506];
  assign o[9505] = i[9505];
  assign o[9504] = i[9504];
  assign o[9503] = i[9503];
  assign o[9502] = i[9502];
  assign o[9501] = i[9501];
  assign o[9500] = i[9500];
  assign o[9499] = i[9499];
  assign o[9498] = i[9498];
  assign o[9497] = i[9497];
  assign o[9496] = i[9496];
  assign o[9495] = i[9495];
  assign o[9494] = i[9494];
  assign o[9493] = i[9493];
  assign o[9492] = i[9492];
  assign o[9491] = i[9491];
  assign o[9490] = i[9490];
  assign o[9489] = i[9489];
  assign o[9488] = i[9488];
  assign o[9487] = i[9487];
  assign o[9486] = i[9486];
  assign o[9485] = i[9485];
  assign o[9484] = i[9484];
  assign o[9483] = i[9483];
  assign o[9482] = i[9482];
  assign o[9481] = i[9481];
  assign o[9480] = i[9480];
  assign o[9479] = i[9479];
  assign o[9478] = i[9478];
  assign o[9477] = i[9477];
  assign o[9476] = i[9476];
  assign o[9475] = i[9475];
  assign o[9474] = i[9474];
  assign o[9473] = i[9473];
  assign o[9472] = i[9472];
  assign o[9471] = i[9471];
  assign o[9470] = i[9470];
  assign o[9469] = i[9469];
  assign o[9468] = i[9468];
  assign o[9467] = i[9467];
  assign o[9466] = i[9466];
  assign o[9465] = i[9465];
  assign o[9464] = i[9464];
  assign o[9463] = i[9463];
  assign o[9462] = i[9462];
  assign o[9461] = i[9461];
  assign o[9460] = i[9460];
  assign o[9459] = i[9459];
  assign o[9458] = i[9458];
  assign o[9457] = i[9457];
  assign o[9456] = i[9456];
  assign o[9455] = i[9455];
  assign o[9454] = i[9454];
  assign o[9453] = i[9453];
  assign o[9452] = i[9452];
  assign o[9451] = i[9451];
  assign o[9450] = i[9450];
  assign o[9449] = i[9449];
  assign o[9448] = i[9448];
  assign o[9447] = i[9447];
  assign o[9446] = i[9446];
  assign o[9445] = i[9445];
  assign o[9444] = i[9444];
  assign o[9443] = i[9443];
  assign o[9442] = i[9442];
  assign o[9441] = i[9441];
  assign o[9440] = i[9440];
  assign o[9439] = i[9439];
  assign o[9438] = i[9438];
  assign o[9437] = i[9437];
  assign o[9436] = i[9436];
  assign o[9435] = i[9435];
  assign o[9434] = i[9434];
  assign o[9433] = i[9433];
  assign o[9432] = i[9432];
  assign o[9431] = i[9431];
  assign o[9430] = i[9430];
  assign o[9429] = i[9429];
  assign o[9428] = i[9428];
  assign o[9427] = i[9427];
  assign o[9426] = i[9426];
  assign o[9425] = i[9425];
  assign o[9424] = i[9424];
  assign o[9423] = i[9423];
  assign o[9422] = i[9422];
  assign o[9421] = i[9421];
  assign o[9420] = i[9420];
  assign o[9419] = i[9419];
  assign o[9418] = i[9418];
  assign o[9417] = i[9417];
  assign o[9416] = i[9416];
  assign o[9415] = i[9415];
  assign o[9414] = i[9414];
  assign o[9413] = i[9413];
  assign o[9412] = i[9412];
  assign o[9411] = i[9411];
  assign o[9410] = i[9410];
  assign o[9409] = i[9409];
  assign o[9408] = i[9408];
  assign o[9407] = i[9407];
  assign o[9406] = i[9406];
  assign o[9405] = i[9405];
  assign o[9404] = i[9404];
  assign o[9403] = i[9403];
  assign o[9402] = i[9402];
  assign o[9401] = i[9401];
  assign o[9400] = i[9400];
  assign o[9399] = i[9399];
  assign o[9398] = i[9398];
  assign o[9397] = i[9397];
  assign o[9396] = i[9396];
  assign o[9395] = i[9395];
  assign o[9394] = i[9394];
  assign o[9393] = i[9393];
  assign o[9392] = i[9392];
  assign o[9391] = i[9391];
  assign o[9390] = i[9390];
  assign o[9389] = i[9389];
  assign o[9388] = i[9388];
  assign o[9387] = i[9387];
  assign o[9386] = i[9386];
  assign o[9385] = i[9385];
  assign o[9384] = i[9384];
  assign o[9383] = i[9383];
  assign o[9382] = i[9382];
  assign o[9381] = i[9381];
  assign o[9380] = i[9380];
  assign o[9379] = i[9379];
  assign o[9378] = i[9378];
  assign o[9377] = i[9377];
  assign o[9376] = i[9376];
  assign o[9375] = i[9375];
  assign o[9374] = i[9374];
  assign o[9373] = i[9373];
  assign o[9372] = i[9372];
  assign o[9371] = i[9371];
  assign o[9370] = i[9370];
  assign o[9369] = i[9369];
  assign o[9368] = i[9368];
  assign o[9367] = i[9367];
  assign o[9366] = i[9366];
  assign o[9365] = i[9365];
  assign o[9364] = i[9364];
  assign o[9363] = i[9363];
  assign o[9362] = i[9362];
  assign o[9361] = i[9361];
  assign o[9360] = i[9360];
  assign o[9359] = i[9359];
  assign o[9358] = i[9358];
  assign o[9357] = i[9357];
  assign o[9356] = i[9356];
  assign o[9355] = i[9355];
  assign o[9354] = i[9354];
  assign o[9353] = i[9353];
  assign o[9352] = i[9352];
  assign o[9351] = i[9351];
  assign o[9350] = i[9350];
  assign o[9349] = i[9349];
  assign o[9348] = i[9348];
  assign o[9347] = i[9347];
  assign o[9346] = i[9346];
  assign o[9345] = i[9345];
  assign o[9344] = i[9344];
  assign o[9343] = i[9343];
  assign o[9342] = i[9342];
  assign o[9341] = i[9341];
  assign o[9340] = i[9340];
  assign o[9339] = i[9339];
  assign o[9338] = i[9338];
  assign o[9337] = i[9337];
  assign o[9336] = i[9336];
  assign o[9335] = i[9335];
  assign o[9334] = i[9334];
  assign o[9333] = i[9333];
  assign o[9332] = i[9332];
  assign o[9331] = i[9331];
  assign o[9330] = i[9330];
  assign o[9329] = i[9329];
  assign o[9328] = i[9328];
  assign o[9327] = i[9327];
  assign o[9326] = i[9326];
  assign o[9325] = i[9325];
  assign o[9324] = i[9324];
  assign o[9323] = i[9323];
  assign o[9322] = i[9322];
  assign o[9321] = i[9321];
  assign o[9320] = i[9320];
  assign o[9319] = i[9319];
  assign o[9318] = i[9318];
  assign o[9317] = i[9317];
  assign o[9316] = i[9316];
  assign o[9315] = i[9315];
  assign o[9314] = i[9314];
  assign o[9313] = i[9313];
  assign o[9312] = i[9312];
  assign o[9311] = i[9311];
  assign o[9310] = i[9310];
  assign o[9309] = i[9309];
  assign o[9308] = i[9308];
  assign o[9307] = i[9307];
  assign o[9306] = i[9306];
  assign o[9305] = i[9305];
  assign o[9304] = i[9304];
  assign o[9303] = i[9303];
  assign o[9302] = i[9302];
  assign o[9301] = i[9301];
  assign o[9300] = i[9300];
  assign o[9299] = i[9299];
  assign o[9298] = i[9298];
  assign o[9297] = i[9297];
  assign o[9296] = i[9296];
  assign o[9295] = i[9295];
  assign o[9294] = i[9294];
  assign o[9293] = i[9293];
  assign o[9292] = i[9292];
  assign o[9291] = i[9291];
  assign o[9290] = i[9290];
  assign o[9289] = i[9289];
  assign o[9288] = i[9288];
  assign o[9287] = i[9287];
  assign o[9286] = i[9286];
  assign o[9285] = i[9285];
  assign o[9284] = i[9284];
  assign o[9283] = i[9283];
  assign o[9282] = i[9282];
  assign o[9281] = i[9281];
  assign o[9280] = i[9280];
  assign o[9279] = i[9279];
  assign o[9278] = i[9278];
  assign o[9277] = i[9277];
  assign o[9276] = i[9276];
  assign o[9275] = i[9275];
  assign o[9274] = i[9274];
  assign o[9273] = i[9273];
  assign o[9272] = i[9272];
  assign o[9271] = i[9271];
  assign o[9270] = i[9270];
  assign o[9269] = i[9269];
  assign o[9268] = i[9268];
  assign o[9267] = i[9267];
  assign o[9266] = i[9266];
  assign o[9265] = i[9265];
  assign o[9264] = i[9264];
  assign o[9263] = i[9263];
  assign o[9262] = i[9262];
  assign o[9261] = i[9261];
  assign o[9260] = i[9260];
  assign o[9259] = i[9259];
  assign o[9258] = i[9258];
  assign o[9257] = i[9257];
  assign o[9256] = i[9256];
  assign o[9255] = i[9255];
  assign o[9254] = i[9254];
  assign o[9253] = i[9253];
  assign o[9252] = i[9252];
  assign o[9251] = i[9251];
  assign o[9250] = i[9250];
  assign o[9249] = i[9249];
  assign o[9248] = i[9248];
  assign o[9247] = i[9247];
  assign o[9246] = i[9246];
  assign o[9245] = i[9245];
  assign o[9244] = i[9244];
  assign o[9243] = i[9243];
  assign o[9242] = i[9242];
  assign o[9241] = i[9241];
  assign o[9240] = i[9240];
  assign o[9239] = i[9239];
  assign o[9238] = i[9238];
  assign o[9237] = i[9237];
  assign o[9236] = i[9236];
  assign o[9235] = i[9235];
  assign o[9234] = i[9234];
  assign o[9233] = i[9233];
  assign o[9232] = i[9232];
  assign o[9231] = i[9231];
  assign o[9230] = i[9230];
  assign o[9229] = i[9229];
  assign o[9228] = i[9228];
  assign o[9227] = i[9227];
  assign o[9226] = i[9226];
  assign o[9225] = i[9225];
  assign o[9224] = i[9224];
  assign o[9223] = i[9223];
  assign o[9222] = i[9222];
  assign o[9221] = i[9221];
  assign o[9220] = i[9220];
  assign o[9219] = i[9219];
  assign o[9218] = i[9218];
  assign o[9217] = i[9217];
  assign o[9216] = i[9216];
  assign o[9215] = i[9215];
  assign o[9214] = i[9214];
  assign o[9213] = i[9213];
  assign o[9212] = i[9212];
  assign o[9211] = i[9211];
  assign o[9210] = i[9210];
  assign o[9209] = i[9209];
  assign o[9208] = i[9208];
  assign o[9207] = i[9207];
  assign o[9206] = i[9206];
  assign o[9205] = i[9205];
  assign o[9204] = i[9204];
  assign o[9203] = i[9203];
  assign o[9202] = i[9202];
  assign o[9201] = i[9201];
  assign o[9200] = i[9200];
  assign o[9199] = i[9199];
  assign o[9198] = i[9198];
  assign o[9197] = i[9197];
  assign o[9196] = i[9196];
  assign o[9195] = i[9195];
  assign o[9194] = i[9194];
  assign o[9193] = i[9193];
  assign o[9192] = i[9192];
  assign o[9191] = i[9191];
  assign o[9190] = i[9190];
  assign o[9189] = i[9189];
  assign o[9188] = i[9188];
  assign o[9187] = i[9187];
  assign o[9186] = i[9186];
  assign o[9185] = i[9185];
  assign o[9184] = i[9184];
  assign o[9183] = i[9183];
  assign o[9182] = i[9182];
  assign o[9181] = i[9181];
  assign o[9180] = i[9180];
  assign o[9179] = i[9179];
  assign o[9178] = i[9178];
  assign o[9177] = i[9177];
  assign o[9176] = i[9176];
  assign o[9175] = i[9175];
  assign o[9174] = i[9174];
  assign o[9173] = i[9173];
  assign o[9172] = i[9172];
  assign o[9171] = i[9171];
  assign o[9170] = i[9170];
  assign o[9169] = i[9169];
  assign o[9168] = i[9168];
  assign o[9167] = i[9167];
  assign o[9166] = i[9166];
  assign o[9165] = i[9165];
  assign o[9164] = i[9164];
  assign o[9163] = i[9163];
  assign o[9162] = i[9162];
  assign o[9161] = i[9161];
  assign o[9160] = i[9160];
  assign o[9159] = i[9159];
  assign o[9158] = i[9158];
  assign o[9157] = i[9157];
  assign o[9156] = i[9156];
  assign o[9155] = i[9155];
  assign o[9154] = i[9154];
  assign o[9153] = i[9153];
  assign o[9152] = i[9152];
  assign o[9151] = i[9151];
  assign o[9150] = i[9150];
  assign o[9149] = i[9149];
  assign o[9148] = i[9148];
  assign o[9147] = i[9147];
  assign o[9146] = i[9146];
  assign o[9145] = i[9145];
  assign o[9144] = i[9144];
  assign o[9143] = i[9143];
  assign o[9142] = i[9142];
  assign o[9141] = i[9141];
  assign o[9140] = i[9140];
  assign o[9139] = i[9139];
  assign o[9138] = i[9138];
  assign o[9137] = i[9137];
  assign o[9136] = i[9136];
  assign o[9135] = i[9135];
  assign o[9134] = i[9134];
  assign o[9133] = i[9133];
  assign o[9132] = i[9132];
  assign o[9131] = i[9131];
  assign o[9130] = i[9130];
  assign o[9129] = i[9129];
  assign o[9128] = i[9128];
  assign o[9127] = i[9127];
  assign o[9126] = i[9126];
  assign o[9125] = i[9125];
  assign o[9124] = i[9124];
  assign o[9123] = i[9123];
  assign o[9122] = i[9122];
  assign o[9121] = i[9121];
  assign o[9120] = i[9120];
  assign o[9119] = i[9119];
  assign o[9118] = i[9118];
  assign o[9117] = i[9117];
  assign o[9116] = i[9116];
  assign o[9115] = i[9115];
  assign o[9114] = i[9114];
  assign o[9113] = i[9113];
  assign o[9112] = i[9112];
  assign o[9111] = i[9111];
  assign o[9110] = i[9110];
  assign o[9109] = i[9109];
  assign o[9108] = i[9108];
  assign o[9107] = i[9107];
  assign o[9106] = i[9106];
  assign o[9105] = i[9105];
  assign o[9104] = i[9104];
  assign o[9103] = i[9103];
  assign o[9102] = i[9102];
  assign o[9101] = i[9101];
  assign o[9100] = i[9100];
  assign o[9099] = i[9099];
  assign o[9098] = i[9098];
  assign o[9097] = i[9097];
  assign o[9096] = i[9096];
  assign o[9095] = i[9095];
  assign o[9094] = i[9094];
  assign o[9093] = i[9093];
  assign o[9092] = i[9092];
  assign o[9091] = i[9091];
  assign o[9090] = i[9090];
  assign o[9089] = i[9089];
  assign o[9088] = i[9088];
  assign o[9087] = i[9087];
  assign o[9086] = i[9086];
  assign o[9085] = i[9085];
  assign o[9084] = i[9084];
  assign o[9083] = i[9083];
  assign o[9082] = i[9082];
  assign o[9081] = i[9081];
  assign o[9080] = i[9080];
  assign o[9079] = i[9079];
  assign o[9078] = i[9078];
  assign o[9077] = i[9077];
  assign o[9076] = i[9076];
  assign o[9075] = i[9075];
  assign o[9074] = i[9074];
  assign o[9073] = i[9073];
  assign o[9072] = i[9072];
  assign o[9071] = i[9071];
  assign o[9070] = i[9070];
  assign o[9069] = i[9069];
  assign o[9068] = i[9068];
  assign o[9067] = i[9067];
  assign o[9066] = i[9066];
  assign o[9065] = i[9065];
  assign o[9064] = i[9064];
  assign o[9063] = i[9063];
  assign o[9062] = i[9062];
  assign o[9061] = i[9061];
  assign o[9060] = i[9060];
  assign o[9059] = i[9059];
  assign o[9058] = i[9058];
  assign o[9057] = i[9057];
  assign o[9056] = i[9056];
  assign o[9055] = i[9055];
  assign o[9054] = i[9054];
  assign o[9053] = i[9053];
  assign o[9052] = i[9052];
  assign o[9051] = i[9051];
  assign o[9050] = i[9050];
  assign o[9049] = i[9049];
  assign o[9048] = i[9048];
  assign o[9047] = i[9047];
  assign o[9046] = i[9046];
  assign o[9045] = i[9045];
  assign o[9044] = i[9044];
  assign o[9043] = i[9043];
  assign o[9042] = i[9042];
  assign o[9041] = i[9041];
  assign o[9040] = i[9040];
  assign o[9039] = i[9039];
  assign o[9038] = i[9038];
  assign o[9037] = i[9037];
  assign o[9036] = i[9036];
  assign o[9035] = i[9035];
  assign o[9034] = i[9034];
  assign o[9033] = i[9033];
  assign o[9032] = i[9032];
  assign o[9031] = i[9031];
  assign o[9030] = i[9030];
  assign o[9029] = i[9029];
  assign o[9028] = i[9028];
  assign o[9027] = i[9027];
  assign o[9026] = i[9026];
  assign o[9025] = i[9025];
  assign o[9024] = i[9024];
  assign o[9023] = i[9023];
  assign o[9022] = i[9022];
  assign o[9021] = i[9021];
  assign o[9020] = i[9020];
  assign o[9019] = i[9019];
  assign o[9018] = i[9018];
  assign o[9017] = i[9017];
  assign o[9016] = i[9016];
  assign o[9015] = i[9015];
  assign o[9014] = i[9014];
  assign o[9013] = i[9013];
  assign o[9012] = i[9012];
  assign o[9011] = i[9011];
  assign o[9010] = i[9010];
  assign o[9009] = i[9009];
  assign o[9008] = i[9008];
  assign o[9007] = i[9007];
  assign o[9006] = i[9006];
  assign o[9005] = i[9005];
  assign o[9004] = i[9004];
  assign o[9003] = i[9003];
  assign o[9002] = i[9002];
  assign o[9001] = i[9001];
  assign o[9000] = i[9000];
  assign o[8999] = i[8999];
  assign o[8998] = i[8998];
  assign o[8997] = i[8997];
  assign o[8996] = i[8996];
  assign o[8995] = i[8995];
  assign o[8994] = i[8994];
  assign o[8993] = i[8993];
  assign o[8992] = i[8992];
  assign o[8991] = i[8991];
  assign o[8990] = i[8990];
  assign o[8989] = i[8989];
  assign o[8988] = i[8988];
  assign o[8987] = i[8987];
  assign o[8986] = i[8986];
  assign o[8985] = i[8985];
  assign o[8984] = i[8984];
  assign o[8983] = i[8983];
  assign o[8982] = i[8982];
  assign o[8981] = i[8981];
  assign o[8980] = i[8980];
  assign o[8979] = i[8979];
  assign o[8978] = i[8978];
  assign o[8977] = i[8977];
  assign o[8976] = i[8976];
  assign o[8975] = i[8975];
  assign o[8974] = i[8974];
  assign o[8973] = i[8973];
  assign o[8972] = i[8972];
  assign o[8971] = i[8971];
  assign o[8970] = i[8970];
  assign o[8969] = i[8969];
  assign o[8968] = i[8968];
  assign o[8967] = i[8967];
  assign o[8966] = i[8966];
  assign o[8965] = i[8965];
  assign o[8964] = i[8964];
  assign o[8963] = i[8963];
  assign o[8962] = i[8962];
  assign o[8961] = i[8961];
  assign o[8960] = i[8960];
  assign o[8959] = i[8959];
  assign o[8958] = i[8958];
  assign o[8957] = i[8957];
  assign o[8956] = i[8956];
  assign o[8955] = i[8955];
  assign o[8954] = i[8954];
  assign o[8953] = i[8953];
  assign o[8952] = i[8952];
  assign o[8951] = i[8951];
  assign o[8950] = i[8950];
  assign o[8949] = i[8949];
  assign o[8948] = i[8948];
  assign o[8947] = i[8947];
  assign o[8946] = i[8946];
  assign o[8945] = i[8945];
  assign o[8944] = i[8944];
  assign o[8943] = i[8943];
  assign o[8942] = i[8942];
  assign o[8941] = i[8941];
  assign o[8940] = i[8940];
  assign o[8939] = i[8939];
  assign o[8938] = i[8938];
  assign o[8937] = i[8937];
  assign o[8936] = i[8936];
  assign o[8935] = i[8935];
  assign o[8934] = i[8934];
  assign o[8933] = i[8933];
  assign o[8932] = i[8932];
  assign o[8931] = i[8931];
  assign o[8930] = i[8930];
  assign o[8929] = i[8929];
  assign o[8928] = i[8928];
  assign o[8927] = i[8927];
  assign o[8926] = i[8926];
  assign o[8925] = i[8925];
  assign o[8924] = i[8924];
  assign o[8923] = i[8923];
  assign o[8922] = i[8922];
  assign o[8921] = i[8921];
  assign o[8920] = i[8920];
  assign o[8919] = i[8919];
  assign o[8918] = i[8918];
  assign o[8917] = i[8917];
  assign o[8916] = i[8916];
  assign o[8915] = i[8915];
  assign o[8914] = i[8914];
  assign o[8913] = i[8913];
  assign o[8912] = i[8912];
  assign o[8911] = i[8911];
  assign o[8910] = i[8910];
  assign o[8909] = i[8909];
  assign o[8908] = i[8908];
  assign o[8907] = i[8907];
  assign o[8906] = i[8906];
  assign o[8905] = i[8905];
  assign o[8904] = i[8904];
  assign o[8903] = i[8903];
  assign o[8902] = i[8902];
  assign o[8901] = i[8901];
  assign o[8900] = i[8900];
  assign o[8899] = i[8899];
  assign o[8898] = i[8898];
  assign o[8897] = i[8897];
  assign o[8896] = i[8896];
  assign o[8895] = i[8895];
  assign o[8894] = i[8894];
  assign o[8893] = i[8893];
  assign o[8892] = i[8892];
  assign o[8891] = i[8891];
  assign o[8890] = i[8890];
  assign o[8889] = i[8889];
  assign o[8888] = i[8888];
  assign o[8887] = i[8887];
  assign o[8886] = i[8886];
  assign o[8885] = i[8885];
  assign o[8884] = i[8884];
  assign o[8883] = i[8883];
  assign o[8882] = i[8882];
  assign o[8881] = i[8881];
  assign o[8880] = i[8880];
  assign o[8879] = i[8879];
  assign o[8878] = i[8878];
  assign o[8877] = i[8877];
  assign o[8876] = i[8876];
  assign o[8875] = i[8875];
  assign o[8874] = i[8874];
  assign o[8873] = i[8873];
  assign o[8872] = i[8872];
  assign o[8871] = i[8871];
  assign o[8870] = i[8870];
  assign o[8869] = i[8869];
  assign o[8868] = i[8868];
  assign o[8867] = i[8867];
  assign o[8866] = i[8866];
  assign o[8865] = i[8865];
  assign o[8864] = i[8864];
  assign o[8863] = i[8863];
  assign o[8862] = i[8862];
  assign o[8861] = i[8861];
  assign o[8860] = i[8860];
  assign o[8859] = i[8859];
  assign o[8858] = i[8858];
  assign o[8857] = i[8857];
  assign o[8856] = i[8856];
  assign o[8855] = i[8855];
  assign o[8854] = i[8854];
  assign o[8853] = i[8853];
  assign o[8852] = i[8852];
  assign o[8851] = i[8851];
  assign o[8850] = i[8850];
  assign o[8849] = i[8849];
  assign o[8848] = i[8848];
  assign o[8847] = i[8847];
  assign o[8846] = i[8846];
  assign o[8845] = i[8845];
  assign o[8844] = i[8844];
  assign o[8843] = i[8843];
  assign o[8842] = i[8842];
  assign o[8841] = i[8841];
  assign o[8840] = i[8840];
  assign o[8839] = i[8839];
  assign o[8838] = i[8838];
  assign o[8837] = i[8837];
  assign o[8836] = i[8836];
  assign o[8835] = i[8835];
  assign o[8834] = i[8834];
  assign o[8833] = i[8833];
  assign o[8832] = i[8832];
  assign o[8831] = i[8831];
  assign o[8830] = i[8830];
  assign o[8829] = i[8829];
  assign o[8828] = i[8828];
  assign o[8827] = i[8827];
  assign o[8826] = i[8826];
  assign o[8825] = i[8825];
  assign o[8824] = i[8824];
  assign o[8823] = i[8823];
  assign o[8822] = i[8822];
  assign o[8821] = i[8821];
  assign o[8820] = i[8820];
  assign o[8819] = i[8819];
  assign o[8818] = i[8818];
  assign o[8817] = i[8817];
  assign o[8816] = i[8816];
  assign o[8815] = i[8815];
  assign o[8814] = i[8814];
  assign o[8813] = i[8813];
  assign o[8812] = i[8812];
  assign o[8811] = i[8811];
  assign o[8810] = i[8810];
  assign o[8809] = i[8809];
  assign o[8808] = i[8808];
  assign o[8807] = i[8807];
  assign o[8806] = i[8806];
  assign o[8805] = i[8805];
  assign o[8804] = i[8804];
  assign o[8803] = i[8803];
  assign o[8802] = i[8802];
  assign o[8801] = i[8801];
  assign o[8800] = i[8800];
  assign o[8799] = i[8799];
  assign o[8798] = i[8798];
  assign o[8797] = i[8797];
  assign o[8796] = i[8796];
  assign o[8795] = i[8795];
  assign o[8794] = i[8794];
  assign o[8793] = i[8793];
  assign o[8792] = i[8792];
  assign o[8791] = i[8791];
  assign o[8790] = i[8790];
  assign o[8789] = i[8789];
  assign o[8788] = i[8788];
  assign o[8787] = i[8787];
  assign o[8786] = i[8786];
  assign o[8785] = i[8785];
  assign o[8784] = i[8784];
  assign o[8783] = i[8783];
  assign o[8782] = i[8782];
  assign o[8781] = i[8781];
  assign o[8780] = i[8780];
  assign o[8779] = i[8779];
  assign o[8778] = i[8778];
  assign o[8777] = i[8777];
  assign o[8776] = i[8776];
  assign o[8775] = i[8775];
  assign o[8774] = i[8774];
  assign o[8773] = i[8773];
  assign o[8772] = i[8772];
  assign o[8771] = i[8771];
  assign o[8770] = i[8770];
  assign o[8769] = i[8769];
  assign o[8768] = i[8768];
  assign o[8767] = i[8767];
  assign o[8766] = i[8766];
  assign o[8765] = i[8765];
  assign o[8764] = i[8764];
  assign o[8763] = i[8763];
  assign o[8762] = i[8762];
  assign o[8761] = i[8761];
  assign o[8760] = i[8760];
  assign o[8759] = i[8759];
  assign o[8758] = i[8758];
  assign o[8757] = i[8757];
  assign o[8756] = i[8756];
  assign o[8755] = i[8755];
  assign o[8754] = i[8754];
  assign o[8753] = i[8753];
  assign o[8752] = i[8752];
  assign o[8751] = i[8751];
  assign o[8750] = i[8750];
  assign o[8749] = i[8749];
  assign o[8748] = i[8748];
  assign o[8747] = i[8747];
  assign o[8746] = i[8746];
  assign o[8745] = i[8745];
  assign o[8744] = i[8744];
  assign o[8743] = i[8743];
  assign o[8742] = i[8742];
  assign o[8741] = i[8741];
  assign o[8740] = i[8740];
  assign o[8739] = i[8739];
  assign o[8738] = i[8738];
  assign o[8737] = i[8737];
  assign o[8736] = i[8736];
  assign o[8735] = i[8735];
  assign o[8734] = i[8734];
  assign o[8733] = i[8733];
  assign o[8732] = i[8732];
  assign o[8731] = i[8731];
  assign o[8730] = i[8730];
  assign o[8729] = i[8729];
  assign o[8728] = i[8728];
  assign o[8727] = i[8727];
  assign o[8726] = i[8726];
  assign o[8725] = i[8725];
  assign o[8724] = i[8724];
  assign o[8723] = i[8723];
  assign o[8722] = i[8722];
  assign o[8721] = i[8721];
  assign o[8720] = i[8720];
  assign o[8719] = i[8719];
  assign o[8718] = i[8718];
  assign o[8717] = i[8717];
  assign o[8716] = i[8716];
  assign o[8715] = i[8715];
  assign o[8714] = i[8714];
  assign o[8713] = i[8713];
  assign o[8712] = i[8712];
  assign o[8711] = i[8711];
  assign o[8710] = i[8710];
  assign o[8709] = i[8709];
  assign o[8708] = i[8708];
  assign o[8707] = i[8707];
  assign o[8706] = i[8706];
  assign o[8705] = i[8705];
  assign o[8704] = i[8704];
  assign o[8703] = i[8703];
  assign o[8702] = i[8702];
  assign o[8701] = i[8701];
  assign o[8700] = i[8700];
  assign o[8699] = i[8699];
  assign o[8698] = i[8698];
  assign o[8697] = i[8697];
  assign o[8696] = i[8696];
  assign o[8695] = i[8695];
  assign o[8694] = i[8694];
  assign o[8693] = i[8693];
  assign o[8692] = i[8692];
  assign o[8691] = i[8691];
  assign o[8690] = i[8690];
  assign o[8689] = i[8689];
  assign o[8688] = i[8688];
  assign o[8687] = i[8687];
  assign o[8686] = i[8686];
  assign o[8685] = i[8685];
  assign o[8684] = i[8684];
  assign o[8683] = i[8683];
  assign o[8682] = i[8682];
  assign o[8681] = i[8681];
  assign o[8680] = i[8680];
  assign o[8679] = i[8679];
  assign o[8678] = i[8678];
  assign o[8677] = i[8677];
  assign o[8676] = i[8676];
  assign o[8675] = i[8675];
  assign o[8674] = i[8674];
  assign o[8673] = i[8673];
  assign o[8672] = i[8672];
  assign o[8671] = i[8671];
  assign o[8670] = i[8670];
  assign o[8669] = i[8669];
  assign o[8668] = i[8668];
  assign o[8667] = i[8667];
  assign o[8666] = i[8666];
  assign o[8665] = i[8665];
  assign o[8664] = i[8664];
  assign o[8663] = i[8663];
  assign o[8662] = i[8662];
  assign o[8661] = i[8661];
  assign o[8660] = i[8660];
  assign o[8659] = i[8659];
  assign o[8658] = i[8658];
  assign o[8657] = i[8657];
  assign o[8656] = i[8656];
  assign o[8655] = i[8655];
  assign o[8654] = i[8654];
  assign o[8653] = i[8653];
  assign o[8652] = i[8652];
  assign o[8651] = i[8651];
  assign o[8650] = i[8650];
  assign o[8649] = i[8649];
  assign o[8648] = i[8648];
  assign o[8647] = i[8647];
  assign o[8646] = i[8646];
  assign o[8645] = i[8645];
  assign o[8644] = i[8644];
  assign o[8643] = i[8643];
  assign o[8642] = i[8642];
  assign o[8641] = i[8641];
  assign o[8640] = i[8640];
  assign o[8639] = i[8639];
  assign o[8638] = i[8638];
  assign o[8637] = i[8637];
  assign o[8636] = i[8636];
  assign o[8635] = i[8635];
  assign o[8634] = i[8634];
  assign o[8633] = i[8633];
  assign o[8632] = i[8632];
  assign o[8631] = i[8631];
  assign o[8630] = i[8630];
  assign o[8629] = i[8629];
  assign o[8628] = i[8628];
  assign o[8627] = i[8627];
  assign o[8626] = i[8626];
  assign o[8625] = i[8625];
  assign o[8624] = i[8624];
  assign o[8623] = i[8623];
  assign o[8622] = i[8622];
  assign o[8621] = i[8621];
  assign o[8620] = i[8620];
  assign o[8619] = i[8619];
  assign o[8618] = i[8618];
  assign o[8617] = i[8617];
  assign o[8616] = i[8616];
  assign o[8615] = i[8615];
  assign o[8614] = i[8614];
  assign o[8613] = i[8613];
  assign o[8612] = i[8612];
  assign o[8611] = i[8611];
  assign o[8610] = i[8610];
  assign o[8609] = i[8609];
  assign o[8608] = i[8608];
  assign o[8607] = i[8607];
  assign o[8606] = i[8606];
  assign o[8605] = i[8605];
  assign o[8604] = i[8604];
  assign o[8603] = i[8603];
  assign o[8602] = i[8602];
  assign o[8601] = i[8601];
  assign o[8600] = i[8600];
  assign o[8599] = i[8599];
  assign o[8598] = i[8598];
  assign o[8597] = i[8597];
  assign o[8596] = i[8596];
  assign o[8595] = i[8595];
  assign o[8594] = i[8594];
  assign o[8593] = i[8593];
  assign o[8592] = i[8592];
  assign o[8591] = i[8591];
  assign o[8590] = i[8590];
  assign o[8589] = i[8589];
  assign o[8588] = i[8588];
  assign o[8587] = i[8587];
  assign o[8586] = i[8586];
  assign o[8585] = i[8585];
  assign o[8584] = i[8584];
  assign o[8583] = i[8583];
  assign o[8582] = i[8582];
  assign o[8581] = i[8581];
  assign o[8580] = i[8580];
  assign o[8579] = i[8579];
  assign o[8578] = i[8578];
  assign o[8577] = i[8577];
  assign o[8576] = i[8576];
  assign o[8575] = i[8575];
  assign o[8574] = i[8574];
  assign o[8573] = i[8573];
  assign o[8572] = i[8572];
  assign o[8571] = i[8571];
  assign o[8570] = i[8570];
  assign o[8569] = i[8569];
  assign o[8568] = i[8568];
  assign o[8567] = i[8567];
  assign o[8566] = i[8566];
  assign o[8565] = i[8565];
  assign o[8564] = i[8564];
  assign o[8563] = i[8563];
  assign o[8562] = i[8562];
  assign o[8561] = i[8561];
  assign o[8560] = i[8560];
  assign o[8559] = i[8559];
  assign o[8558] = i[8558];
  assign o[8557] = i[8557];
  assign o[8556] = i[8556];
  assign o[8555] = i[8555];
  assign o[8554] = i[8554];
  assign o[8553] = i[8553];
  assign o[8552] = i[8552];
  assign o[8551] = i[8551];
  assign o[8550] = i[8550];
  assign o[8549] = i[8549];
  assign o[8548] = i[8548];
  assign o[8547] = i[8547];
  assign o[8546] = i[8546];
  assign o[8545] = i[8545];
  assign o[8544] = i[8544];
  assign o[8543] = i[8543];
  assign o[8542] = i[8542];
  assign o[8541] = i[8541];
  assign o[8540] = i[8540];
  assign o[8539] = i[8539];
  assign o[8538] = i[8538];
  assign o[8537] = i[8537];
  assign o[8536] = i[8536];
  assign o[8535] = i[8535];
  assign o[8534] = i[8534];
  assign o[8533] = i[8533];
  assign o[8532] = i[8532];
  assign o[8531] = i[8531];
  assign o[8530] = i[8530];
  assign o[8529] = i[8529];
  assign o[8528] = i[8528];
  assign o[8527] = i[8527];
  assign o[8526] = i[8526];
  assign o[8525] = i[8525];
  assign o[8524] = i[8524];
  assign o[8523] = i[8523];
  assign o[8522] = i[8522];
  assign o[8521] = i[8521];
  assign o[8520] = i[8520];
  assign o[8519] = i[8519];
  assign o[8518] = i[8518];
  assign o[8517] = i[8517];
  assign o[8516] = i[8516];
  assign o[8515] = i[8515];
  assign o[8514] = i[8514];
  assign o[8513] = i[8513];
  assign o[8512] = i[8512];
  assign o[8511] = i[8511];
  assign o[8510] = i[8510];
  assign o[8509] = i[8509];
  assign o[8508] = i[8508];
  assign o[8507] = i[8507];
  assign o[8506] = i[8506];
  assign o[8505] = i[8505];
  assign o[8504] = i[8504];
  assign o[8503] = i[8503];
  assign o[8502] = i[8502];
  assign o[8501] = i[8501];
  assign o[8500] = i[8500];
  assign o[8499] = i[8499];
  assign o[8498] = i[8498];
  assign o[8497] = i[8497];
  assign o[8496] = i[8496];
  assign o[8495] = i[8495];
  assign o[8494] = i[8494];
  assign o[8493] = i[8493];
  assign o[8492] = i[8492];
  assign o[8491] = i[8491];
  assign o[8490] = i[8490];
  assign o[8489] = i[8489];
  assign o[8488] = i[8488];
  assign o[8487] = i[8487];
  assign o[8486] = i[8486];
  assign o[8485] = i[8485];
  assign o[8484] = i[8484];
  assign o[8483] = i[8483];
  assign o[8482] = i[8482];
  assign o[8481] = i[8481];
  assign o[8480] = i[8480];
  assign o[8479] = i[8479];
  assign o[8478] = i[8478];
  assign o[8477] = i[8477];
  assign o[8476] = i[8476];
  assign o[8475] = i[8475];
  assign o[8474] = i[8474];
  assign o[8473] = i[8473];
  assign o[8472] = i[8472];
  assign o[8471] = i[8471];
  assign o[8470] = i[8470];
  assign o[8469] = i[8469];
  assign o[8468] = i[8468];
  assign o[8467] = i[8467];
  assign o[8466] = i[8466];
  assign o[8465] = i[8465];
  assign o[8464] = i[8464];
  assign o[8463] = i[8463];
  assign o[8462] = i[8462];
  assign o[8461] = i[8461];
  assign o[8460] = i[8460];
  assign o[8459] = i[8459];
  assign o[8458] = i[8458];
  assign o[8457] = i[8457];
  assign o[8456] = i[8456];
  assign o[8455] = i[8455];
  assign o[8454] = i[8454];
  assign o[8453] = i[8453];
  assign o[8452] = i[8452];
  assign o[8451] = i[8451];
  assign o[8450] = i[8450];
  assign o[8449] = i[8449];
  assign o[8448] = i[8448];
  assign o[8447] = i[8447];
  assign o[8446] = i[8446];
  assign o[8445] = i[8445];
  assign o[8444] = i[8444];
  assign o[8443] = i[8443];
  assign o[8442] = i[8442];
  assign o[8441] = i[8441];
  assign o[8440] = i[8440];
  assign o[8439] = i[8439];
  assign o[8438] = i[8438];
  assign o[8437] = i[8437];
  assign o[8436] = i[8436];
  assign o[8435] = i[8435];
  assign o[8434] = i[8434];
  assign o[8433] = i[8433];
  assign o[8432] = i[8432];
  assign o[8431] = i[8431];
  assign o[8430] = i[8430];
  assign o[8429] = i[8429];
  assign o[8428] = i[8428];
  assign o[8427] = i[8427];
  assign o[8426] = i[8426];
  assign o[8425] = i[8425];
  assign o[8424] = i[8424];
  assign o[8423] = i[8423];
  assign o[8422] = i[8422];
  assign o[8421] = i[8421];
  assign o[8420] = i[8420];
  assign o[8419] = i[8419];
  assign o[8418] = i[8418];
  assign o[8417] = i[8417];
  assign o[8416] = i[8416];
  assign o[8415] = i[8415];
  assign o[8414] = i[8414];
  assign o[8413] = i[8413];
  assign o[8412] = i[8412];
  assign o[8411] = i[8411];
  assign o[8410] = i[8410];
  assign o[8409] = i[8409];
  assign o[8408] = i[8408];
  assign o[8407] = i[8407];
  assign o[8406] = i[8406];
  assign o[8405] = i[8405];
  assign o[8404] = i[8404];
  assign o[8403] = i[8403];
  assign o[8402] = i[8402];
  assign o[8401] = i[8401];
  assign o[8400] = i[8400];
  assign o[8399] = i[8399];
  assign o[8398] = i[8398];
  assign o[8397] = i[8397];
  assign o[8396] = i[8396];
  assign o[8395] = i[8395];
  assign o[8394] = i[8394];
  assign o[8393] = i[8393];
  assign o[8392] = i[8392];
  assign o[8391] = i[8391];
  assign o[8390] = i[8390];
  assign o[8389] = i[8389];
  assign o[8388] = i[8388];
  assign o[8387] = i[8387];
  assign o[8386] = i[8386];
  assign o[8385] = i[8385];
  assign o[8384] = i[8384];
  assign o[8383] = i[8383];
  assign o[8382] = i[8382];
  assign o[8381] = i[8381];
  assign o[8380] = i[8380];
  assign o[8379] = i[8379];
  assign o[8378] = i[8378];
  assign o[8377] = i[8377];
  assign o[8376] = i[8376];
  assign o[8375] = i[8375];
  assign o[8374] = i[8374];
  assign o[8373] = i[8373];
  assign o[8372] = i[8372];
  assign o[8371] = i[8371];
  assign o[8370] = i[8370];
  assign o[8369] = i[8369];
  assign o[8368] = i[8368];
  assign o[8367] = i[8367];
  assign o[8366] = i[8366];
  assign o[8365] = i[8365];
  assign o[8364] = i[8364];
  assign o[8363] = i[8363];
  assign o[8362] = i[8362];
  assign o[8361] = i[8361];
  assign o[8360] = i[8360];
  assign o[8359] = i[8359];
  assign o[8358] = i[8358];
  assign o[8357] = i[8357];
  assign o[8356] = i[8356];
  assign o[8355] = i[8355];
  assign o[8354] = i[8354];
  assign o[8353] = i[8353];
  assign o[8352] = i[8352];
  assign o[8351] = i[8351];
  assign o[8350] = i[8350];
  assign o[8349] = i[8349];
  assign o[8348] = i[8348];
  assign o[8347] = i[8347];
  assign o[8346] = i[8346];
  assign o[8345] = i[8345];
  assign o[8344] = i[8344];
  assign o[8343] = i[8343];
  assign o[8342] = i[8342];
  assign o[8341] = i[8341];
  assign o[8340] = i[8340];
  assign o[8339] = i[8339];
  assign o[8338] = i[8338];
  assign o[8337] = i[8337];
  assign o[8336] = i[8336];
  assign o[8335] = i[8335];
  assign o[8334] = i[8334];
  assign o[8333] = i[8333];
  assign o[8332] = i[8332];
  assign o[8331] = i[8331];
  assign o[8330] = i[8330];
  assign o[8329] = i[8329];
  assign o[8328] = i[8328];
  assign o[8327] = i[8327];
  assign o[8326] = i[8326];
  assign o[8325] = i[8325];
  assign o[8324] = i[8324];
  assign o[8323] = i[8323];
  assign o[8322] = i[8322];
  assign o[8321] = i[8321];
  assign o[8320] = i[8320];
  assign o[8319] = i[8319];
  assign o[8318] = i[8318];
  assign o[8317] = i[8317];
  assign o[8316] = i[8316];
  assign o[8315] = i[8315];
  assign o[8314] = i[8314];
  assign o[8313] = i[8313];
  assign o[8312] = i[8312];
  assign o[8311] = i[8311];
  assign o[8310] = i[8310];
  assign o[8309] = i[8309];
  assign o[8308] = i[8308];
  assign o[8307] = i[8307];
  assign o[8306] = i[8306];
  assign o[8305] = i[8305];
  assign o[8304] = i[8304];
  assign o[8303] = i[8303];
  assign o[8302] = i[8302];
  assign o[8301] = i[8301];
  assign o[8300] = i[8300];
  assign o[8299] = i[8299];
  assign o[8298] = i[8298];
  assign o[8297] = i[8297];
  assign o[8296] = i[8296];
  assign o[8295] = i[8295];
  assign o[8294] = i[8294];
  assign o[8293] = i[8293];
  assign o[8292] = i[8292];
  assign o[8291] = i[8291];
  assign o[8290] = i[8290];
  assign o[8289] = i[8289];
  assign o[8288] = i[8288];
  assign o[8287] = i[8287];
  assign o[8286] = i[8286];
  assign o[8285] = i[8285];
  assign o[8284] = i[8284];
  assign o[8283] = i[8283];
  assign o[8282] = i[8282];
  assign o[8281] = i[8281];
  assign o[8280] = i[8280];
  assign o[8279] = i[8279];
  assign o[8278] = i[8278];
  assign o[8277] = i[8277];
  assign o[8276] = i[8276];
  assign o[8275] = i[8275];
  assign o[8274] = i[8274];
  assign o[8273] = i[8273];
  assign o[8272] = i[8272];
  assign o[8271] = i[8271];
  assign o[8270] = i[8270];
  assign o[8269] = i[8269];
  assign o[8268] = i[8268];
  assign o[8267] = i[8267];
  assign o[8266] = i[8266];
  assign o[8265] = i[8265];
  assign o[8264] = i[8264];
  assign o[8263] = i[8263];
  assign o[8262] = i[8262];
  assign o[8261] = i[8261];
  assign o[8260] = i[8260];
  assign o[8259] = i[8259];
  assign o[8258] = i[8258];
  assign o[8257] = i[8257];
  assign o[8256] = i[8256];
  assign o[8255] = i[8255];
  assign o[8254] = i[8254];
  assign o[8253] = i[8253];
  assign o[8252] = i[8252];
  assign o[8251] = i[8251];
  assign o[8250] = i[8250];
  assign o[8249] = i[8249];
  assign o[8248] = i[8248];
  assign o[8247] = i[8247];
  assign o[8246] = i[8246];
  assign o[8245] = i[8245];
  assign o[8244] = i[8244];
  assign o[8243] = i[8243];
  assign o[8242] = i[8242];
  assign o[8241] = i[8241];
  assign o[8240] = i[8240];
  assign o[8239] = i[8239];
  assign o[8238] = i[8238];
  assign o[8237] = i[8237];
  assign o[8236] = i[8236];
  assign o[8235] = i[8235];
  assign o[8234] = i[8234];
  assign o[8233] = i[8233];
  assign o[8232] = i[8232];
  assign o[8231] = i[8231];
  assign o[8230] = i[8230];
  assign o[8229] = i[8229];
  assign o[8228] = i[8228];
  assign o[8227] = i[8227];
  assign o[8226] = i[8226];
  assign o[8225] = i[8225];
  assign o[8224] = i[8224];
  assign o[8223] = i[8223];
  assign o[8222] = i[8222];
  assign o[8221] = i[8221];
  assign o[8220] = i[8220];
  assign o[8219] = i[8219];
  assign o[8218] = i[8218];
  assign o[8217] = i[8217];
  assign o[8216] = i[8216];
  assign o[8215] = i[8215];
  assign o[8214] = i[8214];
  assign o[8213] = i[8213];
  assign o[8212] = i[8212];
  assign o[8211] = i[8211];
  assign o[8210] = i[8210];
  assign o[8209] = i[8209];
  assign o[8208] = i[8208];
  assign o[8207] = i[8207];
  assign o[8206] = i[8206];
  assign o[8205] = i[8205];
  assign o[8204] = i[8204];
  assign o[8203] = i[8203];
  assign o[8202] = i[8202];
  assign o[8201] = i[8201];
  assign o[8200] = i[8200];
  assign o[8199] = i[8199];
  assign o[8198] = i[8198];
  assign o[8197] = i[8197];
  assign o[8196] = i[8196];
  assign o[8195] = i[8195];
  assign o[8194] = i[8194];
  assign o[8193] = i[8193];
  assign o[8192] = i[8192];
  assign o[8191] = i[8191];
  assign o[8190] = i[8190];
  assign o[8189] = i[8189];
  assign o[8188] = i[8188];
  assign o[8187] = i[8187];
  assign o[8186] = i[8186];
  assign o[8185] = i[8185];
  assign o[8184] = i[8184];
  assign o[8183] = i[8183];
  assign o[8182] = i[8182];
  assign o[8181] = i[8181];
  assign o[8180] = i[8180];
  assign o[8179] = i[8179];
  assign o[8178] = i[8178];
  assign o[8177] = i[8177];
  assign o[8176] = i[8176];
  assign o[8175] = i[8175];
  assign o[8174] = i[8174];
  assign o[8173] = i[8173];
  assign o[8172] = i[8172];
  assign o[8171] = i[8171];
  assign o[8170] = i[8170];
  assign o[8169] = i[8169];
  assign o[8168] = i[8168];
  assign o[8167] = i[8167];
  assign o[8166] = i[8166];
  assign o[8165] = i[8165];
  assign o[8164] = i[8164];
  assign o[8163] = i[8163];
  assign o[8162] = i[8162];
  assign o[8161] = i[8161];
  assign o[8160] = i[8160];
  assign o[8159] = i[8159];
  assign o[8158] = i[8158];
  assign o[8157] = i[8157];
  assign o[8156] = i[8156];
  assign o[8155] = i[8155];
  assign o[8154] = i[8154];
  assign o[8153] = i[8153];
  assign o[8152] = i[8152];
  assign o[8151] = i[8151];
  assign o[8150] = i[8150];
  assign o[8149] = i[8149];
  assign o[8148] = i[8148];
  assign o[8147] = i[8147];
  assign o[8146] = i[8146];
  assign o[8145] = i[8145];
  assign o[8144] = i[8144];
  assign o[8143] = i[8143];
  assign o[8142] = i[8142];
  assign o[8141] = i[8141];
  assign o[8140] = i[8140];
  assign o[8139] = i[8139];
  assign o[8138] = i[8138];
  assign o[8137] = i[8137];
  assign o[8136] = i[8136];
  assign o[8135] = i[8135];
  assign o[8134] = i[8134];
  assign o[8133] = i[8133];
  assign o[8132] = i[8132];
  assign o[8131] = i[8131];
  assign o[8130] = i[8130];
  assign o[8129] = i[8129];
  assign o[8128] = i[8128];
  assign o[8127] = i[8127];
  assign o[8126] = i[8126];
  assign o[8125] = i[8125];
  assign o[8124] = i[8124];
  assign o[8123] = i[8123];
  assign o[8122] = i[8122];
  assign o[8121] = i[8121];
  assign o[8120] = i[8120];
  assign o[8119] = i[8119];
  assign o[8118] = i[8118];
  assign o[8117] = i[8117];
  assign o[8116] = i[8116];
  assign o[8115] = i[8115];
  assign o[8114] = i[8114];
  assign o[8113] = i[8113];
  assign o[8112] = i[8112];
  assign o[8111] = i[8111];
  assign o[8110] = i[8110];
  assign o[8109] = i[8109];
  assign o[8108] = i[8108];
  assign o[8107] = i[8107];
  assign o[8106] = i[8106];
  assign o[8105] = i[8105];
  assign o[8104] = i[8104];
  assign o[8103] = i[8103];
  assign o[8102] = i[8102];
  assign o[8101] = i[8101];
  assign o[8100] = i[8100];
  assign o[8099] = i[8099];
  assign o[8098] = i[8098];
  assign o[8097] = i[8097];
  assign o[8096] = i[8096];
  assign o[8095] = i[8095];
  assign o[8094] = i[8094];
  assign o[8093] = i[8093];
  assign o[8092] = i[8092];
  assign o[8091] = i[8091];
  assign o[8090] = i[8090];
  assign o[8089] = i[8089];
  assign o[8088] = i[8088];
  assign o[8087] = i[8087];
  assign o[8086] = i[8086];
  assign o[8085] = i[8085];
  assign o[8084] = i[8084];
  assign o[8083] = i[8083];
  assign o[8082] = i[8082];
  assign o[8081] = i[8081];
  assign o[8080] = i[8080];
  assign o[8079] = i[8079];
  assign o[8078] = i[8078];
  assign o[8077] = i[8077];
  assign o[8076] = i[8076];
  assign o[8075] = i[8075];
  assign o[8074] = i[8074];
  assign o[8073] = i[8073];
  assign o[8072] = i[8072];
  assign o[8071] = i[8071];
  assign o[8070] = i[8070];
  assign o[8069] = i[8069];
  assign o[8068] = i[8068];
  assign o[8067] = i[8067];
  assign o[8066] = i[8066];
  assign o[8065] = i[8065];
  assign o[8064] = i[8064];
  assign o[8063] = i[8063];
  assign o[8062] = i[8062];
  assign o[8061] = i[8061];
  assign o[8060] = i[8060];
  assign o[8059] = i[8059];
  assign o[8058] = i[8058];
  assign o[8057] = i[8057];
  assign o[8056] = i[8056];
  assign o[8055] = i[8055];
  assign o[8054] = i[8054];
  assign o[8053] = i[8053];
  assign o[8052] = i[8052];
  assign o[8051] = i[8051];
  assign o[8050] = i[8050];
  assign o[8049] = i[8049];
  assign o[8048] = i[8048];
  assign o[8047] = i[8047];
  assign o[8046] = i[8046];
  assign o[8045] = i[8045];
  assign o[8044] = i[8044];
  assign o[8043] = i[8043];
  assign o[8042] = i[8042];
  assign o[8041] = i[8041];
  assign o[8040] = i[8040];
  assign o[8039] = i[8039];
  assign o[8038] = i[8038];
  assign o[8037] = i[8037];
  assign o[8036] = i[8036];
  assign o[8035] = i[8035];
  assign o[8034] = i[8034];
  assign o[8033] = i[8033];
  assign o[8032] = i[8032];
  assign o[8031] = i[8031];
  assign o[8030] = i[8030];
  assign o[8029] = i[8029];
  assign o[8028] = i[8028];
  assign o[8027] = i[8027];
  assign o[8026] = i[8026];
  assign o[8025] = i[8025];
  assign o[8024] = i[8024];
  assign o[8023] = i[8023];
  assign o[8022] = i[8022];
  assign o[8021] = i[8021];
  assign o[8020] = i[8020];
  assign o[8019] = i[8019];
  assign o[8018] = i[8018];
  assign o[8017] = i[8017];
  assign o[8016] = i[8016];
  assign o[8015] = i[8015];
  assign o[8014] = i[8014];
  assign o[8013] = i[8013];
  assign o[8012] = i[8012];
  assign o[8011] = i[8011];
  assign o[8010] = i[8010];
  assign o[8009] = i[8009];
  assign o[8008] = i[8008];
  assign o[8007] = i[8007];
  assign o[8006] = i[8006];
  assign o[8005] = i[8005];
  assign o[8004] = i[8004];
  assign o[8003] = i[8003];
  assign o[8002] = i[8002];
  assign o[8001] = i[8001];
  assign o[8000] = i[8000];
  assign o[7999] = i[7999];
  assign o[7998] = i[7998];
  assign o[7997] = i[7997];
  assign o[7996] = i[7996];
  assign o[7995] = i[7995];
  assign o[7994] = i[7994];
  assign o[7993] = i[7993];
  assign o[7992] = i[7992];
  assign o[7991] = i[7991];
  assign o[7990] = i[7990];
  assign o[7989] = i[7989];
  assign o[7988] = i[7988];
  assign o[7987] = i[7987];
  assign o[7986] = i[7986];
  assign o[7985] = i[7985];
  assign o[7984] = i[7984];
  assign o[7983] = i[7983];
  assign o[7982] = i[7982];
  assign o[7981] = i[7981];
  assign o[7980] = i[7980];
  assign o[7979] = i[7979];
  assign o[7978] = i[7978];
  assign o[7977] = i[7977];
  assign o[7976] = i[7976];
  assign o[7975] = i[7975];
  assign o[7974] = i[7974];
  assign o[7973] = i[7973];
  assign o[7972] = i[7972];
  assign o[7971] = i[7971];
  assign o[7970] = i[7970];
  assign o[7969] = i[7969];
  assign o[7968] = i[7968];
  assign o[7967] = i[7967];
  assign o[7966] = i[7966];
  assign o[7965] = i[7965];
  assign o[7964] = i[7964];
  assign o[7963] = i[7963];
  assign o[7962] = i[7962];
  assign o[7961] = i[7961];
  assign o[7960] = i[7960];
  assign o[7959] = i[7959];
  assign o[7958] = i[7958];
  assign o[7957] = i[7957];
  assign o[7956] = i[7956];
  assign o[7955] = i[7955];
  assign o[7954] = i[7954];
  assign o[7953] = i[7953];
  assign o[7952] = i[7952];
  assign o[7951] = i[7951];
  assign o[7950] = i[7950];
  assign o[7949] = i[7949];
  assign o[7948] = i[7948];
  assign o[7947] = i[7947];
  assign o[7946] = i[7946];
  assign o[7945] = i[7945];
  assign o[7944] = i[7944];
  assign o[7943] = i[7943];
  assign o[7942] = i[7942];
  assign o[7941] = i[7941];
  assign o[7940] = i[7940];
  assign o[7939] = i[7939];
  assign o[7938] = i[7938];
  assign o[7937] = i[7937];
  assign o[7936] = i[7936];
  assign o[7935] = i[7935];
  assign o[7934] = i[7934];
  assign o[7933] = i[7933];
  assign o[7932] = i[7932];
  assign o[7931] = i[7931];
  assign o[7930] = i[7930];
  assign o[7929] = i[7929];
  assign o[7928] = i[7928];
  assign o[7927] = i[7927];
  assign o[7926] = i[7926];
  assign o[7925] = i[7925];
  assign o[7924] = i[7924];
  assign o[7923] = i[7923];
  assign o[7922] = i[7922];
  assign o[7921] = i[7921];
  assign o[7920] = i[7920];
  assign o[7919] = i[7919];
  assign o[7918] = i[7918];
  assign o[7917] = i[7917];
  assign o[7916] = i[7916];
  assign o[7915] = i[7915];
  assign o[7914] = i[7914];
  assign o[7913] = i[7913];
  assign o[7912] = i[7912];
  assign o[7911] = i[7911];
  assign o[7910] = i[7910];
  assign o[7909] = i[7909];
  assign o[7908] = i[7908];
  assign o[7907] = i[7907];
  assign o[7906] = i[7906];
  assign o[7905] = i[7905];
  assign o[7904] = i[7904];
  assign o[7903] = i[7903];
  assign o[7902] = i[7902];
  assign o[7901] = i[7901];
  assign o[7900] = i[7900];
  assign o[7899] = i[7899];
  assign o[7898] = i[7898];
  assign o[7897] = i[7897];
  assign o[7896] = i[7896];
  assign o[7895] = i[7895];
  assign o[7894] = i[7894];
  assign o[7893] = i[7893];
  assign o[7892] = i[7892];
  assign o[7891] = i[7891];
  assign o[7890] = i[7890];
  assign o[7889] = i[7889];
  assign o[7888] = i[7888];
  assign o[7887] = i[7887];
  assign o[7886] = i[7886];
  assign o[7885] = i[7885];
  assign o[7884] = i[7884];
  assign o[7883] = i[7883];
  assign o[7882] = i[7882];
  assign o[7881] = i[7881];
  assign o[7880] = i[7880];
  assign o[7879] = i[7879];
  assign o[7878] = i[7878];
  assign o[7877] = i[7877];
  assign o[7876] = i[7876];
  assign o[7875] = i[7875];
  assign o[7874] = i[7874];
  assign o[7873] = i[7873];
  assign o[7872] = i[7872];
  assign o[7871] = i[7871];
  assign o[7870] = i[7870];
  assign o[7869] = i[7869];
  assign o[7868] = i[7868];
  assign o[7867] = i[7867];
  assign o[7866] = i[7866];
  assign o[7865] = i[7865];
  assign o[7864] = i[7864];
  assign o[7863] = i[7863];
  assign o[7862] = i[7862];
  assign o[7861] = i[7861];
  assign o[7860] = i[7860];
  assign o[7859] = i[7859];
  assign o[7858] = i[7858];
  assign o[7857] = i[7857];
  assign o[7856] = i[7856];
  assign o[7855] = i[7855];
  assign o[7854] = i[7854];
  assign o[7853] = i[7853];
  assign o[7852] = i[7852];
  assign o[7851] = i[7851];
  assign o[7850] = i[7850];
  assign o[7849] = i[7849];
  assign o[7848] = i[7848];
  assign o[7847] = i[7847];
  assign o[7846] = i[7846];
  assign o[7845] = i[7845];
  assign o[7844] = i[7844];
  assign o[7843] = i[7843];
  assign o[7842] = i[7842];
  assign o[7841] = i[7841];
  assign o[7840] = i[7840];
  assign o[7839] = i[7839];
  assign o[7838] = i[7838];
  assign o[7837] = i[7837];
  assign o[7836] = i[7836];
  assign o[7835] = i[7835];
  assign o[7834] = i[7834];
  assign o[7833] = i[7833];
  assign o[7832] = i[7832];
  assign o[7831] = i[7831];
  assign o[7830] = i[7830];
  assign o[7829] = i[7829];
  assign o[7828] = i[7828];
  assign o[7827] = i[7827];
  assign o[7826] = i[7826];
  assign o[7825] = i[7825];
  assign o[7824] = i[7824];
  assign o[7823] = i[7823];
  assign o[7822] = i[7822];
  assign o[7821] = i[7821];
  assign o[7820] = i[7820];
  assign o[7819] = i[7819];
  assign o[7818] = i[7818];
  assign o[7817] = i[7817];
  assign o[7816] = i[7816];
  assign o[7815] = i[7815];
  assign o[7814] = i[7814];
  assign o[7813] = i[7813];
  assign o[7812] = i[7812];
  assign o[7811] = i[7811];
  assign o[7810] = i[7810];
  assign o[7809] = i[7809];
  assign o[7808] = i[7808];
  assign o[7807] = i[7807];
  assign o[7806] = i[7806];
  assign o[7805] = i[7805];
  assign o[7804] = i[7804];
  assign o[7803] = i[7803];
  assign o[7802] = i[7802];
  assign o[7801] = i[7801];
  assign o[7800] = i[7800];
  assign o[7799] = i[7799];
  assign o[7798] = i[7798];
  assign o[7797] = i[7797];
  assign o[7796] = i[7796];
  assign o[7795] = i[7795];
  assign o[7794] = i[7794];
  assign o[7793] = i[7793];
  assign o[7792] = i[7792];
  assign o[7791] = i[7791];
  assign o[7790] = i[7790];
  assign o[7789] = i[7789];
  assign o[7788] = i[7788];
  assign o[7787] = i[7787];
  assign o[7786] = i[7786];
  assign o[7785] = i[7785];
  assign o[7784] = i[7784];
  assign o[7783] = i[7783];
  assign o[7782] = i[7782];
  assign o[7781] = i[7781];
  assign o[7780] = i[7780];
  assign o[7779] = i[7779];
  assign o[7778] = i[7778];
  assign o[7777] = i[7777];
  assign o[7776] = i[7776];
  assign o[7775] = i[7775];
  assign o[7774] = i[7774];
  assign o[7773] = i[7773];
  assign o[7772] = i[7772];
  assign o[7771] = i[7771];
  assign o[7770] = i[7770];
  assign o[7769] = i[7769];
  assign o[7768] = i[7768];
  assign o[7767] = i[7767];
  assign o[7766] = i[7766];
  assign o[7765] = i[7765];
  assign o[7764] = i[7764];
  assign o[7763] = i[7763];
  assign o[7762] = i[7762];
  assign o[7761] = i[7761];
  assign o[7760] = i[7760];
  assign o[7759] = i[7759];
  assign o[7758] = i[7758];
  assign o[7757] = i[7757];
  assign o[7756] = i[7756];
  assign o[7755] = i[7755];
  assign o[7754] = i[7754];
  assign o[7753] = i[7753];
  assign o[7752] = i[7752];
  assign o[7751] = i[7751];
  assign o[7750] = i[7750];
  assign o[7749] = i[7749];
  assign o[7748] = i[7748];
  assign o[7747] = i[7747];
  assign o[7746] = i[7746];
  assign o[7745] = i[7745];
  assign o[7744] = i[7744];
  assign o[7743] = i[7743];
  assign o[7742] = i[7742];
  assign o[7741] = i[7741];
  assign o[7740] = i[7740];
  assign o[7739] = i[7739];
  assign o[7738] = i[7738];
  assign o[7737] = i[7737];
  assign o[7736] = i[7736];
  assign o[7735] = i[7735];
  assign o[7734] = i[7734];
  assign o[7733] = i[7733];
  assign o[7732] = i[7732];
  assign o[7731] = i[7731];
  assign o[7730] = i[7730];
  assign o[7729] = i[7729];
  assign o[7728] = i[7728];
  assign o[7727] = i[7727];
  assign o[7726] = i[7726];
  assign o[7725] = i[7725];
  assign o[7724] = i[7724];
  assign o[7723] = i[7723];
  assign o[7722] = i[7722];
  assign o[7721] = i[7721];
  assign o[7720] = i[7720];
  assign o[7719] = i[7719];
  assign o[7718] = i[7718];
  assign o[7717] = i[7717];
  assign o[7716] = i[7716];
  assign o[7715] = i[7715];
  assign o[7714] = i[7714];
  assign o[7713] = i[7713];
  assign o[7712] = i[7712];
  assign o[7711] = i[7711];
  assign o[7710] = i[7710];
  assign o[7709] = i[7709];
  assign o[7708] = i[7708];
  assign o[7707] = i[7707];
  assign o[7706] = i[7706];
  assign o[7705] = i[7705];
  assign o[7704] = i[7704];
  assign o[7703] = i[7703];
  assign o[7702] = i[7702];
  assign o[7701] = i[7701];
  assign o[7700] = i[7700];
  assign o[7699] = i[7699];
  assign o[7698] = i[7698];
  assign o[7697] = i[7697];
  assign o[7696] = i[7696];
  assign o[7695] = i[7695];
  assign o[7694] = i[7694];
  assign o[7693] = i[7693];
  assign o[7692] = i[7692];
  assign o[7691] = i[7691];
  assign o[7690] = i[7690];
  assign o[7689] = i[7689];
  assign o[7688] = i[7688];
  assign o[7687] = i[7687];
  assign o[7686] = i[7686];
  assign o[7685] = i[7685];
  assign o[7684] = i[7684];
  assign o[7683] = i[7683];
  assign o[7682] = i[7682];
  assign o[7681] = i[7681];
  assign o[7680] = i[7680];
  assign o[7679] = i[7679];
  assign o[7678] = i[7678];
  assign o[7677] = i[7677];
  assign o[7676] = i[7676];
  assign o[7675] = i[7675];
  assign o[7674] = i[7674];
  assign o[7673] = i[7673];
  assign o[7672] = i[7672];
  assign o[7671] = i[7671];
  assign o[7670] = i[7670];
  assign o[7669] = i[7669];
  assign o[7668] = i[7668];
  assign o[7667] = i[7667];
  assign o[7666] = i[7666];
  assign o[7665] = i[7665];
  assign o[7664] = i[7664];
  assign o[7663] = i[7663];
  assign o[7662] = i[7662];
  assign o[7661] = i[7661];
  assign o[7660] = i[7660];
  assign o[7659] = i[7659];
  assign o[7658] = i[7658];
  assign o[7657] = i[7657];
  assign o[7656] = i[7656];
  assign o[7655] = i[7655];
  assign o[7654] = i[7654];
  assign o[7653] = i[7653];
  assign o[7652] = i[7652];
  assign o[7651] = i[7651];
  assign o[7650] = i[7650];
  assign o[7649] = i[7649];
  assign o[7648] = i[7648];
  assign o[7647] = i[7647];
  assign o[7646] = i[7646];
  assign o[7645] = i[7645];
  assign o[7644] = i[7644];
  assign o[7643] = i[7643];
  assign o[7642] = i[7642];
  assign o[7641] = i[7641];
  assign o[7640] = i[7640];
  assign o[7639] = i[7639];
  assign o[7638] = i[7638];
  assign o[7637] = i[7637];
  assign o[7636] = i[7636];
  assign o[7635] = i[7635];
  assign o[7634] = i[7634];
  assign o[7633] = i[7633];
  assign o[7632] = i[7632];
  assign o[7631] = i[7631];
  assign o[7630] = i[7630];
  assign o[7629] = i[7629];
  assign o[7628] = i[7628];
  assign o[7627] = i[7627];
  assign o[7626] = i[7626];
  assign o[7625] = i[7625];
  assign o[7624] = i[7624];
  assign o[7623] = i[7623];
  assign o[7622] = i[7622];
  assign o[7621] = i[7621];
  assign o[7620] = i[7620];
  assign o[7619] = i[7619];
  assign o[7618] = i[7618];
  assign o[7617] = i[7617];
  assign o[7616] = i[7616];
  assign o[7615] = i[7615];
  assign o[7614] = i[7614];
  assign o[7613] = i[7613];
  assign o[7612] = i[7612];
  assign o[7611] = i[7611];
  assign o[7610] = i[7610];
  assign o[7609] = i[7609];
  assign o[7608] = i[7608];
  assign o[7607] = i[7607];
  assign o[7606] = i[7606];
  assign o[7605] = i[7605];
  assign o[7604] = i[7604];
  assign o[7603] = i[7603];
  assign o[7602] = i[7602];
  assign o[7601] = i[7601];
  assign o[7600] = i[7600];
  assign o[7599] = i[7599];
  assign o[7598] = i[7598];
  assign o[7597] = i[7597];
  assign o[7596] = i[7596];
  assign o[7595] = i[7595];
  assign o[7594] = i[7594];
  assign o[7593] = i[7593];
  assign o[7592] = i[7592];
  assign o[7591] = i[7591];
  assign o[7590] = i[7590];
  assign o[7589] = i[7589];
  assign o[7588] = i[7588];
  assign o[7587] = i[7587];
  assign o[7586] = i[7586];
  assign o[7585] = i[7585];
  assign o[7584] = i[7584];
  assign o[7583] = i[7583];
  assign o[7582] = i[7582];
  assign o[7581] = i[7581];
  assign o[7580] = i[7580];
  assign o[7579] = i[7579];
  assign o[7578] = i[7578];
  assign o[7577] = i[7577];
  assign o[7576] = i[7576];
  assign o[7575] = i[7575];
  assign o[7574] = i[7574];
  assign o[7573] = i[7573];
  assign o[7572] = i[7572];
  assign o[7571] = i[7571];
  assign o[7570] = i[7570];
  assign o[7569] = i[7569];
  assign o[7568] = i[7568];
  assign o[7567] = i[7567];
  assign o[7566] = i[7566];
  assign o[7565] = i[7565];
  assign o[7564] = i[7564];
  assign o[7563] = i[7563];
  assign o[7562] = i[7562];
  assign o[7561] = i[7561];
  assign o[7560] = i[7560];
  assign o[7559] = i[7559];
  assign o[7558] = i[7558];
  assign o[7557] = i[7557];
  assign o[7556] = i[7556];
  assign o[7555] = i[7555];
  assign o[7554] = i[7554];
  assign o[7553] = i[7553];
  assign o[7552] = i[7552];
  assign o[7551] = i[7551];
  assign o[7550] = i[7550];
  assign o[7549] = i[7549];
  assign o[7548] = i[7548];
  assign o[7547] = i[7547];
  assign o[7546] = i[7546];
  assign o[7545] = i[7545];
  assign o[7544] = i[7544];
  assign o[7543] = i[7543];
  assign o[7542] = i[7542];
  assign o[7541] = i[7541];
  assign o[7540] = i[7540];
  assign o[7539] = i[7539];
  assign o[7538] = i[7538];
  assign o[7537] = i[7537];
  assign o[7536] = i[7536];
  assign o[7535] = i[7535];
  assign o[7534] = i[7534];
  assign o[7533] = i[7533];
  assign o[7532] = i[7532];
  assign o[7531] = i[7531];
  assign o[7530] = i[7530];
  assign o[7529] = i[7529];
  assign o[7528] = i[7528];
  assign o[7527] = i[7527];
  assign o[7526] = i[7526];
  assign o[7525] = i[7525];
  assign o[7524] = i[7524];
  assign o[7523] = i[7523];
  assign o[7522] = i[7522];
  assign o[7521] = i[7521];
  assign o[7520] = i[7520];
  assign o[7519] = i[7519];
  assign o[7518] = i[7518];
  assign o[7517] = i[7517];
  assign o[7516] = i[7516];
  assign o[7515] = i[7515];
  assign o[7514] = i[7514];
  assign o[7513] = i[7513];
  assign o[7512] = i[7512];
  assign o[7511] = i[7511];
  assign o[7510] = i[7510];
  assign o[7509] = i[7509];
  assign o[7508] = i[7508];
  assign o[7507] = i[7507];
  assign o[7506] = i[7506];
  assign o[7505] = i[7505];
  assign o[7504] = i[7504];
  assign o[7503] = i[7503];
  assign o[7502] = i[7502];
  assign o[7501] = i[7501];
  assign o[7500] = i[7500];
  assign o[7499] = i[7499];
  assign o[7498] = i[7498];
  assign o[7497] = i[7497];
  assign o[7496] = i[7496];
  assign o[7495] = i[7495];
  assign o[7494] = i[7494];
  assign o[7493] = i[7493];
  assign o[7492] = i[7492];
  assign o[7491] = i[7491];
  assign o[7490] = i[7490];
  assign o[7489] = i[7489];
  assign o[7488] = i[7488];
  assign o[7487] = i[7487];
  assign o[7486] = i[7486];
  assign o[7485] = i[7485];
  assign o[7484] = i[7484];
  assign o[7483] = i[7483];
  assign o[7482] = i[7482];
  assign o[7481] = i[7481];
  assign o[7480] = i[7480];
  assign o[7479] = i[7479];
  assign o[7478] = i[7478];
  assign o[7477] = i[7477];
  assign o[7476] = i[7476];
  assign o[7475] = i[7475];
  assign o[7474] = i[7474];
  assign o[7473] = i[7473];
  assign o[7472] = i[7472];
  assign o[7471] = i[7471];
  assign o[7470] = i[7470];
  assign o[7469] = i[7469];
  assign o[7468] = i[7468];
  assign o[7467] = i[7467];
  assign o[7466] = i[7466];
  assign o[7465] = i[7465];
  assign o[7464] = i[7464];
  assign o[7463] = i[7463];
  assign o[7462] = i[7462];
  assign o[7461] = i[7461];
  assign o[7460] = i[7460];
  assign o[7459] = i[7459];
  assign o[7458] = i[7458];
  assign o[7457] = i[7457];
  assign o[7456] = i[7456];
  assign o[7455] = i[7455];
  assign o[7454] = i[7454];
  assign o[7453] = i[7453];
  assign o[7452] = i[7452];
  assign o[7451] = i[7451];
  assign o[7450] = i[7450];
  assign o[7449] = i[7449];
  assign o[7448] = i[7448];
  assign o[7447] = i[7447];
  assign o[7446] = i[7446];
  assign o[7445] = i[7445];
  assign o[7444] = i[7444];
  assign o[7443] = i[7443];
  assign o[7442] = i[7442];
  assign o[7441] = i[7441];
  assign o[7440] = i[7440];
  assign o[7439] = i[7439];
  assign o[7438] = i[7438];
  assign o[7437] = i[7437];
  assign o[7436] = i[7436];
  assign o[7435] = i[7435];
  assign o[7434] = i[7434];
  assign o[7433] = i[7433];
  assign o[7432] = i[7432];
  assign o[7431] = i[7431];
  assign o[7430] = i[7430];
  assign o[7429] = i[7429];
  assign o[7428] = i[7428];
  assign o[7427] = i[7427];
  assign o[7426] = i[7426];
  assign o[7425] = i[7425];
  assign o[7424] = i[7424];
  assign o[7423] = i[7423];
  assign o[7422] = i[7422];
  assign o[7421] = i[7421];
  assign o[7420] = i[7420];
  assign o[7419] = i[7419];
  assign o[7418] = i[7418];
  assign o[7417] = i[7417];
  assign o[7416] = i[7416];
  assign o[7415] = i[7415];
  assign o[7414] = i[7414];
  assign o[7413] = i[7413];
  assign o[7412] = i[7412];
  assign o[7411] = i[7411];
  assign o[7410] = i[7410];
  assign o[7409] = i[7409];
  assign o[7408] = i[7408];
  assign o[7407] = i[7407];
  assign o[7406] = i[7406];
  assign o[7405] = i[7405];
  assign o[7404] = i[7404];
  assign o[7403] = i[7403];
  assign o[7402] = i[7402];
  assign o[7401] = i[7401];
  assign o[7400] = i[7400];
  assign o[7399] = i[7399];
  assign o[7398] = i[7398];
  assign o[7397] = i[7397];
  assign o[7396] = i[7396];
  assign o[7395] = i[7395];
  assign o[7394] = i[7394];
  assign o[7393] = i[7393];
  assign o[7392] = i[7392];
  assign o[7391] = i[7391];
  assign o[7390] = i[7390];
  assign o[7389] = i[7389];
  assign o[7388] = i[7388];
  assign o[7387] = i[7387];
  assign o[7386] = i[7386];
  assign o[7385] = i[7385];
  assign o[7384] = i[7384];
  assign o[7383] = i[7383];
  assign o[7382] = i[7382];
  assign o[7381] = i[7381];
  assign o[7380] = i[7380];
  assign o[7379] = i[7379];
  assign o[7378] = i[7378];
  assign o[7377] = i[7377];
  assign o[7376] = i[7376];
  assign o[7375] = i[7375];
  assign o[7374] = i[7374];
  assign o[7373] = i[7373];
  assign o[7372] = i[7372];
  assign o[7371] = i[7371];
  assign o[7370] = i[7370];
  assign o[7369] = i[7369];
  assign o[7368] = i[7368];
  assign o[7367] = i[7367];
  assign o[7366] = i[7366];
  assign o[7365] = i[7365];
  assign o[7364] = i[7364];
  assign o[7363] = i[7363];
  assign o[7362] = i[7362];
  assign o[7361] = i[7361];
  assign o[7360] = i[7360];
  assign o[7359] = i[7359];
  assign o[7358] = i[7358];
  assign o[7357] = i[7357];
  assign o[7356] = i[7356];
  assign o[7355] = i[7355];
  assign o[7354] = i[7354];
  assign o[7353] = i[7353];
  assign o[7352] = i[7352];
  assign o[7351] = i[7351];
  assign o[7350] = i[7350];
  assign o[7349] = i[7349];
  assign o[7348] = i[7348];
  assign o[7347] = i[7347];
  assign o[7346] = i[7346];
  assign o[7345] = i[7345];
  assign o[7344] = i[7344];
  assign o[7343] = i[7343];
  assign o[7342] = i[7342];
  assign o[7341] = i[7341];
  assign o[7340] = i[7340];
  assign o[7339] = i[7339];
  assign o[7338] = i[7338];
  assign o[7337] = i[7337];
  assign o[7336] = i[7336];
  assign o[7335] = i[7335];
  assign o[7334] = i[7334];
  assign o[7333] = i[7333];
  assign o[7332] = i[7332];
  assign o[7331] = i[7331];
  assign o[7330] = i[7330];
  assign o[7329] = i[7329];
  assign o[7328] = i[7328];
  assign o[7327] = i[7327];
  assign o[7326] = i[7326];
  assign o[7325] = i[7325];
  assign o[7324] = i[7324];
  assign o[7323] = i[7323];
  assign o[7322] = i[7322];
  assign o[7321] = i[7321];
  assign o[7320] = i[7320];
  assign o[7319] = i[7319];
  assign o[7318] = i[7318];
  assign o[7317] = i[7317];
  assign o[7316] = i[7316];
  assign o[7315] = i[7315];
  assign o[7314] = i[7314];
  assign o[7313] = i[7313];
  assign o[7312] = i[7312];
  assign o[7311] = i[7311];
  assign o[7310] = i[7310];
  assign o[7309] = i[7309];
  assign o[7308] = i[7308];
  assign o[7307] = i[7307];
  assign o[7306] = i[7306];
  assign o[7305] = i[7305];
  assign o[7304] = i[7304];
  assign o[7303] = i[7303];
  assign o[7302] = i[7302];
  assign o[7301] = i[7301];
  assign o[7300] = i[7300];
  assign o[7299] = i[7299];
  assign o[7298] = i[7298];
  assign o[7297] = i[7297];
  assign o[7296] = i[7296];
  assign o[7295] = i[7295];
  assign o[7294] = i[7294];
  assign o[7293] = i[7293];
  assign o[7292] = i[7292];
  assign o[7291] = i[7291];
  assign o[7290] = i[7290];
  assign o[7289] = i[7289];
  assign o[7288] = i[7288];
  assign o[7287] = i[7287];
  assign o[7286] = i[7286];
  assign o[7285] = i[7285];
  assign o[7284] = i[7284];
  assign o[7283] = i[7283];
  assign o[7282] = i[7282];
  assign o[7281] = i[7281];
  assign o[7280] = i[7280];
  assign o[7279] = i[7279];
  assign o[7278] = i[7278];
  assign o[7277] = i[7277];
  assign o[7276] = i[7276];
  assign o[7275] = i[7275];
  assign o[7274] = i[7274];
  assign o[7273] = i[7273];
  assign o[7272] = i[7272];
  assign o[7271] = i[7271];
  assign o[7270] = i[7270];
  assign o[7269] = i[7269];
  assign o[7268] = i[7268];
  assign o[7267] = i[7267];
  assign o[7266] = i[7266];
  assign o[7265] = i[7265];
  assign o[7264] = i[7264];
  assign o[7263] = i[7263];
  assign o[7262] = i[7262];
  assign o[7261] = i[7261];
  assign o[7260] = i[7260];
  assign o[7259] = i[7259];
  assign o[7258] = i[7258];
  assign o[7257] = i[7257];
  assign o[7256] = i[7256];
  assign o[7255] = i[7255];
  assign o[7254] = i[7254];
  assign o[7253] = i[7253];
  assign o[7252] = i[7252];
  assign o[7251] = i[7251];
  assign o[7250] = i[7250];
  assign o[7249] = i[7249];
  assign o[7248] = i[7248];
  assign o[7247] = i[7247];
  assign o[7246] = i[7246];
  assign o[7245] = i[7245];
  assign o[7244] = i[7244];
  assign o[7243] = i[7243];
  assign o[7242] = i[7242];
  assign o[7241] = i[7241];
  assign o[7240] = i[7240];
  assign o[7239] = i[7239];
  assign o[7238] = i[7238];
  assign o[7237] = i[7237];
  assign o[7236] = i[7236];
  assign o[7235] = i[7235];
  assign o[7234] = i[7234];
  assign o[7233] = i[7233];
  assign o[7232] = i[7232];
  assign o[7231] = i[7231];
  assign o[7230] = i[7230];
  assign o[7229] = i[7229];
  assign o[7228] = i[7228];
  assign o[7227] = i[7227];
  assign o[7226] = i[7226];
  assign o[7225] = i[7225];
  assign o[7224] = i[7224];
  assign o[7223] = i[7223];
  assign o[7222] = i[7222];
  assign o[7221] = i[7221];
  assign o[7220] = i[7220];
  assign o[7219] = i[7219];
  assign o[7218] = i[7218];
  assign o[7217] = i[7217];
  assign o[7216] = i[7216];
  assign o[7215] = i[7215];
  assign o[7214] = i[7214];
  assign o[7213] = i[7213];
  assign o[7212] = i[7212];
  assign o[7211] = i[7211];
  assign o[7210] = i[7210];
  assign o[7209] = i[7209];
  assign o[7208] = i[7208];
  assign o[7207] = i[7207];
  assign o[7206] = i[7206];
  assign o[7205] = i[7205];
  assign o[7204] = i[7204];
  assign o[7203] = i[7203];
  assign o[7202] = i[7202];
  assign o[7201] = i[7201];
  assign o[7200] = i[7200];
  assign o[7199] = i[7199];
  assign o[7198] = i[7198];
  assign o[7197] = i[7197];
  assign o[7196] = i[7196];
  assign o[7195] = i[7195];
  assign o[7194] = i[7194];
  assign o[7193] = i[7193];
  assign o[7192] = i[7192];
  assign o[7191] = i[7191];
  assign o[7190] = i[7190];
  assign o[7189] = i[7189];
  assign o[7188] = i[7188];
  assign o[7187] = i[7187];
  assign o[7186] = i[7186];
  assign o[7185] = i[7185];
  assign o[7184] = i[7184];
  assign o[7183] = i[7183];
  assign o[7182] = i[7182];
  assign o[7181] = i[7181];
  assign o[7180] = i[7180];
  assign o[7179] = i[7179];
  assign o[7178] = i[7178];
  assign o[7177] = i[7177];
  assign o[7176] = i[7176];
  assign o[7175] = i[7175];
  assign o[7174] = i[7174];
  assign o[7173] = i[7173];
  assign o[7172] = i[7172];
  assign o[7171] = i[7171];
  assign o[7170] = i[7170];
  assign o[7169] = i[7169];
  assign o[7168] = i[7168];
  assign o[7167] = i[7167];
  assign o[7166] = i[7166];
  assign o[7165] = i[7165];
  assign o[7164] = i[7164];
  assign o[7163] = i[7163];
  assign o[7162] = i[7162];
  assign o[7161] = i[7161];
  assign o[7160] = i[7160];
  assign o[7159] = i[7159];
  assign o[7158] = i[7158];
  assign o[7157] = i[7157];
  assign o[7156] = i[7156];
  assign o[7155] = i[7155];
  assign o[7154] = i[7154];
  assign o[7153] = i[7153];
  assign o[7152] = i[7152];
  assign o[7151] = i[7151];
  assign o[7150] = i[7150];
  assign o[7149] = i[7149];
  assign o[7148] = i[7148];
  assign o[7147] = i[7147];
  assign o[7146] = i[7146];
  assign o[7145] = i[7145];
  assign o[7144] = i[7144];
  assign o[7143] = i[7143];
  assign o[7142] = i[7142];
  assign o[7141] = i[7141];
  assign o[7140] = i[7140];
  assign o[7139] = i[7139];
  assign o[7138] = i[7138];
  assign o[7137] = i[7137];
  assign o[7136] = i[7136];
  assign o[7135] = i[7135];
  assign o[7134] = i[7134];
  assign o[7133] = i[7133];
  assign o[7132] = i[7132];
  assign o[7131] = i[7131];
  assign o[7130] = i[7130];
  assign o[7129] = i[7129];
  assign o[7128] = i[7128];
  assign o[7127] = i[7127];
  assign o[7126] = i[7126];
  assign o[7125] = i[7125];
  assign o[7124] = i[7124];
  assign o[7123] = i[7123];
  assign o[7122] = i[7122];
  assign o[7121] = i[7121];
  assign o[7120] = i[7120];
  assign o[7119] = i[7119];
  assign o[7118] = i[7118];
  assign o[7117] = i[7117];
  assign o[7116] = i[7116];
  assign o[7115] = i[7115];
  assign o[7114] = i[7114];
  assign o[7113] = i[7113];
  assign o[7112] = i[7112];
  assign o[7111] = i[7111];
  assign o[7110] = i[7110];
  assign o[7109] = i[7109];
  assign o[7108] = i[7108];
  assign o[7107] = i[7107];
  assign o[7106] = i[7106];
  assign o[7105] = i[7105];
  assign o[7104] = i[7104];
  assign o[7103] = i[7103];
  assign o[7102] = i[7102];
  assign o[7101] = i[7101];
  assign o[7100] = i[7100];
  assign o[7099] = i[7099];
  assign o[7098] = i[7098];
  assign o[7097] = i[7097];
  assign o[7096] = i[7096];
  assign o[7095] = i[7095];
  assign o[7094] = i[7094];
  assign o[7093] = i[7093];
  assign o[7092] = i[7092];
  assign o[7091] = i[7091];
  assign o[7090] = i[7090];
  assign o[7089] = i[7089];
  assign o[7088] = i[7088];
  assign o[7087] = i[7087];
  assign o[7086] = i[7086];
  assign o[7085] = i[7085];
  assign o[7084] = i[7084];
  assign o[7083] = i[7083];
  assign o[7082] = i[7082];
  assign o[7081] = i[7081];
  assign o[7080] = i[7080];
  assign o[7079] = i[7079];
  assign o[7078] = i[7078];
  assign o[7077] = i[7077];
  assign o[7076] = i[7076];
  assign o[7075] = i[7075];
  assign o[7074] = i[7074];
  assign o[7073] = i[7073];
  assign o[7072] = i[7072];
  assign o[7071] = i[7071];
  assign o[7070] = i[7070];
  assign o[7069] = i[7069];
  assign o[7068] = i[7068];
  assign o[7067] = i[7067];
  assign o[7066] = i[7066];
  assign o[7065] = i[7065];
  assign o[7064] = i[7064];
  assign o[7063] = i[7063];
  assign o[7062] = i[7062];
  assign o[7061] = i[7061];
  assign o[7060] = i[7060];
  assign o[7059] = i[7059];
  assign o[7058] = i[7058];
  assign o[7057] = i[7057];
  assign o[7056] = i[7056];
  assign o[7055] = i[7055];
  assign o[7054] = i[7054];
  assign o[7053] = i[7053];
  assign o[7052] = i[7052];
  assign o[7051] = i[7051];
  assign o[7050] = i[7050];
  assign o[7049] = i[7049];
  assign o[7048] = i[7048];
  assign o[7047] = i[7047];
  assign o[7046] = i[7046];
  assign o[7045] = i[7045];
  assign o[7044] = i[7044];
  assign o[7043] = i[7043];
  assign o[7042] = i[7042];
  assign o[7041] = i[7041];
  assign o[7040] = i[7040];
  assign o[7039] = i[7039];
  assign o[7038] = i[7038];
  assign o[7037] = i[7037];
  assign o[7036] = i[7036];
  assign o[7035] = i[7035];
  assign o[7034] = i[7034];
  assign o[7033] = i[7033];
  assign o[7032] = i[7032];
  assign o[7031] = i[7031];
  assign o[7030] = i[7030];
  assign o[7029] = i[7029];
  assign o[7028] = i[7028];
  assign o[7027] = i[7027];
  assign o[7026] = i[7026];
  assign o[7025] = i[7025];
  assign o[7024] = i[7024];
  assign o[7023] = i[7023];
  assign o[7022] = i[7022];
  assign o[7021] = i[7021];
  assign o[7020] = i[7020];
  assign o[7019] = i[7019];
  assign o[7018] = i[7018];
  assign o[7017] = i[7017];
  assign o[7016] = i[7016];
  assign o[7015] = i[7015];
  assign o[7014] = i[7014];
  assign o[7013] = i[7013];
  assign o[7012] = i[7012];
  assign o[7011] = i[7011];
  assign o[7010] = i[7010];
  assign o[7009] = i[7009];
  assign o[7008] = i[7008];
  assign o[7007] = i[7007];
  assign o[7006] = i[7006];
  assign o[7005] = i[7005];
  assign o[7004] = i[7004];
  assign o[7003] = i[7003];
  assign o[7002] = i[7002];
  assign o[7001] = i[7001];
  assign o[7000] = i[7000];
  assign o[6999] = i[6999];
  assign o[6998] = i[6998];
  assign o[6997] = i[6997];
  assign o[6996] = i[6996];
  assign o[6995] = i[6995];
  assign o[6994] = i[6994];
  assign o[6993] = i[6993];
  assign o[6992] = i[6992];
  assign o[6991] = i[6991];
  assign o[6990] = i[6990];
  assign o[6989] = i[6989];
  assign o[6988] = i[6988];
  assign o[6987] = i[6987];
  assign o[6986] = i[6986];
  assign o[6985] = i[6985];
  assign o[6984] = i[6984];
  assign o[6983] = i[6983];
  assign o[6982] = i[6982];
  assign o[6981] = i[6981];
  assign o[6980] = i[6980];
  assign o[6979] = i[6979];
  assign o[6978] = i[6978];
  assign o[6977] = i[6977];
  assign o[6976] = i[6976];
  assign o[6975] = i[6975];
  assign o[6974] = i[6974];
  assign o[6973] = i[6973];
  assign o[6972] = i[6972];
  assign o[6971] = i[6971];
  assign o[6970] = i[6970];
  assign o[6969] = i[6969];
  assign o[6968] = i[6968];
  assign o[6967] = i[6967];
  assign o[6966] = i[6966];
  assign o[6965] = i[6965];
  assign o[6964] = i[6964];
  assign o[6963] = i[6963];
  assign o[6962] = i[6962];
  assign o[6961] = i[6961];
  assign o[6960] = i[6960];
  assign o[6959] = i[6959];
  assign o[6958] = i[6958];
  assign o[6957] = i[6957];
  assign o[6956] = i[6956];
  assign o[6955] = i[6955];
  assign o[6954] = i[6954];
  assign o[6953] = i[6953];
  assign o[6952] = i[6952];
  assign o[6951] = i[6951];
  assign o[6950] = i[6950];
  assign o[6949] = i[6949];
  assign o[6948] = i[6948];
  assign o[6947] = i[6947];
  assign o[6946] = i[6946];
  assign o[6945] = i[6945];
  assign o[6944] = i[6944];
  assign o[6943] = i[6943];
  assign o[6942] = i[6942];
  assign o[6941] = i[6941];
  assign o[6940] = i[6940];
  assign o[6939] = i[6939];
  assign o[6938] = i[6938];
  assign o[6937] = i[6937];
  assign o[6936] = i[6936];
  assign o[6935] = i[6935];
  assign o[6934] = i[6934];
  assign o[6933] = i[6933];
  assign o[6932] = i[6932];
  assign o[6931] = i[6931];
  assign o[6930] = i[6930];
  assign o[6929] = i[6929];
  assign o[6928] = i[6928];
  assign o[6927] = i[6927];
  assign o[6926] = i[6926];
  assign o[6925] = i[6925];
  assign o[6924] = i[6924];
  assign o[6923] = i[6923];
  assign o[6922] = i[6922];
  assign o[6921] = i[6921];
  assign o[6920] = i[6920];
  assign o[6919] = i[6919];
  assign o[6918] = i[6918];
  assign o[6917] = i[6917];
  assign o[6916] = i[6916];
  assign o[6915] = i[6915];
  assign o[6914] = i[6914];
  assign o[6913] = i[6913];
  assign o[6912] = i[6912];
  assign o[6911] = i[6911];
  assign o[6910] = i[6910];
  assign o[6909] = i[6909];
  assign o[6908] = i[6908];
  assign o[6907] = i[6907];
  assign o[6906] = i[6906];
  assign o[6905] = i[6905];
  assign o[6904] = i[6904];
  assign o[6903] = i[6903];
  assign o[6902] = i[6902];
  assign o[6901] = i[6901];
  assign o[6900] = i[6900];
  assign o[6899] = i[6899];
  assign o[6898] = i[6898];
  assign o[6897] = i[6897];
  assign o[6896] = i[6896];
  assign o[6895] = i[6895];
  assign o[6894] = i[6894];
  assign o[6893] = i[6893];
  assign o[6892] = i[6892];
  assign o[6891] = i[6891];
  assign o[6890] = i[6890];
  assign o[6889] = i[6889];
  assign o[6888] = i[6888];
  assign o[6887] = i[6887];
  assign o[6886] = i[6886];
  assign o[6885] = i[6885];
  assign o[6884] = i[6884];
  assign o[6883] = i[6883];
  assign o[6882] = i[6882];
  assign o[6881] = i[6881];
  assign o[6880] = i[6880];
  assign o[6879] = i[6879];
  assign o[6878] = i[6878];
  assign o[6877] = i[6877];
  assign o[6876] = i[6876];
  assign o[6875] = i[6875];
  assign o[6874] = i[6874];
  assign o[6873] = i[6873];
  assign o[6872] = i[6872];
  assign o[6871] = i[6871];
  assign o[6870] = i[6870];
  assign o[6869] = i[6869];
  assign o[6868] = i[6868];
  assign o[6867] = i[6867];
  assign o[6866] = i[6866];
  assign o[6865] = i[6865];
  assign o[6864] = i[6864];
  assign o[6863] = i[6863];
  assign o[6862] = i[6862];
  assign o[6861] = i[6861];
  assign o[6860] = i[6860];
  assign o[6859] = i[6859];
  assign o[6858] = i[6858];
  assign o[6857] = i[6857];
  assign o[6856] = i[6856];
  assign o[6855] = i[6855];
  assign o[6854] = i[6854];
  assign o[6853] = i[6853];
  assign o[6852] = i[6852];
  assign o[6851] = i[6851];
  assign o[6850] = i[6850];
  assign o[6849] = i[6849];
  assign o[6848] = i[6848];
  assign o[6847] = i[6847];
  assign o[6846] = i[6846];
  assign o[6845] = i[6845];
  assign o[6844] = i[6844];
  assign o[6843] = i[6843];
  assign o[6842] = i[6842];
  assign o[6841] = i[6841];
  assign o[6840] = i[6840];
  assign o[6839] = i[6839];
  assign o[6838] = i[6838];
  assign o[6837] = i[6837];
  assign o[6836] = i[6836];
  assign o[6835] = i[6835];
  assign o[6834] = i[6834];
  assign o[6833] = i[6833];
  assign o[6832] = i[6832];
  assign o[6831] = i[6831];
  assign o[6830] = i[6830];
  assign o[6829] = i[6829];
  assign o[6828] = i[6828];
  assign o[6827] = i[6827];
  assign o[6826] = i[6826];
  assign o[6825] = i[6825];
  assign o[6824] = i[6824];
  assign o[6823] = i[6823];
  assign o[6822] = i[6822];
  assign o[6821] = i[6821];
  assign o[6820] = i[6820];
  assign o[6819] = i[6819];
  assign o[6818] = i[6818];
  assign o[6817] = i[6817];
  assign o[6816] = i[6816];
  assign o[6815] = i[6815];
  assign o[6814] = i[6814];
  assign o[6813] = i[6813];
  assign o[6812] = i[6812];
  assign o[6811] = i[6811];
  assign o[6810] = i[6810];
  assign o[6809] = i[6809];
  assign o[6808] = i[6808];
  assign o[6807] = i[6807];
  assign o[6806] = i[6806];
  assign o[6805] = i[6805];
  assign o[6804] = i[6804];
  assign o[6803] = i[6803];
  assign o[6802] = i[6802];
  assign o[6801] = i[6801];
  assign o[6800] = i[6800];
  assign o[6799] = i[6799];
  assign o[6798] = i[6798];
  assign o[6797] = i[6797];
  assign o[6796] = i[6796];
  assign o[6795] = i[6795];
  assign o[6794] = i[6794];
  assign o[6793] = i[6793];
  assign o[6792] = i[6792];
  assign o[6791] = i[6791];
  assign o[6790] = i[6790];
  assign o[6789] = i[6789];
  assign o[6788] = i[6788];
  assign o[6787] = i[6787];
  assign o[6786] = i[6786];
  assign o[6785] = i[6785];
  assign o[6784] = i[6784];
  assign o[6783] = i[6783];
  assign o[6782] = i[6782];
  assign o[6781] = i[6781];
  assign o[6780] = i[6780];
  assign o[6779] = i[6779];
  assign o[6778] = i[6778];
  assign o[6777] = i[6777];
  assign o[6776] = i[6776];
  assign o[6775] = i[6775];
  assign o[6774] = i[6774];
  assign o[6773] = i[6773];
  assign o[6772] = i[6772];
  assign o[6771] = i[6771];
  assign o[6770] = i[6770];
  assign o[6769] = i[6769];
  assign o[6768] = i[6768];
  assign o[6767] = i[6767];
  assign o[6766] = i[6766];
  assign o[6765] = i[6765];
  assign o[6764] = i[6764];
  assign o[6763] = i[6763];
  assign o[6762] = i[6762];
  assign o[6761] = i[6761];
  assign o[6760] = i[6760];
  assign o[6759] = i[6759];
  assign o[6758] = i[6758];
  assign o[6757] = i[6757];
  assign o[6756] = i[6756];
  assign o[6755] = i[6755];
  assign o[6754] = i[6754];
  assign o[6753] = i[6753];
  assign o[6752] = i[6752];
  assign o[6751] = i[6751];
  assign o[6750] = i[6750];
  assign o[6749] = i[6749];
  assign o[6748] = i[6748];
  assign o[6747] = i[6747];
  assign o[6746] = i[6746];
  assign o[6745] = i[6745];
  assign o[6744] = i[6744];
  assign o[6743] = i[6743];
  assign o[6742] = i[6742];
  assign o[6741] = i[6741];
  assign o[6740] = i[6740];
  assign o[6739] = i[6739];
  assign o[6738] = i[6738];
  assign o[6737] = i[6737];
  assign o[6736] = i[6736];
  assign o[6735] = i[6735];
  assign o[6734] = i[6734];
  assign o[6733] = i[6733];
  assign o[6732] = i[6732];
  assign o[6731] = i[6731];
  assign o[6730] = i[6730];
  assign o[6729] = i[6729];
  assign o[6728] = i[6728];
  assign o[6727] = i[6727];
  assign o[6726] = i[6726];
  assign o[6725] = i[6725];
  assign o[6724] = i[6724];
  assign o[6723] = i[6723];
  assign o[6722] = i[6722];
  assign o[6721] = i[6721];
  assign o[6720] = i[6720];
  assign o[6719] = i[6719];
  assign o[6718] = i[6718];
  assign o[6717] = i[6717];
  assign o[6716] = i[6716];
  assign o[6715] = i[6715];
  assign o[6714] = i[6714];
  assign o[6713] = i[6713];
  assign o[6712] = i[6712];
  assign o[6711] = i[6711];
  assign o[6710] = i[6710];
  assign o[6709] = i[6709];
  assign o[6708] = i[6708];
  assign o[6707] = i[6707];
  assign o[6706] = i[6706];
  assign o[6705] = i[6705];
  assign o[6704] = i[6704];
  assign o[6703] = i[6703];
  assign o[6702] = i[6702];
  assign o[6701] = i[6701];
  assign o[6700] = i[6700];
  assign o[6699] = i[6699];
  assign o[6698] = i[6698];
  assign o[6697] = i[6697];
  assign o[6696] = i[6696];
  assign o[6695] = i[6695];
  assign o[6694] = i[6694];
  assign o[6693] = i[6693];
  assign o[6692] = i[6692];
  assign o[6691] = i[6691];
  assign o[6690] = i[6690];
  assign o[6689] = i[6689];
  assign o[6688] = i[6688];
  assign o[6687] = i[6687];
  assign o[6686] = i[6686];
  assign o[6685] = i[6685];
  assign o[6684] = i[6684];
  assign o[6683] = i[6683];
  assign o[6682] = i[6682];
  assign o[6681] = i[6681];
  assign o[6680] = i[6680];
  assign o[6679] = i[6679];
  assign o[6678] = i[6678];
  assign o[6677] = i[6677];
  assign o[6676] = i[6676];
  assign o[6675] = i[6675];
  assign o[6674] = i[6674];
  assign o[6673] = i[6673];
  assign o[6672] = i[6672];
  assign o[6671] = i[6671];
  assign o[6670] = i[6670];
  assign o[6669] = i[6669];
  assign o[6668] = i[6668];
  assign o[6667] = i[6667];
  assign o[6666] = i[6666];
  assign o[6665] = i[6665];
  assign o[6664] = i[6664];
  assign o[6663] = i[6663];
  assign o[6662] = i[6662];
  assign o[6661] = i[6661];
  assign o[6660] = i[6660];
  assign o[6659] = i[6659];
  assign o[6658] = i[6658];
  assign o[6657] = i[6657];
  assign o[6656] = i[6656];
  assign o[6655] = i[6655];
  assign o[6654] = i[6654];
  assign o[6653] = i[6653];
  assign o[6652] = i[6652];
  assign o[6651] = i[6651];
  assign o[6650] = i[6650];
  assign o[6649] = i[6649];
  assign o[6648] = i[6648];
  assign o[6647] = i[6647];
  assign o[6646] = i[6646];
  assign o[6645] = i[6645];
  assign o[6644] = i[6644];
  assign o[6643] = i[6643];
  assign o[6642] = i[6642];
  assign o[6641] = i[6641];
  assign o[6640] = i[6640];
  assign o[6639] = i[6639];
  assign o[6638] = i[6638];
  assign o[6637] = i[6637];
  assign o[6636] = i[6636];
  assign o[6635] = i[6635];
  assign o[6634] = i[6634];
  assign o[6633] = i[6633];
  assign o[6632] = i[6632];
  assign o[6631] = i[6631];
  assign o[6630] = i[6630];
  assign o[6629] = i[6629];
  assign o[6628] = i[6628];
  assign o[6627] = i[6627];
  assign o[6626] = i[6626];
  assign o[6625] = i[6625];
  assign o[6624] = i[6624];
  assign o[6623] = i[6623];
  assign o[6622] = i[6622];
  assign o[6621] = i[6621];
  assign o[6620] = i[6620];
  assign o[6619] = i[6619];
  assign o[6618] = i[6618];
  assign o[6617] = i[6617];
  assign o[6616] = i[6616];
  assign o[6615] = i[6615];
  assign o[6614] = i[6614];
  assign o[6613] = i[6613];
  assign o[6612] = i[6612];
  assign o[6611] = i[6611];
  assign o[6610] = i[6610];
  assign o[6609] = i[6609];
  assign o[6608] = i[6608];
  assign o[6607] = i[6607];
  assign o[6606] = i[6606];
  assign o[6605] = i[6605];
  assign o[6604] = i[6604];
  assign o[6603] = i[6603];
  assign o[6602] = i[6602];
  assign o[6601] = i[6601];
  assign o[6600] = i[6600];
  assign o[6599] = i[6599];
  assign o[6598] = i[6598];
  assign o[6597] = i[6597];
  assign o[6596] = i[6596];
  assign o[6595] = i[6595];
  assign o[6594] = i[6594];
  assign o[6593] = i[6593];
  assign o[6592] = i[6592];
  assign o[6591] = i[6591];
  assign o[6590] = i[6590];
  assign o[6589] = i[6589];
  assign o[6588] = i[6588];
  assign o[6587] = i[6587];
  assign o[6586] = i[6586];
  assign o[6585] = i[6585];
  assign o[6584] = i[6584];
  assign o[6583] = i[6583];
  assign o[6582] = i[6582];
  assign o[6581] = i[6581];
  assign o[6580] = i[6580];
  assign o[6579] = i[6579];
  assign o[6578] = i[6578];
  assign o[6577] = i[6577];
  assign o[6576] = i[6576];
  assign o[6575] = i[6575];
  assign o[6574] = i[6574];
  assign o[6573] = i[6573];
  assign o[6572] = i[6572];
  assign o[6571] = i[6571];
  assign o[6570] = i[6570];
  assign o[6569] = i[6569];
  assign o[6568] = i[6568];
  assign o[6567] = i[6567];
  assign o[6566] = i[6566];
  assign o[6565] = i[6565];
  assign o[6564] = i[6564];
  assign o[6563] = i[6563];
  assign o[6562] = i[6562];
  assign o[6561] = i[6561];
  assign o[6560] = i[6560];
  assign o[6559] = i[6559];
  assign o[6558] = i[6558];
  assign o[6557] = i[6557];
  assign o[6556] = i[6556];
  assign o[6555] = i[6555];
  assign o[6554] = i[6554];
  assign o[6553] = i[6553];
  assign o[6552] = i[6552];
  assign o[6551] = i[6551];
  assign o[6550] = i[6550];
  assign o[6549] = i[6549];
  assign o[6548] = i[6548];
  assign o[6547] = i[6547];
  assign o[6546] = i[6546];
  assign o[6545] = i[6545];
  assign o[6544] = i[6544];
  assign o[6543] = i[6543];
  assign o[6542] = i[6542];
  assign o[6541] = i[6541];
  assign o[6540] = i[6540];
  assign o[6539] = i[6539];
  assign o[6538] = i[6538];
  assign o[6537] = i[6537];
  assign o[6536] = i[6536];
  assign o[6535] = i[6535];
  assign o[6534] = i[6534];
  assign o[6533] = i[6533];
  assign o[6532] = i[6532];
  assign o[6531] = i[6531];
  assign o[6530] = i[6530];
  assign o[6529] = i[6529];
  assign o[6528] = i[6528];
  assign o[6527] = i[6527];
  assign o[6526] = i[6526];
  assign o[6525] = i[6525];
  assign o[6524] = i[6524];
  assign o[6523] = i[6523];
  assign o[6522] = i[6522];
  assign o[6521] = i[6521];
  assign o[6520] = i[6520];
  assign o[6519] = i[6519];
  assign o[6518] = i[6518];
  assign o[6517] = i[6517];
  assign o[6516] = i[6516];
  assign o[6515] = i[6515];
  assign o[6514] = i[6514];
  assign o[6513] = i[6513];
  assign o[6512] = i[6512];
  assign o[6511] = i[6511];
  assign o[6510] = i[6510];
  assign o[6509] = i[6509];
  assign o[6508] = i[6508];
  assign o[6507] = i[6507];
  assign o[6506] = i[6506];
  assign o[6505] = i[6505];
  assign o[6504] = i[6504];
  assign o[6503] = i[6503];
  assign o[6502] = i[6502];
  assign o[6501] = i[6501];
  assign o[6500] = i[6500];
  assign o[6499] = i[6499];
  assign o[6498] = i[6498];
  assign o[6497] = i[6497];
  assign o[6496] = i[6496];
  assign o[6495] = i[6495];
  assign o[6494] = i[6494];
  assign o[6493] = i[6493];
  assign o[6492] = i[6492];
  assign o[6491] = i[6491];
  assign o[6490] = i[6490];
  assign o[6489] = i[6489];
  assign o[6488] = i[6488];
  assign o[6487] = i[6487];
  assign o[6486] = i[6486];
  assign o[6485] = i[6485];
  assign o[6484] = i[6484];
  assign o[6483] = i[6483];
  assign o[6482] = i[6482];
  assign o[6481] = i[6481];
  assign o[6480] = i[6480];
  assign o[6479] = i[6479];
  assign o[6478] = i[6478];
  assign o[6477] = i[6477];
  assign o[6476] = i[6476];
  assign o[6475] = i[6475];
  assign o[6474] = i[6474];
  assign o[6473] = i[6473];
  assign o[6472] = i[6472];
  assign o[6471] = i[6471];
  assign o[6470] = i[6470];
  assign o[6469] = i[6469];
  assign o[6468] = i[6468];
  assign o[6467] = i[6467];
  assign o[6466] = i[6466];
  assign o[6465] = i[6465];
  assign o[6464] = i[6464];
  assign o[6463] = i[6463];
  assign o[6462] = i[6462];
  assign o[6461] = i[6461];
  assign o[6460] = i[6460];
  assign o[6459] = i[6459];
  assign o[6458] = i[6458];
  assign o[6457] = i[6457];
  assign o[6456] = i[6456];
  assign o[6455] = i[6455];
  assign o[6454] = i[6454];
  assign o[6453] = i[6453];
  assign o[6452] = i[6452];
  assign o[6451] = i[6451];
  assign o[6450] = i[6450];
  assign o[6449] = i[6449];
  assign o[6448] = i[6448];
  assign o[6447] = i[6447];
  assign o[6446] = i[6446];
  assign o[6445] = i[6445];
  assign o[6444] = i[6444];
  assign o[6443] = i[6443];
  assign o[6442] = i[6442];
  assign o[6441] = i[6441];
  assign o[6440] = i[6440];
  assign o[6439] = i[6439];
  assign o[6438] = i[6438];
  assign o[6437] = i[6437];
  assign o[6436] = i[6436];
  assign o[6435] = i[6435];
  assign o[6434] = i[6434];
  assign o[6433] = i[6433];
  assign o[6432] = i[6432];
  assign o[6431] = i[6431];
  assign o[6430] = i[6430];
  assign o[6429] = i[6429];
  assign o[6428] = i[6428];
  assign o[6427] = i[6427];
  assign o[6426] = i[6426];
  assign o[6425] = i[6425];
  assign o[6424] = i[6424];
  assign o[6423] = i[6423];
  assign o[6422] = i[6422];
  assign o[6421] = i[6421];
  assign o[6420] = i[6420];
  assign o[6419] = i[6419];
  assign o[6418] = i[6418];
  assign o[6417] = i[6417];
  assign o[6416] = i[6416];
  assign o[6415] = i[6415];
  assign o[6414] = i[6414];
  assign o[6413] = i[6413];
  assign o[6412] = i[6412];
  assign o[6411] = i[6411];
  assign o[6410] = i[6410];
  assign o[6409] = i[6409];
  assign o[6408] = i[6408];
  assign o[6407] = i[6407];
  assign o[6406] = i[6406];
  assign o[6405] = i[6405];
  assign o[6404] = i[6404];
  assign o[6403] = i[6403];
  assign o[6402] = i[6402];
  assign o[6401] = i[6401];
  assign o[6400] = i[6400];
  assign o[6399] = i[6399];
  assign o[6398] = i[6398];
  assign o[6397] = i[6397];
  assign o[6396] = i[6396];
  assign o[6395] = i[6395];
  assign o[6394] = i[6394];
  assign o[6393] = i[6393];
  assign o[6392] = i[6392];
  assign o[6391] = i[6391];
  assign o[6390] = i[6390];
  assign o[6389] = i[6389];
  assign o[6388] = i[6388];
  assign o[6387] = i[6387];
  assign o[6386] = i[6386];
  assign o[6385] = i[6385];
  assign o[6384] = i[6384];
  assign o[6383] = i[6383];
  assign o[6382] = i[6382];
  assign o[6381] = i[6381];
  assign o[6380] = i[6380];
  assign o[6379] = i[6379];
  assign o[6378] = i[6378];
  assign o[6377] = i[6377];
  assign o[6376] = i[6376];
  assign o[6375] = i[6375];
  assign o[6374] = i[6374];
  assign o[6373] = i[6373];
  assign o[6372] = i[6372];
  assign o[6371] = i[6371];
  assign o[6370] = i[6370];
  assign o[6369] = i[6369];
  assign o[6368] = i[6368];
  assign o[6367] = i[6367];
  assign o[6366] = i[6366];
  assign o[6365] = i[6365];
  assign o[6364] = i[6364];
  assign o[6363] = i[6363];
  assign o[6362] = i[6362];
  assign o[6361] = i[6361];
  assign o[6360] = i[6360];
  assign o[6359] = i[6359];
  assign o[6358] = i[6358];
  assign o[6357] = i[6357];
  assign o[6356] = i[6356];
  assign o[6355] = i[6355];
  assign o[6354] = i[6354];
  assign o[6353] = i[6353];
  assign o[6352] = i[6352];
  assign o[6351] = i[6351];
  assign o[6350] = i[6350];
  assign o[6349] = i[6349];
  assign o[6348] = i[6348];
  assign o[6347] = i[6347];
  assign o[6346] = i[6346];
  assign o[6345] = i[6345];
  assign o[6344] = i[6344];
  assign o[6343] = i[6343];
  assign o[6342] = i[6342];
  assign o[6341] = i[6341];
  assign o[6340] = i[6340];
  assign o[6339] = i[6339];
  assign o[6338] = i[6338];
  assign o[6337] = i[6337];
  assign o[6336] = i[6336];
  assign o[6335] = i[6335];
  assign o[6334] = i[6334];
  assign o[6333] = i[6333];
  assign o[6332] = i[6332];
  assign o[6331] = i[6331];
  assign o[6330] = i[6330];
  assign o[6329] = i[6329];
  assign o[6328] = i[6328];
  assign o[6327] = i[6327];
  assign o[6326] = i[6326];
  assign o[6325] = i[6325];
  assign o[6324] = i[6324];
  assign o[6323] = i[6323];
  assign o[6322] = i[6322];
  assign o[6321] = i[6321];
  assign o[6320] = i[6320];
  assign o[6319] = i[6319];
  assign o[6318] = i[6318];
  assign o[6317] = i[6317];
  assign o[6316] = i[6316];
  assign o[6315] = i[6315];
  assign o[6314] = i[6314];
  assign o[6313] = i[6313];
  assign o[6312] = i[6312];
  assign o[6311] = i[6311];
  assign o[6310] = i[6310];
  assign o[6309] = i[6309];
  assign o[6308] = i[6308];
  assign o[6307] = i[6307];
  assign o[6306] = i[6306];
  assign o[6305] = i[6305];
  assign o[6304] = i[6304];
  assign o[6303] = i[6303];
  assign o[6302] = i[6302];
  assign o[6301] = i[6301];
  assign o[6300] = i[6300];
  assign o[6299] = i[6299];
  assign o[6298] = i[6298];
  assign o[6297] = i[6297];
  assign o[6296] = i[6296];
  assign o[6295] = i[6295];
  assign o[6294] = i[6294];
  assign o[6293] = i[6293];
  assign o[6292] = i[6292];
  assign o[6291] = i[6291];
  assign o[6290] = i[6290];
  assign o[6289] = i[6289];
  assign o[6288] = i[6288];
  assign o[6287] = i[6287];
  assign o[6286] = i[6286];
  assign o[6285] = i[6285];
  assign o[6284] = i[6284];
  assign o[6283] = i[6283];
  assign o[6282] = i[6282];
  assign o[6281] = i[6281];
  assign o[6280] = i[6280];
  assign o[6279] = i[6279];
  assign o[6278] = i[6278];
  assign o[6277] = i[6277];
  assign o[6276] = i[6276];
  assign o[6275] = i[6275];
  assign o[6274] = i[6274];
  assign o[6273] = i[6273];
  assign o[6272] = i[6272];
  assign o[6271] = i[6271];
  assign o[6270] = i[6270];
  assign o[6269] = i[6269];
  assign o[6268] = i[6268];
  assign o[6267] = i[6267];
  assign o[6266] = i[6266];
  assign o[6265] = i[6265];
  assign o[6264] = i[6264];
  assign o[6263] = i[6263];
  assign o[6262] = i[6262];
  assign o[6261] = i[6261];
  assign o[6260] = i[6260];
  assign o[6259] = i[6259];
  assign o[6258] = i[6258];
  assign o[6257] = i[6257];
  assign o[6256] = i[6256];
  assign o[6255] = i[6255];
  assign o[6254] = i[6254];
  assign o[6253] = i[6253];
  assign o[6252] = i[6252];
  assign o[6251] = i[6251];
  assign o[6250] = i[6250];
  assign o[6249] = i[6249];
  assign o[6248] = i[6248];
  assign o[6247] = i[6247];
  assign o[6246] = i[6246];
  assign o[6245] = i[6245];
  assign o[6244] = i[6244];
  assign o[6243] = i[6243];
  assign o[6242] = i[6242];
  assign o[6241] = i[6241];
  assign o[6240] = i[6240];
  assign o[6239] = i[6239];
  assign o[6238] = i[6238];
  assign o[6237] = i[6237];
  assign o[6236] = i[6236];
  assign o[6235] = i[6235];
  assign o[6234] = i[6234];
  assign o[6233] = i[6233];
  assign o[6232] = i[6232];
  assign o[6231] = i[6231];
  assign o[6230] = i[6230];
  assign o[6229] = i[6229];
  assign o[6228] = i[6228];
  assign o[6227] = i[6227];
  assign o[6226] = i[6226];
  assign o[6225] = i[6225];
  assign o[6224] = i[6224];
  assign o[6223] = i[6223];
  assign o[6222] = i[6222];
  assign o[6221] = i[6221];
  assign o[6220] = i[6220];
  assign o[6219] = i[6219];
  assign o[6218] = i[6218];
  assign o[6217] = i[6217];
  assign o[6216] = i[6216];
  assign o[6215] = i[6215];
  assign o[6214] = i[6214];
  assign o[6213] = i[6213];
  assign o[6212] = i[6212];
  assign o[6211] = i[6211];
  assign o[6210] = i[6210];
  assign o[6209] = i[6209];
  assign o[6208] = i[6208];
  assign o[6207] = i[6207];
  assign o[6206] = i[6206];
  assign o[6205] = i[6205];
  assign o[6204] = i[6204];
  assign o[6203] = i[6203];
  assign o[6202] = i[6202];
  assign o[6201] = i[6201];
  assign o[6200] = i[6200];
  assign o[6199] = i[6199];
  assign o[6198] = i[6198];
  assign o[6197] = i[6197];
  assign o[6196] = i[6196];
  assign o[6195] = i[6195];
  assign o[6194] = i[6194];
  assign o[6193] = i[6193];
  assign o[6192] = i[6192];
  assign o[6191] = i[6191];
  assign o[6190] = i[6190];
  assign o[6189] = i[6189];
  assign o[6188] = i[6188];
  assign o[6187] = i[6187];
  assign o[6186] = i[6186];
  assign o[6185] = i[6185];
  assign o[6184] = i[6184];
  assign o[6183] = i[6183];
  assign o[6182] = i[6182];
  assign o[6181] = i[6181];
  assign o[6180] = i[6180];
  assign o[6179] = i[6179];
  assign o[6178] = i[6178];
  assign o[6177] = i[6177];
  assign o[6176] = i[6176];
  assign o[6175] = i[6175];
  assign o[6174] = i[6174];
  assign o[6173] = i[6173];
  assign o[6172] = i[6172];
  assign o[6171] = i[6171];
  assign o[6170] = i[6170];
  assign o[6169] = i[6169];
  assign o[6168] = i[6168];
  assign o[6167] = i[6167];
  assign o[6166] = i[6166];
  assign o[6165] = i[6165];
  assign o[6164] = i[6164];
  assign o[6163] = i[6163];
  assign o[6162] = i[6162];
  assign o[6161] = i[6161];
  assign o[6160] = i[6160];
  assign o[6159] = i[6159];
  assign o[6158] = i[6158];
  assign o[6157] = i[6157];
  assign o[6156] = i[6156];
  assign o[6155] = i[6155];
  assign o[6154] = i[6154];
  assign o[6153] = i[6153];
  assign o[6152] = i[6152];
  assign o[6151] = i[6151];
  assign o[6150] = i[6150];
  assign o[6149] = i[6149];
  assign o[6148] = i[6148];
  assign o[6147] = i[6147];
  assign o[6146] = i[6146];
  assign o[6145] = i[6145];
  assign o[6144] = i[6144];
  assign o[6143] = i[6143];
  assign o[6142] = i[6142];
  assign o[6141] = i[6141];
  assign o[6140] = i[6140];
  assign o[6139] = i[6139];
  assign o[6138] = i[6138];
  assign o[6137] = i[6137];
  assign o[6136] = i[6136];
  assign o[6135] = i[6135];
  assign o[6134] = i[6134];
  assign o[6133] = i[6133];
  assign o[6132] = i[6132];
  assign o[6131] = i[6131];
  assign o[6130] = i[6130];
  assign o[6129] = i[6129];
  assign o[6128] = i[6128];
  assign o[6127] = i[6127];
  assign o[6126] = i[6126];
  assign o[6125] = i[6125];
  assign o[6124] = i[6124];
  assign o[6123] = i[6123];
  assign o[6122] = i[6122];
  assign o[6121] = i[6121];
  assign o[6120] = i[6120];
  assign o[6119] = i[6119];
  assign o[6118] = i[6118];
  assign o[6117] = i[6117];
  assign o[6116] = i[6116];
  assign o[6115] = i[6115];
  assign o[6114] = i[6114];
  assign o[6113] = i[6113];
  assign o[6112] = i[6112];
  assign o[6111] = i[6111];
  assign o[6110] = i[6110];
  assign o[6109] = i[6109];
  assign o[6108] = i[6108];
  assign o[6107] = i[6107];
  assign o[6106] = i[6106];
  assign o[6105] = i[6105];
  assign o[6104] = i[6104];
  assign o[6103] = i[6103];
  assign o[6102] = i[6102];
  assign o[6101] = i[6101];
  assign o[6100] = i[6100];
  assign o[6099] = i[6099];
  assign o[6098] = i[6098];
  assign o[6097] = i[6097];
  assign o[6096] = i[6096];
  assign o[6095] = i[6095];
  assign o[6094] = i[6094];
  assign o[6093] = i[6093];
  assign o[6092] = i[6092];
  assign o[6091] = i[6091];
  assign o[6090] = i[6090];
  assign o[6089] = i[6089];
  assign o[6088] = i[6088];
  assign o[6087] = i[6087];
  assign o[6086] = i[6086];
  assign o[6085] = i[6085];
  assign o[6084] = i[6084];
  assign o[6083] = i[6083];
  assign o[6082] = i[6082];
  assign o[6081] = i[6081];
  assign o[6080] = i[6080];
  assign o[6079] = i[6079];
  assign o[6078] = i[6078];
  assign o[6077] = i[6077];
  assign o[6076] = i[6076];
  assign o[6075] = i[6075];
  assign o[6074] = i[6074];
  assign o[6073] = i[6073];
  assign o[6072] = i[6072];
  assign o[6071] = i[6071];
  assign o[6070] = i[6070];
  assign o[6069] = i[6069];
  assign o[6068] = i[6068];
  assign o[6067] = i[6067];
  assign o[6066] = i[6066];
  assign o[6065] = i[6065];
  assign o[6064] = i[6064];
  assign o[6063] = i[6063];
  assign o[6062] = i[6062];
  assign o[6061] = i[6061];
  assign o[6060] = i[6060];
  assign o[6059] = i[6059];
  assign o[6058] = i[6058];
  assign o[6057] = i[6057];
  assign o[6056] = i[6056];
  assign o[6055] = i[6055];
  assign o[6054] = i[6054];
  assign o[6053] = i[6053];
  assign o[6052] = i[6052];
  assign o[6051] = i[6051];
  assign o[6050] = i[6050];
  assign o[6049] = i[6049];
  assign o[6048] = i[6048];
  assign o[6047] = i[6047];
  assign o[6046] = i[6046];
  assign o[6045] = i[6045];
  assign o[6044] = i[6044];
  assign o[6043] = i[6043];
  assign o[6042] = i[6042];
  assign o[6041] = i[6041];
  assign o[6040] = i[6040];
  assign o[6039] = i[6039];
  assign o[6038] = i[6038];
  assign o[6037] = i[6037];
  assign o[6036] = i[6036];
  assign o[6035] = i[6035];
  assign o[6034] = i[6034];
  assign o[6033] = i[6033];
  assign o[6032] = i[6032];
  assign o[6031] = i[6031];
  assign o[6030] = i[6030];
  assign o[6029] = i[6029];
  assign o[6028] = i[6028];
  assign o[6027] = i[6027];
  assign o[6026] = i[6026];
  assign o[6025] = i[6025];
  assign o[6024] = i[6024];
  assign o[6023] = i[6023];
  assign o[6022] = i[6022];
  assign o[6021] = i[6021];
  assign o[6020] = i[6020];
  assign o[6019] = i[6019];
  assign o[6018] = i[6018];
  assign o[6017] = i[6017];
  assign o[6016] = i[6016];
  assign o[6015] = i[6015];
  assign o[6014] = i[6014];
  assign o[6013] = i[6013];
  assign o[6012] = i[6012];
  assign o[6011] = i[6011];
  assign o[6010] = i[6010];
  assign o[6009] = i[6009];
  assign o[6008] = i[6008];
  assign o[6007] = i[6007];
  assign o[6006] = i[6006];
  assign o[6005] = i[6005];
  assign o[6004] = i[6004];
  assign o[6003] = i[6003];
  assign o[6002] = i[6002];
  assign o[6001] = i[6001];
  assign o[6000] = i[6000];
  assign o[5999] = i[5999];
  assign o[5998] = i[5998];
  assign o[5997] = i[5997];
  assign o[5996] = i[5996];
  assign o[5995] = i[5995];
  assign o[5994] = i[5994];
  assign o[5993] = i[5993];
  assign o[5992] = i[5992];
  assign o[5991] = i[5991];
  assign o[5990] = i[5990];
  assign o[5989] = i[5989];
  assign o[5988] = i[5988];
  assign o[5987] = i[5987];
  assign o[5986] = i[5986];
  assign o[5985] = i[5985];
  assign o[5984] = i[5984];
  assign o[5983] = i[5983];
  assign o[5982] = i[5982];
  assign o[5981] = i[5981];
  assign o[5980] = i[5980];
  assign o[5979] = i[5979];
  assign o[5978] = i[5978];
  assign o[5977] = i[5977];
  assign o[5976] = i[5976];
  assign o[5975] = i[5975];
  assign o[5974] = i[5974];
  assign o[5973] = i[5973];
  assign o[5972] = i[5972];
  assign o[5971] = i[5971];
  assign o[5970] = i[5970];
  assign o[5969] = i[5969];
  assign o[5968] = i[5968];
  assign o[5967] = i[5967];
  assign o[5966] = i[5966];
  assign o[5965] = i[5965];
  assign o[5964] = i[5964];
  assign o[5963] = i[5963];
  assign o[5962] = i[5962];
  assign o[5961] = i[5961];
  assign o[5960] = i[5960];
  assign o[5959] = i[5959];
  assign o[5958] = i[5958];
  assign o[5957] = i[5957];
  assign o[5956] = i[5956];
  assign o[5955] = i[5955];
  assign o[5954] = i[5954];
  assign o[5953] = i[5953];
  assign o[5952] = i[5952];
  assign o[5951] = i[5951];
  assign o[5950] = i[5950];
  assign o[5949] = i[5949];
  assign o[5948] = i[5948];
  assign o[5947] = i[5947];
  assign o[5946] = i[5946];
  assign o[5945] = i[5945];
  assign o[5944] = i[5944];
  assign o[5943] = i[5943];
  assign o[5942] = i[5942];
  assign o[5941] = i[5941];
  assign o[5940] = i[5940];
  assign o[5939] = i[5939];
  assign o[5938] = i[5938];
  assign o[5937] = i[5937];
  assign o[5936] = i[5936];
  assign o[5935] = i[5935];
  assign o[5934] = i[5934];
  assign o[5933] = i[5933];
  assign o[5932] = i[5932];
  assign o[5931] = i[5931];
  assign o[5930] = i[5930];
  assign o[5929] = i[5929];
  assign o[5928] = i[5928];
  assign o[5927] = i[5927];
  assign o[5926] = i[5926];
  assign o[5925] = i[5925];
  assign o[5924] = i[5924];
  assign o[5923] = i[5923];
  assign o[5922] = i[5922];
  assign o[5921] = i[5921];
  assign o[5920] = i[5920];
  assign o[5919] = i[5919];
  assign o[5918] = i[5918];
  assign o[5917] = i[5917];
  assign o[5916] = i[5916];
  assign o[5915] = i[5915];
  assign o[5914] = i[5914];
  assign o[5913] = i[5913];
  assign o[5912] = i[5912];
  assign o[5911] = i[5911];
  assign o[5910] = i[5910];
  assign o[5909] = i[5909];
  assign o[5908] = i[5908];
  assign o[5907] = i[5907];
  assign o[5906] = i[5906];
  assign o[5905] = i[5905];
  assign o[5904] = i[5904];
  assign o[5903] = i[5903];
  assign o[5902] = i[5902];
  assign o[5901] = i[5901];
  assign o[5900] = i[5900];
  assign o[5899] = i[5899];
  assign o[5898] = i[5898];
  assign o[5897] = i[5897];
  assign o[5896] = i[5896];
  assign o[5895] = i[5895];
  assign o[5894] = i[5894];
  assign o[5893] = i[5893];
  assign o[5892] = i[5892];
  assign o[5891] = i[5891];
  assign o[5890] = i[5890];
  assign o[5889] = i[5889];
  assign o[5888] = i[5888];
  assign o[5887] = i[5887];
  assign o[5886] = i[5886];
  assign o[5885] = i[5885];
  assign o[5884] = i[5884];
  assign o[5883] = i[5883];
  assign o[5882] = i[5882];
  assign o[5881] = i[5881];
  assign o[5880] = i[5880];
  assign o[5879] = i[5879];
  assign o[5878] = i[5878];
  assign o[5877] = i[5877];
  assign o[5876] = i[5876];
  assign o[5875] = i[5875];
  assign o[5874] = i[5874];
  assign o[5873] = i[5873];
  assign o[5872] = i[5872];
  assign o[5871] = i[5871];
  assign o[5870] = i[5870];
  assign o[5869] = i[5869];
  assign o[5868] = i[5868];
  assign o[5867] = i[5867];
  assign o[5866] = i[5866];
  assign o[5865] = i[5865];
  assign o[5864] = i[5864];
  assign o[5863] = i[5863];
  assign o[5862] = i[5862];
  assign o[5861] = i[5861];
  assign o[5860] = i[5860];
  assign o[5859] = i[5859];
  assign o[5858] = i[5858];
  assign o[5857] = i[5857];
  assign o[5856] = i[5856];
  assign o[5855] = i[5855];
  assign o[5854] = i[5854];
  assign o[5853] = i[5853];
  assign o[5852] = i[5852];
  assign o[5851] = i[5851];
  assign o[5850] = i[5850];
  assign o[5849] = i[5849];
  assign o[5848] = i[5848];
  assign o[5847] = i[5847];
  assign o[5846] = i[5846];
  assign o[5845] = i[5845];
  assign o[5844] = i[5844];
  assign o[5843] = i[5843];
  assign o[5842] = i[5842];
  assign o[5841] = i[5841];
  assign o[5840] = i[5840];
  assign o[5839] = i[5839];
  assign o[5838] = i[5838];
  assign o[5837] = i[5837];
  assign o[5836] = i[5836];
  assign o[5835] = i[5835];
  assign o[5834] = i[5834];
  assign o[5833] = i[5833];
  assign o[5832] = i[5832];
  assign o[5831] = i[5831];
  assign o[5830] = i[5830];
  assign o[5829] = i[5829];
  assign o[5828] = i[5828];
  assign o[5827] = i[5827];
  assign o[5826] = i[5826];
  assign o[5825] = i[5825];
  assign o[5824] = i[5824];
  assign o[5823] = i[5823];
  assign o[5822] = i[5822];
  assign o[5821] = i[5821];
  assign o[5820] = i[5820];
  assign o[5819] = i[5819];
  assign o[5818] = i[5818];
  assign o[5817] = i[5817];
  assign o[5816] = i[5816];
  assign o[5815] = i[5815];
  assign o[5814] = i[5814];
  assign o[5813] = i[5813];
  assign o[5812] = i[5812];
  assign o[5811] = i[5811];
  assign o[5810] = i[5810];
  assign o[5809] = i[5809];
  assign o[5808] = i[5808];
  assign o[5807] = i[5807];
  assign o[5806] = i[5806];
  assign o[5805] = i[5805];
  assign o[5804] = i[5804];
  assign o[5803] = i[5803];
  assign o[5802] = i[5802];
  assign o[5801] = i[5801];
  assign o[5800] = i[5800];
  assign o[5799] = i[5799];
  assign o[5798] = i[5798];
  assign o[5797] = i[5797];
  assign o[5796] = i[5796];
  assign o[5795] = i[5795];
  assign o[5794] = i[5794];
  assign o[5793] = i[5793];
  assign o[5792] = i[5792];
  assign o[5791] = i[5791];
  assign o[5790] = i[5790];
  assign o[5789] = i[5789];
  assign o[5788] = i[5788];
  assign o[5787] = i[5787];
  assign o[5786] = i[5786];
  assign o[5785] = i[5785];
  assign o[5784] = i[5784];
  assign o[5783] = i[5783];
  assign o[5782] = i[5782];
  assign o[5781] = i[5781];
  assign o[5780] = i[5780];
  assign o[5779] = i[5779];
  assign o[5778] = i[5778];
  assign o[5777] = i[5777];
  assign o[5776] = i[5776];
  assign o[5775] = i[5775];
  assign o[5774] = i[5774];
  assign o[5773] = i[5773];
  assign o[5772] = i[5772];
  assign o[5771] = i[5771];
  assign o[5770] = i[5770];
  assign o[5769] = i[5769];
  assign o[5768] = i[5768];
  assign o[5767] = i[5767];
  assign o[5766] = i[5766];
  assign o[5765] = i[5765];
  assign o[5764] = i[5764];
  assign o[5763] = i[5763];
  assign o[5762] = i[5762];
  assign o[5761] = i[5761];
  assign o[5760] = i[5760];
  assign o[5759] = i[5759];
  assign o[5758] = i[5758];
  assign o[5757] = i[5757];
  assign o[5756] = i[5756];
  assign o[5755] = i[5755];
  assign o[5754] = i[5754];
  assign o[5753] = i[5753];
  assign o[5752] = i[5752];
  assign o[5751] = i[5751];
  assign o[5750] = i[5750];
  assign o[5749] = i[5749];
  assign o[5748] = i[5748];
  assign o[5747] = i[5747];
  assign o[5746] = i[5746];
  assign o[5745] = i[5745];
  assign o[5744] = i[5744];
  assign o[5743] = i[5743];
  assign o[5742] = i[5742];
  assign o[5741] = i[5741];
  assign o[5740] = i[5740];
  assign o[5739] = i[5739];
  assign o[5738] = i[5738];
  assign o[5737] = i[5737];
  assign o[5736] = i[5736];
  assign o[5735] = i[5735];
  assign o[5734] = i[5734];
  assign o[5733] = i[5733];
  assign o[5732] = i[5732];
  assign o[5731] = i[5731];
  assign o[5730] = i[5730];
  assign o[5729] = i[5729];
  assign o[5728] = i[5728];
  assign o[5727] = i[5727];
  assign o[5726] = i[5726];
  assign o[5725] = i[5725];
  assign o[5724] = i[5724];
  assign o[5723] = i[5723];
  assign o[5722] = i[5722];
  assign o[5721] = i[5721];
  assign o[5720] = i[5720];
  assign o[5719] = i[5719];
  assign o[5718] = i[5718];
  assign o[5717] = i[5717];
  assign o[5716] = i[5716];
  assign o[5715] = i[5715];
  assign o[5714] = i[5714];
  assign o[5713] = i[5713];
  assign o[5712] = i[5712];
  assign o[5711] = i[5711];
  assign o[5710] = i[5710];
  assign o[5709] = i[5709];
  assign o[5708] = i[5708];
  assign o[5707] = i[5707];
  assign o[5706] = i[5706];
  assign o[5705] = i[5705];
  assign o[5704] = i[5704];
  assign o[5703] = i[5703];
  assign o[5702] = i[5702];
  assign o[5701] = i[5701];
  assign o[5700] = i[5700];
  assign o[5699] = i[5699];
  assign o[5698] = i[5698];
  assign o[5697] = i[5697];
  assign o[5696] = i[5696];
  assign o[5695] = i[5695];
  assign o[5694] = i[5694];
  assign o[5693] = i[5693];
  assign o[5692] = i[5692];
  assign o[5691] = i[5691];
  assign o[5690] = i[5690];
  assign o[5689] = i[5689];
  assign o[5688] = i[5688];
  assign o[5687] = i[5687];
  assign o[5686] = i[5686];
  assign o[5685] = i[5685];
  assign o[5684] = i[5684];
  assign o[5683] = i[5683];
  assign o[5682] = i[5682];
  assign o[5681] = i[5681];
  assign o[5680] = i[5680];
  assign o[5679] = i[5679];
  assign o[5678] = i[5678];
  assign o[5677] = i[5677];
  assign o[5676] = i[5676];
  assign o[5675] = i[5675];
  assign o[5674] = i[5674];
  assign o[5673] = i[5673];
  assign o[5672] = i[5672];
  assign o[5671] = i[5671];
  assign o[5670] = i[5670];
  assign o[5669] = i[5669];
  assign o[5668] = i[5668];
  assign o[5667] = i[5667];
  assign o[5666] = i[5666];
  assign o[5665] = i[5665];
  assign o[5664] = i[5664];
  assign o[5663] = i[5663];
  assign o[5662] = i[5662];
  assign o[5661] = i[5661];
  assign o[5660] = i[5660];
  assign o[5659] = i[5659];
  assign o[5658] = i[5658];
  assign o[5657] = i[5657];
  assign o[5656] = i[5656];
  assign o[5655] = i[5655];
  assign o[5654] = i[5654];
  assign o[5653] = i[5653];
  assign o[5652] = i[5652];
  assign o[5651] = i[5651];
  assign o[5650] = i[5650];
  assign o[5649] = i[5649];
  assign o[5648] = i[5648];
  assign o[5647] = i[5647];
  assign o[5646] = i[5646];
  assign o[5645] = i[5645];
  assign o[5644] = i[5644];
  assign o[5643] = i[5643];
  assign o[5642] = i[5642];
  assign o[5641] = i[5641];
  assign o[5640] = i[5640];
  assign o[5639] = i[5639];
  assign o[5638] = i[5638];
  assign o[5637] = i[5637];
  assign o[5636] = i[5636];
  assign o[5635] = i[5635];
  assign o[5634] = i[5634];
  assign o[5633] = i[5633];
  assign o[5632] = i[5632];
  assign o[5631] = i[5631];
  assign o[5630] = i[5630];
  assign o[5629] = i[5629];
  assign o[5628] = i[5628];
  assign o[5627] = i[5627];
  assign o[5626] = i[5626];
  assign o[5625] = i[5625];
  assign o[5624] = i[5624];
  assign o[5623] = i[5623];
  assign o[5622] = i[5622];
  assign o[5621] = i[5621];
  assign o[5620] = i[5620];
  assign o[5619] = i[5619];
  assign o[5618] = i[5618];
  assign o[5617] = i[5617];
  assign o[5616] = i[5616];
  assign o[5615] = i[5615];
  assign o[5614] = i[5614];
  assign o[5613] = i[5613];
  assign o[5612] = i[5612];
  assign o[5611] = i[5611];
  assign o[5610] = i[5610];
  assign o[5609] = i[5609];
  assign o[5608] = i[5608];
  assign o[5607] = i[5607];
  assign o[5606] = i[5606];
  assign o[5605] = i[5605];
  assign o[5604] = i[5604];
  assign o[5603] = i[5603];
  assign o[5602] = i[5602];
  assign o[5601] = i[5601];
  assign o[5600] = i[5600];
  assign o[5599] = i[5599];
  assign o[5598] = i[5598];
  assign o[5597] = i[5597];
  assign o[5596] = i[5596];
  assign o[5595] = i[5595];
  assign o[5594] = i[5594];
  assign o[5593] = i[5593];
  assign o[5592] = i[5592];
  assign o[5591] = i[5591];
  assign o[5590] = i[5590];
  assign o[5589] = i[5589];
  assign o[5588] = i[5588];
  assign o[5587] = i[5587];
  assign o[5586] = i[5586];
  assign o[5585] = i[5585];
  assign o[5584] = i[5584];
  assign o[5583] = i[5583];
  assign o[5582] = i[5582];
  assign o[5581] = i[5581];
  assign o[5580] = i[5580];
  assign o[5579] = i[5579];
  assign o[5578] = i[5578];
  assign o[5577] = i[5577];
  assign o[5576] = i[5576];
  assign o[5575] = i[5575];
  assign o[5574] = i[5574];
  assign o[5573] = i[5573];
  assign o[5572] = i[5572];
  assign o[5571] = i[5571];
  assign o[5570] = i[5570];
  assign o[5569] = i[5569];
  assign o[5568] = i[5568];
  assign o[5567] = i[5567];
  assign o[5566] = i[5566];
  assign o[5565] = i[5565];
  assign o[5564] = i[5564];
  assign o[5563] = i[5563];
  assign o[5562] = i[5562];
  assign o[5561] = i[5561];
  assign o[5560] = i[5560];
  assign o[5559] = i[5559];
  assign o[5558] = i[5558];
  assign o[5557] = i[5557];
  assign o[5556] = i[5556];
  assign o[5555] = i[5555];
  assign o[5554] = i[5554];
  assign o[5553] = i[5553];
  assign o[5552] = i[5552];
  assign o[5551] = i[5551];
  assign o[5550] = i[5550];
  assign o[5549] = i[5549];
  assign o[5548] = i[5548];
  assign o[5547] = i[5547];
  assign o[5546] = i[5546];
  assign o[5545] = i[5545];
  assign o[5544] = i[5544];
  assign o[5543] = i[5543];
  assign o[5542] = i[5542];
  assign o[5541] = i[5541];
  assign o[5540] = i[5540];
  assign o[5539] = i[5539];
  assign o[5538] = i[5538];
  assign o[5537] = i[5537];
  assign o[5536] = i[5536];
  assign o[5535] = i[5535];
  assign o[5534] = i[5534];
  assign o[5533] = i[5533];
  assign o[5532] = i[5532];
  assign o[5531] = i[5531];
  assign o[5530] = i[5530];
  assign o[5529] = i[5529];
  assign o[5528] = i[5528];
  assign o[5527] = i[5527];
  assign o[5526] = i[5526];
  assign o[5525] = i[5525];
  assign o[5524] = i[5524];
  assign o[5523] = i[5523];
  assign o[5522] = i[5522];
  assign o[5521] = i[5521];
  assign o[5520] = i[5520];
  assign o[5519] = i[5519];
  assign o[5518] = i[5518];
  assign o[5517] = i[5517];
  assign o[5516] = i[5516];
  assign o[5515] = i[5515];
  assign o[5514] = i[5514];
  assign o[5513] = i[5513];
  assign o[5512] = i[5512];
  assign o[5511] = i[5511];
  assign o[5510] = i[5510];
  assign o[5509] = i[5509];
  assign o[5508] = i[5508];
  assign o[5507] = i[5507];
  assign o[5506] = i[5506];
  assign o[5505] = i[5505];
  assign o[5504] = i[5504];
  assign o[5503] = i[5503];
  assign o[5502] = i[5502];
  assign o[5501] = i[5501];
  assign o[5500] = i[5500];
  assign o[5499] = i[5499];
  assign o[5498] = i[5498];
  assign o[5497] = i[5497];
  assign o[5496] = i[5496];
  assign o[5495] = i[5495];
  assign o[5494] = i[5494];
  assign o[5493] = i[5493];
  assign o[5492] = i[5492];
  assign o[5491] = i[5491];
  assign o[5490] = i[5490];
  assign o[5489] = i[5489];
  assign o[5488] = i[5488];
  assign o[5487] = i[5487];
  assign o[5486] = i[5486];
  assign o[5485] = i[5485];
  assign o[5484] = i[5484];
  assign o[5483] = i[5483];
  assign o[5482] = i[5482];
  assign o[5481] = i[5481];
  assign o[5480] = i[5480];
  assign o[5479] = i[5479];
  assign o[5478] = i[5478];
  assign o[5477] = i[5477];
  assign o[5476] = i[5476];
  assign o[5475] = i[5475];
  assign o[5474] = i[5474];
  assign o[5473] = i[5473];
  assign o[5472] = i[5472];
  assign o[5471] = i[5471];
  assign o[5470] = i[5470];
  assign o[5469] = i[5469];
  assign o[5468] = i[5468];
  assign o[5467] = i[5467];
  assign o[5466] = i[5466];
  assign o[5465] = i[5465];
  assign o[5464] = i[5464];
  assign o[5463] = i[5463];
  assign o[5462] = i[5462];
  assign o[5461] = i[5461];
  assign o[5460] = i[5460];
  assign o[5459] = i[5459];
  assign o[5458] = i[5458];
  assign o[5457] = i[5457];
  assign o[5456] = i[5456];
  assign o[5455] = i[5455];
  assign o[5454] = i[5454];
  assign o[5453] = i[5453];
  assign o[5452] = i[5452];
  assign o[5451] = i[5451];
  assign o[5450] = i[5450];
  assign o[5449] = i[5449];
  assign o[5448] = i[5448];
  assign o[5447] = i[5447];
  assign o[5446] = i[5446];
  assign o[5445] = i[5445];
  assign o[5444] = i[5444];
  assign o[5443] = i[5443];
  assign o[5442] = i[5442];
  assign o[5441] = i[5441];
  assign o[5440] = i[5440];
  assign o[5439] = i[5439];
  assign o[5438] = i[5438];
  assign o[5437] = i[5437];
  assign o[5436] = i[5436];
  assign o[5435] = i[5435];
  assign o[5434] = i[5434];
  assign o[5433] = i[5433];
  assign o[5432] = i[5432];
  assign o[5431] = i[5431];
  assign o[5430] = i[5430];
  assign o[5429] = i[5429];
  assign o[5428] = i[5428];
  assign o[5427] = i[5427];
  assign o[5426] = i[5426];
  assign o[5425] = i[5425];
  assign o[5424] = i[5424];
  assign o[5423] = i[5423];
  assign o[5422] = i[5422];
  assign o[5421] = i[5421];
  assign o[5420] = i[5420];
  assign o[5419] = i[5419];
  assign o[5418] = i[5418];
  assign o[5417] = i[5417];
  assign o[5416] = i[5416];
  assign o[5415] = i[5415];
  assign o[5414] = i[5414];
  assign o[5413] = i[5413];
  assign o[5412] = i[5412];
  assign o[5411] = i[5411];
  assign o[5410] = i[5410];
  assign o[5409] = i[5409];
  assign o[5408] = i[5408];
  assign o[5407] = i[5407];
  assign o[5406] = i[5406];
  assign o[5405] = i[5405];
  assign o[5404] = i[5404];
  assign o[5403] = i[5403];
  assign o[5402] = i[5402];
  assign o[5401] = i[5401];
  assign o[5400] = i[5400];
  assign o[5399] = i[5399];
  assign o[5398] = i[5398];
  assign o[5397] = i[5397];
  assign o[5396] = i[5396];
  assign o[5395] = i[5395];
  assign o[5394] = i[5394];
  assign o[5393] = i[5393];
  assign o[5392] = i[5392];
  assign o[5391] = i[5391];
  assign o[5390] = i[5390];
  assign o[5389] = i[5389];
  assign o[5388] = i[5388];
  assign o[5387] = i[5387];
  assign o[5386] = i[5386];
  assign o[5385] = i[5385];
  assign o[5384] = i[5384];
  assign o[5383] = i[5383];
  assign o[5382] = i[5382];
  assign o[5381] = i[5381];
  assign o[5380] = i[5380];
  assign o[5379] = i[5379];
  assign o[5378] = i[5378];
  assign o[5377] = i[5377];
  assign o[5376] = i[5376];
  assign o[5375] = i[5375];
  assign o[5374] = i[5374];
  assign o[5373] = i[5373];
  assign o[5372] = i[5372];
  assign o[5371] = i[5371];
  assign o[5370] = i[5370];
  assign o[5369] = i[5369];
  assign o[5368] = i[5368];
  assign o[5367] = i[5367];
  assign o[5366] = i[5366];
  assign o[5365] = i[5365];
  assign o[5364] = i[5364];
  assign o[5363] = i[5363];
  assign o[5362] = i[5362];
  assign o[5361] = i[5361];
  assign o[5360] = i[5360];
  assign o[5359] = i[5359];
  assign o[5358] = i[5358];
  assign o[5357] = i[5357];
  assign o[5356] = i[5356];
  assign o[5355] = i[5355];
  assign o[5354] = i[5354];
  assign o[5353] = i[5353];
  assign o[5352] = i[5352];
  assign o[5351] = i[5351];
  assign o[5350] = i[5350];
  assign o[5349] = i[5349];
  assign o[5348] = i[5348];
  assign o[5347] = i[5347];
  assign o[5346] = i[5346];
  assign o[5345] = i[5345];
  assign o[5344] = i[5344];
  assign o[5343] = i[5343];
  assign o[5342] = i[5342];
  assign o[5341] = i[5341];
  assign o[5340] = i[5340];
  assign o[5339] = i[5339];
  assign o[5338] = i[5338];
  assign o[5337] = i[5337];
  assign o[5336] = i[5336];
  assign o[5335] = i[5335];
  assign o[5334] = i[5334];
  assign o[5333] = i[5333];
  assign o[5332] = i[5332];
  assign o[5331] = i[5331];
  assign o[5330] = i[5330];
  assign o[5329] = i[5329];
  assign o[5328] = i[5328];
  assign o[5327] = i[5327];
  assign o[5326] = i[5326];
  assign o[5325] = i[5325];
  assign o[5324] = i[5324];
  assign o[5323] = i[5323];
  assign o[5322] = i[5322];
  assign o[5321] = i[5321];
  assign o[5320] = i[5320];
  assign o[5319] = i[5319];
  assign o[5318] = i[5318];
  assign o[5317] = i[5317];
  assign o[5316] = i[5316];
  assign o[5315] = i[5315];
  assign o[5314] = i[5314];
  assign o[5313] = i[5313];
  assign o[5312] = i[5312];
  assign o[5311] = i[5311];
  assign o[5310] = i[5310];
  assign o[5309] = i[5309];
  assign o[5308] = i[5308];
  assign o[5307] = i[5307];
  assign o[5306] = i[5306];
  assign o[5305] = i[5305];
  assign o[5304] = i[5304];
  assign o[5303] = i[5303];
  assign o[5302] = i[5302];
  assign o[5301] = i[5301];
  assign o[5300] = i[5300];
  assign o[5299] = i[5299];
  assign o[5298] = i[5298];
  assign o[5297] = i[5297];
  assign o[5296] = i[5296];
  assign o[5295] = i[5295];
  assign o[5294] = i[5294];
  assign o[5293] = i[5293];
  assign o[5292] = i[5292];
  assign o[5291] = i[5291];
  assign o[5290] = i[5290];
  assign o[5289] = i[5289];
  assign o[5288] = i[5288];
  assign o[5287] = i[5287];
  assign o[5286] = i[5286];
  assign o[5285] = i[5285];
  assign o[5284] = i[5284];
  assign o[5283] = i[5283];
  assign o[5282] = i[5282];
  assign o[5281] = i[5281];
  assign o[5280] = i[5280];
  assign o[5279] = i[5279];
  assign o[5278] = i[5278];
  assign o[5277] = i[5277];
  assign o[5276] = i[5276];
  assign o[5275] = i[5275];
  assign o[5274] = i[5274];
  assign o[5273] = i[5273];
  assign o[5272] = i[5272];
  assign o[5271] = i[5271];
  assign o[5270] = i[5270];
  assign o[5269] = i[5269];
  assign o[5268] = i[5268];
  assign o[5267] = i[5267];
  assign o[5266] = i[5266];
  assign o[5265] = i[5265];
  assign o[5264] = i[5264];
  assign o[5263] = i[5263];
  assign o[5262] = i[5262];
  assign o[5261] = i[5261];
  assign o[5260] = i[5260];
  assign o[5259] = i[5259];
  assign o[5258] = i[5258];
  assign o[5257] = i[5257];
  assign o[5256] = i[5256];
  assign o[5255] = i[5255];
  assign o[5254] = i[5254];
  assign o[5253] = i[5253];
  assign o[5252] = i[5252];
  assign o[5251] = i[5251];
  assign o[5250] = i[5250];
  assign o[5249] = i[5249];
  assign o[5248] = i[5248];
  assign o[5247] = i[5247];
  assign o[5246] = i[5246];
  assign o[5245] = i[5245];
  assign o[5244] = i[5244];
  assign o[5243] = i[5243];
  assign o[5242] = i[5242];
  assign o[5241] = i[5241];
  assign o[5240] = i[5240];
  assign o[5239] = i[5239];
  assign o[5238] = i[5238];
  assign o[5237] = i[5237];
  assign o[5236] = i[5236];
  assign o[5235] = i[5235];
  assign o[5234] = i[5234];
  assign o[5233] = i[5233];
  assign o[5232] = i[5232];
  assign o[5231] = i[5231];
  assign o[5230] = i[5230];
  assign o[5229] = i[5229];
  assign o[5228] = i[5228];
  assign o[5227] = i[5227];
  assign o[5226] = i[5226];
  assign o[5225] = i[5225];
  assign o[5224] = i[5224];
  assign o[5223] = i[5223];
  assign o[5222] = i[5222];
  assign o[5221] = i[5221];
  assign o[5220] = i[5220];
  assign o[5219] = i[5219];
  assign o[5218] = i[5218];
  assign o[5217] = i[5217];
  assign o[5216] = i[5216];
  assign o[5215] = i[5215];
  assign o[5214] = i[5214];
  assign o[5213] = i[5213];
  assign o[5212] = i[5212];
  assign o[5211] = i[5211];
  assign o[5210] = i[5210];
  assign o[5209] = i[5209];
  assign o[5208] = i[5208];
  assign o[5207] = i[5207];
  assign o[5206] = i[5206];
  assign o[5205] = i[5205];
  assign o[5204] = i[5204];
  assign o[5203] = i[5203];
  assign o[5202] = i[5202];
  assign o[5201] = i[5201];
  assign o[5200] = i[5200];
  assign o[5199] = i[5199];
  assign o[5198] = i[5198];
  assign o[5197] = i[5197];
  assign o[5196] = i[5196];
  assign o[5195] = i[5195];
  assign o[5194] = i[5194];
  assign o[5193] = i[5193];
  assign o[5192] = i[5192];
  assign o[5191] = i[5191];
  assign o[5190] = i[5190];
  assign o[5189] = i[5189];
  assign o[5188] = i[5188];
  assign o[5187] = i[5187];
  assign o[5186] = i[5186];
  assign o[5185] = i[5185];
  assign o[5184] = i[5184];
  assign o[5183] = i[5183];
  assign o[5182] = i[5182];
  assign o[5181] = i[5181];
  assign o[5180] = i[5180];
  assign o[5179] = i[5179];
  assign o[5178] = i[5178];
  assign o[5177] = i[5177];
  assign o[5176] = i[5176];
  assign o[5175] = i[5175];
  assign o[5174] = i[5174];
  assign o[5173] = i[5173];
  assign o[5172] = i[5172];
  assign o[5171] = i[5171];
  assign o[5170] = i[5170];
  assign o[5169] = i[5169];
  assign o[5168] = i[5168];
  assign o[5167] = i[5167];
  assign o[5166] = i[5166];
  assign o[5165] = i[5165];
  assign o[5164] = i[5164];
  assign o[5163] = i[5163];
  assign o[5162] = i[5162];
  assign o[5161] = i[5161];
  assign o[5160] = i[5160];
  assign o[5159] = i[5159];
  assign o[5158] = i[5158];
  assign o[5157] = i[5157];
  assign o[5156] = i[5156];
  assign o[5155] = i[5155];
  assign o[5154] = i[5154];
  assign o[5153] = i[5153];
  assign o[5152] = i[5152];
  assign o[5151] = i[5151];
  assign o[5150] = i[5150];
  assign o[5149] = i[5149];
  assign o[5148] = i[5148];
  assign o[5147] = i[5147];
  assign o[5146] = i[5146];
  assign o[5145] = i[5145];
  assign o[5144] = i[5144];
  assign o[5143] = i[5143];
  assign o[5142] = i[5142];
  assign o[5141] = i[5141];
  assign o[5140] = i[5140];
  assign o[5139] = i[5139];
  assign o[5138] = i[5138];
  assign o[5137] = i[5137];
  assign o[5136] = i[5136];
  assign o[5135] = i[5135];
  assign o[5134] = i[5134];
  assign o[5133] = i[5133];
  assign o[5132] = i[5132];
  assign o[5131] = i[5131];
  assign o[5130] = i[5130];
  assign o[5129] = i[5129];
  assign o[5128] = i[5128];
  assign o[5127] = i[5127];
  assign o[5126] = i[5126];
  assign o[5125] = i[5125];
  assign o[5124] = i[5124];
  assign o[5123] = i[5123];
  assign o[5122] = i[5122];
  assign o[5121] = i[5121];
  assign o[5120] = i[5120];
  assign o[5119] = i[5119];
  assign o[5118] = i[5118];
  assign o[5117] = i[5117];
  assign o[5116] = i[5116];
  assign o[5115] = i[5115];
  assign o[5114] = i[5114];
  assign o[5113] = i[5113];
  assign o[5112] = i[5112];
  assign o[5111] = i[5111];
  assign o[5110] = i[5110];
  assign o[5109] = i[5109];
  assign o[5108] = i[5108];
  assign o[5107] = i[5107];
  assign o[5106] = i[5106];
  assign o[5105] = i[5105];
  assign o[5104] = i[5104];
  assign o[5103] = i[5103];
  assign o[5102] = i[5102];
  assign o[5101] = i[5101];
  assign o[5100] = i[5100];
  assign o[5099] = i[5099];
  assign o[5098] = i[5098];
  assign o[5097] = i[5097];
  assign o[5096] = i[5096];
  assign o[5095] = i[5095];
  assign o[5094] = i[5094];
  assign o[5093] = i[5093];
  assign o[5092] = i[5092];
  assign o[5091] = i[5091];
  assign o[5090] = i[5090];
  assign o[5089] = i[5089];
  assign o[5088] = i[5088];
  assign o[5087] = i[5087];
  assign o[5086] = i[5086];
  assign o[5085] = i[5085];
  assign o[5084] = i[5084];
  assign o[5083] = i[5083];
  assign o[5082] = i[5082];
  assign o[5081] = i[5081];
  assign o[5080] = i[5080];
  assign o[5079] = i[5079];
  assign o[5078] = i[5078];
  assign o[5077] = i[5077];
  assign o[5076] = i[5076];
  assign o[5075] = i[5075];
  assign o[5074] = i[5074];
  assign o[5073] = i[5073];
  assign o[5072] = i[5072];
  assign o[5071] = i[5071];
  assign o[5070] = i[5070];
  assign o[5069] = i[5069];
  assign o[5068] = i[5068];
  assign o[5067] = i[5067];
  assign o[5066] = i[5066];
  assign o[5065] = i[5065];
  assign o[5064] = i[5064];
  assign o[5063] = i[5063];
  assign o[5062] = i[5062];
  assign o[5061] = i[5061];
  assign o[5060] = i[5060];
  assign o[5059] = i[5059];
  assign o[5058] = i[5058];
  assign o[5057] = i[5057];
  assign o[5056] = i[5056];
  assign o[5055] = i[5055];
  assign o[5054] = i[5054];
  assign o[5053] = i[5053];
  assign o[5052] = i[5052];
  assign o[5051] = i[5051];
  assign o[5050] = i[5050];
  assign o[5049] = i[5049];
  assign o[5048] = i[5048];
  assign o[5047] = i[5047];
  assign o[5046] = i[5046];
  assign o[5045] = i[5045];
  assign o[5044] = i[5044];
  assign o[5043] = i[5043];
  assign o[5042] = i[5042];
  assign o[5041] = i[5041];
  assign o[5040] = i[5040];
  assign o[5039] = i[5039];
  assign o[5038] = i[5038];
  assign o[5037] = i[5037];
  assign o[5036] = i[5036];
  assign o[5035] = i[5035];
  assign o[5034] = i[5034];
  assign o[5033] = i[5033];
  assign o[5032] = i[5032];
  assign o[5031] = i[5031];
  assign o[5030] = i[5030];
  assign o[5029] = i[5029];
  assign o[5028] = i[5028];
  assign o[5027] = i[5027];
  assign o[5026] = i[5026];
  assign o[5025] = i[5025];
  assign o[5024] = i[5024];
  assign o[5023] = i[5023];
  assign o[5022] = i[5022];
  assign o[5021] = i[5021];
  assign o[5020] = i[5020];
  assign o[5019] = i[5019];
  assign o[5018] = i[5018];
  assign o[5017] = i[5017];
  assign o[5016] = i[5016];
  assign o[5015] = i[5015];
  assign o[5014] = i[5014];
  assign o[5013] = i[5013];
  assign o[5012] = i[5012];
  assign o[5011] = i[5011];
  assign o[5010] = i[5010];
  assign o[5009] = i[5009];
  assign o[5008] = i[5008];
  assign o[5007] = i[5007];
  assign o[5006] = i[5006];
  assign o[5005] = i[5005];
  assign o[5004] = i[5004];
  assign o[5003] = i[5003];
  assign o[5002] = i[5002];
  assign o[5001] = i[5001];
  assign o[5000] = i[5000];
  assign o[4999] = i[4999];
  assign o[4998] = i[4998];
  assign o[4997] = i[4997];
  assign o[4996] = i[4996];
  assign o[4995] = i[4995];
  assign o[4994] = i[4994];
  assign o[4993] = i[4993];
  assign o[4992] = i[4992];
  assign o[4991] = i[4991];
  assign o[4990] = i[4990];
  assign o[4989] = i[4989];
  assign o[4988] = i[4988];
  assign o[4987] = i[4987];
  assign o[4986] = i[4986];
  assign o[4985] = i[4985];
  assign o[4984] = i[4984];
  assign o[4983] = i[4983];
  assign o[4982] = i[4982];
  assign o[4981] = i[4981];
  assign o[4980] = i[4980];
  assign o[4979] = i[4979];
  assign o[4978] = i[4978];
  assign o[4977] = i[4977];
  assign o[4976] = i[4976];
  assign o[4975] = i[4975];
  assign o[4974] = i[4974];
  assign o[4973] = i[4973];
  assign o[4972] = i[4972];
  assign o[4971] = i[4971];
  assign o[4970] = i[4970];
  assign o[4969] = i[4969];
  assign o[4968] = i[4968];
  assign o[4967] = i[4967];
  assign o[4966] = i[4966];
  assign o[4965] = i[4965];
  assign o[4964] = i[4964];
  assign o[4963] = i[4963];
  assign o[4962] = i[4962];
  assign o[4961] = i[4961];
  assign o[4960] = i[4960];
  assign o[4959] = i[4959];
  assign o[4958] = i[4958];
  assign o[4957] = i[4957];
  assign o[4956] = i[4956];
  assign o[4955] = i[4955];
  assign o[4954] = i[4954];
  assign o[4953] = i[4953];
  assign o[4952] = i[4952];
  assign o[4951] = i[4951];
  assign o[4950] = i[4950];
  assign o[4949] = i[4949];
  assign o[4948] = i[4948];
  assign o[4947] = i[4947];
  assign o[4946] = i[4946];
  assign o[4945] = i[4945];
  assign o[4944] = i[4944];
  assign o[4943] = i[4943];
  assign o[4942] = i[4942];
  assign o[4941] = i[4941];
  assign o[4940] = i[4940];
  assign o[4939] = i[4939];
  assign o[4938] = i[4938];
  assign o[4937] = i[4937];
  assign o[4936] = i[4936];
  assign o[4935] = i[4935];
  assign o[4934] = i[4934];
  assign o[4933] = i[4933];
  assign o[4932] = i[4932];
  assign o[4931] = i[4931];
  assign o[4930] = i[4930];
  assign o[4929] = i[4929];
  assign o[4928] = i[4928];
  assign o[4927] = i[4927];
  assign o[4926] = i[4926];
  assign o[4925] = i[4925];
  assign o[4924] = i[4924];
  assign o[4923] = i[4923];
  assign o[4922] = i[4922];
  assign o[4921] = i[4921];
  assign o[4920] = i[4920];
  assign o[4919] = i[4919];
  assign o[4918] = i[4918];
  assign o[4917] = i[4917];
  assign o[4916] = i[4916];
  assign o[4915] = i[4915];
  assign o[4914] = i[4914];
  assign o[4913] = i[4913];
  assign o[4912] = i[4912];
  assign o[4911] = i[4911];
  assign o[4910] = i[4910];
  assign o[4909] = i[4909];
  assign o[4908] = i[4908];
  assign o[4907] = i[4907];
  assign o[4906] = i[4906];
  assign o[4905] = i[4905];
  assign o[4904] = i[4904];
  assign o[4903] = i[4903];
  assign o[4902] = i[4902];
  assign o[4901] = i[4901];
  assign o[4900] = i[4900];
  assign o[4899] = i[4899];
  assign o[4898] = i[4898];
  assign o[4897] = i[4897];
  assign o[4896] = i[4896];
  assign o[4895] = i[4895];
  assign o[4894] = i[4894];
  assign o[4893] = i[4893];
  assign o[4892] = i[4892];
  assign o[4891] = i[4891];
  assign o[4890] = i[4890];
  assign o[4889] = i[4889];
  assign o[4888] = i[4888];
  assign o[4887] = i[4887];
  assign o[4886] = i[4886];
  assign o[4885] = i[4885];
  assign o[4884] = i[4884];
  assign o[4883] = i[4883];
  assign o[4882] = i[4882];
  assign o[4881] = i[4881];
  assign o[4880] = i[4880];
  assign o[4879] = i[4879];
  assign o[4878] = i[4878];
  assign o[4877] = i[4877];
  assign o[4876] = i[4876];
  assign o[4875] = i[4875];
  assign o[4874] = i[4874];
  assign o[4873] = i[4873];
  assign o[4872] = i[4872];
  assign o[4871] = i[4871];
  assign o[4870] = i[4870];
  assign o[4869] = i[4869];
  assign o[4868] = i[4868];
  assign o[4867] = i[4867];
  assign o[4866] = i[4866];
  assign o[4865] = i[4865];
  assign o[4864] = i[4864];
  assign o[4863] = i[4863];
  assign o[4862] = i[4862];
  assign o[4861] = i[4861];
  assign o[4860] = i[4860];
  assign o[4859] = i[4859];
  assign o[4858] = i[4858];
  assign o[4857] = i[4857];
  assign o[4856] = i[4856];
  assign o[4855] = i[4855];
  assign o[4854] = i[4854];
  assign o[4853] = i[4853];
  assign o[4852] = i[4852];
  assign o[4851] = i[4851];
  assign o[4850] = i[4850];
  assign o[4849] = i[4849];
  assign o[4848] = i[4848];
  assign o[4847] = i[4847];
  assign o[4846] = i[4846];
  assign o[4845] = i[4845];
  assign o[4844] = i[4844];
  assign o[4843] = i[4843];
  assign o[4842] = i[4842];
  assign o[4841] = i[4841];
  assign o[4840] = i[4840];
  assign o[4839] = i[4839];
  assign o[4838] = i[4838];
  assign o[4837] = i[4837];
  assign o[4836] = i[4836];
  assign o[4835] = i[4835];
  assign o[4834] = i[4834];
  assign o[4833] = i[4833];
  assign o[4832] = i[4832];
  assign o[4831] = i[4831];
  assign o[4830] = i[4830];
  assign o[4829] = i[4829];
  assign o[4828] = i[4828];
  assign o[4827] = i[4827];
  assign o[4826] = i[4826];
  assign o[4825] = i[4825];
  assign o[4824] = i[4824];
  assign o[4823] = i[4823];
  assign o[4822] = i[4822];
  assign o[4821] = i[4821];
  assign o[4820] = i[4820];
  assign o[4819] = i[4819];
  assign o[4818] = i[4818];
  assign o[4817] = i[4817];
  assign o[4816] = i[4816];
  assign o[4815] = i[4815];
  assign o[4814] = i[4814];
  assign o[4813] = i[4813];
  assign o[4812] = i[4812];
  assign o[4811] = i[4811];
  assign o[4810] = i[4810];
  assign o[4809] = i[4809];
  assign o[4808] = i[4808];
  assign o[4807] = i[4807];
  assign o[4806] = i[4806];
  assign o[4805] = i[4805];
  assign o[4804] = i[4804];
  assign o[4803] = i[4803];
  assign o[4802] = i[4802];
  assign o[4801] = i[4801];
  assign o[4800] = i[4800];
  assign o[4799] = i[4799];
  assign o[4798] = i[4798];
  assign o[4797] = i[4797];
  assign o[4796] = i[4796];
  assign o[4795] = i[4795];
  assign o[4794] = i[4794];
  assign o[4793] = i[4793];
  assign o[4792] = i[4792];
  assign o[4791] = i[4791];
  assign o[4790] = i[4790];
  assign o[4789] = i[4789];
  assign o[4788] = i[4788];
  assign o[4787] = i[4787];
  assign o[4786] = i[4786];
  assign o[4785] = i[4785];
  assign o[4784] = i[4784];
  assign o[4783] = i[4783];
  assign o[4782] = i[4782];
  assign o[4781] = i[4781];
  assign o[4780] = i[4780];
  assign o[4779] = i[4779];
  assign o[4778] = i[4778];
  assign o[4777] = i[4777];
  assign o[4776] = i[4776];
  assign o[4775] = i[4775];
  assign o[4774] = i[4774];
  assign o[4773] = i[4773];
  assign o[4772] = i[4772];
  assign o[4771] = i[4771];
  assign o[4770] = i[4770];
  assign o[4769] = i[4769];
  assign o[4768] = i[4768];
  assign o[4767] = i[4767];
  assign o[4766] = i[4766];
  assign o[4765] = i[4765];
  assign o[4764] = i[4764];
  assign o[4763] = i[4763];
  assign o[4762] = i[4762];
  assign o[4761] = i[4761];
  assign o[4760] = i[4760];
  assign o[4759] = i[4759];
  assign o[4758] = i[4758];
  assign o[4757] = i[4757];
  assign o[4756] = i[4756];
  assign o[4755] = i[4755];
  assign o[4754] = i[4754];
  assign o[4753] = i[4753];
  assign o[4752] = i[4752];
  assign o[4751] = i[4751];
  assign o[4750] = i[4750];
  assign o[4749] = i[4749];
  assign o[4748] = i[4748];
  assign o[4747] = i[4747];
  assign o[4746] = i[4746];
  assign o[4745] = i[4745];
  assign o[4744] = i[4744];
  assign o[4743] = i[4743];
  assign o[4742] = i[4742];
  assign o[4741] = i[4741];
  assign o[4740] = i[4740];
  assign o[4739] = i[4739];
  assign o[4738] = i[4738];
  assign o[4737] = i[4737];
  assign o[4736] = i[4736];
  assign o[4735] = i[4735];
  assign o[4734] = i[4734];
  assign o[4733] = i[4733];
  assign o[4732] = i[4732];
  assign o[4731] = i[4731];
  assign o[4730] = i[4730];
  assign o[4729] = i[4729];
  assign o[4728] = i[4728];
  assign o[4727] = i[4727];
  assign o[4726] = i[4726];
  assign o[4725] = i[4725];
  assign o[4724] = i[4724];
  assign o[4723] = i[4723];
  assign o[4722] = i[4722];
  assign o[4721] = i[4721];
  assign o[4720] = i[4720];
  assign o[4719] = i[4719];
  assign o[4718] = i[4718];
  assign o[4717] = i[4717];
  assign o[4716] = i[4716];
  assign o[4715] = i[4715];
  assign o[4714] = i[4714];
  assign o[4713] = i[4713];
  assign o[4712] = i[4712];
  assign o[4711] = i[4711];
  assign o[4710] = i[4710];
  assign o[4709] = i[4709];
  assign o[4708] = i[4708];
  assign o[4707] = i[4707];
  assign o[4706] = i[4706];
  assign o[4705] = i[4705];
  assign o[4704] = i[4704];
  assign o[4703] = i[4703];
  assign o[4702] = i[4702];
  assign o[4701] = i[4701];
  assign o[4700] = i[4700];
  assign o[4699] = i[4699];
  assign o[4698] = i[4698];
  assign o[4697] = i[4697];
  assign o[4696] = i[4696];
  assign o[4695] = i[4695];
  assign o[4694] = i[4694];
  assign o[4693] = i[4693];
  assign o[4692] = i[4692];
  assign o[4691] = i[4691];
  assign o[4690] = i[4690];
  assign o[4689] = i[4689];
  assign o[4688] = i[4688];
  assign o[4687] = i[4687];
  assign o[4686] = i[4686];
  assign o[4685] = i[4685];
  assign o[4684] = i[4684];
  assign o[4683] = i[4683];
  assign o[4682] = i[4682];
  assign o[4681] = i[4681];
  assign o[4680] = i[4680];
  assign o[4679] = i[4679];
  assign o[4678] = i[4678];
  assign o[4677] = i[4677];
  assign o[4676] = i[4676];
  assign o[4675] = i[4675];
  assign o[4674] = i[4674];
  assign o[4673] = i[4673];
  assign o[4672] = i[4672];
  assign o[4671] = i[4671];
  assign o[4670] = i[4670];
  assign o[4669] = i[4669];
  assign o[4668] = i[4668];
  assign o[4667] = i[4667];
  assign o[4666] = i[4666];
  assign o[4665] = i[4665];
  assign o[4664] = i[4664];
  assign o[4663] = i[4663];
  assign o[4662] = i[4662];
  assign o[4661] = i[4661];
  assign o[4660] = i[4660];
  assign o[4659] = i[4659];
  assign o[4658] = i[4658];
  assign o[4657] = i[4657];
  assign o[4656] = i[4656];
  assign o[4655] = i[4655];
  assign o[4654] = i[4654];
  assign o[4653] = i[4653];
  assign o[4652] = i[4652];
  assign o[4651] = i[4651];
  assign o[4650] = i[4650];
  assign o[4649] = i[4649];
  assign o[4648] = i[4648];
  assign o[4647] = i[4647];
  assign o[4646] = i[4646];
  assign o[4645] = i[4645];
  assign o[4644] = i[4644];
  assign o[4643] = i[4643];
  assign o[4642] = i[4642];
  assign o[4641] = i[4641];
  assign o[4640] = i[4640];
  assign o[4639] = i[4639];
  assign o[4638] = i[4638];
  assign o[4637] = i[4637];
  assign o[4636] = i[4636];
  assign o[4635] = i[4635];
  assign o[4634] = i[4634];
  assign o[4633] = i[4633];
  assign o[4632] = i[4632];
  assign o[4631] = i[4631];
  assign o[4630] = i[4630];
  assign o[4629] = i[4629];
  assign o[4628] = i[4628];
  assign o[4627] = i[4627];
  assign o[4626] = i[4626];
  assign o[4625] = i[4625];
  assign o[4624] = i[4624];
  assign o[4623] = i[4623];
  assign o[4622] = i[4622];
  assign o[4621] = i[4621];
  assign o[4620] = i[4620];
  assign o[4619] = i[4619];
  assign o[4618] = i[4618];
  assign o[4617] = i[4617];
  assign o[4616] = i[4616];
  assign o[4615] = i[4615];
  assign o[4614] = i[4614];
  assign o[4613] = i[4613];
  assign o[4612] = i[4612];
  assign o[4611] = i[4611];
  assign o[4610] = i[4610];
  assign o[4609] = i[4609];
  assign o[4608] = i[4608];
  assign o[4607] = i[4607];
  assign o[4606] = i[4606];
  assign o[4605] = i[4605];
  assign o[4604] = i[4604];
  assign o[4603] = i[4603];
  assign o[4602] = i[4602];
  assign o[4601] = i[4601];
  assign o[4600] = i[4600];
  assign o[4599] = i[4599];
  assign o[4598] = i[4598];
  assign o[4597] = i[4597];
  assign o[4596] = i[4596];
  assign o[4595] = i[4595];
  assign o[4594] = i[4594];
  assign o[4593] = i[4593];
  assign o[4592] = i[4592];
  assign o[4591] = i[4591];
  assign o[4590] = i[4590];
  assign o[4589] = i[4589];
  assign o[4588] = i[4588];
  assign o[4587] = i[4587];
  assign o[4586] = i[4586];
  assign o[4585] = i[4585];
  assign o[4584] = i[4584];
  assign o[4583] = i[4583];
  assign o[4582] = i[4582];
  assign o[4581] = i[4581];
  assign o[4580] = i[4580];
  assign o[4579] = i[4579];
  assign o[4578] = i[4578];
  assign o[4577] = i[4577];
  assign o[4576] = i[4576];
  assign o[4575] = i[4575];
  assign o[4574] = i[4574];
  assign o[4573] = i[4573];
  assign o[4572] = i[4572];
  assign o[4571] = i[4571];
  assign o[4570] = i[4570];
  assign o[4569] = i[4569];
  assign o[4568] = i[4568];
  assign o[4567] = i[4567];
  assign o[4566] = i[4566];
  assign o[4565] = i[4565];
  assign o[4564] = i[4564];
  assign o[4563] = i[4563];
  assign o[4562] = i[4562];
  assign o[4561] = i[4561];
  assign o[4560] = i[4560];
  assign o[4559] = i[4559];
  assign o[4558] = i[4558];
  assign o[4557] = i[4557];
  assign o[4556] = i[4556];
  assign o[4555] = i[4555];
  assign o[4554] = i[4554];
  assign o[4553] = i[4553];
  assign o[4552] = i[4552];
  assign o[4551] = i[4551];
  assign o[4550] = i[4550];
  assign o[4549] = i[4549];
  assign o[4548] = i[4548];
  assign o[4547] = i[4547];
  assign o[4546] = i[4546];
  assign o[4545] = i[4545];
  assign o[4544] = i[4544];
  assign o[4543] = i[4543];
  assign o[4542] = i[4542];
  assign o[4541] = i[4541];
  assign o[4540] = i[4540];
  assign o[4539] = i[4539];
  assign o[4538] = i[4538];
  assign o[4537] = i[4537];
  assign o[4536] = i[4536];
  assign o[4535] = i[4535];
  assign o[4534] = i[4534];
  assign o[4533] = i[4533];
  assign o[4532] = i[4532];
  assign o[4531] = i[4531];
  assign o[4530] = i[4530];
  assign o[4529] = i[4529];
  assign o[4528] = i[4528];
  assign o[4527] = i[4527];
  assign o[4526] = i[4526];
  assign o[4525] = i[4525];
  assign o[4524] = i[4524];
  assign o[4523] = i[4523];
  assign o[4522] = i[4522];
  assign o[4521] = i[4521];
  assign o[4520] = i[4520];
  assign o[4519] = i[4519];
  assign o[4518] = i[4518];
  assign o[4517] = i[4517];
  assign o[4516] = i[4516];
  assign o[4515] = i[4515];
  assign o[4514] = i[4514];
  assign o[4513] = i[4513];
  assign o[4512] = i[4512];
  assign o[4511] = i[4511];
  assign o[4510] = i[4510];
  assign o[4509] = i[4509];
  assign o[4508] = i[4508];
  assign o[4507] = i[4507];
  assign o[4506] = i[4506];
  assign o[4505] = i[4505];
  assign o[4504] = i[4504];
  assign o[4503] = i[4503];
  assign o[4502] = i[4502];
  assign o[4501] = i[4501];
  assign o[4500] = i[4500];
  assign o[4499] = i[4499];
  assign o[4498] = i[4498];
  assign o[4497] = i[4497];
  assign o[4496] = i[4496];
  assign o[4495] = i[4495];
  assign o[4494] = i[4494];
  assign o[4493] = i[4493];
  assign o[4492] = i[4492];
  assign o[4491] = i[4491];
  assign o[4490] = i[4490];
  assign o[4489] = i[4489];
  assign o[4488] = i[4488];
  assign o[4487] = i[4487];
  assign o[4486] = i[4486];
  assign o[4485] = i[4485];
  assign o[4484] = i[4484];
  assign o[4483] = i[4483];
  assign o[4482] = i[4482];
  assign o[4481] = i[4481];
  assign o[4480] = i[4480];
  assign o[4479] = i[4479];
  assign o[4478] = i[4478];
  assign o[4477] = i[4477];
  assign o[4476] = i[4476];
  assign o[4475] = i[4475];
  assign o[4474] = i[4474];
  assign o[4473] = i[4473];
  assign o[4472] = i[4472];
  assign o[4471] = i[4471];
  assign o[4470] = i[4470];
  assign o[4469] = i[4469];
  assign o[4468] = i[4468];
  assign o[4467] = i[4467];
  assign o[4466] = i[4466];
  assign o[4465] = i[4465];
  assign o[4464] = i[4464];
  assign o[4463] = i[4463];
  assign o[4462] = i[4462];
  assign o[4461] = i[4461];
  assign o[4460] = i[4460];
  assign o[4459] = i[4459];
  assign o[4458] = i[4458];
  assign o[4457] = i[4457];
  assign o[4456] = i[4456];
  assign o[4455] = i[4455];
  assign o[4454] = i[4454];
  assign o[4453] = i[4453];
  assign o[4452] = i[4452];
  assign o[4451] = i[4451];
  assign o[4450] = i[4450];
  assign o[4449] = i[4449];
  assign o[4448] = i[4448];
  assign o[4447] = i[4447];
  assign o[4446] = i[4446];
  assign o[4445] = i[4445];
  assign o[4444] = i[4444];
  assign o[4443] = i[4443];
  assign o[4442] = i[4442];
  assign o[4441] = i[4441];
  assign o[4440] = i[4440];
  assign o[4439] = i[4439];
  assign o[4438] = i[4438];
  assign o[4437] = i[4437];
  assign o[4436] = i[4436];
  assign o[4435] = i[4435];
  assign o[4434] = i[4434];
  assign o[4433] = i[4433];
  assign o[4432] = i[4432];
  assign o[4431] = i[4431];
  assign o[4430] = i[4430];
  assign o[4429] = i[4429];
  assign o[4428] = i[4428];
  assign o[4427] = i[4427];
  assign o[4426] = i[4426];
  assign o[4425] = i[4425];
  assign o[4424] = i[4424];
  assign o[4423] = i[4423];
  assign o[4422] = i[4422];
  assign o[4421] = i[4421];
  assign o[4420] = i[4420];
  assign o[4419] = i[4419];
  assign o[4418] = i[4418];
  assign o[4417] = i[4417];
  assign o[4416] = i[4416];
  assign o[4415] = i[4415];
  assign o[4414] = i[4414];
  assign o[4413] = i[4413];
  assign o[4412] = i[4412];
  assign o[4411] = i[4411];
  assign o[4410] = i[4410];
  assign o[4409] = i[4409];
  assign o[4408] = i[4408];
  assign o[4407] = i[4407];
  assign o[4406] = i[4406];
  assign o[4405] = i[4405];
  assign o[4404] = i[4404];
  assign o[4403] = i[4403];
  assign o[4402] = i[4402];
  assign o[4401] = i[4401];
  assign o[4400] = i[4400];
  assign o[4399] = i[4399];
  assign o[4398] = i[4398];
  assign o[4397] = i[4397];
  assign o[4396] = i[4396];
  assign o[4395] = i[4395];
  assign o[4394] = i[4394];
  assign o[4393] = i[4393];
  assign o[4392] = i[4392];
  assign o[4391] = i[4391];
  assign o[4390] = i[4390];
  assign o[4389] = i[4389];
  assign o[4388] = i[4388];
  assign o[4387] = i[4387];
  assign o[4386] = i[4386];
  assign o[4385] = i[4385];
  assign o[4384] = i[4384];
  assign o[4383] = i[4383];
  assign o[4382] = i[4382];
  assign o[4381] = i[4381];
  assign o[4380] = i[4380];
  assign o[4379] = i[4379];
  assign o[4378] = i[4378];
  assign o[4377] = i[4377];
  assign o[4376] = i[4376];
  assign o[4375] = i[4375];
  assign o[4374] = i[4374];
  assign o[4373] = i[4373];
  assign o[4372] = i[4372];
  assign o[4371] = i[4371];
  assign o[4370] = i[4370];
  assign o[4369] = i[4369];
  assign o[4368] = i[4368];
  assign o[4367] = i[4367];
  assign o[4366] = i[4366];
  assign o[4365] = i[4365];
  assign o[4364] = i[4364];
  assign o[4363] = i[4363];
  assign o[4362] = i[4362];
  assign o[4361] = i[4361];
  assign o[4360] = i[4360];
  assign o[4359] = i[4359];
  assign o[4358] = i[4358];
  assign o[4357] = i[4357];
  assign o[4356] = i[4356];
  assign o[4355] = i[4355];
  assign o[4354] = i[4354];
  assign o[4353] = i[4353];
  assign o[4352] = i[4352];
  assign o[4351] = i[4351];
  assign o[4350] = i[4350];
  assign o[4349] = i[4349];
  assign o[4348] = i[4348];
  assign o[4347] = i[4347];
  assign o[4346] = i[4346];
  assign o[4345] = i[4345];
  assign o[4344] = i[4344];
  assign o[4343] = i[4343];
  assign o[4342] = i[4342];
  assign o[4341] = i[4341];
  assign o[4340] = i[4340];
  assign o[4339] = i[4339];
  assign o[4338] = i[4338];
  assign o[4337] = i[4337];
  assign o[4336] = i[4336];
  assign o[4335] = i[4335];
  assign o[4334] = i[4334];
  assign o[4333] = i[4333];
  assign o[4332] = i[4332];
  assign o[4331] = i[4331];
  assign o[4330] = i[4330];
  assign o[4329] = i[4329];
  assign o[4328] = i[4328];
  assign o[4327] = i[4327];
  assign o[4326] = i[4326];
  assign o[4325] = i[4325];
  assign o[4324] = i[4324];
  assign o[4323] = i[4323];
  assign o[4322] = i[4322];
  assign o[4321] = i[4321];
  assign o[4320] = i[4320];
  assign o[4319] = i[4319];
  assign o[4318] = i[4318];
  assign o[4317] = i[4317];
  assign o[4316] = i[4316];
  assign o[4315] = i[4315];
  assign o[4314] = i[4314];
  assign o[4313] = i[4313];
  assign o[4312] = i[4312];
  assign o[4311] = i[4311];
  assign o[4310] = i[4310];
  assign o[4309] = i[4309];
  assign o[4308] = i[4308];
  assign o[4307] = i[4307];
  assign o[4306] = i[4306];
  assign o[4305] = i[4305];
  assign o[4304] = i[4304];
  assign o[4303] = i[4303];
  assign o[4302] = i[4302];
  assign o[4301] = i[4301];
  assign o[4300] = i[4300];
  assign o[4299] = i[4299];
  assign o[4298] = i[4298];
  assign o[4297] = i[4297];
  assign o[4296] = i[4296];
  assign o[4295] = i[4295];
  assign o[4294] = i[4294];
  assign o[4293] = i[4293];
  assign o[4292] = i[4292];
  assign o[4291] = i[4291];
  assign o[4290] = i[4290];
  assign o[4289] = i[4289];
  assign o[4288] = i[4288];
  assign o[4287] = i[4287];
  assign o[4286] = i[4286];
  assign o[4285] = i[4285];
  assign o[4284] = i[4284];
  assign o[4283] = i[4283];
  assign o[4282] = i[4282];
  assign o[4281] = i[4281];
  assign o[4280] = i[4280];
  assign o[4279] = i[4279];
  assign o[4278] = i[4278];
  assign o[4277] = i[4277];
  assign o[4276] = i[4276];
  assign o[4275] = i[4275];
  assign o[4274] = i[4274];
  assign o[4273] = i[4273];
  assign o[4272] = i[4272];
  assign o[4271] = i[4271];
  assign o[4270] = i[4270];
  assign o[4269] = i[4269];
  assign o[4268] = i[4268];
  assign o[4267] = i[4267];
  assign o[4266] = i[4266];
  assign o[4265] = i[4265];
  assign o[4264] = i[4264];
  assign o[4263] = i[4263];
  assign o[4262] = i[4262];
  assign o[4261] = i[4261];
  assign o[4260] = i[4260];
  assign o[4259] = i[4259];
  assign o[4258] = i[4258];
  assign o[4257] = i[4257];
  assign o[4256] = i[4256];
  assign o[4255] = i[4255];
  assign o[4254] = i[4254];
  assign o[4253] = i[4253];
  assign o[4252] = i[4252];
  assign o[4251] = i[4251];
  assign o[4250] = i[4250];
  assign o[4249] = i[4249];
  assign o[4248] = i[4248];
  assign o[4247] = i[4247];
  assign o[4246] = i[4246];
  assign o[4245] = i[4245];
  assign o[4244] = i[4244];
  assign o[4243] = i[4243];
  assign o[4242] = i[4242];
  assign o[4241] = i[4241];
  assign o[4240] = i[4240];
  assign o[4239] = i[4239];
  assign o[4238] = i[4238];
  assign o[4237] = i[4237];
  assign o[4236] = i[4236];
  assign o[4235] = i[4235];
  assign o[4234] = i[4234];
  assign o[4233] = i[4233];
  assign o[4232] = i[4232];
  assign o[4231] = i[4231];
  assign o[4230] = i[4230];
  assign o[4229] = i[4229];
  assign o[4228] = i[4228];
  assign o[4227] = i[4227];
  assign o[4226] = i[4226];
  assign o[4225] = i[4225];
  assign o[4224] = i[4224];
  assign o[4223] = i[4223];
  assign o[4222] = i[4222];
  assign o[4221] = i[4221];
  assign o[4220] = i[4220];
  assign o[4219] = i[4219];
  assign o[4218] = i[4218];
  assign o[4217] = i[4217];
  assign o[4216] = i[4216];
  assign o[4215] = i[4215];
  assign o[4214] = i[4214];
  assign o[4213] = i[4213];
  assign o[4212] = i[4212];
  assign o[4211] = i[4211];
  assign o[4210] = i[4210];
  assign o[4209] = i[4209];
  assign o[4208] = i[4208];
  assign o[4207] = i[4207];
  assign o[4206] = i[4206];
  assign o[4205] = i[4205];
  assign o[4204] = i[4204];
  assign o[4203] = i[4203];
  assign o[4202] = i[4202];
  assign o[4201] = i[4201];
  assign o[4200] = i[4200];
  assign o[4199] = i[4199];
  assign o[4198] = i[4198];
  assign o[4197] = i[4197];
  assign o[4196] = i[4196];
  assign o[4195] = i[4195];
  assign o[4194] = i[4194];
  assign o[4193] = i[4193];
  assign o[4192] = i[4192];
  assign o[4191] = i[4191];
  assign o[4190] = i[4190];
  assign o[4189] = i[4189];
  assign o[4188] = i[4188];
  assign o[4187] = i[4187];
  assign o[4186] = i[4186];
  assign o[4185] = i[4185];
  assign o[4184] = i[4184];
  assign o[4183] = i[4183];
  assign o[4182] = i[4182];
  assign o[4181] = i[4181];
  assign o[4180] = i[4180];
  assign o[4179] = i[4179];
  assign o[4178] = i[4178];
  assign o[4177] = i[4177];
  assign o[4176] = i[4176];
  assign o[4175] = i[4175];
  assign o[4174] = i[4174];
  assign o[4173] = i[4173];
  assign o[4172] = i[4172];
  assign o[4171] = i[4171];
  assign o[4170] = i[4170];
  assign o[4169] = i[4169];
  assign o[4168] = i[4168];
  assign o[4167] = i[4167];
  assign o[4166] = i[4166];
  assign o[4165] = i[4165];
  assign o[4164] = i[4164];
  assign o[4163] = i[4163];
  assign o[4162] = i[4162];
  assign o[4161] = i[4161];
  assign o[4160] = i[4160];
  assign o[4159] = i[4159];
  assign o[4158] = i[4158];
  assign o[4157] = i[4157];
  assign o[4156] = i[4156];
  assign o[4155] = i[4155];
  assign o[4154] = i[4154];
  assign o[4153] = i[4153];
  assign o[4152] = i[4152];
  assign o[4151] = i[4151];
  assign o[4150] = i[4150];
  assign o[4149] = i[4149];
  assign o[4148] = i[4148];
  assign o[4147] = i[4147];
  assign o[4146] = i[4146];
  assign o[4145] = i[4145];
  assign o[4144] = i[4144];
  assign o[4143] = i[4143];
  assign o[4142] = i[4142];
  assign o[4141] = i[4141];
  assign o[4140] = i[4140];
  assign o[4139] = i[4139];
  assign o[4138] = i[4138];
  assign o[4137] = i[4137];
  assign o[4136] = i[4136];
  assign o[4135] = i[4135];
  assign o[4134] = i[4134];
  assign o[4133] = i[4133];
  assign o[4132] = i[4132];
  assign o[4131] = i[4131];
  assign o[4130] = i[4130];
  assign o[4129] = i[4129];
  assign o[4128] = i[4128];
  assign o[4127] = i[4127];
  assign o[4126] = i[4126];
  assign o[4125] = i[4125];
  assign o[4124] = i[4124];
  assign o[4123] = i[4123];
  assign o[4122] = i[4122];
  assign o[4121] = i[4121];
  assign o[4120] = i[4120];
  assign o[4119] = i[4119];
  assign o[4118] = i[4118];
  assign o[4117] = i[4117];
  assign o[4116] = i[4116];
  assign o[4115] = i[4115];
  assign o[4114] = i[4114];
  assign o[4113] = i[4113];
  assign o[4112] = i[4112];
  assign o[4111] = i[4111];
  assign o[4110] = i[4110];
  assign o[4109] = i[4109];
  assign o[4108] = i[4108];
  assign o[4107] = i[4107];
  assign o[4106] = i[4106];
  assign o[4105] = i[4105];
  assign o[4104] = i[4104];
  assign o[4103] = i[4103];
  assign o[4102] = i[4102];
  assign o[4101] = i[4101];
  assign o[4100] = i[4100];
  assign o[4099] = i[4099];
  assign o[4098] = i[4098];
  assign o[4097] = i[4097];
  assign o[4096] = i[4096];
  assign o[4095] = i[4095];
  assign o[4094] = i[4094];
  assign o[4093] = i[4093];
  assign o[4092] = i[4092];
  assign o[4091] = i[4091];
  assign o[4090] = i[4090];
  assign o[4089] = i[4089];
  assign o[4088] = i[4088];
  assign o[4087] = i[4087];
  assign o[4086] = i[4086];
  assign o[4085] = i[4085];
  assign o[4084] = i[4084];
  assign o[4083] = i[4083];
  assign o[4082] = i[4082];
  assign o[4081] = i[4081];
  assign o[4080] = i[4080];
  assign o[4079] = i[4079];
  assign o[4078] = i[4078];
  assign o[4077] = i[4077];
  assign o[4076] = i[4076];
  assign o[4075] = i[4075];
  assign o[4074] = i[4074];
  assign o[4073] = i[4073];
  assign o[4072] = i[4072];
  assign o[4071] = i[4071];
  assign o[4070] = i[4070];
  assign o[4069] = i[4069];
  assign o[4068] = i[4068];
  assign o[4067] = i[4067];
  assign o[4066] = i[4066];
  assign o[4065] = i[4065];
  assign o[4064] = i[4064];
  assign o[4063] = i[4063];
  assign o[4062] = i[4062];
  assign o[4061] = i[4061];
  assign o[4060] = i[4060];
  assign o[4059] = i[4059];
  assign o[4058] = i[4058];
  assign o[4057] = i[4057];
  assign o[4056] = i[4056];
  assign o[4055] = i[4055];
  assign o[4054] = i[4054];
  assign o[4053] = i[4053];
  assign o[4052] = i[4052];
  assign o[4051] = i[4051];
  assign o[4050] = i[4050];
  assign o[4049] = i[4049];
  assign o[4048] = i[4048];
  assign o[4047] = i[4047];
  assign o[4046] = i[4046];
  assign o[4045] = i[4045];
  assign o[4044] = i[4044];
  assign o[4043] = i[4043];
  assign o[4042] = i[4042];
  assign o[4041] = i[4041];
  assign o[4040] = i[4040];
  assign o[4039] = i[4039];
  assign o[4038] = i[4038];
  assign o[4037] = i[4037];
  assign o[4036] = i[4036];
  assign o[4035] = i[4035];
  assign o[4034] = i[4034];
  assign o[4033] = i[4033];
  assign o[4032] = i[4032];
  assign o[4031] = i[4031];
  assign o[4030] = i[4030];
  assign o[4029] = i[4029];
  assign o[4028] = i[4028];
  assign o[4027] = i[4027];
  assign o[4026] = i[4026];
  assign o[4025] = i[4025];
  assign o[4024] = i[4024];
  assign o[4023] = i[4023];
  assign o[4022] = i[4022];
  assign o[4021] = i[4021];
  assign o[4020] = i[4020];
  assign o[4019] = i[4019];
  assign o[4018] = i[4018];
  assign o[4017] = i[4017];
  assign o[4016] = i[4016];
  assign o[4015] = i[4015];
  assign o[4014] = i[4014];
  assign o[4013] = i[4013];
  assign o[4012] = i[4012];
  assign o[4011] = i[4011];
  assign o[4010] = i[4010];
  assign o[4009] = i[4009];
  assign o[4008] = i[4008];
  assign o[4007] = i[4007];
  assign o[4006] = i[4006];
  assign o[4005] = i[4005];
  assign o[4004] = i[4004];
  assign o[4003] = i[4003];
  assign o[4002] = i[4002];
  assign o[4001] = i[4001];
  assign o[4000] = i[4000];
  assign o[3999] = i[3999];
  assign o[3998] = i[3998];
  assign o[3997] = i[3997];
  assign o[3996] = i[3996];
  assign o[3995] = i[3995];
  assign o[3994] = i[3994];
  assign o[3993] = i[3993];
  assign o[3992] = i[3992];
  assign o[3991] = i[3991];
  assign o[3990] = i[3990];
  assign o[3989] = i[3989];
  assign o[3988] = i[3988];
  assign o[3987] = i[3987];
  assign o[3986] = i[3986];
  assign o[3985] = i[3985];
  assign o[3984] = i[3984];
  assign o[3983] = i[3983];
  assign o[3982] = i[3982];
  assign o[3981] = i[3981];
  assign o[3980] = i[3980];
  assign o[3979] = i[3979];
  assign o[3978] = i[3978];
  assign o[3977] = i[3977];
  assign o[3976] = i[3976];
  assign o[3975] = i[3975];
  assign o[3974] = i[3974];
  assign o[3973] = i[3973];
  assign o[3972] = i[3972];
  assign o[3971] = i[3971];
  assign o[3970] = i[3970];
  assign o[3969] = i[3969];
  assign o[3968] = i[3968];
  assign o[3967] = i[3967];
  assign o[3966] = i[3966];
  assign o[3965] = i[3965];
  assign o[3964] = i[3964];
  assign o[3963] = i[3963];
  assign o[3962] = i[3962];
  assign o[3961] = i[3961];
  assign o[3960] = i[3960];
  assign o[3959] = i[3959];
  assign o[3958] = i[3958];
  assign o[3957] = i[3957];
  assign o[3956] = i[3956];
  assign o[3955] = i[3955];
  assign o[3954] = i[3954];
  assign o[3953] = i[3953];
  assign o[3952] = i[3952];
  assign o[3951] = i[3951];
  assign o[3950] = i[3950];
  assign o[3949] = i[3949];
  assign o[3948] = i[3948];
  assign o[3947] = i[3947];
  assign o[3946] = i[3946];
  assign o[3945] = i[3945];
  assign o[3944] = i[3944];
  assign o[3943] = i[3943];
  assign o[3942] = i[3942];
  assign o[3941] = i[3941];
  assign o[3940] = i[3940];
  assign o[3939] = i[3939];
  assign o[3938] = i[3938];
  assign o[3937] = i[3937];
  assign o[3936] = i[3936];
  assign o[3935] = i[3935];
  assign o[3934] = i[3934];
  assign o[3933] = i[3933];
  assign o[3932] = i[3932];
  assign o[3931] = i[3931];
  assign o[3930] = i[3930];
  assign o[3929] = i[3929];
  assign o[3928] = i[3928];
  assign o[3927] = i[3927];
  assign o[3926] = i[3926];
  assign o[3925] = i[3925];
  assign o[3924] = i[3924];
  assign o[3923] = i[3923];
  assign o[3922] = i[3922];
  assign o[3921] = i[3921];
  assign o[3920] = i[3920];
  assign o[3919] = i[3919];
  assign o[3918] = i[3918];
  assign o[3917] = i[3917];
  assign o[3916] = i[3916];
  assign o[3915] = i[3915];
  assign o[3914] = i[3914];
  assign o[3913] = i[3913];
  assign o[3912] = i[3912];
  assign o[3911] = i[3911];
  assign o[3910] = i[3910];
  assign o[3909] = i[3909];
  assign o[3908] = i[3908];
  assign o[3907] = i[3907];
  assign o[3906] = i[3906];
  assign o[3905] = i[3905];
  assign o[3904] = i[3904];
  assign o[3903] = i[3903];
  assign o[3902] = i[3902];
  assign o[3901] = i[3901];
  assign o[3900] = i[3900];
  assign o[3899] = i[3899];
  assign o[3898] = i[3898];
  assign o[3897] = i[3897];
  assign o[3896] = i[3896];
  assign o[3895] = i[3895];
  assign o[3894] = i[3894];
  assign o[3893] = i[3893];
  assign o[3892] = i[3892];
  assign o[3891] = i[3891];
  assign o[3890] = i[3890];
  assign o[3889] = i[3889];
  assign o[3888] = i[3888];
  assign o[3887] = i[3887];
  assign o[3886] = i[3886];
  assign o[3885] = i[3885];
  assign o[3884] = i[3884];
  assign o[3883] = i[3883];
  assign o[3882] = i[3882];
  assign o[3881] = i[3881];
  assign o[3880] = i[3880];
  assign o[3879] = i[3879];
  assign o[3878] = i[3878];
  assign o[3877] = i[3877];
  assign o[3876] = i[3876];
  assign o[3875] = i[3875];
  assign o[3874] = i[3874];
  assign o[3873] = i[3873];
  assign o[3872] = i[3872];
  assign o[3871] = i[3871];
  assign o[3870] = i[3870];
  assign o[3869] = i[3869];
  assign o[3868] = i[3868];
  assign o[3867] = i[3867];
  assign o[3866] = i[3866];
  assign o[3865] = i[3865];
  assign o[3864] = i[3864];
  assign o[3863] = i[3863];
  assign o[3862] = i[3862];
  assign o[3861] = i[3861];
  assign o[3860] = i[3860];
  assign o[3859] = i[3859];
  assign o[3858] = i[3858];
  assign o[3857] = i[3857];
  assign o[3856] = i[3856];
  assign o[3855] = i[3855];
  assign o[3854] = i[3854];
  assign o[3853] = i[3853];
  assign o[3852] = i[3852];
  assign o[3851] = i[3851];
  assign o[3850] = i[3850];
  assign o[3849] = i[3849];
  assign o[3848] = i[3848];
  assign o[3847] = i[3847];
  assign o[3846] = i[3846];
  assign o[3845] = i[3845];
  assign o[3844] = i[3844];
  assign o[3843] = i[3843];
  assign o[3842] = i[3842];
  assign o[3841] = i[3841];
  assign o[3840] = i[3840];
  assign o[3839] = i[3839];
  assign o[3838] = i[3838];
  assign o[3837] = i[3837];
  assign o[3836] = i[3836];
  assign o[3835] = i[3835];
  assign o[3834] = i[3834];
  assign o[3833] = i[3833];
  assign o[3832] = i[3832];
  assign o[3831] = i[3831];
  assign o[3830] = i[3830];
  assign o[3829] = i[3829];
  assign o[3828] = i[3828];
  assign o[3827] = i[3827];
  assign o[3826] = i[3826];
  assign o[3825] = i[3825];
  assign o[3824] = i[3824];
  assign o[3823] = i[3823];
  assign o[3822] = i[3822];
  assign o[3821] = i[3821];
  assign o[3820] = i[3820];
  assign o[3819] = i[3819];
  assign o[3818] = i[3818];
  assign o[3817] = i[3817];
  assign o[3816] = i[3816];
  assign o[3815] = i[3815];
  assign o[3814] = i[3814];
  assign o[3813] = i[3813];
  assign o[3812] = i[3812];
  assign o[3811] = i[3811];
  assign o[3810] = i[3810];
  assign o[3809] = i[3809];
  assign o[3808] = i[3808];
  assign o[3807] = i[3807];
  assign o[3806] = i[3806];
  assign o[3805] = i[3805];
  assign o[3804] = i[3804];
  assign o[3803] = i[3803];
  assign o[3802] = i[3802];
  assign o[3801] = i[3801];
  assign o[3800] = i[3800];
  assign o[3799] = i[3799];
  assign o[3798] = i[3798];
  assign o[3797] = i[3797];
  assign o[3796] = i[3796];
  assign o[3795] = i[3795];
  assign o[3794] = i[3794];
  assign o[3793] = i[3793];
  assign o[3792] = i[3792];
  assign o[3791] = i[3791];
  assign o[3790] = i[3790];
  assign o[3789] = i[3789];
  assign o[3788] = i[3788];
  assign o[3787] = i[3787];
  assign o[3786] = i[3786];
  assign o[3785] = i[3785];
  assign o[3784] = i[3784];
  assign o[3783] = i[3783];
  assign o[3782] = i[3782];
  assign o[3781] = i[3781];
  assign o[3780] = i[3780];
  assign o[3779] = i[3779];
  assign o[3778] = i[3778];
  assign o[3777] = i[3777];
  assign o[3776] = i[3776];
  assign o[3775] = i[3775];
  assign o[3774] = i[3774];
  assign o[3773] = i[3773];
  assign o[3772] = i[3772];
  assign o[3771] = i[3771];
  assign o[3770] = i[3770];
  assign o[3769] = i[3769];
  assign o[3768] = i[3768];
  assign o[3767] = i[3767];
  assign o[3766] = i[3766];
  assign o[3765] = i[3765];
  assign o[3764] = i[3764];
  assign o[3763] = i[3763];
  assign o[3762] = i[3762];
  assign o[3761] = i[3761];
  assign o[3760] = i[3760];
  assign o[3759] = i[3759];
  assign o[3758] = i[3758];
  assign o[3757] = i[3757];
  assign o[3756] = i[3756];
  assign o[3755] = i[3755];
  assign o[3754] = i[3754];
  assign o[3753] = i[3753];
  assign o[3752] = i[3752];
  assign o[3751] = i[3751];
  assign o[3750] = i[3750];
  assign o[3749] = i[3749];
  assign o[3748] = i[3748];
  assign o[3747] = i[3747];
  assign o[3746] = i[3746];
  assign o[3745] = i[3745];
  assign o[3744] = i[3744];
  assign o[3743] = i[3743];
  assign o[3742] = i[3742];
  assign o[3741] = i[3741];
  assign o[3740] = i[3740];
  assign o[3739] = i[3739];
  assign o[3738] = i[3738];
  assign o[3737] = i[3737];
  assign o[3736] = i[3736];
  assign o[3735] = i[3735];
  assign o[3734] = i[3734];
  assign o[3733] = i[3733];
  assign o[3732] = i[3732];
  assign o[3731] = i[3731];
  assign o[3730] = i[3730];
  assign o[3729] = i[3729];
  assign o[3728] = i[3728];
  assign o[3727] = i[3727];
  assign o[3726] = i[3726];
  assign o[3725] = i[3725];
  assign o[3724] = i[3724];
  assign o[3723] = i[3723];
  assign o[3722] = i[3722];
  assign o[3721] = i[3721];
  assign o[3720] = i[3720];
  assign o[3719] = i[3719];
  assign o[3718] = i[3718];
  assign o[3717] = i[3717];
  assign o[3716] = i[3716];
  assign o[3715] = i[3715];
  assign o[3714] = i[3714];
  assign o[3713] = i[3713];
  assign o[3712] = i[3712];
  assign o[3711] = i[3711];
  assign o[3710] = i[3710];
  assign o[3709] = i[3709];
  assign o[3708] = i[3708];
  assign o[3707] = i[3707];
  assign o[3706] = i[3706];
  assign o[3705] = i[3705];
  assign o[3704] = i[3704];
  assign o[3703] = i[3703];
  assign o[3702] = i[3702];
  assign o[3701] = i[3701];
  assign o[3700] = i[3700];
  assign o[3699] = i[3699];
  assign o[3698] = i[3698];
  assign o[3697] = i[3697];
  assign o[3696] = i[3696];
  assign o[3695] = i[3695];
  assign o[3694] = i[3694];
  assign o[3693] = i[3693];
  assign o[3692] = i[3692];
  assign o[3691] = i[3691];
  assign o[3690] = i[3690];
  assign o[3689] = i[3689];
  assign o[3688] = i[3688];
  assign o[3687] = i[3687];
  assign o[3686] = i[3686];
  assign o[3685] = i[3685];
  assign o[3684] = i[3684];
  assign o[3683] = i[3683];
  assign o[3682] = i[3682];
  assign o[3681] = i[3681];
  assign o[3680] = i[3680];
  assign o[3679] = i[3679];
  assign o[3678] = i[3678];
  assign o[3677] = i[3677];
  assign o[3676] = i[3676];
  assign o[3675] = i[3675];
  assign o[3674] = i[3674];
  assign o[3673] = i[3673];
  assign o[3672] = i[3672];
  assign o[3671] = i[3671];
  assign o[3670] = i[3670];
  assign o[3669] = i[3669];
  assign o[3668] = i[3668];
  assign o[3667] = i[3667];
  assign o[3666] = i[3666];
  assign o[3665] = i[3665];
  assign o[3664] = i[3664];
  assign o[3663] = i[3663];
  assign o[3662] = i[3662];
  assign o[3661] = i[3661];
  assign o[3660] = i[3660];
  assign o[3659] = i[3659];
  assign o[3658] = i[3658];
  assign o[3657] = i[3657];
  assign o[3656] = i[3656];
  assign o[3655] = i[3655];
  assign o[3654] = i[3654];
  assign o[3653] = i[3653];
  assign o[3652] = i[3652];
  assign o[3651] = i[3651];
  assign o[3650] = i[3650];
  assign o[3649] = i[3649];
  assign o[3648] = i[3648];
  assign o[3647] = i[3647];
  assign o[3646] = i[3646];
  assign o[3645] = i[3645];
  assign o[3644] = i[3644];
  assign o[3643] = i[3643];
  assign o[3642] = i[3642];
  assign o[3641] = i[3641];
  assign o[3640] = i[3640];
  assign o[3639] = i[3639];
  assign o[3638] = i[3638];
  assign o[3637] = i[3637];
  assign o[3636] = i[3636];
  assign o[3635] = i[3635];
  assign o[3634] = i[3634];
  assign o[3633] = i[3633];
  assign o[3632] = i[3632];
  assign o[3631] = i[3631];
  assign o[3630] = i[3630];
  assign o[3629] = i[3629];
  assign o[3628] = i[3628];
  assign o[3627] = i[3627];
  assign o[3626] = i[3626];
  assign o[3625] = i[3625];
  assign o[3624] = i[3624];
  assign o[3623] = i[3623];
  assign o[3622] = i[3622];
  assign o[3621] = i[3621];
  assign o[3620] = i[3620];
  assign o[3619] = i[3619];
  assign o[3618] = i[3618];
  assign o[3617] = i[3617];
  assign o[3616] = i[3616];
  assign o[3615] = i[3615];
  assign o[3614] = i[3614];
  assign o[3613] = i[3613];
  assign o[3612] = i[3612];
  assign o[3611] = i[3611];
  assign o[3610] = i[3610];
  assign o[3609] = i[3609];
  assign o[3608] = i[3608];
  assign o[3607] = i[3607];
  assign o[3606] = i[3606];
  assign o[3605] = i[3605];
  assign o[3604] = i[3604];
  assign o[3603] = i[3603];
  assign o[3602] = i[3602];
  assign o[3601] = i[3601];
  assign o[3600] = i[3600];
  assign o[3599] = i[3599];
  assign o[3598] = i[3598];
  assign o[3597] = i[3597];
  assign o[3596] = i[3596];
  assign o[3595] = i[3595];
  assign o[3594] = i[3594];
  assign o[3593] = i[3593];
  assign o[3592] = i[3592];
  assign o[3591] = i[3591];
  assign o[3590] = i[3590];
  assign o[3589] = i[3589];
  assign o[3588] = i[3588];
  assign o[3587] = i[3587];
  assign o[3586] = i[3586];
  assign o[3585] = i[3585];
  assign o[3584] = i[3584];
  assign o[3583] = i[3583];
  assign o[3582] = i[3582];
  assign o[3581] = i[3581];
  assign o[3580] = i[3580];
  assign o[3579] = i[3579];
  assign o[3578] = i[3578];
  assign o[3577] = i[3577];
  assign o[3576] = i[3576];
  assign o[3575] = i[3575];
  assign o[3574] = i[3574];
  assign o[3573] = i[3573];
  assign o[3572] = i[3572];
  assign o[3571] = i[3571];
  assign o[3570] = i[3570];
  assign o[3569] = i[3569];
  assign o[3568] = i[3568];
  assign o[3567] = i[3567];
  assign o[3566] = i[3566];
  assign o[3565] = i[3565];
  assign o[3564] = i[3564];
  assign o[3563] = i[3563];
  assign o[3562] = i[3562];
  assign o[3561] = i[3561];
  assign o[3560] = i[3560];
  assign o[3559] = i[3559];
  assign o[3558] = i[3558];
  assign o[3557] = i[3557];
  assign o[3556] = i[3556];
  assign o[3555] = i[3555];
  assign o[3554] = i[3554];
  assign o[3553] = i[3553];
  assign o[3552] = i[3552];
  assign o[3551] = i[3551];
  assign o[3550] = i[3550];
  assign o[3549] = i[3549];
  assign o[3548] = i[3548];
  assign o[3547] = i[3547];
  assign o[3546] = i[3546];
  assign o[3545] = i[3545];
  assign o[3544] = i[3544];
  assign o[3543] = i[3543];
  assign o[3542] = i[3542];
  assign o[3541] = i[3541];
  assign o[3540] = i[3540];
  assign o[3539] = i[3539];
  assign o[3538] = i[3538];
  assign o[3537] = i[3537];
  assign o[3536] = i[3536];
  assign o[3535] = i[3535];
  assign o[3534] = i[3534];
  assign o[3533] = i[3533];
  assign o[3532] = i[3532];
  assign o[3531] = i[3531];
  assign o[3530] = i[3530];
  assign o[3529] = i[3529];
  assign o[3528] = i[3528];
  assign o[3527] = i[3527];
  assign o[3526] = i[3526];
  assign o[3525] = i[3525];
  assign o[3524] = i[3524];
  assign o[3523] = i[3523];
  assign o[3522] = i[3522];
  assign o[3521] = i[3521];
  assign o[3520] = i[3520];
  assign o[3519] = i[3519];
  assign o[3518] = i[3518];
  assign o[3517] = i[3517];
  assign o[3516] = i[3516];
  assign o[3515] = i[3515];
  assign o[3514] = i[3514];
  assign o[3513] = i[3513];
  assign o[3512] = i[3512];
  assign o[3511] = i[3511];
  assign o[3510] = i[3510];
  assign o[3509] = i[3509];
  assign o[3508] = i[3508];
  assign o[3507] = i[3507];
  assign o[3506] = i[3506];
  assign o[3505] = i[3505];
  assign o[3504] = i[3504];
  assign o[3503] = i[3503];
  assign o[3502] = i[3502];
  assign o[3501] = i[3501];
  assign o[3500] = i[3500];
  assign o[3499] = i[3499];
  assign o[3498] = i[3498];
  assign o[3497] = i[3497];
  assign o[3496] = i[3496];
  assign o[3495] = i[3495];
  assign o[3494] = i[3494];
  assign o[3493] = i[3493];
  assign o[3492] = i[3492];
  assign o[3491] = i[3491];
  assign o[3490] = i[3490];
  assign o[3489] = i[3489];
  assign o[3488] = i[3488];
  assign o[3487] = i[3487];
  assign o[3486] = i[3486];
  assign o[3485] = i[3485];
  assign o[3484] = i[3484];
  assign o[3483] = i[3483];
  assign o[3482] = i[3482];
  assign o[3481] = i[3481];
  assign o[3480] = i[3480];
  assign o[3479] = i[3479];
  assign o[3478] = i[3478];
  assign o[3477] = i[3477];
  assign o[3476] = i[3476];
  assign o[3475] = i[3475];
  assign o[3474] = i[3474];
  assign o[3473] = i[3473];
  assign o[3472] = i[3472];
  assign o[3471] = i[3471];
  assign o[3470] = i[3470];
  assign o[3469] = i[3469];
  assign o[3468] = i[3468];
  assign o[3467] = i[3467];
  assign o[3466] = i[3466];
  assign o[3465] = i[3465];
  assign o[3464] = i[3464];
  assign o[3463] = i[3463];
  assign o[3462] = i[3462];
  assign o[3461] = i[3461];
  assign o[3460] = i[3460];
  assign o[3459] = i[3459];
  assign o[3458] = i[3458];
  assign o[3457] = i[3457];
  assign o[3456] = i[3456];
  assign o[3455] = i[3455];
  assign o[3454] = i[3454];
  assign o[3453] = i[3453];
  assign o[3452] = i[3452];
  assign o[3451] = i[3451];
  assign o[3450] = i[3450];
  assign o[3449] = i[3449];
  assign o[3448] = i[3448];
  assign o[3447] = i[3447];
  assign o[3446] = i[3446];
  assign o[3445] = i[3445];
  assign o[3444] = i[3444];
  assign o[3443] = i[3443];
  assign o[3442] = i[3442];
  assign o[3441] = i[3441];
  assign o[3440] = i[3440];
  assign o[3439] = i[3439];
  assign o[3438] = i[3438];
  assign o[3437] = i[3437];
  assign o[3436] = i[3436];
  assign o[3435] = i[3435];
  assign o[3434] = i[3434];
  assign o[3433] = i[3433];
  assign o[3432] = i[3432];
  assign o[3431] = i[3431];
  assign o[3430] = i[3430];
  assign o[3429] = i[3429];
  assign o[3428] = i[3428];
  assign o[3427] = i[3427];
  assign o[3426] = i[3426];
  assign o[3425] = i[3425];
  assign o[3424] = i[3424];
  assign o[3423] = i[3423];
  assign o[3422] = i[3422];
  assign o[3421] = i[3421];
  assign o[3420] = i[3420];
  assign o[3419] = i[3419];
  assign o[3418] = i[3418];
  assign o[3417] = i[3417];
  assign o[3416] = i[3416];
  assign o[3415] = i[3415];
  assign o[3414] = i[3414];
  assign o[3413] = i[3413];
  assign o[3412] = i[3412];
  assign o[3411] = i[3411];
  assign o[3410] = i[3410];
  assign o[3409] = i[3409];
  assign o[3408] = i[3408];
  assign o[3407] = i[3407];
  assign o[3406] = i[3406];
  assign o[3405] = i[3405];
  assign o[3404] = i[3404];
  assign o[3403] = i[3403];
  assign o[3402] = i[3402];
  assign o[3401] = i[3401];
  assign o[3400] = i[3400];
  assign o[3399] = i[3399];
  assign o[3398] = i[3398];
  assign o[3397] = i[3397];
  assign o[3396] = i[3396];
  assign o[3395] = i[3395];
  assign o[3394] = i[3394];
  assign o[3393] = i[3393];
  assign o[3392] = i[3392];
  assign o[3391] = i[3391];
  assign o[3390] = i[3390];
  assign o[3389] = i[3389];
  assign o[3388] = i[3388];
  assign o[3387] = i[3387];
  assign o[3386] = i[3386];
  assign o[3385] = i[3385];
  assign o[3384] = i[3384];
  assign o[3383] = i[3383];
  assign o[3382] = i[3382];
  assign o[3381] = i[3381];
  assign o[3380] = i[3380];
  assign o[3379] = i[3379];
  assign o[3378] = i[3378];
  assign o[3377] = i[3377];
  assign o[3376] = i[3376];
  assign o[3375] = i[3375];
  assign o[3374] = i[3374];
  assign o[3373] = i[3373];
  assign o[3372] = i[3372];
  assign o[3371] = i[3371];
  assign o[3370] = i[3370];
  assign o[3369] = i[3369];
  assign o[3368] = i[3368];
  assign o[3367] = i[3367];
  assign o[3366] = i[3366];
  assign o[3365] = i[3365];
  assign o[3364] = i[3364];
  assign o[3363] = i[3363];
  assign o[3362] = i[3362];
  assign o[3361] = i[3361];
  assign o[3360] = i[3360];
  assign o[3359] = i[3359];
  assign o[3358] = i[3358];
  assign o[3357] = i[3357];
  assign o[3356] = i[3356];
  assign o[3355] = i[3355];
  assign o[3354] = i[3354];
  assign o[3353] = i[3353];
  assign o[3352] = i[3352];
  assign o[3351] = i[3351];
  assign o[3350] = i[3350];
  assign o[3349] = i[3349];
  assign o[3348] = i[3348];
  assign o[3347] = i[3347];
  assign o[3346] = i[3346];
  assign o[3345] = i[3345];
  assign o[3344] = i[3344];
  assign o[3343] = i[3343];
  assign o[3342] = i[3342];
  assign o[3341] = i[3341];
  assign o[3340] = i[3340];
  assign o[3339] = i[3339];
  assign o[3338] = i[3338];
  assign o[3337] = i[3337];
  assign o[3336] = i[3336];
  assign o[3335] = i[3335];
  assign o[3334] = i[3334];
  assign o[3333] = i[3333];
  assign o[3332] = i[3332];
  assign o[3331] = i[3331];
  assign o[3330] = i[3330];
  assign o[3329] = i[3329];
  assign o[3328] = i[3328];
  assign o[3327] = i[3327];
  assign o[3326] = i[3326];
  assign o[3325] = i[3325];
  assign o[3324] = i[3324];
  assign o[3323] = i[3323];
  assign o[3322] = i[3322];
  assign o[3321] = i[3321];
  assign o[3320] = i[3320];
  assign o[3319] = i[3319];
  assign o[3318] = i[3318];
  assign o[3317] = i[3317];
  assign o[3316] = i[3316];
  assign o[3315] = i[3315];
  assign o[3314] = i[3314];
  assign o[3313] = i[3313];
  assign o[3312] = i[3312];
  assign o[3311] = i[3311];
  assign o[3310] = i[3310];
  assign o[3309] = i[3309];
  assign o[3308] = i[3308];
  assign o[3307] = i[3307];
  assign o[3306] = i[3306];
  assign o[3305] = i[3305];
  assign o[3304] = i[3304];
  assign o[3303] = i[3303];
  assign o[3302] = i[3302];
  assign o[3301] = i[3301];
  assign o[3300] = i[3300];
  assign o[3299] = i[3299];
  assign o[3298] = i[3298];
  assign o[3297] = i[3297];
  assign o[3296] = i[3296];
  assign o[3295] = i[3295];
  assign o[3294] = i[3294];
  assign o[3293] = i[3293];
  assign o[3292] = i[3292];
  assign o[3291] = i[3291];
  assign o[3290] = i[3290];
  assign o[3289] = i[3289];
  assign o[3288] = i[3288];
  assign o[3287] = i[3287];
  assign o[3286] = i[3286];
  assign o[3285] = i[3285];
  assign o[3284] = i[3284];
  assign o[3283] = i[3283];
  assign o[3282] = i[3282];
  assign o[3281] = i[3281];
  assign o[3280] = i[3280];
  assign o[3279] = i[3279];
  assign o[3278] = i[3278];
  assign o[3277] = i[3277];
  assign o[3276] = i[3276];
  assign o[3275] = i[3275];
  assign o[3274] = i[3274];
  assign o[3273] = i[3273];
  assign o[3272] = i[3272];
  assign o[3271] = i[3271];
  assign o[3270] = i[3270];
  assign o[3269] = i[3269];
  assign o[3268] = i[3268];
  assign o[3267] = i[3267];
  assign o[3266] = i[3266];
  assign o[3265] = i[3265];
  assign o[3264] = i[3264];
  assign o[3263] = i[3263];
  assign o[3262] = i[3262];
  assign o[3261] = i[3261];
  assign o[3260] = i[3260];
  assign o[3259] = i[3259];
  assign o[3258] = i[3258];
  assign o[3257] = i[3257];
  assign o[3256] = i[3256];
  assign o[3255] = i[3255];
  assign o[3254] = i[3254];
  assign o[3253] = i[3253];
  assign o[3252] = i[3252];
  assign o[3251] = i[3251];
  assign o[3250] = i[3250];
  assign o[3249] = i[3249];
  assign o[3248] = i[3248];
  assign o[3247] = i[3247];
  assign o[3246] = i[3246];
  assign o[3245] = i[3245];
  assign o[3244] = i[3244];
  assign o[3243] = i[3243];
  assign o[3242] = i[3242];
  assign o[3241] = i[3241];
  assign o[3240] = i[3240];
  assign o[3239] = i[3239];
  assign o[3238] = i[3238];
  assign o[3237] = i[3237];
  assign o[3236] = i[3236];
  assign o[3235] = i[3235];
  assign o[3234] = i[3234];
  assign o[3233] = i[3233];
  assign o[3232] = i[3232];
  assign o[3231] = i[3231];
  assign o[3230] = i[3230];
  assign o[3229] = i[3229];
  assign o[3228] = i[3228];
  assign o[3227] = i[3227];
  assign o[3226] = i[3226];
  assign o[3225] = i[3225];
  assign o[3224] = i[3224];
  assign o[3223] = i[3223];
  assign o[3222] = i[3222];
  assign o[3221] = i[3221];
  assign o[3220] = i[3220];
  assign o[3219] = i[3219];
  assign o[3218] = i[3218];
  assign o[3217] = i[3217];
  assign o[3216] = i[3216];
  assign o[3215] = i[3215];
  assign o[3214] = i[3214];
  assign o[3213] = i[3213];
  assign o[3212] = i[3212];
  assign o[3211] = i[3211];
  assign o[3210] = i[3210];
  assign o[3209] = i[3209];
  assign o[3208] = i[3208];
  assign o[3207] = i[3207];
  assign o[3206] = i[3206];
  assign o[3205] = i[3205];
  assign o[3204] = i[3204];
  assign o[3203] = i[3203];
  assign o[3202] = i[3202];
  assign o[3201] = i[3201];
  assign o[3200] = i[3200];
  assign o[3199] = i[3199];
  assign o[3198] = i[3198];
  assign o[3197] = i[3197];
  assign o[3196] = i[3196];
  assign o[3195] = i[3195];
  assign o[3194] = i[3194];
  assign o[3193] = i[3193];
  assign o[3192] = i[3192];
  assign o[3191] = i[3191];
  assign o[3190] = i[3190];
  assign o[3189] = i[3189];
  assign o[3188] = i[3188];
  assign o[3187] = i[3187];
  assign o[3186] = i[3186];
  assign o[3185] = i[3185];
  assign o[3184] = i[3184];
  assign o[3183] = i[3183];
  assign o[3182] = i[3182];
  assign o[3181] = i[3181];
  assign o[3180] = i[3180];
  assign o[3179] = i[3179];
  assign o[3178] = i[3178];
  assign o[3177] = i[3177];
  assign o[3176] = i[3176];
  assign o[3175] = i[3175];
  assign o[3174] = i[3174];
  assign o[3173] = i[3173];
  assign o[3172] = i[3172];
  assign o[3171] = i[3171];
  assign o[3170] = i[3170];
  assign o[3169] = i[3169];
  assign o[3168] = i[3168];
  assign o[3167] = i[3167];
  assign o[3166] = i[3166];
  assign o[3165] = i[3165];
  assign o[3164] = i[3164];
  assign o[3163] = i[3163];
  assign o[3162] = i[3162];
  assign o[3161] = i[3161];
  assign o[3160] = i[3160];
  assign o[3159] = i[3159];
  assign o[3158] = i[3158];
  assign o[3157] = i[3157];
  assign o[3156] = i[3156];
  assign o[3155] = i[3155];
  assign o[3154] = i[3154];
  assign o[3153] = i[3153];
  assign o[3152] = i[3152];
  assign o[3151] = i[3151];
  assign o[3150] = i[3150];
  assign o[3149] = i[3149];
  assign o[3148] = i[3148];
  assign o[3147] = i[3147];
  assign o[3146] = i[3146];
  assign o[3145] = i[3145];
  assign o[3144] = i[3144];
  assign o[3143] = i[3143];
  assign o[3142] = i[3142];
  assign o[3141] = i[3141];
  assign o[3140] = i[3140];
  assign o[3139] = i[3139];
  assign o[3138] = i[3138];
  assign o[3137] = i[3137];
  assign o[3136] = i[3136];
  assign o[3135] = i[3135];
  assign o[3134] = i[3134];
  assign o[3133] = i[3133];
  assign o[3132] = i[3132];
  assign o[3131] = i[3131];
  assign o[3130] = i[3130];
  assign o[3129] = i[3129];
  assign o[3128] = i[3128];
  assign o[3127] = i[3127];
  assign o[3126] = i[3126];
  assign o[3125] = i[3125];
  assign o[3124] = i[3124];
  assign o[3123] = i[3123];
  assign o[3122] = i[3122];
  assign o[3121] = i[3121];
  assign o[3120] = i[3120];
  assign o[3119] = i[3119];
  assign o[3118] = i[3118];
  assign o[3117] = i[3117];
  assign o[3116] = i[3116];
  assign o[3115] = i[3115];
  assign o[3114] = i[3114];
  assign o[3113] = i[3113];
  assign o[3112] = i[3112];
  assign o[3111] = i[3111];
  assign o[3110] = i[3110];
  assign o[3109] = i[3109];
  assign o[3108] = i[3108];
  assign o[3107] = i[3107];
  assign o[3106] = i[3106];
  assign o[3105] = i[3105];
  assign o[3104] = i[3104];
  assign o[3103] = i[3103];
  assign o[3102] = i[3102];
  assign o[3101] = i[3101];
  assign o[3100] = i[3100];
  assign o[3099] = i[3099];
  assign o[3098] = i[3098];
  assign o[3097] = i[3097];
  assign o[3096] = i[3096];
  assign o[3095] = i[3095];
  assign o[3094] = i[3094];
  assign o[3093] = i[3093];
  assign o[3092] = i[3092];
  assign o[3091] = i[3091];
  assign o[3090] = i[3090];
  assign o[3089] = i[3089];
  assign o[3088] = i[3088];
  assign o[3087] = i[3087];
  assign o[3086] = i[3086];
  assign o[3085] = i[3085];
  assign o[3084] = i[3084];
  assign o[3083] = i[3083];
  assign o[3082] = i[3082];
  assign o[3081] = i[3081];
  assign o[3080] = i[3080];
  assign o[3079] = i[3079];
  assign o[3078] = i[3078];
  assign o[3077] = i[3077];
  assign o[3076] = i[3076];
  assign o[3075] = i[3075];
  assign o[3074] = i[3074];
  assign o[3073] = i[3073];
  assign o[3072] = i[3072];
  assign o[3071] = i[3071];
  assign o[3070] = i[3070];
  assign o[3069] = i[3069];
  assign o[3068] = i[3068];
  assign o[3067] = i[3067];
  assign o[3066] = i[3066];
  assign o[3065] = i[3065];
  assign o[3064] = i[3064];
  assign o[3063] = i[3063];
  assign o[3062] = i[3062];
  assign o[3061] = i[3061];
  assign o[3060] = i[3060];
  assign o[3059] = i[3059];
  assign o[3058] = i[3058];
  assign o[3057] = i[3057];
  assign o[3056] = i[3056];
  assign o[3055] = i[3055];
  assign o[3054] = i[3054];
  assign o[3053] = i[3053];
  assign o[3052] = i[3052];
  assign o[3051] = i[3051];
  assign o[3050] = i[3050];
  assign o[3049] = i[3049];
  assign o[3048] = i[3048];
  assign o[3047] = i[3047];
  assign o[3046] = i[3046];
  assign o[3045] = i[3045];
  assign o[3044] = i[3044];
  assign o[3043] = i[3043];
  assign o[3042] = i[3042];
  assign o[3041] = i[3041];
  assign o[3040] = i[3040];
  assign o[3039] = i[3039];
  assign o[3038] = i[3038];
  assign o[3037] = i[3037];
  assign o[3036] = i[3036];
  assign o[3035] = i[3035];
  assign o[3034] = i[3034];
  assign o[3033] = i[3033];
  assign o[3032] = i[3032];
  assign o[3031] = i[3031];
  assign o[3030] = i[3030];
  assign o[3029] = i[3029];
  assign o[3028] = i[3028];
  assign o[3027] = i[3027];
  assign o[3026] = i[3026];
  assign o[3025] = i[3025];
  assign o[3024] = i[3024];
  assign o[3023] = i[3023];
  assign o[3022] = i[3022];
  assign o[3021] = i[3021];
  assign o[3020] = i[3020];
  assign o[3019] = i[3019];
  assign o[3018] = i[3018];
  assign o[3017] = i[3017];
  assign o[3016] = i[3016];
  assign o[3015] = i[3015];
  assign o[3014] = i[3014];
  assign o[3013] = i[3013];
  assign o[3012] = i[3012];
  assign o[3011] = i[3011];
  assign o[3010] = i[3010];
  assign o[3009] = i[3009];
  assign o[3008] = i[3008];
  assign o[3007] = i[3007];
  assign o[3006] = i[3006];
  assign o[3005] = i[3005];
  assign o[3004] = i[3004];
  assign o[3003] = i[3003];
  assign o[3002] = i[3002];
  assign o[3001] = i[3001];
  assign o[3000] = i[3000];
  assign o[2999] = i[2999];
  assign o[2998] = i[2998];
  assign o[2997] = i[2997];
  assign o[2996] = i[2996];
  assign o[2995] = i[2995];
  assign o[2994] = i[2994];
  assign o[2993] = i[2993];
  assign o[2992] = i[2992];
  assign o[2991] = i[2991];
  assign o[2990] = i[2990];
  assign o[2989] = i[2989];
  assign o[2988] = i[2988];
  assign o[2987] = i[2987];
  assign o[2986] = i[2986];
  assign o[2985] = i[2985];
  assign o[2984] = i[2984];
  assign o[2983] = i[2983];
  assign o[2982] = i[2982];
  assign o[2981] = i[2981];
  assign o[2980] = i[2980];
  assign o[2979] = i[2979];
  assign o[2978] = i[2978];
  assign o[2977] = i[2977];
  assign o[2976] = i[2976];
  assign o[2975] = i[2975];
  assign o[2974] = i[2974];
  assign o[2973] = i[2973];
  assign o[2972] = i[2972];
  assign o[2971] = i[2971];
  assign o[2970] = i[2970];
  assign o[2969] = i[2969];
  assign o[2968] = i[2968];
  assign o[2967] = i[2967];
  assign o[2966] = i[2966];
  assign o[2965] = i[2965];
  assign o[2964] = i[2964];
  assign o[2963] = i[2963];
  assign o[2962] = i[2962];
  assign o[2961] = i[2961];
  assign o[2960] = i[2960];
  assign o[2959] = i[2959];
  assign o[2958] = i[2958];
  assign o[2957] = i[2957];
  assign o[2956] = i[2956];
  assign o[2955] = i[2955];
  assign o[2954] = i[2954];
  assign o[2953] = i[2953];
  assign o[2952] = i[2952];
  assign o[2951] = i[2951];
  assign o[2950] = i[2950];
  assign o[2949] = i[2949];
  assign o[2948] = i[2948];
  assign o[2947] = i[2947];
  assign o[2946] = i[2946];
  assign o[2945] = i[2945];
  assign o[2944] = i[2944];
  assign o[2943] = i[2943];
  assign o[2942] = i[2942];
  assign o[2941] = i[2941];
  assign o[2940] = i[2940];
  assign o[2939] = i[2939];
  assign o[2938] = i[2938];
  assign o[2937] = i[2937];
  assign o[2936] = i[2936];
  assign o[2935] = i[2935];
  assign o[2934] = i[2934];
  assign o[2933] = i[2933];
  assign o[2932] = i[2932];
  assign o[2931] = i[2931];
  assign o[2930] = i[2930];
  assign o[2929] = i[2929];
  assign o[2928] = i[2928];
  assign o[2927] = i[2927];
  assign o[2926] = i[2926];
  assign o[2925] = i[2925];
  assign o[2924] = i[2924];
  assign o[2923] = i[2923];
  assign o[2922] = i[2922];
  assign o[2921] = i[2921];
  assign o[2920] = i[2920];
  assign o[2919] = i[2919];
  assign o[2918] = i[2918];
  assign o[2917] = i[2917];
  assign o[2916] = i[2916];
  assign o[2915] = i[2915];
  assign o[2914] = i[2914];
  assign o[2913] = i[2913];
  assign o[2912] = i[2912];
  assign o[2911] = i[2911];
  assign o[2910] = i[2910];
  assign o[2909] = i[2909];
  assign o[2908] = i[2908];
  assign o[2907] = i[2907];
  assign o[2906] = i[2906];
  assign o[2905] = i[2905];
  assign o[2904] = i[2904];
  assign o[2903] = i[2903];
  assign o[2902] = i[2902];
  assign o[2901] = i[2901];
  assign o[2900] = i[2900];
  assign o[2899] = i[2899];
  assign o[2898] = i[2898];
  assign o[2897] = i[2897];
  assign o[2896] = i[2896];
  assign o[2895] = i[2895];
  assign o[2894] = i[2894];
  assign o[2893] = i[2893];
  assign o[2892] = i[2892];
  assign o[2891] = i[2891];
  assign o[2890] = i[2890];
  assign o[2889] = i[2889];
  assign o[2888] = i[2888];
  assign o[2887] = i[2887];
  assign o[2886] = i[2886];
  assign o[2885] = i[2885];
  assign o[2884] = i[2884];
  assign o[2883] = i[2883];
  assign o[2882] = i[2882];
  assign o[2881] = i[2881];
  assign o[2880] = i[2880];
  assign o[2879] = i[2879];
  assign o[2878] = i[2878];
  assign o[2877] = i[2877];
  assign o[2876] = i[2876];
  assign o[2875] = i[2875];
  assign o[2874] = i[2874];
  assign o[2873] = i[2873];
  assign o[2872] = i[2872];
  assign o[2871] = i[2871];
  assign o[2870] = i[2870];
  assign o[2869] = i[2869];
  assign o[2868] = i[2868];
  assign o[2867] = i[2867];
  assign o[2866] = i[2866];
  assign o[2865] = i[2865];
  assign o[2864] = i[2864];
  assign o[2863] = i[2863];
  assign o[2862] = i[2862];
  assign o[2861] = i[2861];
  assign o[2860] = i[2860];
  assign o[2859] = i[2859];
  assign o[2858] = i[2858];
  assign o[2857] = i[2857];
  assign o[2856] = i[2856];
  assign o[2855] = i[2855];
  assign o[2854] = i[2854];
  assign o[2853] = i[2853];
  assign o[2852] = i[2852];
  assign o[2851] = i[2851];
  assign o[2850] = i[2850];
  assign o[2849] = i[2849];
  assign o[2848] = i[2848];
  assign o[2847] = i[2847];
  assign o[2846] = i[2846];
  assign o[2845] = i[2845];
  assign o[2844] = i[2844];
  assign o[2843] = i[2843];
  assign o[2842] = i[2842];
  assign o[2841] = i[2841];
  assign o[2840] = i[2840];
  assign o[2839] = i[2839];
  assign o[2838] = i[2838];
  assign o[2837] = i[2837];
  assign o[2836] = i[2836];
  assign o[2835] = i[2835];
  assign o[2834] = i[2834];
  assign o[2833] = i[2833];
  assign o[2832] = i[2832];
  assign o[2831] = i[2831];
  assign o[2830] = i[2830];
  assign o[2829] = i[2829];
  assign o[2828] = i[2828];
  assign o[2827] = i[2827];
  assign o[2826] = i[2826];
  assign o[2825] = i[2825];
  assign o[2824] = i[2824];
  assign o[2823] = i[2823];
  assign o[2822] = i[2822];
  assign o[2821] = i[2821];
  assign o[2820] = i[2820];
  assign o[2819] = i[2819];
  assign o[2818] = i[2818];
  assign o[2817] = i[2817];
  assign o[2816] = i[2816];
  assign o[2815] = i[2815];
  assign o[2814] = i[2814];
  assign o[2813] = i[2813];
  assign o[2812] = i[2812];
  assign o[2811] = i[2811];
  assign o[2810] = i[2810];
  assign o[2809] = i[2809];
  assign o[2808] = i[2808];
  assign o[2807] = i[2807];
  assign o[2806] = i[2806];
  assign o[2805] = i[2805];
  assign o[2804] = i[2804];
  assign o[2803] = i[2803];
  assign o[2802] = i[2802];
  assign o[2801] = i[2801];
  assign o[2800] = i[2800];
  assign o[2799] = i[2799];
  assign o[2798] = i[2798];
  assign o[2797] = i[2797];
  assign o[2796] = i[2796];
  assign o[2795] = i[2795];
  assign o[2794] = i[2794];
  assign o[2793] = i[2793];
  assign o[2792] = i[2792];
  assign o[2791] = i[2791];
  assign o[2790] = i[2790];
  assign o[2789] = i[2789];
  assign o[2788] = i[2788];
  assign o[2787] = i[2787];
  assign o[2786] = i[2786];
  assign o[2785] = i[2785];
  assign o[2784] = i[2784];
  assign o[2783] = i[2783];
  assign o[2782] = i[2782];
  assign o[2781] = i[2781];
  assign o[2780] = i[2780];
  assign o[2779] = i[2779];
  assign o[2778] = i[2778];
  assign o[2777] = i[2777];
  assign o[2776] = i[2776];
  assign o[2775] = i[2775];
  assign o[2774] = i[2774];
  assign o[2773] = i[2773];
  assign o[2772] = i[2772];
  assign o[2771] = i[2771];
  assign o[2770] = i[2770];
  assign o[2769] = i[2769];
  assign o[2768] = i[2768];
  assign o[2767] = i[2767];
  assign o[2766] = i[2766];
  assign o[2765] = i[2765];
  assign o[2764] = i[2764];
  assign o[2763] = i[2763];
  assign o[2762] = i[2762];
  assign o[2761] = i[2761];
  assign o[2760] = i[2760];
  assign o[2759] = i[2759];
  assign o[2758] = i[2758];
  assign o[2757] = i[2757];
  assign o[2756] = i[2756];
  assign o[2755] = i[2755];
  assign o[2754] = i[2754];
  assign o[2753] = i[2753];
  assign o[2752] = i[2752];
  assign o[2751] = i[2751];
  assign o[2750] = i[2750];
  assign o[2749] = i[2749];
  assign o[2748] = i[2748];
  assign o[2747] = i[2747];
  assign o[2746] = i[2746];
  assign o[2745] = i[2745];
  assign o[2744] = i[2744];
  assign o[2743] = i[2743];
  assign o[2742] = i[2742];
  assign o[2741] = i[2741];
  assign o[2740] = i[2740];
  assign o[2739] = i[2739];
  assign o[2738] = i[2738];
  assign o[2737] = i[2737];
  assign o[2736] = i[2736];
  assign o[2735] = i[2735];
  assign o[2734] = i[2734];
  assign o[2733] = i[2733];
  assign o[2732] = i[2732];
  assign o[2731] = i[2731];
  assign o[2730] = i[2730];
  assign o[2729] = i[2729];
  assign o[2728] = i[2728];
  assign o[2727] = i[2727];
  assign o[2726] = i[2726];
  assign o[2725] = i[2725];
  assign o[2724] = i[2724];
  assign o[2723] = i[2723];
  assign o[2722] = i[2722];
  assign o[2721] = i[2721];
  assign o[2720] = i[2720];
  assign o[2719] = i[2719];
  assign o[2718] = i[2718];
  assign o[2717] = i[2717];
  assign o[2716] = i[2716];
  assign o[2715] = i[2715];
  assign o[2714] = i[2714];
  assign o[2713] = i[2713];
  assign o[2712] = i[2712];
  assign o[2711] = i[2711];
  assign o[2710] = i[2710];
  assign o[2709] = i[2709];
  assign o[2708] = i[2708];
  assign o[2707] = i[2707];
  assign o[2706] = i[2706];
  assign o[2705] = i[2705];
  assign o[2704] = i[2704];
  assign o[2703] = i[2703];
  assign o[2702] = i[2702];
  assign o[2701] = i[2701];
  assign o[2700] = i[2700];
  assign o[2699] = i[2699];
  assign o[2698] = i[2698];
  assign o[2697] = i[2697];
  assign o[2696] = i[2696];
  assign o[2695] = i[2695];
  assign o[2694] = i[2694];
  assign o[2693] = i[2693];
  assign o[2692] = i[2692];
  assign o[2691] = i[2691];
  assign o[2690] = i[2690];
  assign o[2689] = i[2689];
  assign o[2688] = i[2688];
  assign o[2687] = i[2687];
  assign o[2686] = i[2686];
  assign o[2685] = i[2685];
  assign o[2684] = i[2684];
  assign o[2683] = i[2683];
  assign o[2682] = i[2682];
  assign o[2681] = i[2681];
  assign o[2680] = i[2680];
  assign o[2679] = i[2679];
  assign o[2678] = i[2678];
  assign o[2677] = i[2677];
  assign o[2676] = i[2676];
  assign o[2675] = i[2675];
  assign o[2674] = i[2674];
  assign o[2673] = i[2673];
  assign o[2672] = i[2672];
  assign o[2671] = i[2671];
  assign o[2670] = i[2670];
  assign o[2669] = i[2669];
  assign o[2668] = i[2668];
  assign o[2667] = i[2667];
  assign o[2666] = i[2666];
  assign o[2665] = i[2665];
  assign o[2664] = i[2664];
  assign o[2663] = i[2663];
  assign o[2662] = i[2662];
  assign o[2661] = i[2661];
  assign o[2660] = i[2660];
  assign o[2659] = i[2659];
  assign o[2658] = i[2658];
  assign o[2657] = i[2657];
  assign o[2656] = i[2656];
  assign o[2655] = i[2655];
  assign o[2654] = i[2654];
  assign o[2653] = i[2653];
  assign o[2652] = i[2652];
  assign o[2651] = i[2651];
  assign o[2650] = i[2650];
  assign o[2649] = i[2649];
  assign o[2648] = i[2648];
  assign o[2647] = i[2647];
  assign o[2646] = i[2646];
  assign o[2645] = i[2645];
  assign o[2644] = i[2644];
  assign o[2643] = i[2643];
  assign o[2642] = i[2642];
  assign o[2641] = i[2641];
  assign o[2640] = i[2640];
  assign o[2639] = i[2639];
  assign o[2638] = i[2638];
  assign o[2637] = i[2637];
  assign o[2636] = i[2636];
  assign o[2635] = i[2635];
  assign o[2634] = i[2634];
  assign o[2633] = i[2633];
  assign o[2632] = i[2632];
  assign o[2631] = i[2631];
  assign o[2630] = i[2630];
  assign o[2629] = i[2629];
  assign o[2628] = i[2628];
  assign o[2627] = i[2627];
  assign o[2626] = i[2626];
  assign o[2625] = i[2625];
  assign o[2624] = i[2624];
  assign o[2623] = i[2623];
  assign o[2622] = i[2622];
  assign o[2621] = i[2621];
  assign o[2620] = i[2620];
  assign o[2619] = i[2619];
  assign o[2618] = i[2618];
  assign o[2617] = i[2617];
  assign o[2616] = i[2616];
  assign o[2615] = i[2615];
  assign o[2614] = i[2614];
  assign o[2613] = i[2613];
  assign o[2612] = i[2612];
  assign o[2611] = i[2611];
  assign o[2610] = i[2610];
  assign o[2609] = i[2609];
  assign o[2608] = i[2608];
  assign o[2607] = i[2607];
  assign o[2606] = i[2606];
  assign o[2605] = i[2605];
  assign o[2604] = i[2604];
  assign o[2603] = i[2603];
  assign o[2602] = i[2602];
  assign o[2601] = i[2601];
  assign o[2600] = i[2600];
  assign o[2599] = i[2599];
  assign o[2598] = i[2598];
  assign o[2597] = i[2597];
  assign o[2596] = i[2596];
  assign o[2595] = i[2595];
  assign o[2594] = i[2594];
  assign o[2593] = i[2593];
  assign o[2592] = i[2592];
  assign o[2591] = i[2591];
  assign o[2590] = i[2590];
  assign o[2589] = i[2589];
  assign o[2588] = i[2588];
  assign o[2587] = i[2587];
  assign o[2586] = i[2586];
  assign o[2585] = i[2585];
  assign o[2584] = i[2584];
  assign o[2583] = i[2583];
  assign o[2582] = i[2582];
  assign o[2581] = i[2581];
  assign o[2580] = i[2580];
  assign o[2579] = i[2579];
  assign o[2578] = i[2578];
  assign o[2577] = i[2577];
  assign o[2576] = i[2576];
  assign o[2575] = i[2575];
  assign o[2574] = i[2574];
  assign o[2573] = i[2573];
  assign o[2572] = i[2572];
  assign o[2571] = i[2571];
  assign o[2570] = i[2570];
  assign o[2569] = i[2569];
  assign o[2568] = i[2568];
  assign o[2567] = i[2567];
  assign o[2566] = i[2566];
  assign o[2565] = i[2565];
  assign o[2564] = i[2564];
  assign o[2563] = i[2563];
  assign o[2562] = i[2562];
  assign o[2561] = i[2561];
  assign o[2560] = i[2560];
  assign o[2559] = i[2559];
  assign o[2558] = i[2558];
  assign o[2557] = i[2557];
  assign o[2556] = i[2556];
  assign o[2555] = i[2555];
  assign o[2554] = i[2554];
  assign o[2553] = i[2553];
  assign o[2552] = i[2552];
  assign o[2551] = i[2551];
  assign o[2550] = i[2550];
  assign o[2549] = i[2549];
  assign o[2548] = i[2548];
  assign o[2547] = i[2547];
  assign o[2546] = i[2546];
  assign o[2545] = i[2545];
  assign o[2544] = i[2544];
  assign o[2543] = i[2543];
  assign o[2542] = i[2542];
  assign o[2541] = i[2541];
  assign o[2540] = i[2540];
  assign o[2539] = i[2539];
  assign o[2538] = i[2538];
  assign o[2537] = i[2537];
  assign o[2536] = i[2536];
  assign o[2535] = i[2535];
  assign o[2534] = i[2534];
  assign o[2533] = i[2533];
  assign o[2532] = i[2532];
  assign o[2531] = i[2531];
  assign o[2530] = i[2530];
  assign o[2529] = i[2529];
  assign o[2528] = i[2528];
  assign o[2527] = i[2527];
  assign o[2526] = i[2526];
  assign o[2525] = i[2525];
  assign o[2524] = i[2524];
  assign o[2523] = i[2523];
  assign o[2522] = i[2522];
  assign o[2521] = i[2521];
  assign o[2520] = i[2520];
  assign o[2519] = i[2519];
  assign o[2518] = i[2518];
  assign o[2517] = i[2517];
  assign o[2516] = i[2516];
  assign o[2515] = i[2515];
  assign o[2514] = i[2514];
  assign o[2513] = i[2513];
  assign o[2512] = i[2512];
  assign o[2511] = i[2511];
  assign o[2510] = i[2510];
  assign o[2509] = i[2509];
  assign o[2508] = i[2508];
  assign o[2507] = i[2507];
  assign o[2506] = i[2506];
  assign o[2505] = i[2505];
  assign o[2504] = i[2504];
  assign o[2503] = i[2503];
  assign o[2502] = i[2502];
  assign o[2501] = i[2501];
  assign o[2500] = i[2500];
  assign o[2499] = i[2499];
  assign o[2498] = i[2498];
  assign o[2497] = i[2497];
  assign o[2496] = i[2496];
  assign o[2495] = i[2495];
  assign o[2494] = i[2494];
  assign o[2493] = i[2493];
  assign o[2492] = i[2492];
  assign o[2491] = i[2491];
  assign o[2490] = i[2490];
  assign o[2489] = i[2489];
  assign o[2488] = i[2488];
  assign o[2487] = i[2487];
  assign o[2486] = i[2486];
  assign o[2485] = i[2485];
  assign o[2484] = i[2484];
  assign o[2483] = i[2483];
  assign o[2482] = i[2482];
  assign o[2481] = i[2481];
  assign o[2480] = i[2480];
  assign o[2479] = i[2479];
  assign o[2478] = i[2478];
  assign o[2477] = i[2477];
  assign o[2476] = i[2476];
  assign o[2475] = i[2475];
  assign o[2474] = i[2474];
  assign o[2473] = i[2473];
  assign o[2472] = i[2472];
  assign o[2471] = i[2471];
  assign o[2470] = i[2470];
  assign o[2469] = i[2469];
  assign o[2468] = i[2468];
  assign o[2467] = i[2467];
  assign o[2466] = i[2466];
  assign o[2465] = i[2465];
  assign o[2464] = i[2464];
  assign o[2463] = i[2463];
  assign o[2462] = i[2462];
  assign o[2461] = i[2461];
  assign o[2460] = i[2460];
  assign o[2459] = i[2459];
  assign o[2458] = i[2458];
  assign o[2457] = i[2457];
  assign o[2456] = i[2456];
  assign o[2455] = i[2455];
  assign o[2454] = i[2454];
  assign o[2453] = i[2453];
  assign o[2452] = i[2452];
  assign o[2451] = i[2451];
  assign o[2450] = i[2450];
  assign o[2449] = i[2449];
  assign o[2448] = i[2448];
  assign o[2447] = i[2447];
  assign o[2446] = i[2446];
  assign o[2445] = i[2445];
  assign o[2444] = i[2444];
  assign o[2443] = i[2443];
  assign o[2442] = i[2442];
  assign o[2441] = i[2441];
  assign o[2440] = i[2440];
  assign o[2439] = i[2439];
  assign o[2438] = i[2438];
  assign o[2437] = i[2437];
  assign o[2436] = i[2436];
  assign o[2435] = i[2435];
  assign o[2434] = i[2434];
  assign o[2433] = i[2433];
  assign o[2432] = i[2432];
  assign o[2431] = i[2431];
  assign o[2430] = i[2430];
  assign o[2429] = i[2429];
  assign o[2428] = i[2428];
  assign o[2427] = i[2427];
  assign o[2426] = i[2426];
  assign o[2425] = i[2425];
  assign o[2424] = i[2424];
  assign o[2423] = i[2423];
  assign o[2422] = i[2422];
  assign o[2421] = i[2421];
  assign o[2420] = i[2420];
  assign o[2419] = i[2419];
  assign o[2418] = i[2418];
  assign o[2417] = i[2417];
  assign o[2416] = i[2416];
  assign o[2415] = i[2415];
  assign o[2414] = i[2414];
  assign o[2413] = i[2413];
  assign o[2412] = i[2412];
  assign o[2411] = i[2411];
  assign o[2410] = i[2410];
  assign o[2409] = i[2409];
  assign o[2408] = i[2408];
  assign o[2407] = i[2407];
  assign o[2406] = i[2406];
  assign o[2405] = i[2405];
  assign o[2404] = i[2404];
  assign o[2403] = i[2403];
  assign o[2402] = i[2402];
  assign o[2401] = i[2401];
  assign o[2400] = i[2400];
  assign o[2399] = i[2399];
  assign o[2398] = i[2398];
  assign o[2397] = i[2397];
  assign o[2396] = i[2396];
  assign o[2395] = i[2395];
  assign o[2394] = i[2394];
  assign o[2393] = i[2393];
  assign o[2392] = i[2392];
  assign o[2391] = i[2391];
  assign o[2390] = i[2390];
  assign o[2389] = i[2389];
  assign o[2388] = i[2388];
  assign o[2387] = i[2387];
  assign o[2386] = i[2386];
  assign o[2385] = i[2385];
  assign o[2384] = i[2384];
  assign o[2383] = i[2383];
  assign o[2382] = i[2382];
  assign o[2381] = i[2381];
  assign o[2380] = i[2380];
  assign o[2379] = i[2379];
  assign o[2378] = i[2378];
  assign o[2377] = i[2377];
  assign o[2376] = i[2376];
  assign o[2375] = i[2375];
  assign o[2374] = i[2374];
  assign o[2373] = i[2373];
  assign o[2372] = i[2372];
  assign o[2371] = i[2371];
  assign o[2370] = i[2370];
  assign o[2369] = i[2369];
  assign o[2368] = i[2368];
  assign o[2367] = i[2367];
  assign o[2366] = i[2366];
  assign o[2365] = i[2365];
  assign o[2364] = i[2364];
  assign o[2363] = i[2363];
  assign o[2362] = i[2362];
  assign o[2361] = i[2361];
  assign o[2360] = i[2360];
  assign o[2359] = i[2359];
  assign o[2358] = i[2358];
  assign o[2357] = i[2357];
  assign o[2356] = i[2356];
  assign o[2355] = i[2355];
  assign o[2354] = i[2354];
  assign o[2353] = i[2353];
  assign o[2352] = i[2352];
  assign o[2351] = i[2351];
  assign o[2350] = i[2350];
  assign o[2349] = i[2349];
  assign o[2348] = i[2348];
  assign o[2347] = i[2347];
  assign o[2346] = i[2346];
  assign o[2345] = i[2345];
  assign o[2344] = i[2344];
  assign o[2343] = i[2343];
  assign o[2342] = i[2342];
  assign o[2341] = i[2341];
  assign o[2340] = i[2340];
  assign o[2339] = i[2339];
  assign o[2338] = i[2338];
  assign o[2337] = i[2337];
  assign o[2336] = i[2336];
  assign o[2335] = i[2335];
  assign o[2334] = i[2334];
  assign o[2333] = i[2333];
  assign o[2332] = i[2332];
  assign o[2331] = i[2331];
  assign o[2330] = i[2330];
  assign o[2329] = i[2329];
  assign o[2328] = i[2328];
  assign o[2327] = i[2327];
  assign o[2326] = i[2326];
  assign o[2325] = i[2325];
  assign o[2324] = i[2324];
  assign o[2323] = i[2323];
  assign o[2322] = i[2322];
  assign o[2321] = i[2321];
  assign o[2320] = i[2320];
  assign o[2319] = i[2319];
  assign o[2318] = i[2318];
  assign o[2317] = i[2317];
  assign o[2316] = i[2316];
  assign o[2315] = i[2315];
  assign o[2314] = i[2314];
  assign o[2313] = i[2313];
  assign o[2312] = i[2312];
  assign o[2311] = i[2311];
  assign o[2310] = i[2310];
  assign o[2309] = i[2309];
  assign o[2308] = i[2308];
  assign o[2307] = i[2307];
  assign o[2306] = i[2306];
  assign o[2305] = i[2305];
  assign o[2304] = i[2304];
  assign o[2303] = i[2303];
  assign o[2302] = i[2302];
  assign o[2301] = i[2301];
  assign o[2300] = i[2300];
  assign o[2299] = i[2299];
  assign o[2298] = i[2298];
  assign o[2297] = i[2297];
  assign o[2296] = i[2296];
  assign o[2295] = i[2295];
  assign o[2294] = i[2294];
  assign o[2293] = i[2293];
  assign o[2292] = i[2292];
  assign o[2291] = i[2291];
  assign o[2290] = i[2290];
  assign o[2289] = i[2289];
  assign o[2288] = i[2288];
  assign o[2287] = i[2287];
  assign o[2286] = i[2286];
  assign o[2285] = i[2285];
  assign o[2284] = i[2284];
  assign o[2283] = i[2283];
  assign o[2282] = i[2282];
  assign o[2281] = i[2281];
  assign o[2280] = i[2280];
  assign o[2279] = i[2279];
  assign o[2278] = i[2278];
  assign o[2277] = i[2277];
  assign o[2276] = i[2276];
  assign o[2275] = i[2275];
  assign o[2274] = i[2274];
  assign o[2273] = i[2273];
  assign o[2272] = i[2272];
  assign o[2271] = i[2271];
  assign o[2270] = i[2270];
  assign o[2269] = i[2269];
  assign o[2268] = i[2268];
  assign o[2267] = i[2267];
  assign o[2266] = i[2266];
  assign o[2265] = i[2265];
  assign o[2264] = i[2264];
  assign o[2263] = i[2263];
  assign o[2262] = i[2262];
  assign o[2261] = i[2261];
  assign o[2260] = i[2260];
  assign o[2259] = i[2259];
  assign o[2258] = i[2258];
  assign o[2257] = i[2257];
  assign o[2256] = i[2256];
  assign o[2255] = i[2255];
  assign o[2254] = i[2254];
  assign o[2253] = i[2253];
  assign o[2252] = i[2252];
  assign o[2251] = i[2251];
  assign o[2250] = i[2250];
  assign o[2249] = i[2249];
  assign o[2248] = i[2248];
  assign o[2247] = i[2247];
  assign o[2246] = i[2246];
  assign o[2245] = i[2245];
  assign o[2244] = i[2244];
  assign o[2243] = i[2243];
  assign o[2242] = i[2242];
  assign o[2241] = i[2241];
  assign o[2240] = i[2240];
  assign o[2239] = i[2239];
  assign o[2238] = i[2238];
  assign o[2237] = i[2237];
  assign o[2236] = i[2236];
  assign o[2235] = i[2235];
  assign o[2234] = i[2234];
  assign o[2233] = i[2233];
  assign o[2232] = i[2232];
  assign o[2231] = i[2231];
  assign o[2230] = i[2230];
  assign o[2229] = i[2229];
  assign o[2228] = i[2228];
  assign o[2227] = i[2227];
  assign o[2226] = i[2226];
  assign o[2225] = i[2225];
  assign o[2224] = i[2224];
  assign o[2223] = i[2223];
  assign o[2222] = i[2222];
  assign o[2221] = i[2221];
  assign o[2220] = i[2220];
  assign o[2219] = i[2219];
  assign o[2218] = i[2218];
  assign o[2217] = i[2217];
  assign o[2216] = i[2216];
  assign o[2215] = i[2215];
  assign o[2214] = i[2214];
  assign o[2213] = i[2213];
  assign o[2212] = i[2212];
  assign o[2211] = i[2211];
  assign o[2210] = i[2210];
  assign o[2209] = i[2209];
  assign o[2208] = i[2208];
  assign o[2207] = i[2207];
  assign o[2206] = i[2206];
  assign o[2205] = i[2205];
  assign o[2204] = i[2204];
  assign o[2203] = i[2203];
  assign o[2202] = i[2202];
  assign o[2201] = i[2201];
  assign o[2200] = i[2200];
  assign o[2199] = i[2199];
  assign o[2198] = i[2198];
  assign o[2197] = i[2197];
  assign o[2196] = i[2196];
  assign o[2195] = i[2195];
  assign o[2194] = i[2194];
  assign o[2193] = i[2193];
  assign o[2192] = i[2192];
  assign o[2191] = i[2191];
  assign o[2190] = i[2190];
  assign o[2189] = i[2189];
  assign o[2188] = i[2188];
  assign o[2187] = i[2187];
  assign o[2186] = i[2186];
  assign o[2185] = i[2185];
  assign o[2184] = i[2184];
  assign o[2183] = i[2183];
  assign o[2182] = i[2182];
  assign o[2181] = i[2181];
  assign o[2180] = i[2180];
  assign o[2179] = i[2179];
  assign o[2178] = i[2178];
  assign o[2177] = i[2177];
  assign o[2176] = i[2176];
  assign o[2175] = i[2175];
  assign o[2174] = i[2174];
  assign o[2173] = i[2173];
  assign o[2172] = i[2172];
  assign o[2171] = i[2171];
  assign o[2170] = i[2170];
  assign o[2169] = i[2169];
  assign o[2168] = i[2168];
  assign o[2167] = i[2167];
  assign o[2166] = i[2166];
  assign o[2165] = i[2165];
  assign o[2164] = i[2164];
  assign o[2163] = i[2163];
  assign o[2162] = i[2162];
  assign o[2161] = i[2161];
  assign o[2160] = i[2160];
  assign o[2159] = i[2159];
  assign o[2158] = i[2158];
  assign o[2157] = i[2157];
  assign o[2156] = i[2156];
  assign o[2155] = i[2155];
  assign o[2154] = i[2154];
  assign o[2153] = i[2153];
  assign o[2152] = i[2152];
  assign o[2151] = i[2151];
  assign o[2150] = i[2150];
  assign o[2149] = i[2149];
  assign o[2148] = i[2148];
  assign o[2147] = i[2147];
  assign o[2146] = i[2146];
  assign o[2145] = i[2145];
  assign o[2144] = i[2144];
  assign o[2143] = i[2143];
  assign o[2142] = i[2142];
  assign o[2141] = i[2141];
  assign o[2140] = i[2140];
  assign o[2139] = i[2139];
  assign o[2138] = i[2138];
  assign o[2137] = i[2137];
  assign o[2136] = i[2136];
  assign o[2135] = i[2135];
  assign o[2134] = i[2134];
  assign o[2133] = i[2133];
  assign o[2132] = i[2132];
  assign o[2131] = i[2131];
  assign o[2130] = i[2130];
  assign o[2129] = i[2129];
  assign o[2128] = i[2128];
  assign o[2127] = i[2127];
  assign o[2126] = i[2126];
  assign o[2125] = i[2125];
  assign o[2124] = i[2124];
  assign o[2123] = i[2123];
  assign o[2122] = i[2122];
  assign o[2121] = i[2121];
  assign o[2120] = i[2120];
  assign o[2119] = i[2119];
  assign o[2118] = i[2118];
  assign o[2117] = i[2117];
  assign o[2116] = i[2116];
  assign o[2115] = i[2115];
  assign o[2114] = i[2114];
  assign o[2113] = i[2113];
  assign o[2112] = i[2112];
  assign o[2111] = i[2111];
  assign o[2110] = i[2110];
  assign o[2109] = i[2109];
  assign o[2108] = i[2108];
  assign o[2107] = i[2107];
  assign o[2106] = i[2106];
  assign o[2105] = i[2105];
  assign o[2104] = i[2104];
  assign o[2103] = i[2103];
  assign o[2102] = i[2102];
  assign o[2101] = i[2101];
  assign o[2100] = i[2100];
  assign o[2099] = i[2099];
  assign o[2098] = i[2098];
  assign o[2097] = i[2097];
  assign o[2096] = i[2096];
  assign o[2095] = i[2095];
  assign o[2094] = i[2094];
  assign o[2093] = i[2093];
  assign o[2092] = i[2092];
  assign o[2091] = i[2091];
  assign o[2090] = i[2090];
  assign o[2089] = i[2089];
  assign o[2088] = i[2088];
  assign o[2087] = i[2087];
  assign o[2086] = i[2086];
  assign o[2085] = i[2085];
  assign o[2084] = i[2084];
  assign o[2083] = i[2083];
  assign o[2082] = i[2082];
  assign o[2081] = i[2081];
  assign o[2080] = i[2080];
  assign o[2079] = i[2079];
  assign o[2078] = i[2078];
  assign o[2077] = i[2077];
  assign o[2076] = i[2076];
  assign o[2075] = i[2075];
  assign o[2074] = i[2074];
  assign o[2073] = i[2073];
  assign o[2072] = i[2072];
  assign o[2071] = i[2071];
  assign o[2070] = i[2070];
  assign o[2069] = i[2069];
  assign o[2068] = i[2068];
  assign o[2067] = i[2067];
  assign o[2066] = i[2066];
  assign o[2065] = i[2065];
  assign o[2064] = i[2064];
  assign o[2063] = i[2063];
  assign o[2062] = i[2062];
  assign o[2061] = i[2061];
  assign o[2060] = i[2060];
  assign o[2059] = i[2059];
  assign o[2058] = i[2058];
  assign o[2057] = i[2057];
  assign o[2056] = i[2056];
  assign o[2055] = i[2055];
  assign o[2054] = i[2054];
  assign o[2053] = i[2053];
  assign o[2052] = i[2052];
  assign o[2051] = i[2051];
  assign o[2050] = i[2050];
  assign o[2049] = i[2049];
  assign o[2048] = i[2048];
  assign o[2047] = i[2047];
  assign o[2046] = i[2046];
  assign o[2045] = i[2045];
  assign o[2044] = i[2044];
  assign o[2043] = i[2043];
  assign o[2042] = i[2042];
  assign o[2041] = i[2041];
  assign o[2040] = i[2040];
  assign o[2039] = i[2039];
  assign o[2038] = i[2038];
  assign o[2037] = i[2037];
  assign o[2036] = i[2036];
  assign o[2035] = i[2035];
  assign o[2034] = i[2034];
  assign o[2033] = i[2033];
  assign o[2032] = i[2032];
  assign o[2031] = i[2031];
  assign o[2030] = i[2030];
  assign o[2029] = i[2029];
  assign o[2028] = i[2028];
  assign o[2027] = i[2027];
  assign o[2026] = i[2026];
  assign o[2025] = i[2025];
  assign o[2024] = i[2024];
  assign o[2023] = i[2023];
  assign o[2022] = i[2022];
  assign o[2021] = i[2021];
  assign o[2020] = i[2020];
  assign o[2019] = i[2019];
  assign o[2018] = i[2018];
  assign o[2017] = i[2017];
  assign o[2016] = i[2016];
  assign o[2015] = i[2015];
  assign o[2014] = i[2014];
  assign o[2013] = i[2013];
  assign o[2012] = i[2012];
  assign o[2011] = i[2011];
  assign o[2010] = i[2010];
  assign o[2009] = i[2009];
  assign o[2008] = i[2008];
  assign o[2007] = i[2007];
  assign o[2006] = i[2006];
  assign o[2005] = i[2005];
  assign o[2004] = i[2004];
  assign o[2003] = i[2003];
  assign o[2002] = i[2002];
  assign o[2001] = i[2001];
  assign o[2000] = i[2000];
  assign o[1999] = i[1999];
  assign o[1998] = i[1998];
  assign o[1997] = i[1997];
  assign o[1996] = i[1996];
  assign o[1995] = i[1995];
  assign o[1994] = i[1994];
  assign o[1993] = i[1993];
  assign o[1992] = i[1992];
  assign o[1991] = i[1991];
  assign o[1990] = i[1990];
  assign o[1989] = i[1989];
  assign o[1988] = i[1988];
  assign o[1987] = i[1987];
  assign o[1986] = i[1986];
  assign o[1985] = i[1985];
  assign o[1984] = i[1984];
  assign o[1983] = i[1983];
  assign o[1982] = i[1982];
  assign o[1981] = i[1981];
  assign o[1980] = i[1980];
  assign o[1979] = i[1979];
  assign o[1978] = i[1978];
  assign o[1977] = i[1977];
  assign o[1976] = i[1976];
  assign o[1975] = i[1975];
  assign o[1974] = i[1974];
  assign o[1973] = i[1973];
  assign o[1972] = i[1972];
  assign o[1971] = i[1971];
  assign o[1970] = i[1970];
  assign o[1969] = i[1969];
  assign o[1968] = i[1968];
  assign o[1967] = i[1967];
  assign o[1966] = i[1966];
  assign o[1965] = i[1965];
  assign o[1964] = i[1964];
  assign o[1963] = i[1963];
  assign o[1962] = i[1962];
  assign o[1961] = i[1961];
  assign o[1960] = i[1960];
  assign o[1959] = i[1959];
  assign o[1958] = i[1958];
  assign o[1957] = i[1957];
  assign o[1956] = i[1956];
  assign o[1955] = i[1955];
  assign o[1954] = i[1954];
  assign o[1953] = i[1953];
  assign o[1952] = i[1952];
  assign o[1951] = i[1951];
  assign o[1950] = i[1950];
  assign o[1949] = i[1949];
  assign o[1948] = i[1948];
  assign o[1947] = i[1947];
  assign o[1946] = i[1946];
  assign o[1945] = i[1945];
  assign o[1944] = i[1944];
  assign o[1943] = i[1943];
  assign o[1942] = i[1942];
  assign o[1941] = i[1941];
  assign o[1940] = i[1940];
  assign o[1939] = i[1939];
  assign o[1938] = i[1938];
  assign o[1937] = i[1937];
  assign o[1936] = i[1936];
  assign o[1935] = i[1935];
  assign o[1934] = i[1934];
  assign o[1933] = i[1933];
  assign o[1932] = i[1932];
  assign o[1931] = i[1931];
  assign o[1930] = i[1930];
  assign o[1929] = i[1929];
  assign o[1928] = i[1928];
  assign o[1927] = i[1927];
  assign o[1926] = i[1926];
  assign o[1925] = i[1925];
  assign o[1924] = i[1924];
  assign o[1923] = i[1923];
  assign o[1922] = i[1922];
  assign o[1921] = i[1921];
  assign o[1920] = i[1920];
  assign o[1919] = i[1919];
  assign o[1918] = i[1918];
  assign o[1917] = i[1917];
  assign o[1916] = i[1916];
  assign o[1915] = i[1915];
  assign o[1914] = i[1914];
  assign o[1913] = i[1913];
  assign o[1912] = i[1912];
  assign o[1911] = i[1911];
  assign o[1910] = i[1910];
  assign o[1909] = i[1909];
  assign o[1908] = i[1908];
  assign o[1907] = i[1907];
  assign o[1906] = i[1906];
  assign o[1905] = i[1905];
  assign o[1904] = i[1904];
  assign o[1903] = i[1903];
  assign o[1902] = i[1902];
  assign o[1901] = i[1901];
  assign o[1900] = i[1900];
  assign o[1899] = i[1899];
  assign o[1898] = i[1898];
  assign o[1897] = i[1897];
  assign o[1896] = i[1896];
  assign o[1895] = i[1895];
  assign o[1894] = i[1894];
  assign o[1893] = i[1893];
  assign o[1892] = i[1892];
  assign o[1891] = i[1891];
  assign o[1890] = i[1890];
  assign o[1889] = i[1889];
  assign o[1888] = i[1888];
  assign o[1887] = i[1887];
  assign o[1886] = i[1886];
  assign o[1885] = i[1885];
  assign o[1884] = i[1884];
  assign o[1883] = i[1883];
  assign o[1882] = i[1882];
  assign o[1881] = i[1881];
  assign o[1880] = i[1880];
  assign o[1879] = i[1879];
  assign o[1878] = i[1878];
  assign o[1877] = i[1877];
  assign o[1876] = i[1876];
  assign o[1875] = i[1875];
  assign o[1874] = i[1874];
  assign o[1873] = i[1873];
  assign o[1872] = i[1872];
  assign o[1871] = i[1871];
  assign o[1870] = i[1870];
  assign o[1869] = i[1869];
  assign o[1868] = i[1868];
  assign o[1867] = i[1867];
  assign o[1866] = i[1866];
  assign o[1865] = i[1865];
  assign o[1864] = i[1864];
  assign o[1863] = i[1863];
  assign o[1862] = i[1862];
  assign o[1861] = i[1861];
  assign o[1860] = i[1860];
  assign o[1859] = i[1859];
  assign o[1858] = i[1858];
  assign o[1857] = i[1857];
  assign o[1856] = i[1856];
  assign o[1855] = i[1855];
  assign o[1854] = i[1854];
  assign o[1853] = i[1853];
  assign o[1852] = i[1852];
  assign o[1851] = i[1851];
  assign o[1850] = i[1850];
  assign o[1849] = i[1849];
  assign o[1848] = i[1848];
  assign o[1847] = i[1847];
  assign o[1846] = i[1846];
  assign o[1845] = i[1845];
  assign o[1844] = i[1844];
  assign o[1843] = i[1843];
  assign o[1842] = i[1842];
  assign o[1841] = i[1841];
  assign o[1840] = i[1840];
  assign o[1839] = i[1839];
  assign o[1838] = i[1838];
  assign o[1837] = i[1837];
  assign o[1836] = i[1836];
  assign o[1835] = i[1835];
  assign o[1834] = i[1834];
  assign o[1833] = i[1833];
  assign o[1832] = i[1832];
  assign o[1831] = i[1831];
  assign o[1830] = i[1830];
  assign o[1829] = i[1829];
  assign o[1828] = i[1828];
  assign o[1827] = i[1827];
  assign o[1826] = i[1826];
  assign o[1825] = i[1825];
  assign o[1824] = i[1824];
  assign o[1823] = i[1823];
  assign o[1822] = i[1822];
  assign o[1821] = i[1821];
  assign o[1820] = i[1820];
  assign o[1819] = i[1819];
  assign o[1818] = i[1818];
  assign o[1817] = i[1817];
  assign o[1816] = i[1816];
  assign o[1815] = i[1815];
  assign o[1814] = i[1814];
  assign o[1813] = i[1813];
  assign o[1812] = i[1812];
  assign o[1811] = i[1811];
  assign o[1810] = i[1810];
  assign o[1809] = i[1809];
  assign o[1808] = i[1808];
  assign o[1807] = i[1807];
  assign o[1806] = i[1806];
  assign o[1805] = i[1805];
  assign o[1804] = i[1804];
  assign o[1803] = i[1803];
  assign o[1802] = i[1802];
  assign o[1801] = i[1801];
  assign o[1800] = i[1800];
  assign o[1799] = i[1799];
  assign o[1798] = i[1798];
  assign o[1797] = i[1797];
  assign o[1796] = i[1796];
  assign o[1795] = i[1795];
  assign o[1794] = i[1794];
  assign o[1793] = i[1793];
  assign o[1792] = i[1792];
  assign o[1791] = i[1791];
  assign o[1790] = i[1790];
  assign o[1789] = i[1789];
  assign o[1788] = i[1788];
  assign o[1787] = i[1787];
  assign o[1786] = i[1786];
  assign o[1785] = i[1785];
  assign o[1784] = i[1784];
  assign o[1783] = i[1783];
  assign o[1782] = i[1782];
  assign o[1781] = i[1781];
  assign o[1780] = i[1780];
  assign o[1779] = i[1779];
  assign o[1778] = i[1778];
  assign o[1777] = i[1777];
  assign o[1776] = i[1776];
  assign o[1775] = i[1775];
  assign o[1774] = i[1774];
  assign o[1773] = i[1773];
  assign o[1772] = i[1772];
  assign o[1771] = i[1771];
  assign o[1770] = i[1770];
  assign o[1769] = i[1769];
  assign o[1768] = i[1768];
  assign o[1767] = i[1767];
  assign o[1766] = i[1766];
  assign o[1765] = i[1765];
  assign o[1764] = i[1764];
  assign o[1763] = i[1763];
  assign o[1762] = i[1762];
  assign o[1761] = i[1761];
  assign o[1760] = i[1760];
  assign o[1759] = i[1759];
  assign o[1758] = i[1758];
  assign o[1757] = i[1757];
  assign o[1756] = i[1756];
  assign o[1755] = i[1755];
  assign o[1754] = i[1754];
  assign o[1753] = i[1753];
  assign o[1752] = i[1752];
  assign o[1751] = i[1751];
  assign o[1750] = i[1750];
  assign o[1749] = i[1749];
  assign o[1748] = i[1748];
  assign o[1747] = i[1747];
  assign o[1746] = i[1746];
  assign o[1745] = i[1745];
  assign o[1744] = i[1744];
  assign o[1743] = i[1743];
  assign o[1742] = i[1742];
  assign o[1741] = i[1741];
  assign o[1740] = i[1740];
  assign o[1739] = i[1739];
  assign o[1738] = i[1738];
  assign o[1737] = i[1737];
  assign o[1736] = i[1736];
  assign o[1735] = i[1735];
  assign o[1734] = i[1734];
  assign o[1733] = i[1733];
  assign o[1732] = i[1732];
  assign o[1731] = i[1731];
  assign o[1730] = i[1730];
  assign o[1729] = i[1729];
  assign o[1728] = i[1728];
  assign o[1727] = i[1727];
  assign o[1726] = i[1726];
  assign o[1725] = i[1725];
  assign o[1724] = i[1724];
  assign o[1723] = i[1723];
  assign o[1722] = i[1722];
  assign o[1721] = i[1721];
  assign o[1720] = i[1720];
  assign o[1719] = i[1719];
  assign o[1718] = i[1718];
  assign o[1717] = i[1717];
  assign o[1716] = i[1716];
  assign o[1715] = i[1715];
  assign o[1714] = i[1714];
  assign o[1713] = i[1713];
  assign o[1712] = i[1712];
  assign o[1711] = i[1711];
  assign o[1710] = i[1710];
  assign o[1709] = i[1709];
  assign o[1708] = i[1708];
  assign o[1707] = i[1707];
  assign o[1706] = i[1706];
  assign o[1705] = i[1705];
  assign o[1704] = i[1704];
  assign o[1703] = i[1703];
  assign o[1702] = i[1702];
  assign o[1701] = i[1701];
  assign o[1700] = i[1700];
  assign o[1699] = i[1699];
  assign o[1698] = i[1698];
  assign o[1697] = i[1697];
  assign o[1696] = i[1696];
  assign o[1695] = i[1695];
  assign o[1694] = i[1694];
  assign o[1693] = i[1693];
  assign o[1692] = i[1692];
  assign o[1691] = i[1691];
  assign o[1690] = i[1690];
  assign o[1689] = i[1689];
  assign o[1688] = i[1688];
  assign o[1687] = i[1687];
  assign o[1686] = i[1686];
  assign o[1685] = i[1685];
  assign o[1684] = i[1684];
  assign o[1683] = i[1683];
  assign o[1682] = i[1682];
  assign o[1681] = i[1681];
  assign o[1680] = i[1680];
  assign o[1679] = i[1679];
  assign o[1678] = i[1678];
  assign o[1677] = i[1677];
  assign o[1676] = i[1676];
  assign o[1675] = i[1675];
  assign o[1674] = i[1674];
  assign o[1673] = i[1673];
  assign o[1672] = i[1672];
  assign o[1671] = i[1671];
  assign o[1670] = i[1670];
  assign o[1669] = i[1669];
  assign o[1668] = i[1668];
  assign o[1667] = i[1667];
  assign o[1666] = i[1666];
  assign o[1665] = i[1665];
  assign o[1664] = i[1664];
  assign o[1663] = i[1663];
  assign o[1662] = i[1662];
  assign o[1661] = i[1661];
  assign o[1660] = i[1660];
  assign o[1659] = i[1659];
  assign o[1658] = i[1658];
  assign o[1657] = i[1657];
  assign o[1656] = i[1656];
  assign o[1655] = i[1655];
  assign o[1654] = i[1654];
  assign o[1653] = i[1653];
  assign o[1652] = i[1652];
  assign o[1651] = i[1651];
  assign o[1650] = i[1650];
  assign o[1649] = i[1649];
  assign o[1648] = i[1648];
  assign o[1647] = i[1647];
  assign o[1646] = i[1646];
  assign o[1645] = i[1645];
  assign o[1644] = i[1644];
  assign o[1643] = i[1643];
  assign o[1642] = i[1642];
  assign o[1641] = i[1641];
  assign o[1640] = i[1640];
  assign o[1639] = i[1639];
  assign o[1638] = i[1638];
  assign o[1637] = i[1637];
  assign o[1636] = i[1636];
  assign o[1635] = i[1635];
  assign o[1634] = i[1634];
  assign o[1633] = i[1633];
  assign o[1632] = i[1632];
  assign o[1631] = i[1631];
  assign o[1630] = i[1630];
  assign o[1629] = i[1629];
  assign o[1628] = i[1628];
  assign o[1627] = i[1627];
  assign o[1626] = i[1626];
  assign o[1625] = i[1625];
  assign o[1624] = i[1624];
  assign o[1623] = i[1623];
  assign o[1622] = i[1622];
  assign o[1621] = i[1621];
  assign o[1620] = i[1620];
  assign o[1619] = i[1619];
  assign o[1618] = i[1618];
  assign o[1617] = i[1617];
  assign o[1616] = i[1616];
  assign o[1615] = i[1615];
  assign o[1614] = i[1614];
  assign o[1613] = i[1613];
  assign o[1612] = i[1612];
  assign o[1611] = i[1611];
  assign o[1610] = i[1610];
  assign o[1609] = i[1609];
  assign o[1608] = i[1608];
  assign o[1607] = i[1607];
  assign o[1606] = i[1606];
  assign o[1605] = i[1605];
  assign o[1604] = i[1604];
  assign o[1603] = i[1603];
  assign o[1602] = i[1602];
  assign o[1601] = i[1601];
  assign o[1600] = i[1600];
  assign o[1599] = i[1599];
  assign o[1598] = i[1598];
  assign o[1597] = i[1597];
  assign o[1596] = i[1596];
  assign o[1595] = i[1595];
  assign o[1594] = i[1594];
  assign o[1593] = i[1593];
  assign o[1592] = i[1592];
  assign o[1591] = i[1591];
  assign o[1590] = i[1590];
  assign o[1589] = i[1589];
  assign o[1588] = i[1588];
  assign o[1587] = i[1587];
  assign o[1586] = i[1586];
  assign o[1585] = i[1585];
  assign o[1584] = i[1584];
  assign o[1583] = i[1583];
  assign o[1582] = i[1582];
  assign o[1581] = i[1581];
  assign o[1580] = i[1580];
  assign o[1579] = i[1579];
  assign o[1578] = i[1578];
  assign o[1577] = i[1577];
  assign o[1576] = i[1576];
  assign o[1575] = i[1575];
  assign o[1574] = i[1574];
  assign o[1573] = i[1573];
  assign o[1572] = i[1572];
  assign o[1571] = i[1571];
  assign o[1570] = i[1570];
  assign o[1569] = i[1569];
  assign o[1568] = i[1568];
  assign o[1567] = i[1567];
  assign o[1566] = i[1566];
  assign o[1565] = i[1565];
  assign o[1564] = i[1564];
  assign o[1563] = i[1563];
  assign o[1562] = i[1562];
  assign o[1561] = i[1561];
  assign o[1560] = i[1560];
  assign o[1559] = i[1559];
  assign o[1558] = i[1558];
  assign o[1557] = i[1557];
  assign o[1556] = i[1556];
  assign o[1555] = i[1555];
  assign o[1554] = i[1554];
  assign o[1553] = i[1553];
  assign o[1552] = i[1552];
  assign o[1551] = i[1551];
  assign o[1550] = i[1550];
  assign o[1549] = i[1549];
  assign o[1548] = i[1548];
  assign o[1547] = i[1547];
  assign o[1546] = i[1546];
  assign o[1545] = i[1545];
  assign o[1544] = i[1544];
  assign o[1543] = i[1543];
  assign o[1542] = i[1542];
  assign o[1541] = i[1541];
  assign o[1540] = i[1540];
  assign o[1539] = i[1539];
  assign o[1538] = i[1538];
  assign o[1537] = i[1537];
  assign o[1536] = i[1536];
  assign o[1535] = i[1535];
  assign o[1534] = i[1534];
  assign o[1533] = i[1533];
  assign o[1532] = i[1532];
  assign o[1531] = i[1531];
  assign o[1530] = i[1530];
  assign o[1529] = i[1529];
  assign o[1528] = i[1528];
  assign o[1527] = i[1527];
  assign o[1526] = i[1526];
  assign o[1525] = i[1525];
  assign o[1524] = i[1524];
  assign o[1523] = i[1523];
  assign o[1522] = i[1522];
  assign o[1521] = i[1521];
  assign o[1520] = i[1520];
  assign o[1519] = i[1519];
  assign o[1518] = i[1518];
  assign o[1517] = i[1517];
  assign o[1516] = i[1516];
  assign o[1515] = i[1515];
  assign o[1514] = i[1514];
  assign o[1513] = i[1513];
  assign o[1512] = i[1512];
  assign o[1511] = i[1511];
  assign o[1510] = i[1510];
  assign o[1509] = i[1509];
  assign o[1508] = i[1508];
  assign o[1507] = i[1507];
  assign o[1506] = i[1506];
  assign o[1505] = i[1505];
  assign o[1504] = i[1504];
  assign o[1503] = i[1503];
  assign o[1502] = i[1502];
  assign o[1501] = i[1501];
  assign o[1500] = i[1500];
  assign o[1499] = i[1499];
  assign o[1498] = i[1498];
  assign o[1497] = i[1497];
  assign o[1496] = i[1496];
  assign o[1495] = i[1495];
  assign o[1494] = i[1494];
  assign o[1493] = i[1493];
  assign o[1492] = i[1492];
  assign o[1491] = i[1491];
  assign o[1490] = i[1490];
  assign o[1489] = i[1489];
  assign o[1488] = i[1488];
  assign o[1487] = i[1487];
  assign o[1486] = i[1486];
  assign o[1485] = i[1485];
  assign o[1484] = i[1484];
  assign o[1483] = i[1483];
  assign o[1482] = i[1482];
  assign o[1481] = i[1481];
  assign o[1480] = i[1480];
  assign o[1479] = i[1479];
  assign o[1478] = i[1478];
  assign o[1477] = i[1477];
  assign o[1476] = i[1476];
  assign o[1475] = i[1475];
  assign o[1474] = i[1474];
  assign o[1473] = i[1473];
  assign o[1472] = i[1472];
  assign o[1471] = i[1471];
  assign o[1470] = i[1470];
  assign o[1469] = i[1469];
  assign o[1468] = i[1468];
  assign o[1467] = i[1467];
  assign o[1466] = i[1466];
  assign o[1465] = i[1465];
  assign o[1464] = i[1464];
  assign o[1463] = i[1463];
  assign o[1462] = i[1462];
  assign o[1461] = i[1461];
  assign o[1460] = i[1460];
  assign o[1459] = i[1459];
  assign o[1458] = i[1458];
  assign o[1457] = i[1457];
  assign o[1456] = i[1456];
  assign o[1455] = i[1455];
  assign o[1454] = i[1454];
  assign o[1453] = i[1453];
  assign o[1452] = i[1452];
  assign o[1451] = i[1451];
  assign o[1450] = i[1450];
  assign o[1449] = i[1449];
  assign o[1448] = i[1448];
  assign o[1447] = i[1447];
  assign o[1446] = i[1446];
  assign o[1445] = i[1445];
  assign o[1444] = i[1444];
  assign o[1443] = i[1443];
  assign o[1442] = i[1442];
  assign o[1441] = i[1441];
  assign o[1440] = i[1440];
  assign o[1439] = i[1439];
  assign o[1438] = i[1438];
  assign o[1437] = i[1437];
  assign o[1436] = i[1436];
  assign o[1435] = i[1435];
  assign o[1434] = i[1434];
  assign o[1433] = i[1433];
  assign o[1432] = i[1432];
  assign o[1431] = i[1431];
  assign o[1430] = i[1430];
  assign o[1429] = i[1429];
  assign o[1428] = i[1428];
  assign o[1427] = i[1427];
  assign o[1426] = i[1426];
  assign o[1425] = i[1425];
  assign o[1424] = i[1424];
  assign o[1423] = i[1423];
  assign o[1422] = i[1422];
  assign o[1421] = i[1421];
  assign o[1420] = i[1420];
  assign o[1419] = i[1419];
  assign o[1418] = i[1418];
  assign o[1417] = i[1417];
  assign o[1416] = i[1416];
  assign o[1415] = i[1415];
  assign o[1414] = i[1414];
  assign o[1413] = i[1413];
  assign o[1412] = i[1412];
  assign o[1411] = i[1411];
  assign o[1410] = i[1410];
  assign o[1409] = i[1409];
  assign o[1408] = i[1408];
  assign o[1407] = i[1407];
  assign o[1406] = i[1406];
  assign o[1405] = i[1405];
  assign o[1404] = i[1404];
  assign o[1403] = i[1403];
  assign o[1402] = i[1402];
  assign o[1401] = i[1401];
  assign o[1400] = i[1400];
  assign o[1399] = i[1399];
  assign o[1398] = i[1398];
  assign o[1397] = i[1397];
  assign o[1396] = i[1396];
  assign o[1395] = i[1395];
  assign o[1394] = i[1394];
  assign o[1393] = i[1393];
  assign o[1392] = i[1392];
  assign o[1391] = i[1391];
  assign o[1390] = i[1390];
  assign o[1389] = i[1389];
  assign o[1388] = i[1388];
  assign o[1387] = i[1387];
  assign o[1386] = i[1386];
  assign o[1385] = i[1385];
  assign o[1384] = i[1384];
  assign o[1383] = i[1383];
  assign o[1382] = i[1382];
  assign o[1381] = i[1381];
  assign o[1380] = i[1380];
  assign o[1379] = i[1379];
  assign o[1378] = i[1378];
  assign o[1377] = i[1377];
  assign o[1376] = i[1376];
  assign o[1375] = i[1375];
  assign o[1374] = i[1374];
  assign o[1373] = i[1373];
  assign o[1372] = i[1372];
  assign o[1371] = i[1371];
  assign o[1370] = i[1370];
  assign o[1369] = i[1369];
  assign o[1368] = i[1368];
  assign o[1367] = i[1367];
  assign o[1366] = i[1366];
  assign o[1365] = i[1365];
  assign o[1364] = i[1364];
  assign o[1363] = i[1363];
  assign o[1362] = i[1362];
  assign o[1361] = i[1361];
  assign o[1360] = i[1360];
  assign o[1359] = i[1359];
  assign o[1358] = i[1358];
  assign o[1357] = i[1357];
  assign o[1356] = i[1356];
  assign o[1355] = i[1355];
  assign o[1354] = i[1354];
  assign o[1353] = i[1353];
  assign o[1352] = i[1352];
  assign o[1351] = i[1351];
  assign o[1350] = i[1350];
  assign o[1349] = i[1349];
  assign o[1348] = i[1348];
  assign o[1347] = i[1347];
  assign o[1346] = i[1346];
  assign o[1345] = i[1345];
  assign o[1344] = i[1344];
  assign o[1343] = i[1343];
  assign o[1342] = i[1342];
  assign o[1341] = i[1341];
  assign o[1340] = i[1340];
  assign o[1339] = i[1339];
  assign o[1338] = i[1338];
  assign o[1337] = i[1337];
  assign o[1336] = i[1336];
  assign o[1335] = i[1335];
  assign o[1334] = i[1334];
  assign o[1333] = i[1333];
  assign o[1332] = i[1332];
  assign o[1331] = i[1331];
  assign o[1330] = i[1330];
  assign o[1329] = i[1329];
  assign o[1328] = i[1328];
  assign o[1327] = i[1327];
  assign o[1326] = i[1326];
  assign o[1325] = i[1325];
  assign o[1324] = i[1324];
  assign o[1323] = i[1323];
  assign o[1322] = i[1322];
  assign o[1321] = i[1321];
  assign o[1320] = i[1320];
  assign o[1319] = i[1319];
  assign o[1318] = i[1318];
  assign o[1317] = i[1317];
  assign o[1316] = i[1316];
  assign o[1315] = i[1315];
  assign o[1314] = i[1314];
  assign o[1313] = i[1313];
  assign o[1312] = i[1312];
  assign o[1311] = i[1311];
  assign o[1310] = i[1310];
  assign o[1309] = i[1309];
  assign o[1308] = i[1308];
  assign o[1307] = i[1307];
  assign o[1306] = i[1306];
  assign o[1305] = i[1305];
  assign o[1304] = i[1304];
  assign o[1303] = i[1303];
  assign o[1302] = i[1302];
  assign o[1301] = i[1301];
  assign o[1300] = i[1300];
  assign o[1299] = i[1299];
  assign o[1298] = i[1298];
  assign o[1297] = i[1297];
  assign o[1296] = i[1296];
  assign o[1295] = i[1295];
  assign o[1294] = i[1294];
  assign o[1293] = i[1293];
  assign o[1292] = i[1292];
  assign o[1291] = i[1291];
  assign o[1290] = i[1290];
  assign o[1289] = i[1289];
  assign o[1288] = i[1288];
  assign o[1287] = i[1287];
  assign o[1286] = i[1286];
  assign o[1285] = i[1285];
  assign o[1284] = i[1284];
  assign o[1283] = i[1283];
  assign o[1282] = i[1282];
  assign o[1281] = i[1281];
  assign o[1280] = i[1280];
  assign o[1279] = i[1279];
  assign o[1278] = i[1278];
  assign o[1277] = i[1277];
  assign o[1276] = i[1276];
  assign o[1275] = i[1275];
  assign o[1274] = i[1274];
  assign o[1273] = i[1273];
  assign o[1272] = i[1272];
  assign o[1271] = i[1271];
  assign o[1270] = i[1270];
  assign o[1269] = i[1269];
  assign o[1268] = i[1268];
  assign o[1267] = i[1267];
  assign o[1266] = i[1266];
  assign o[1265] = i[1265];
  assign o[1264] = i[1264];
  assign o[1263] = i[1263];
  assign o[1262] = i[1262];
  assign o[1261] = i[1261];
  assign o[1260] = i[1260];
  assign o[1259] = i[1259];
  assign o[1258] = i[1258];
  assign o[1257] = i[1257];
  assign o[1256] = i[1256];
  assign o[1255] = i[1255];
  assign o[1254] = i[1254];
  assign o[1253] = i[1253];
  assign o[1252] = i[1252];
  assign o[1251] = i[1251];
  assign o[1250] = i[1250];
  assign o[1249] = i[1249];
  assign o[1248] = i[1248];
  assign o[1247] = i[1247];
  assign o[1246] = i[1246];
  assign o[1245] = i[1245];
  assign o[1244] = i[1244];
  assign o[1243] = i[1243];
  assign o[1242] = i[1242];
  assign o[1241] = i[1241];
  assign o[1240] = i[1240];
  assign o[1239] = i[1239];
  assign o[1238] = i[1238];
  assign o[1237] = i[1237];
  assign o[1236] = i[1236];
  assign o[1235] = i[1235];
  assign o[1234] = i[1234];
  assign o[1233] = i[1233];
  assign o[1232] = i[1232];
  assign o[1231] = i[1231];
  assign o[1230] = i[1230];
  assign o[1229] = i[1229];
  assign o[1228] = i[1228];
  assign o[1227] = i[1227];
  assign o[1226] = i[1226];
  assign o[1225] = i[1225];
  assign o[1224] = i[1224];
  assign o[1223] = i[1223];
  assign o[1222] = i[1222];
  assign o[1221] = i[1221];
  assign o[1220] = i[1220];
  assign o[1219] = i[1219];
  assign o[1218] = i[1218];
  assign o[1217] = i[1217];
  assign o[1216] = i[1216];
  assign o[1215] = i[1215];
  assign o[1214] = i[1214];
  assign o[1213] = i[1213];
  assign o[1212] = i[1212];
  assign o[1211] = i[1211];
  assign o[1210] = i[1210];
  assign o[1209] = i[1209];
  assign o[1208] = i[1208];
  assign o[1207] = i[1207];
  assign o[1206] = i[1206];
  assign o[1205] = i[1205];
  assign o[1204] = i[1204];
  assign o[1203] = i[1203];
  assign o[1202] = i[1202];
  assign o[1201] = i[1201];
  assign o[1200] = i[1200];
  assign o[1199] = i[1199];
  assign o[1198] = i[1198];
  assign o[1197] = i[1197];
  assign o[1196] = i[1196];
  assign o[1195] = i[1195];
  assign o[1194] = i[1194];
  assign o[1193] = i[1193];
  assign o[1192] = i[1192];
  assign o[1191] = i[1191];
  assign o[1190] = i[1190];
  assign o[1189] = i[1189];
  assign o[1188] = i[1188];
  assign o[1187] = i[1187];
  assign o[1186] = i[1186];
  assign o[1185] = i[1185];
  assign o[1184] = i[1184];
  assign o[1183] = i[1183];
  assign o[1182] = i[1182];
  assign o[1181] = i[1181];
  assign o[1180] = i[1180];
  assign o[1179] = i[1179];
  assign o[1178] = i[1178];
  assign o[1177] = i[1177];
  assign o[1176] = i[1176];
  assign o[1175] = i[1175];
  assign o[1174] = i[1174];
  assign o[1173] = i[1173];
  assign o[1172] = i[1172];
  assign o[1171] = i[1171];
  assign o[1170] = i[1170];
  assign o[1169] = i[1169];
  assign o[1168] = i[1168];
  assign o[1167] = i[1167];
  assign o[1166] = i[1166];
  assign o[1165] = i[1165];
  assign o[1164] = i[1164];
  assign o[1163] = i[1163];
  assign o[1162] = i[1162];
  assign o[1161] = i[1161];
  assign o[1160] = i[1160];
  assign o[1159] = i[1159];
  assign o[1158] = i[1158];
  assign o[1157] = i[1157];
  assign o[1156] = i[1156];
  assign o[1155] = i[1155];
  assign o[1154] = i[1154];
  assign o[1153] = i[1153];
  assign o[1152] = i[1152];
  assign o[1151] = i[1151];
  assign o[1150] = i[1150];
  assign o[1149] = i[1149];
  assign o[1148] = i[1148];
  assign o[1147] = i[1147];
  assign o[1146] = i[1146];
  assign o[1145] = i[1145];
  assign o[1144] = i[1144];
  assign o[1143] = i[1143];
  assign o[1142] = i[1142];
  assign o[1141] = i[1141];
  assign o[1140] = i[1140];
  assign o[1139] = i[1139];
  assign o[1138] = i[1138];
  assign o[1137] = i[1137];
  assign o[1136] = i[1136];
  assign o[1135] = i[1135];
  assign o[1134] = i[1134];
  assign o[1133] = i[1133];
  assign o[1132] = i[1132];
  assign o[1131] = i[1131];
  assign o[1130] = i[1130];
  assign o[1129] = i[1129];
  assign o[1128] = i[1128];
  assign o[1127] = i[1127];
  assign o[1126] = i[1126];
  assign o[1125] = i[1125];
  assign o[1124] = i[1124];
  assign o[1123] = i[1123];
  assign o[1122] = i[1122];
  assign o[1121] = i[1121];
  assign o[1120] = i[1120];
  assign o[1119] = i[1119];
  assign o[1118] = i[1118];
  assign o[1117] = i[1117];
  assign o[1116] = i[1116];
  assign o[1115] = i[1115];
  assign o[1114] = i[1114];
  assign o[1113] = i[1113];
  assign o[1112] = i[1112];
  assign o[1111] = i[1111];
  assign o[1110] = i[1110];
  assign o[1109] = i[1109];
  assign o[1108] = i[1108];
  assign o[1107] = i[1107];
  assign o[1106] = i[1106];
  assign o[1105] = i[1105];
  assign o[1104] = i[1104];
  assign o[1103] = i[1103];
  assign o[1102] = i[1102];
  assign o[1101] = i[1101];
  assign o[1100] = i[1100];
  assign o[1099] = i[1099];
  assign o[1098] = i[1098];
  assign o[1097] = i[1097];
  assign o[1096] = i[1096];
  assign o[1095] = i[1095];
  assign o[1094] = i[1094];
  assign o[1093] = i[1093];
  assign o[1092] = i[1092];
  assign o[1091] = i[1091];
  assign o[1090] = i[1090];
  assign o[1089] = i[1089];
  assign o[1088] = i[1088];
  assign o[1087] = i[1087];
  assign o[1086] = i[1086];
  assign o[1085] = i[1085];
  assign o[1084] = i[1084];
  assign o[1083] = i[1083];
  assign o[1082] = i[1082];
  assign o[1081] = i[1081];
  assign o[1080] = i[1080];
  assign o[1079] = i[1079];
  assign o[1078] = i[1078];
  assign o[1077] = i[1077];
  assign o[1076] = i[1076];
  assign o[1075] = i[1075];
  assign o[1074] = i[1074];
  assign o[1073] = i[1073];
  assign o[1072] = i[1072];
  assign o[1071] = i[1071];
  assign o[1070] = i[1070];
  assign o[1069] = i[1069];
  assign o[1068] = i[1068];
  assign o[1067] = i[1067];
  assign o[1066] = i[1066];
  assign o[1065] = i[1065];
  assign o[1064] = i[1064];
  assign o[1063] = i[1063];
  assign o[1062] = i[1062];
  assign o[1061] = i[1061];
  assign o[1060] = i[1060];
  assign o[1059] = i[1059];
  assign o[1058] = i[1058];
  assign o[1057] = i[1057];
  assign o[1056] = i[1056];
  assign o[1055] = i[1055];
  assign o[1054] = i[1054];
  assign o[1053] = i[1053];
  assign o[1052] = i[1052];
  assign o[1051] = i[1051];
  assign o[1050] = i[1050];
  assign o[1049] = i[1049];
  assign o[1048] = i[1048];
  assign o[1047] = i[1047];
  assign o[1046] = i[1046];
  assign o[1045] = i[1045];
  assign o[1044] = i[1044];
  assign o[1043] = i[1043];
  assign o[1042] = i[1042];
  assign o[1041] = i[1041];
  assign o[1040] = i[1040];
  assign o[1039] = i[1039];
  assign o[1038] = i[1038];
  assign o[1037] = i[1037];
  assign o[1036] = i[1036];
  assign o[1035] = i[1035];
  assign o[1034] = i[1034];
  assign o[1033] = i[1033];
  assign o[1032] = i[1032];
  assign o[1031] = i[1031];
  assign o[1030] = i[1030];
  assign o[1029] = i[1029];
  assign o[1028] = i[1028];
  assign o[1027] = i[1027];
  assign o[1026] = i[1026];
  assign o[1025] = i[1025];
  assign o[1024] = i[1024];
  assign o[1023] = i[1023];
  assign o[1022] = i[1022];
  assign o[1021] = i[1021];
  assign o[1020] = i[1020];
  assign o[1019] = i[1019];
  assign o[1018] = i[1018];
  assign o[1017] = i[1017];
  assign o[1016] = i[1016];
  assign o[1015] = i[1015];
  assign o[1014] = i[1014];
  assign o[1013] = i[1013];
  assign o[1012] = i[1012];
  assign o[1011] = i[1011];
  assign o[1010] = i[1010];
  assign o[1009] = i[1009];
  assign o[1008] = i[1008];
  assign o[1007] = i[1007];
  assign o[1006] = i[1006];
  assign o[1005] = i[1005];
  assign o[1004] = i[1004];
  assign o[1003] = i[1003];
  assign o[1002] = i[1002];
  assign o[1001] = i[1001];
  assign o[1000] = i[1000];
  assign o[999] = i[999];
  assign o[998] = i[998];
  assign o[997] = i[997];
  assign o[996] = i[996];
  assign o[995] = i[995];
  assign o[994] = i[994];
  assign o[993] = i[993];
  assign o[992] = i[992];
  assign o[991] = i[991];
  assign o[990] = i[990];
  assign o[989] = i[989];
  assign o[988] = i[988];
  assign o[987] = i[987];
  assign o[986] = i[986];
  assign o[985] = i[985];
  assign o[984] = i[984];
  assign o[983] = i[983];
  assign o[982] = i[982];
  assign o[981] = i[981];
  assign o[980] = i[980];
  assign o[979] = i[979];
  assign o[978] = i[978];
  assign o[977] = i[977];
  assign o[976] = i[976];
  assign o[975] = i[975];
  assign o[974] = i[974];
  assign o[973] = i[973];
  assign o[972] = i[972];
  assign o[971] = i[971];
  assign o[970] = i[970];
  assign o[969] = i[969];
  assign o[968] = i[968];
  assign o[967] = i[967];
  assign o[966] = i[966];
  assign o[965] = i[965];
  assign o[964] = i[964];
  assign o[963] = i[963];
  assign o[962] = i[962];
  assign o[961] = i[961];
  assign o[960] = i[960];
  assign o[959] = i[959];
  assign o[958] = i[958];
  assign o[957] = i[957];
  assign o[956] = i[956];
  assign o[955] = i[955];
  assign o[954] = i[954];
  assign o[953] = i[953];
  assign o[952] = i[952];
  assign o[951] = i[951];
  assign o[950] = i[950];
  assign o[949] = i[949];
  assign o[948] = i[948];
  assign o[947] = i[947];
  assign o[946] = i[946];
  assign o[945] = i[945];
  assign o[944] = i[944];
  assign o[943] = i[943];
  assign o[942] = i[942];
  assign o[941] = i[941];
  assign o[940] = i[940];
  assign o[939] = i[939];
  assign o[938] = i[938];
  assign o[937] = i[937];
  assign o[936] = i[936];
  assign o[935] = i[935];
  assign o[934] = i[934];
  assign o[933] = i[933];
  assign o[932] = i[932];
  assign o[931] = i[931];
  assign o[930] = i[930];
  assign o[929] = i[929];
  assign o[928] = i[928];
  assign o[927] = i[927];
  assign o[926] = i[926];
  assign o[925] = i[925];
  assign o[924] = i[924];
  assign o[923] = i[923];
  assign o[922] = i[922];
  assign o[921] = i[921];
  assign o[920] = i[920];
  assign o[919] = i[919];
  assign o[918] = i[918];
  assign o[917] = i[917];
  assign o[916] = i[916];
  assign o[915] = i[915];
  assign o[914] = i[914];
  assign o[913] = i[913];
  assign o[912] = i[912];
  assign o[911] = i[911];
  assign o[910] = i[910];
  assign o[909] = i[909];
  assign o[908] = i[908];
  assign o[907] = i[907];
  assign o[906] = i[906];
  assign o[905] = i[905];
  assign o[904] = i[904];
  assign o[903] = i[903];
  assign o[902] = i[902];
  assign o[901] = i[901];
  assign o[900] = i[900];
  assign o[899] = i[899];
  assign o[898] = i[898];
  assign o[897] = i[897];
  assign o[896] = i[896];
  assign o[895] = i[895];
  assign o[894] = i[894];
  assign o[893] = i[893];
  assign o[892] = i[892];
  assign o[891] = i[891];
  assign o[890] = i[890];
  assign o[889] = i[889];
  assign o[888] = i[888];
  assign o[887] = i[887];
  assign o[886] = i[886];
  assign o[885] = i[885];
  assign o[884] = i[884];
  assign o[883] = i[883];
  assign o[882] = i[882];
  assign o[881] = i[881];
  assign o[880] = i[880];
  assign o[879] = i[879];
  assign o[878] = i[878];
  assign o[877] = i[877];
  assign o[876] = i[876];
  assign o[875] = i[875];
  assign o[874] = i[874];
  assign o[873] = i[873];
  assign o[872] = i[872];
  assign o[871] = i[871];
  assign o[870] = i[870];
  assign o[869] = i[869];
  assign o[868] = i[868];
  assign o[867] = i[867];
  assign o[866] = i[866];
  assign o[865] = i[865];
  assign o[864] = i[864];
  assign o[863] = i[863];
  assign o[862] = i[862];
  assign o[861] = i[861];
  assign o[860] = i[860];
  assign o[859] = i[859];
  assign o[858] = i[858];
  assign o[857] = i[857];
  assign o[856] = i[856];
  assign o[855] = i[855];
  assign o[854] = i[854];
  assign o[853] = i[853];
  assign o[852] = i[852];
  assign o[851] = i[851];
  assign o[850] = i[850];
  assign o[849] = i[849];
  assign o[848] = i[848];
  assign o[847] = i[847];
  assign o[846] = i[846];
  assign o[845] = i[845];
  assign o[844] = i[844];
  assign o[843] = i[843];
  assign o[842] = i[842];
  assign o[841] = i[841];
  assign o[840] = i[840];
  assign o[839] = i[839];
  assign o[838] = i[838];
  assign o[837] = i[837];
  assign o[836] = i[836];
  assign o[835] = i[835];
  assign o[834] = i[834];
  assign o[833] = i[833];
  assign o[832] = i[832];
  assign o[831] = i[831];
  assign o[830] = i[830];
  assign o[829] = i[829];
  assign o[828] = i[828];
  assign o[827] = i[827];
  assign o[826] = i[826];
  assign o[825] = i[825];
  assign o[824] = i[824];
  assign o[823] = i[823];
  assign o[822] = i[822];
  assign o[821] = i[821];
  assign o[820] = i[820];
  assign o[819] = i[819];
  assign o[818] = i[818];
  assign o[817] = i[817];
  assign o[816] = i[816];
  assign o[815] = i[815];
  assign o[814] = i[814];
  assign o[813] = i[813];
  assign o[812] = i[812];
  assign o[811] = i[811];
  assign o[810] = i[810];
  assign o[809] = i[809];
  assign o[808] = i[808];
  assign o[807] = i[807];
  assign o[806] = i[806];
  assign o[805] = i[805];
  assign o[804] = i[804];
  assign o[803] = i[803];
  assign o[802] = i[802];
  assign o[801] = i[801];
  assign o[800] = i[800];
  assign o[799] = i[799];
  assign o[798] = i[798];
  assign o[797] = i[797];
  assign o[796] = i[796];
  assign o[795] = i[795];
  assign o[794] = i[794];
  assign o[793] = i[793];
  assign o[792] = i[792];
  assign o[791] = i[791];
  assign o[790] = i[790];
  assign o[789] = i[789];
  assign o[788] = i[788];
  assign o[787] = i[787];
  assign o[786] = i[786];
  assign o[785] = i[785];
  assign o[784] = i[784];
  assign o[783] = i[783];
  assign o[782] = i[782];
  assign o[781] = i[781];
  assign o[780] = i[780];
  assign o[779] = i[779];
  assign o[778] = i[778];
  assign o[777] = i[777];
  assign o[776] = i[776];
  assign o[775] = i[775];
  assign o[774] = i[774];
  assign o[773] = i[773];
  assign o[772] = i[772];
  assign o[771] = i[771];
  assign o[770] = i[770];
  assign o[769] = i[769];
  assign o[768] = i[768];
  assign o[767] = i[767];
  assign o[766] = i[766];
  assign o[765] = i[765];
  assign o[764] = i[764];
  assign o[763] = i[763];
  assign o[762] = i[762];
  assign o[761] = i[761];
  assign o[760] = i[760];
  assign o[759] = i[759];
  assign o[758] = i[758];
  assign o[757] = i[757];
  assign o[756] = i[756];
  assign o[755] = i[755];
  assign o[754] = i[754];
  assign o[753] = i[753];
  assign o[752] = i[752];
  assign o[751] = i[751];
  assign o[750] = i[750];
  assign o[749] = i[749];
  assign o[748] = i[748];
  assign o[747] = i[747];
  assign o[746] = i[746];
  assign o[745] = i[745];
  assign o[744] = i[744];
  assign o[743] = i[743];
  assign o[742] = i[742];
  assign o[741] = i[741];
  assign o[740] = i[740];
  assign o[739] = i[739];
  assign o[738] = i[738];
  assign o[737] = i[737];
  assign o[736] = i[736];
  assign o[735] = i[735];
  assign o[734] = i[734];
  assign o[733] = i[733];
  assign o[732] = i[732];
  assign o[731] = i[731];
  assign o[730] = i[730];
  assign o[729] = i[729];
  assign o[728] = i[728];
  assign o[727] = i[727];
  assign o[726] = i[726];
  assign o[725] = i[725];
  assign o[724] = i[724];
  assign o[723] = i[723];
  assign o[722] = i[722];
  assign o[721] = i[721];
  assign o[720] = i[720];
  assign o[719] = i[719];
  assign o[718] = i[718];
  assign o[717] = i[717];
  assign o[716] = i[716];
  assign o[715] = i[715];
  assign o[714] = i[714];
  assign o[713] = i[713];
  assign o[712] = i[712];
  assign o[711] = i[711];
  assign o[710] = i[710];
  assign o[709] = i[709];
  assign o[708] = i[708];
  assign o[707] = i[707];
  assign o[706] = i[706];
  assign o[705] = i[705];
  assign o[704] = i[704];
  assign o[703] = i[703];
  assign o[702] = i[702];
  assign o[701] = i[701];
  assign o[700] = i[700];
  assign o[699] = i[699];
  assign o[698] = i[698];
  assign o[697] = i[697];
  assign o[696] = i[696];
  assign o[695] = i[695];
  assign o[694] = i[694];
  assign o[693] = i[693];
  assign o[692] = i[692];
  assign o[691] = i[691];
  assign o[690] = i[690];
  assign o[689] = i[689];
  assign o[688] = i[688];
  assign o[687] = i[687];
  assign o[686] = i[686];
  assign o[685] = i[685];
  assign o[684] = i[684];
  assign o[683] = i[683];
  assign o[682] = i[682];
  assign o[681] = i[681];
  assign o[680] = i[680];
  assign o[679] = i[679];
  assign o[678] = i[678];
  assign o[677] = i[677];
  assign o[676] = i[676];
  assign o[675] = i[675];
  assign o[674] = i[674];
  assign o[673] = i[673];
  assign o[672] = i[672];
  assign o[671] = i[671];
  assign o[670] = i[670];
  assign o[669] = i[669];
  assign o[668] = i[668];
  assign o[667] = i[667];
  assign o[666] = i[666];
  assign o[665] = i[665];
  assign o[664] = i[664];
  assign o[663] = i[663];
  assign o[662] = i[662];
  assign o[661] = i[661];
  assign o[660] = i[660];
  assign o[659] = i[659];
  assign o[658] = i[658];
  assign o[657] = i[657];
  assign o[656] = i[656];
  assign o[655] = i[655];
  assign o[654] = i[654];
  assign o[653] = i[653];
  assign o[652] = i[652];
  assign o[651] = i[651];
  assign o[650] = i[650];
  assign o[649] = i[649];
  assign o[648] = i[648];
  assign o[647] = i[647];
  assign o[646] = i[646];
  assign o[645] = i[645];
  assign o[644] = i[644];
  assign o[643] = i[643];
  assign o[642] = i[642];
  assign o[641] = i[641];
  assign o[640] = i[640];
  assign o[639] = i[639];
  assign o[638] = i[638];
  assign o[637] = i[637];
  assign o[636] = i[636];
  assign o[635] = i[635];
  assign o[634] = i[634];
  assign o[633] = i[633];
  assign o[632] = i[632];
  assign o[631] = i[631];
  assign o[630] = i[630];
  assign o[629] = i[629];
  assign o[628] = i[628];
  assign o[627] = i[627];
  assign o[626] = i[626];
  assign o[625] = i[625];
  assign o[624] = i[624];
  assign o[623] = i[623];
  assign o[622] = i[622];
  assign o[621] = i[621];
  assign o[620] = i[620];
  assign o[619] = i[619];
  assign o[618] = i[618];
  assign o[617] = i[617];
  assign o[616] = i[616];
  assign o[615] = i[615];
  assign o[614] = i[614];
  assign o[613] = i[613];
  assign o[612] = i[612];
  assign o[611] = i[611];
  assign o[610] = i[610];
  assign o[609] = i[609];
  assign o[608] = i[608];
  assign o[607] = i[607];
  assign o[606] = i[606];
  assign o[605] = i[605];
  assign o[604] = i[604];
  assign o[603] = i[603];
  assign o[602] = i[602];
  assign o[601] = i[601];
  assign o[600] = i[600];
  assign o[599] = i[599];
  assign o[598] = i[598];
  assign o[597] = i[597];
  assign o[596] = i[596];
  assign o[595] = i[595];
  assign o[594] = i[594];
  assign o[593] = i[593];
  assign o[592] = i[592];
  assign o[591] = i[591];
  assign o[590] = i[590];
  assign o[589] = i[589];
  assign o[588] = i[588];
  assign o[587] = i[587];
  assign o[586] = i[586];
  assign o[585] = i[585];
  assign o[584] = i[584];
  assign o[583] = i[583];
  assign o[582] = i[582];
  assign o[581] = i[581];
  assign o[580] = i[580];
  assign o[579] = i[579];
  assign o[578] = i[578];
  assign o[577] = i[577];
  assign o[576] = i[576];
  assign o[575] = i[575];
  assign o[574] = i[574];
  assign o[573] = i[573];
  assign o[572] = i[572];
  assign o[571] = i[571];
  assign o[570] = i[570];
  assign o[569] = i[569];
  assign o[568] = i[568];
  assign o[567] = i[567];
  assign o[566] = i[566];
  assign o[565] = i[565];
  assign o[564] = i[564];
  assign o[563] = i[563];
  assign o[562] = i[562];
  assign o[561] = i[561];
  assign o[560] = i[560];
  assign o[559] = i[559];
  assign o[558] = i[558];
  assign o[557] = i[557];
  assign o[556] = i[556];
  assign o[555] = i[555];
  assign o[554] = i[554];
  assign o[553] = i[553];
  assign o[552] = i[552];
  assign o[551] = i[551];
  assign o[550] = i[550];
  assign o[549] = i[549];
  assign o[548] = i[548];
  assign o[547] = i[547];
  assign o[546] = i[546];
  assign o[545] = i[545];
  assign o[544] = i[544];
  assign o[543] = i[543];
  assign o[542] = i[542];
  assign o[541] = i[541];
  assign o[540] = i[540];
  assign o[539] = i[539];
  assign o[538] = i[538];
  assign o[537] = i[537];
  assign o[536] = i[536];
  assign o[535] = i[535];
  assign o[534] = i[534];
  assign o[533] = i[533];
  assign o[532] = i[532];
  assign o[531] = i[531];
  assign o[530] = i[530];
  assign o[529] = i[529];
  assign o[528] = i[528];
  assign o[527] = i[527];
  assign o[526] = i[526];
  assign o[525] = i[525];
  assign o[524] = i[524];
  assign o[523] = i[523];
  assign o[522] = i[522];
  assign o[521] = i[521];
  assign o[520] = i[520];
  assign o[519] = i[519];
  assign o[518] = i[518];
  assign o[517] = i[517];
  assign o[516] = i[516];
  assign o[515] = i[515];
  assign o[514] = i[514];
  assign o[513] = i[513];
  assign o[512] = i[512];
  assign o[511] = i[511];
  assign o[510] = i[510];
  assign o[509] = i[509];
  assign o[508] = i[508];
  assign o[507] = i[507];
  assign o[506] = i[506];
  assign o[505] = i[505];
  assign o[504] = i[504];
  assign o[503] = i[503];
  assign o[502] = i[502];
  assign o[501] = i[501];
  assign o[500] = i[500];
  assign o[499] = i[499];
  assign o[498] = i[498];
  assign o[497] = i[497];
  assign o[496] = i[496];
  assign o[495] = i[495];
  assign o[494] = i[494];
  assign o[493] = i[493];
  assign o[492] = i[492];
  assign o[491] = i[491];
  assign o[490] = i[490];
  assign o[489] = i[489];
  assign o[488] = i[488];
  assign o[487] = i[487];
  assign o[486] = i[486];
  assign o[485] = i[485];
  assign o[484] = i[484];
  assign o[483] = i[483];
  assign o[482] = i[482];
  assign o[481] = i[481];
  assign o[480] = i[480];
  assign o[479] = i[479];
  assign o[478] = i[478];
  assign o[477] = i[477];
  assign o[476] = i[476];
  assign o[475] = i[475];
  assign o[474] = i[474];
  assign o[473] = i[473];
  assign o[472] = i[472];
  assign o[471] = i[471];
  assign o[470] = i[470];
  assign o[469] = i[469];
  assign o[468] = i[468];
  assign o[467] = i[467];
  assign o[466] = i[466];
  assign o[465] = i[465];
  assign o[464] = i[464];
  assign o[463] = i[463];
  assign o[462] = i[462];
  assign o[461] = i[461];
  assign o[460] = i[460];
  assign o[459] = i[459];
  assign o[458] = i[458];
  assign o[457] = i[457];
  assign o[456] = i[456];
  assign o[455] = i[455];
  assign o[454] = i[454];
  assign o[453] = i[453];
  assign o[452] = i[452];
  assign o[451] = i[451];
  assign o[450] = i[450];
  assign o[449] = i[449];
  assign o[448] = i[448];
  assign o[447] = i[447];
  assign o[446] = i[446];
  assign o[445] = i[445];
  assign o[444] = i[444];
  assign o[443] = i[443];
  assign o[442] = i[442];
  assign o[441] = i[441];
  assign o[440] = i[440];
  assign o[439] = i[439];
  assign o[438] = i[438];
  assign o[437] = i[437];
  assign o[436] = i[436];
  assign o[435] = i[435];
  assign o[434] = i[434];
  assign o[433] = i[433];
  assign o[432] = i[432];
  assign o[431] = i[431];
  assign o[430] = i[430];
  assign o[429] = i[429];
  assign o[428] = i[428];
  assign o[427] = i[427];
  assign o[426] = i[426];
  assign o[425] = i[425];
  assign o[424] = i[424];
  assign o[423] = i[423];
  assign o[422] = i[422];
  assign o[421] = i[421];
  assign o[420] = i[420];
  assign o[419] = i[419];
  assign o[418] = i[418];
  assign o[417] = i[417];
  assign o[416] = i[416];
  assign o[415] = i[415];
  assign o[414] = i[414];
  assign o[413] = i[413];
  assign o[412] = i[412];
  assign o[411] = i[411];
  assign o[410] = i[410];
  assign o[409] = i[409];
  assign o[408] = i[408];
  assign o[407] = i[407];
  assign o[406] = i[406];
  assign o[405] = i[405];
  assign o[404] = i[404];
  assign o[403] = i[403];
  assign o[402] = i[402];
  assign o[401] = i[401];
  assign o[400] = i[400];
  assign o[399] = i[399];
  assign o[398] = i[398];
  assign o[397] = i[397];
  assign o[396] = i[396];
  assign o[395] = i[395];
  assign o[394] = i[394];
  assign o[393] = i[393];
  assign o[392] = i[392];
  assign o[391] = i[391];
  assign o[390] = i[390];
  assign o[389] = i[389];
  assign o[388] = i[388];
  assign o[387] = i[387];
  assign o[386] = i[386];
  assign o[385] = i[385];
  assign o[384] = i[384];
  assign o[383] = i[383];
  assign o[382] = i[382];
  assign o[381] = i[381];
  assign o[380] = i[380];
  assign o[379] = i[379];
  assign o[378] = i[378];
  assign o[377] = i[377];
  assign o[376] = i[376];
  assign o[375] = i[375];
  assign o[374] = i[374];
  assign o[373] = i[373];
  assign o[372] = i[372];
  assign o[371] = i[371];
  assign o[370] = i[370];
  assign o[369] = i[369];
  assign o[368] = i[368];
  assign o[367] = i[367];
  assign o[366] = i[366];
  assign o[365] = i[365];
  assign o[364] = i[364];
  assign o[363] = i[363];
  assign o[362] = i[362];
  assign o[361] = i[361];
  assign o[360] = i[360];
  assign o[359] = i[359];
  assign o[358] = i[358];
  assign o[357] = i[357];
  assign o[356] = i[356];
  assign o[355] = i[355];
  assign o[354] = i[354];
  assign o[353] = i[353];
  assign o[352] = i[352];
  assign o[351] = i[351];
  assign o[350] = i[350];
  assign o[349] = i[349];
  assign o[348] = i[348];
  assign o[347] = i[347];
  assign o[346] = i[346];
  assign o[345] = i[345];
  assign o[344] = i[344];
  assign o[343] = i[343];
  assign o[342] = i[342];
  assign o[341] = i[341];
  assign o[340] = i[340];
  assign o[339] = i[339];
  assign o[338] = i[338];
  assign o[337] = i[337];
  assign o[336] = i[336];
  assign o[335] = i[335];
  assign o[334] = i[334];
  assign o[333] = i[333];
  assign o[332] = i[332];
  assign o[331] = i[331];
  assign o[330] = i[330];
  assign o[329] = i[329];
  assign o[328] = i[328];
  assign o[327] = i[327];
  assign o[326] = i[326];
  assign o[325] = i[325];
  assign o[324] = i[324];
  assign o[323] = i[323];
  assign o[322] = i[322];
  assign o[321] = i[321];
  assign o[320] = i[320];
  assign o[319] = i[319];
  assign o[318] = i[318];
  assign o[317] = i[317];
  assign o[316] = i[316];
  assign o[315] = i[315];
  assign o[314] = i[314];
  assign o[313] = i[313];
  assign o[312] = i[312];
  assign o[311] = i[311];
  assign o[310] = i[310];
  assign o[309] = i[309];
  assign o[308] = i[308];
  assign o[307] = i[307];
  assign o[306] = i[306];
  assign o[305] = i[305];
  assign o[304] = i[304];
  assign o[303] = i[303];
  assign o[302] = i[302];
  assign o[301] = i[301];
  assign o[300] = i[300];
  assign o[299] = i[299];
  assign o[298] = i[298];
  assign o[297] = i[297];
  assign o[296] = i[296];
  assign o[295] = i[295];
  assign o[294] = i[294];
  assign o[293] = i[293];
  assign o[292] = i[292];
  assign o[291] = i[291];
  assign o[290] = i[290];
  assign o[289] = i[289];
  assign o[288] = i[288];
  assign o[287] = i[287];
  assign o[286] = i[286];
  assign o[285] = i[285];
  assign o[284] = i[284];
  assign o[283] = i[283];
  assign o[282] = i[282];
  assign o[281] = i[281];
  assign o[280] = i[280];
  assign o[279] = i[279];
  assign o[278] = i[278];
  assign o[277] = i[277];
  assign o[276] = i[276];
  assign o[275] = i[275];
  assign o[274] = i[274];
  assign o[273] = i[273];
  assign o[272] = i[272];
  assign o[271] = i[271];
  assign o[270] = i[270];
  assign o[269] = i[269];
  assign o[268] = i[268];
  assign o[267] = i[267];
  assign o[266] = i[266];
  assign o[265] = i[265];
  assign o[264] = i[264];
  assign o[263] = i[263];
  assign o[262] = i[262];
  assign o[261] = i[261];
  assign o[260] = i[260];
  assign o[259] = i[259];
  assign o[258] = i[258];
  assign o[257] = i[257];
  assign o[256] = i[256];
  assign o[255] = i[255];
  assign o[254] = i[254];
  assign o[253] = i[253];
  assign o[252] = i[252];
  assign o[251] = i[251];
  assign o[250] = i[250];
  assign o[249] = i[249];
  assign o[248] = i[248];
  assign o[247] = i[247];
  assign o[246] = i[246];
  assign o[245] = i[245];
  assign o[244] = i[244];
  assign o[243] = i[243];
  assign o[242] = i[242];
  assign o[241] = i[241];
  assign o[240] = i[240];
  assign o[239] = i[239];
  assign o[238] = i[238];
  assign o[237] = i[237];
  assign o[236] = i[236];
  assign o[235] = i[235];
  assign o[234] = i[234];
  assign o[233] = i[233];
  assign o[232] = i[232];
  assign o[231] = i[231];
  assign o[230] = i[230];
  assign o[229] = i[229];
  assign o[228] = i[228];
  assign o[227] = i[227];
  assign o[226] = i[226];
  assign o[225] = i[225];
  assign o[224] = i[224];
  assign o[223] = i[223];
  assign o[222] = i[222];
  assign o[221] = i[221];
  assign o[220] = i[220];
  assign o[219] = i[219];
  assign o[218] = i[218];
  assign o[217] = i[217];
  assign o[216] = i[216];
  assign o[215] = i[215];
  assign o[214] = i[214];
  assign o[213] = i[213];
  assign o[212] = i[212];
  assign o[211] = i[211];
  assign o[210] = i[210];
  assign o[209] = i[209];
  assign o[208] = i[208];
  assign o[207] = i[207];
  assign o[206] = i[206];
  assign o[205] = i[205];
  assign o[204] = i[204];
  assign o[203] = i[203];
  assign o[202] = i[202];
  assign o[201] = i[201];
  assign o[200] = i[200];
  assign o[199] = i[199];
  assign o[198] = i[198];
  assign o[197] = i[197];
  assign o[196] = i[196];
  assign o[195] = i[195];
  assign o[194] = i[194];
  assign o[193] = i[193];
  assign o[192] = i[192];
  assign o[191] = i[191];
  assign o[190] = i[190];
  assign o[189] = i[189];
  assign o[188] = i[188];
  assign o[187] = i[187];
  assign o[186] = i[186];
  assign o[185] = i[185];
  assign o[184] = i[184];
  assign o[183] = i[183];
  assign o[182] = i[182];
  assign o[181] = i[181];
  assign o[180] = i[180];
  assign o[179] = i[179];
  assign o[178] = i[178];
  assign o[177] = i[177];
  assign o[176] = i[176];
  assign o[175] = i[175];
  assign o[174] = i[174];
  assign o[173] = i[173];
  assign o[172] = i[172];
  assign o[171] = i[171];
  assign o[170] = i[170];
  assign o[169] = i[169];
  assign o[168] = i[168];
  assign o[167] = i[167];
  assign o[166] = i[166];
  assign o[165] = i[165];
  assign o[164] = i[164];
  assign o[163] = i[163];
  assign o[162] = i[162];
  assign o[161] = i[161];
  assign o[160] = i[160];
  assign o[159] = i[159];
  assign o[158] = i[158];
  assign o[157] = i[157];
  assign o[156] = i[156];
  assign o[155] = i[155];
  assign o[154] = i[154];
  assign o[153] = i[153];
  assign o[152] = i[152];
  assign o[151] = i[151];
  assign o[150] = i[150];
  assign o[149] = i[149];
  assign o[148] = i[148];
  assign o[147] = i[147];
  assign o[146] = i[146];
  assign o[145] = i[145];
  assign o[144] = i[144];
  assign o[143] = i[143];
  assign o[142] = i[142];
  assign o[141] = i[141];
  assign o[140] = i[140];
  assign o[139] = i[139];
  assign o[138] = i[138];
  assign o[137] = i[137];
  assign o[136] = i[136];
  assign o[135] = i[135];
  assign o[134] = i[134];
  assign o[133] = i[133];
  assign o[132] = i[132];
  assign o[131] = i[131];
  assign o[130] = i[130];
  assign o[129] = i[129];
  assign o[128] = i[128];
  assign o[127] = i[127];
  assign o[126] = i[126];
  assign o[125] = i[125];
  assign o[124] = i[124];
  assign o[123] = i[123];
  assign o[122] = i[122];
  assign o[121] = i[121];
  assign o[120] = i[120];
  assign o[119] = i[119];
  assign o[118] = i[118];
  assign o[117] = i[117];
  assign o[116] = i[116];
  assign o[115] = i[115];
  assign o[114] = i[114];
  assign o[113] = i[113];
  assign o[112] = i[112];
  assign o[111] = i[111];
  assign o[110] = i[110];
  assign o[109] = i[109];
  assign o[108] = i[108];
  assign o[107] = i[107];
  assign o[106] = i[106];
  assign o[105] = i[105];
  assign o[104] = i[104];
  assign o[103] = i[103];
  assign o[102] = i[102];
  assign o[101] = i[101];
  assign o[100] = i[100];
  assign o[99] = i[99];
  assign o[98] = i[98];
  assign o[97] = i[97];
  assign o[96] = i[96];
  assign o[95] = i[95];
  assign o[94] = i[94];
  assign o[93] = i[93];
  assign o[92] = i[92];
  assign o[91] = i[91];
  assign o[90] = i[90];
  assign o[89] = i[89];
  assign o[88] = i[88];
  assign o[87] = i[87];
  assign o[86] = i[86];
  assign o[85] = i[85];
  assign o[84] = i[84];
  assign o[83] = i[83];
  assign o[82] = i[82];
  assign o[81] = i[81];
  assign o[80] = i[80];
  assign o[79] = i[79];
  assign o[78] = i[78];
  assign o[77] = i[77];
  assign o[76] = i[76];
  assign o[75] = i[75];
  assign o[74] = i[74];
  assign o[73] = i[73];
  assign o[72] = i[72];
  assign o[71] = i[71];
  assign o[70] = i[70];
  assign o[69] = i[69];
  assign o[68] = i[68];
  assign o[67] = i[67];
  assign o[66] = i[66];
  assign o[65] = i[65];
  assign o[64] = i[64];
  assign o[63] = i[63];
  assign o[62] = i[62];
  assign o[61] = i[61];
  assign o[60] = i[60];
  assign o[59] = i[59];
  assign o[58] = i[58];
  assign o[57] = i[57];
  assign o[56] = i[56];
  assign o[55] = i[55];
  assign o[54] = i[54];
  assign o[53] = i[53];
  assign o[52] = i[52];
  assign o[51] = i[51];
  assign o[50] = i[50];
  assign o[49] = i[49];
  assign o[48] = i[48];
  assign o[47] = i[47];
  assign o[46] = i[46];
  assign o[45] = i[45];
  assign o[44] = i[44];
  assign o[43] = i[43];
  assign o[42] = i[42];
  assign o[41] = i[41];
  assign o[40] = i[40];
  assign o[39] = i[39];
  assign o[38] = i[38];
  assign o[37] = i[37];
  assign o[36] = i[36];
  assign o[35] = i[35];
  assign o[34] = i[34];
  assign o[33] = i[33];
  assign o[32] = i[32];
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule

