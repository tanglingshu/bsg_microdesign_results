

module top
(
  clk_i,
  ready_i,
  unlock_i,
  reqs_i,
  grants_o
);

  input [127:0] reqs_i;
  output [127:0] grants_o;
  input clk_i;
  input ready_i;
  input unlock_i;

  bsg_locking_arb_fixed
  wrapper
  (
    .reqs_i(reqs_i),
    .grants_o(grants_o),
    .clk_i(clk_i),
    .ready_i(ready_i),
    .unlock_i(unlock_i)
  );


endmodule



module bsg_dff_reset_en_width_p128
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [127:0] data_i;
  output [127:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134;
  reg [127:0] data_o;
  assign { N5, N3 } = (N0)? { 1'b1, 1'b1 } : 
                      (N134)? { 1'b1, 1'b1 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N0 = reset_i;
  assign { N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N4 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N134)? data_i : 1'b0;
  assign N1 = en_i | reset_i;
  assign N2 = ~N1;
  assign N133 = ~reset_i;
  assign N134 = en_i & N133;

  always @(posedge clk_i) begin
    if(N3) begin
      { data_o[127:29], data_o[0:0] } <= { N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N4 };
    end 
    if(N5) begin
      { data_o[28:1] } <= { N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6 };
    end 
  end


endmodule



module bsg_scan_width_p128_or_p1_lo_to_hi_p0
(
  i,
  o
);

  input [127:0] i;
  output [127:0] o;
  wire [127:0] o;
  wire t_3__127_,t_3__126_,t_3__125_,t_3__124_,t_3__123_,t_3__122_,t_3__121_,t_3__120_,
  t_3__119_,t_3__118_,t_3__117_,t_3__116_,t_3__115_,t_3__114_,t_3__113_,t_3__112_,
  t_3__111_,t_3__110_,t_3__109_,t_3__108_,t_3__107_,t_3__106_,t_3__105_,t_3__104_,
  t_3__103_,t_3__102_,t_3__101_,t_3__100_,t_3__99_,t_3__98_,t_3__97_,t_3__96_,
  t_3__95_,t_3__94_,t_3__93_,t_3__92_,t_3__91_,t_3__90_,t_3__89_,t_3__88_,t_3__87_,
  t_3__86_,t_3__85_,t_3__84_,t_3__83_,t_3__82_,t_3__81_,t_3__80_,t_3__79_,t_3__78_,
  t_3__77_,t_3__76_,t_3__75_,t_3__74_,t_3__73_,t_3__72_,t_3__71_,t_3__70_,t_3__69_,
  t_3__68_,t_3__67_,t_3__66_,t_3__65_,t_3__64_,t_3__63_,t_3__62_,t_3__61_,t_3__60_,
  t_3__59_,t_3__58_,t_3__57_,t_3__56_,t_3__55_,t_3__54_,t_3__53_,t_3__52_,
  t_3__51_,t_3__50_,t_3__49_,t_3__48_,t_3__47_,t_3__46_,t_3__45_,t_3__44_,t_3__43_,
  t_3__42_,t_3__41_,t_3__40_,t_3__39_,t_3__38_,t_3__37_,t_3__36_,t_3__35_,t_3__34_,
  t_3__33_,t_3__32_,t_3__31_,t_3__30_,t_3__29_,t_3__28_,t_3__27_,t_3__26_,t_3__25_,
  t_3__24_,t_3__23_,t_3__22_,t_3__21_,t_3__20_,t_3__19_,t_3__18_,t_3__17_,t_3__16_,
  t_3__15_,t_3__14_,t_3__13_,t_3__12_,t_3__11_,t_3__10_,t_3__9_,t_3__8_,t_3__7_,
  t_3__6_,t_3__5_,t_3__4_,t_3__3_,t_3__2_,t_3__1_,t_3__0_,t_2__127_,t_2__126_,t_2__125_,
  t_2__124_,t_2__123_,t_2__122_,t_2__121_,t_2__120_,t_2__119_,t_2__118_,t_2__117_,
  t_2__116_,t_2__115_,t_2__114_,t_2__113_,t_2__112_,t_2__111_,t_2__110_,t_2__109_,
  t_2__108_,t_2__107_,t_2__106_,t_2__105_,t_2__104_,t_2__103_,t_2__102_,t_2__101_,
  t_2__100_,t_2__99_,t_2__98_,t_2__97_,t_2__96_,t_2__95_,t_2__94_,t_2__93_,
  t_2__92_,t_2__91_,t_2__90_,t_2__89_,t_2__88_,t_2__87_,t_2__86_,t_2__85_,t_2__84_,
  t_2__83_,t_2__82_,t_2__81_,t_2__80_,t_2__79_,t_2__78_,t_2__77_,t_2__76_,t_2__75_,
  t_2__74_,t_2__73_,t_2__72_,t_2__71_,t_2__70_,t_2__69_,t_2__68_,t_2__67_,t_2__66_,
  t_2__65_,t_2__64_,t_2__63_,t_2__62_,t_2__61_,t_2__60_,t_2__59_,t_2__58_,t_2__57_,
  t_2__56_,t_2__55_,t_2__54_,t_2__53_,t_2__52_,t_2__51_,t_2__50_,t_2__49_,t_2__48_,
  t_2__47_,t_2__46_,t_2__45_,t_2__44_,t_2__43_,t_2__42_,t_2__41_,t_2__40_,t_2__39_,
  t_2__38_,t_2__37_,t_2__36_,t_2__35_,t_2__34_,t_2__33_,t_2__32_,t_2__31_,t_2__30_,
  t_2__29_,t_2__28_,t_2__27_,t_2__26_,t_2__25_,t_2__24_,t_2__23_,t_2__22_,
  t_2__21_,t_2__20_,t_2__19_,t_2__18_,t_2__17_,t_2__16_,t_2__15_,t_2__14_,t_2__13_,
  t_2__12_,t_2__11_,t_2__10_,t_2__9_,t_2__8_,t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,
  t_2__2_,t_2__1_,t_2__0_,t_1__127_,t_1__126_,t_1__125_,t_1__124_,t_1__123_,t_1__122_,
  t_1__121_,t_1__120_,t_1__119_,t_1__118_,t_1__117_,t_1__116_,t_1__115_,t_1__114_,
  t_1__113_,t_1__112_,t_1__111_,t_1__110_,t_1__109_,t_1__108_,t_1__107_,t_1__106_,
  t_1__105_,t_1__104_,t_1__103_,t_1__102_,t_1__101_,t_1__100_,t_1__99_,t_1__98_,
  t_1__97_,t_1__96_,t_1__95_,t_1__94_,t_1__93_,t_1__92_,t_1__91_,t_1__90_,t_1__89_,
  t_1__88_,t_1__87_,t_1__86_,t_1__85_,t_1__84_,t_1__83_,t_1__82_,t_1__81_,t_1__80_,
  t_1__79_,t_1__78_,t_1__77_,t_1__76_,t_1__75_,t_1__74_,t_1__73_,t_1__72_,
  t_1__71_,t_1__70_,t_1__69_,t_1__68_,t_1__67_,t_1__66_,t_1__65_,t_1__64_,t_1__63_,
  t_1__62_,t_1__61_,t_1__60_,t_1__59_,t_1__58_,t_1__57_,t_1__56_,t_1__55_,t_1__54_,
  t_1__53_,t_1__52_,t_1__51_,t_1__50_,t_1__49_,t_1__48_,t_1__47_,t_1__46_,t_1__45_,
  t_1__44_,t_1__43_,t_1__42_,t_1__41_,t_1__40_,t_1__39_,t_1__38_,t_1__37_,t_1__36_,
  t_1__35_,t_1__34_,t_1__33_,t_1__32_,t_1__31_,t_1__30_,t_1__29_,t_1__28_,t_1__27_,
  t_1__26_,t_1__25_,t_1__24_,t_1__23_,t_1__22_,t_1__21_,t_1__20_,t_1__19_,t_1__18_,
  t_1__17_,t_1__16_,t_1__15_,t_1__14_,t_1__13_,t_1__12_,t_1__11_,t_1__10_,t_1__9_,
  t_1__8_,t_1__7_,t_1__6_,t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_,t_6__127_,
  t_6__126_,t_6__125_,t_6__124_,t_6__123_,t_6__122_,t_6__121_,t_6__120_,t_6__119_,
  t_6__118_,t_6__117_,t_6__116_,t_6__115_,t_6__114_,t_6__113_,t_6__112_,t_6__111_,
  t_6__110_,t_6__109_,t_6__108_,t_6__107_,t_6__106_,t_6__105_,t_6__104_,t_6__103_,
  t_6__102_,t_6__101_,t_6__100_,t_6__99_,t_6__98_,t_6__97_,t_6__96_,t_6__95_,
  t_6__94_,t_6__93_,t_6__92_,t_6__91_,t_6__90_,t_6__89_,t_6__88_,t_6__87_,t_6__86_,
  t_6__85_,t_6__84_,t_6__83_,t_6__82_,t_6__81_,t_6__80_,t_6__79_,t_6__78_,t_6__77_,
  t_6__76_,t_6__75_,t_6__74_,t_6__73_,t_6__72_,t_6__71_,t_6__70_,t_6__69_,t_6__68_,
  t_6__67_,t_6__66_,t_6__65_,t_6__64_,t_6__63_,t_6__62_,t_6__61_,t_6__60_,t_6__59_,
  t_6__58_,t_6__57_,t_6__56_,t_6__55_,t_6__54_,t_6__53_,t_6__52_,t_6__51_,t_6__50_,
  t_6__49_,t_6__48_,t_6__47_,t_6__46_,t_6__45_,t_6__44_,t_6__43_,t_6__42_,
  t_6__41_,t_6__40_,t_6__39_,t_6__38_,t_6__37_,t_6__36_,t_6__35_,t_6__34_,t_6__33_,
  t_6__32_,t_6__31_,t_6__30_,t_6__29_,t_6__28_,t_6__27_,t_6__26_,t_6__25_,t_6__24_,
  t_6__23_,t_6__22_,t_6__21_,t_6__20_,t_6__19_,t_6__18_,t_6__17_,t_6__16_,t_6__15_,
  t_6__14_,t_6__13_,t_6__12_,t_6__11_,t_6__10_,t_6__9_,t_6__8_,t_6__7_,t_6__6_,t_6__5_,
  t_6__4_,t_6__3_,t_6__2_,t_6__1_,t_6__0_,t_5__127_,t_5__126_,t_5__125_,t_5__124_,
  t_5__123_,t_5__122_,t_5__121_,t_5__120_,t_5__119_,t_5__118_,t_5__117_,t_5__116_,
  t_5__115_,t_5__114_,t_5__113_,t_5__112_,t_5__111_,t_5__110_,t_5__109_,t_5__108_,
  t_5__107_,t_5__106_,t_5__105_,t_5__104_,t_5__103_,t_5__102_,t_5__101_,t_5__100_,
  t_5__99_,t_5__98_,t_5__97_,t_5__96_,t_5__95_,t_5__94_,t_5__93_,t_5__92_,
  t_5__91_,t_5__90_,t_5__89_,t_5__88_,t_5__87_,t_5__86_,t_5__85_,t_5__84_,t_5__83_,
  t_5__82_,t_5__81_,t_5__80_,t_5__79_,t_5__78_,t_5__77_,t_5__76_,t_5__75_,t_5__74_,
  t_5__73_,t_5__72_,t_5__71_,t_5__70_,t_5__69_,t_5__68_,t_5__67_,t_5__66_,t_5__65_,
  t_5__64_,t_5__63_,t_5__62_,t_5__61_,t_5__60_,t_5__59_,t_5__58_,t_5__57_,t_5__56_,
  t_5__55_,t_5__54_,t_5__53_,t_5__52_,t_5__51_,t_5__50_,t_5__49_,t_5__48_,t_5__47_,
  t_5__46_,t_5__45_,t_5__44_,t_5__43_,t_5__42_,t_5__41_,t_5__40_,t_5__39_,t_5__38_,
  t_5__37_,t_5__36_,t_5__35_,t_5__34_,t_5__33_,t_5__32_,t_5__31_,t_5__30_,t_5__29_,
  t_5__28_,t_5__27_,t_5__26_,t_5__25_,t_5__24_,t_5__23_,t_5__22_,t_5__21_,t_5__20_,
  t_5__19_,t_5__18_,t_5__17_,t_5__16_,t_5__15_,t_5__14_,t_5__13_,t_5__12_,
  t_5__11_,t_5__10_,t_5__9_,t_5__8_,t_5__7_,t_5__6_,t_5__5_,t_5__4_,t_5__3_,t_5__2_,
  t_5__1_,t_5__0_,t_4__127_,t_4__126_,t_4__125_,t_4__124_,t_4__123_,t_4__122_,t_4__121_,
  t_4__120_,t_4__119_,t_4__118_,t_4__117_,t_4__116_,t_4__115_,t_4__114_,t_4__113_,
  t_4__112_,t_4__111_,t_4__110_,t_4__109_,t_4__108_,t_4__107_,t_4__106_,t_4__105_,
  t_4__104_,t_4__103_,t_4__102_,t_4__101_,t_4__100_,t_4__99_,t_4__98_,t_4__97_,
  t_4__96_,t_4__95_,t_4__94_,t_4__93_,t_4__92_,t_4__91_,t_4__90_,t_4__89_,t_4__88_,
  t_4__87_,t_4__86_,t_4__85_,t_4__84_,t_4__83_,t_4__82_,t_4__81_,t_4__80_,t_4__79_,
  t_4__78_,t_4__77_,t_4__76_,t_4__75_,t_4__74_,t_4__73_,t_4__72_,t_4__71_,t_4__70_,
  t_4__69_,t_4__68_,t_4__67_,t_4__66_,t_4__65_,t_4__64_,t_4__63_,t_4__62_,
  t_4__61_,t_4__60_,t_4__59_,t_4__58_,t_4__57_,t_4__56_,t_4__55_,t_4__54_,t_4__53_,
  t_4__52_,t_4__51_,t_4__50_,t_4__49_,t_4__48_,t_4__47_,t_4__46_,t_4__45_,t_4__44_,
  t_4__43_,t_4__42_,t_4__41_,t_4__40_,t_4__39_,t_4__38_,t_4__37_,t_4__36_,t_4__35_,
  t_4__34_,t_4__33_,t_4__32_,t_4__31_,t_4__30_,t_4__29_,t_4__28_,t_4__27_,t_4__26_,
  t_4__25_,t_4__24_,t_4__23_,t_4__22_,t_4__21_,t_4__20_,t_4__19_,t_4__18_,t_4__17_,
  t_4__16_,t_4__15_,t_4__14_,t_4__13_,t_4__12_,t_4__11_,t_4__10_,t_4__9_,t_4__8_,
  t_4__7_,t_4__6_,t_4__5_,t_4__4_,t_4__3_,t_4__2_,t_4__1_,t_4__0_;
  assign t_1__127_ = i[127] | 1'b0;
  assign t_1__126_ = i[126] | i[127];
  assign t_1__125_ = i[125] | i[126];
  assign t_1__124_ = i[124] | i[125];
  assign t_1__123_ = i[123] | i[124];
  assign t_1__122_ = i[122] | i[123];
  assign t_1__121_ = i[121] | i[122];
  assign t_1__120_ = i[120] | i[121];
  assign t_1__119_ = i[119] | i[120];
  assign t_1__118_ = i[118] | i[119];
  assign t_1__117_ = i[117] | i[118];
  assign t_1__116_ = i[116] | i[117];
  assign t_1__115_ = i[115] | i[116];
  assign t_1__114_ = i[114] | i[115];
  assign t_1__113_ = i[113] | i[114];
  assign t_1__112_ = i[112] | i[113];
  assign t_1__111_ = i[111] | i[112];
  assign t_1__110_ = i[110] | i[111];
  assign t_1__109_ = i[109] | i[110];
  assign t_1__108_ = i[108] | i[109];
  assign t_1__107_ = i[107] | i[108];
  assign t_1__106_ = i[106] | i[107];
  assign t_1__105_ = i[105] | i[106];
  assign t_1__104_ = i[104] | i[105];
  assign t_1__103_ = i[103] | i[104];
  assign t_1__102_ = i[102] | i[103];
  assign t_1__101_ = i[101] | i[102];
  assign t_1__100_ = i[100] | i[101];
  assign t_1__99_ = i[99] | i[100];
  assign t_1__98_ = i[98] | i[99];
  assign t_1__97_ = i[97] | i[98];
  assign t_1__96_ = i[96] | i[97];
  assign t_1__95_ = i[95] | i[96];
  assign t_1__94_ = i[94] | i[95];
  assign t_1__93_ = i[93] | i[94];
  assign t_1__92_ = i[92] | i[93];
  assign t_1__91_ = i[91] | i[92];
  assign t_1__90_ = i[90] | i[91];
  assign t_1__89_ = i[89] | i[90];
  assign t_1__88_ = i[88] | i[89];
  assign t_1__87_ = i[87] | i[88];
  assign t_1__86_ = i[86] | i[87];
  assign t_1__85_ = i[85] | i[86];
  assign t_1__84_ = i[84] | i[85];
  assign t_1__83_ = i[83] | i[84];
  assign t_1__82_ = i[82] | i[83];
  assign t_1__81_ = i[81] | i[82];
  assign t_1__80_ = i[80] | i[81];
  assign t_1__79_ = i[79] | i[80];
  assign t_1__78_ = i[78] | i[79];
  assign t_1__77_ = i[77] | i[78];
  assign t_1__76_ = i[76] | i[77];
  assign t_1__75_ = i[75] | i[76];
  assign t_1__74_ = i[74] | i[75];
  assign t_1__73_ = i[73] | i[74];
  assign t_1__72_ = i[72] | i[73];
  assign t_1__71_ = i[71] | i[72];
  assign t_1__70_ = i[70] | i[71];
  assign t_1__69_ = i[69] | i[70];
  assign t_1__68_ = i[68] | i[69];
  assign t_1__67_ = i[67] | i[68];
  assign t_1__66_ = i[66] | i[67];
  assign t_1__65_ = i[65] | i[66];
  assign t_1__64_ = i[64] | i[65];
  assign t_1__63_ = i[63] | i[64];
  assign t_1__62_ = i[62] | i[63];
  assign t_1__61_ = i[61] | i[62];
  assign t_1__60_ = i[60] | i[61];
  assign t_1__59_ = i[59] | i[60];
  assign t_1__58_ = i[58] | i[59];
  assign t_1__57_ = i[57] | i[58];
  assign t_1__56_ = i[56] | i[57];
  assign t_1__55_ = i[55] | i[56];
  assign t_1__54_ = i[54] | i[55];
  assign t_1__53_ = i[53] | i[54];
  assign t_1__52_ = i[52] | i[53];
  assign t_1__51_ = i[51] | i[52];
  assign t_1__50_ = i[50] | i[51];
  assign t_1__49_ = i[49] | i[50];
  assign t_1__48_ = i[48] | i[49];
  assign t_1__47_ = i[47] | i[48];
  assign t_1__46_ = i[46] | i[47];
  assign t_1__45_ = i[45] | i[46];
  assign t_1__44_ = i[44] | i[45];
  assign t_1__43_ = i[43] | i[44];
  assign t_1__42_ = i[42] | i[43];
  assign t_1__41_ = i[41] | i[42];
  assign t_1__40_ = i[40] | i[41];
  assign t_1__39_ = i[39] | i[40];
  assign t_1__38_ = i[38] | i[39];
  assign t_1__37_ = i[37] | i[38];
  assign t_1__36_ = i[36] | i[37];
  assign t_1__35_ = i[35] | i[36];
  assign t_1__34_ = i[34] | i[35];
  assign t_1__33_ = i[33] | i[34];
  assign t_1__32_ = i[32] | i[33];
  assign t_1__31_ = i[31] | i[32];
  assign t_1__30_ = i[30] | i[31];
  assign t_1__29_ = i[29] | i[30];
  assign t_1__28_ = i[28] | i[29];
  assign t_1__27_ = i[27] | i[28];
  assign t_1__26_ = i[26] | i[27];
  assign t_1__25_ = i[25] | i[26];
  assign t_1__24_ = i[24] | i[25];
  assign t_1__23_ = i[23] | i[24];
  assign t_1__22_ = i[22] | i[23];
  assign t_1__21_ = i[21] | i[22];
  assign t_1__20_ = i[20] | i[21];
  assign t_1__19_ = i[19] | i[20];
  assign t_1__18_ = i[18] | i[19];
  assign t_1__17_ = i[17] | i[18];
  assign t_1__16_ = i[16] | i[17];
  assign t_1__15_ = i[15] | i[16];
  assign t_1__14_ = i[14] | i[15];
  assign t_1__13_ = i[13] | i[14];
  assign t_1__12_ = i[12] | i[13];
  assign t_1__11_ = i[11] | i[12];
  assign t_1__10_ = i[10] | i[11];
  assign t_1__9_ = i[9] | i[10];
  assign t_1__8_ = i[8] | i[9];
  assign t_1__7_ = i[7] | i[8];
  assign t_1__6_ = i[6] | i[7];
  assign t_1__5_ = i[5] | i[6];
  assign t_1__4_ = i[4] | i[5];
  assign t_1__3_ = i[3] | i[4];
  assign t_1__2_ = i[2] | i[3];
  assign t_1__1_ = i[1] | i[2];
  assign t_1__0_ = i[0] | i[1];
  assign t_2__127_ = t_1__127_ | 1'b0;
  assign t_2__126_ = t_1__126_ | 1'b0;
  assign t_2__125_ = t_1__125_ | t_1__127_;
  assign t_2__124_ = t_1__124_ | t_1__126_;
  assign t_2__123_ = t_1__123_ | t_1__125_;
  assign t_2__122_ = t_1__122_ | t_1__124_;
  assign t_2__121_ = t_1__121_ | t_1__123_;
  assign t_2__120_ = t_1__120_ | t_1__122_;
  assign t_2__119_ = t_1__119_ | t_1__121_;
  assign t_2__118_ = t_1__118_ | t_1__120_;
  assign t_2__117_ = t_1__117_ | t_1__119_;
  assign t_2__116_ = t_1__116_ | t_1__118_;
  assign t_2__115_ = t_1__115_ | t_1__117_;
  assign t_2__114_ = t_1__114_ | t_1__116_;
  assign t_2__113_ = t_1__113_ | t_1__115_;
  assign t_2__112_ = t_1__112_ | t_1__114_;
  assign t_2__111_ = t_1__111_ | t_1__113_;
  assign t_2__110_ = t_1__110_ | t_1__112_;
  assign t_2__109_ = t_1__109_ | t_1__111_;
  assign t_2__108_ = t_1__108_ | t_1__110_;
  assign t_2__107_ = t_1__107_ | t_1__109_;
  assign t_2__106_ = t_1__106_ | t_1__108_;
  assign t_2__105_ = t_1__105_ | t_1__107_;
  assign t_2__104_ = t_1__104_ | t_1__106_;
  assign t_2__103_ = t_1__103_ | t_1__105_;
  assign t_2__102_ = t_1__102_ | t_1__104_;
  assign t_2__101_ = t_1__101_ | t_1__103_;
  assign t_2__100_ = t_1__100_ | t_1__102_;
  assign t_2__99_ = t_1__99_ | t_1__101_;
  assign t_2__98_ = t_1__98_ | t_1__100_;
  assign t_2__97_ = t_1__97_ | t_1__99_;
  assign t_2__96_ = t_1__96_ | t_1__98_;
  assign t_2__95_ = t_1__95_ | t_1__97_;
  assign t_2__94_ = t_1__94_ | t_1__96_;
  assign t_2__93_ = t_1__93_ | t_1__95_;
  assign t_2__92_ = t_1__92_ | t_1__94_;
  assign t_2__91_ = t_1__91_ | t_1__93_;
  assign t_2__90_ = t_1__90_ | t_1__92_;
  assign t_2__89_ = t_1__89_ | t_1__91_;
  assign t_2__88_ = t_1__88_ | t_1__90_;
  assign t_2__87_ = t_1__87_ | t_1__89_;
  assign t_2__86_ = t_1__86_ | t_1__88_;
  assign t_2__85_ = t_1__85_ | t_1__87_;
  assign t_2__84_ = t_1__84_ | t_1__86_;
  assign t_2__83_ = t_1__83_ | t_1__85_;
  assign t_2__82_ = t_1__82_ | t_1__84_;
  assign t_2__81_ = t_1__81_ | t_1__83_;
  assign t_2__80_ = t_1__80_ | t_1__82_;
  assign t_2__79_ = t_1__79_ | t_1__81_;
  assign t_2__78_ = t_1__78_ | t_1__80_;
  assign t_2__77_ = t_1__77_ | t_1__79_;
  assign t_2__76_ = t_1__76_ | t_1__78_;
  assign t_2__75_ = t_1__75_ | t_1__77_;
  assign t_2__74_ = t_1__74_ | t_1__76_;
  assign t_2__73_ = t_1__73_ | t_1__75_;
  assign t_2__72_ = t_1__72_ | t_1__74_;
  assign t_2__71_ = t_1__71_ | t_1__73_;
  assign t_2__70_ = t_1__70_ | t_1__72_;
  assign t_2__69_ = t_1__69_ | t_1__71_;
  assign t_2__68_ = t_1__68_ | t_1__70_;
  assign t_2__67_ = t_1__67_ | t_1__69_;
  assign t_2__66_ = t_1__66_ | t_1__68_;
  assign t_2__65_ = t_1__65_ | t_1__67_;
  assign t_2__64_ = t_1__64_ | t_1__66_;
  assign t_2__63_ = t_1__63_ | t_1__65_;
  assign t_2__62_ = t_1__62_ | t_1__64_;
  assign t_2__61_ = t_1__61_ | t_1__63_;
  assign t_2__60_ = t_1__60_ | t_1__62_;
  assign t_2__59_ = t_1__59_ | t_1__61_;
  assign t_2__58_ = t_1__58_ | t_1__60_;
  assign t_2__57_ = t_1__57_ | t_1__59_;
  assign t_2__56_ = t_1__56_ | t_1__58_;
  assign t_2__55_ = t_1__55_ | t_1__57_;
  assign t_2__54_ = t_1__54_ | t_1__56_;
  assign t_2__53_ = t_1__53_ | t_1__55_;
  assign t_2__52_ = t_1__52_ | t_1__54_;
  assign t_2__51_ = t_1__51_ | t_1__53_;
  assign t_2__50_ = t_1__50_ | t_1__52_;
  assign t_2__49_ = t_1__49_ | t_1__51_;
  assign t_2__48_ = t_1__48_ | t_1__50_;
  assign t_2__47_ = t_1__47_ | t_1__49_;
  assign t_2__46_ = t_1__46_ | t_1__48_;
  assign t_2__45_ = t_1__45_ | t_1__47_;
  assign t_2__44_ = t_1__44_ | t_1__46_;
  assign t_2__43_ = t_1__43_ | t_1__45_;
  assign t_2__42_ = t_1__42_ | t_1__44_;
  assign t_2__41_ = t_1__41_ | t_1__43_;
  assign t_2__40_ = t_1__40_ | t_1__42_;
  assign t_2__39_ = t_1__39_ | t_1__41_;
  assign t_2__38_ = t_1__38_ | t_1__40_;
  assign t_2__37_ = t_1__37_ | t_1__39_;
  assign t_2__36_ = t_1__36_ | t_1__38_;
  assign t_2__35_ = t_1__35_ | t_1__37_;
  assign t_2__34_ = t_1__34_ | t_1__36_;
  assign t_2__33_ = t_1__33_ | t_1__35_;
  assign t_2__32_ = t_1__32_ | t_1__34_;
  assign t_2__31_ = t_1__31_ | t_1__33_;
  assign t_2__30_ = t_1__30_ | t_1__32_;
  assign t_2__29_ = t_1__29_ | t_1__31_;
  assign t_2__28_ = t_1__28_ | t_1__30_;
  assign t_2__27_ = t_1__27_ | t_1__29_;
  assign t_2__26_ = t_1__26_ | t_1__28_;
  assign t_2__25_ = t_1__25_ | t_1__27_;
  assign t_2__24_ = t_1__24_ | t_1__26_;
  assign t_2__23_ = t_1__23_ | t_1__25_;
  assign t_2__22_ = t_1__22_ | t_1__24_;
  assign t_2__21_ = t_1__21_ | t_1__23_;
  assign t_2__20_ = t_1__20_ | t_1__22_;
  assign t_2__19_ = t_1__19_ | t_1__21_;
  assign t_2__18_ = t_1__18_ | t_1__20_;
  assign t_2__17_ = t_1__17_ | t_1__19_;
  assign t_2__16_ = t_1__16_ | t_1__18_;
  assign t_2__15_ = t_1__15_ | t_1__17_;
  assign t_2__14_ = t_1__14_ | t_1__16_;
  assign t_2__13_ = t_1__13_ | t_1__15_;
  assign t_2__12_ = t_1__12_ | t_1__14_;
  assign t_2__11_ = t_1__11_ | t_1__13_;
  assign t_2__10_ = t_1__10_ | t_1__12_;
  assign t_2__9_ = t_1__9_ | t_1__11_;
  assign t_2__8_ = t_1__8_ | t_1__10_;
  assign t_2__7_ = t_1__7_ | t_1__9_;
  assign t_2__6_ = t_1__6_ | t_1__8_;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign t_3__127_ = t_2__127_ | 1'b0;
  assign t_3__126_ = t_2__126_ | 1'b0;
  assign t_3__125_ = t_2__125_ | 1'b0;
  assign t_3__124_ = t_2__124_ | 1'b0;
  assign t_3__123_ = t_2__123_ | t_2__127_;
  assign t_3__122_ = t_2__122_ | t_2__126_;
  assign t_3__121_ = t_2__121_ | t_2__125_;
  assign t_3__120_ = t_2__120_ | t_2__124_;
  assign t_3__119_ = t_2__119_ | t_2__123_;
  assign t_3__118_ = t_2__118_ | t_2__122_;
  assign t_3__117_ = t_2__117_ | t_2__121_;
  assign t_3__116_ = t_2__116_ | t_2__120_;
  assign t_3__115_ = t_2__115_ | t_2__119_;
  assign t_3__114_ = t_2__114_ | t_2__118_;
  assign t_3__113_ = t_2__113_ | t_2__117_;
  assign t_3__112_ = t_2__112_ | t_2__116_;
  assign t_3__111_ = t_2__111_ | t_2__115_;
  assign t_3__110_ = t_2__110_ | t_2__114_;
  assign t_3__109_ = t_2__109_ | t_2__113_;
  assign t_3__108_ = t_2__108_ | t_2__112_;
  assign t_3__107_ = t_2__107_ | t_2__111_;
  assign t_3__106_ = t_2__106_ | t_2__110_;
  assign t_3__105_ = t_2__105_ | t_2__109_;
  assign t_3__104_ = t_2__104_ | t_2__108_;
  assign t_3__103_ = t_2__103_ | t_2__107_;
  assign t_3__102_ = t_2__102_ | t_2__106_;
  assign t_3__101_ = t_2__101_ | t_2__105_;
  assign t_3__100_ = t_2__100_ | t_2__104_;
  assign t_3__99_ = t_2__99_ | t_2__103_;
  assign t_3__98_ = t_2__98_ | t_2__102_;
  assign t_3__97_ = t_2__97_ | t_2__101_;
  assign t_3__96_ = t_2__96_ | t_2__100_;
  assign t_3__95_ = t_2__95_ | t_2__99_;
  assign t_3__94_ = t_2__94_ | t_2__98_;
  assign t_3__93_ = t_2__93_ | t_2__97_;
  assign t_3__92_ = t_2__92_ | t_2__96_;
  assign t_3__91_ = t_2__91_ | t_2__95_;
  assign t_3__90_ = t_2__90_ | t_2__94_;
  assign t_3__89_ = t_2__89_ | t_2__93_;
  assign t_3__88_ = t_2__88_ | t_2__92_;
  assign t_3__87_ = t_2__87_ | t_2__91_;
  assign t_3__86_ = t_2__86_ | t_2__90_;
  assign t_3__85_ = t_2__85_ | t_2__89_;
  assign t_3__84_ = t_2__84_ | t_2__88_;
  assign t_3__83_ = t_2__83_ | t_2__87_;
  assign t_3__82_ = t_2__82_ | t_2__86_;
  assign t_3__81_ = t_2__81_ | t_2__85_;
  assign t_3__80_ = t_2__80_ | t_2__84_;
  assign t_3__79_ = t_2__79_ | t_2__83_;
  assign t_3__78_ = t_2__78_ | t_2__82_;
  assign t_3__77_ = t_2__77_ | t_2__81_;
  assign t_3__76_ = t_2__76_ | t_2__80_;
  assign t_3__75_ = t_2__75_ | t_2__79_;
  assign t_3__74_ = t_2__74_ | t_2__78_;
  assign t_3__73_ = t_2__73_ | t_2__77_;
  assign t_3__72_ = t_2__72_ | t_2__76_;
  assign t_3__71_ = t_2__71_ | t_2__75_;
  assign t_3__70_ = t_2__70_ | t_2__74_;
  assign t_3__69_ = t_2__69_ | t_2__73_;
  assign t_3__68_ = t_2__68_ | t_2__72_;
  assign t_3__67_ = t_2__67_ | t_2__71_;
  assign t_3__66_ = t_2__66_ | t_2__70_;
  assign t_3__65_ = t_2__65_ | t_2__69_;
  assign t_3__64_ = t_2__64_ | t_2__68_;
  assign t_3__63_ = t_2__63_ | t_2__67_;
  assign t_3__62_ = t_2__62_ | t_2__66_;
  assign t_3__61_ = t_2__61_ | t_2__65_;
  assign t_3__60_ = t_2__60_ | t_2__64_;
  assign t_3__59_ = t_2__59_ | t_2__63_;
  assign t_3__58_ = t_2__58_ | t_2__62_;
  assign t_3__57_ = t_2__57_ | t_2__61_;
  assign t_3__56_ = t_2__56_ | t_2__60_;
  assign t_3__55_ = t_2__55_ | t_2__59_;
  assign t_3__54_ = t_2__54_ | t_2__58_;
  assign t_3__53_ = t_2__53_ | t_2__57_;
  assign t_3__52_ = t_2__52_ | t_2__56_;
  assign t_3__51_ = t_2__51_ | t_2__55_;
  assign t_3__50_ = t_2__50_ | t_2__54_;
  assign t_3__49_ = t_2__49_ | t_2__53_;
  assign t_3__48_ = t_2__48_ | t_2__52_;
  assign t_3__47_ = t_2__47_ | t_2__51_;
  assign t_3__46_ = t_2__46_ | t_2__50_;
  assign t_3__45_ = t_2__45_ | t_2__49_;
  assign t_3__44_ = t_2__44_ | t_2__48_;
  assign t_3__43_ = t_2__43_ | t_2__47_;
  assign t_3__42_ = t_2__42_ | t_2__46_;
  assign t_3__41_ = t_2__41_ | t_2__45_;
  assign t_3__40_ = t_2__40_ | t_2__44_;
  assign t_3__39_ = t_2__39_ | t_2__43_;
  assign t_3__38_ = t_2__38_ | t_2__42_;
  assign t_3__37_ = t_2__37_ | t_2__41_;
  assign t_3__36_ = t_2__36_ | t_2__40_;
  assign t_3__35_ = t_2__35_ | t_2__39_;
  assign t_3__34_ = t_2__34_ | t_2__38_;
  assign t_3__33_ = t_2__33_ | t_2__37_;
  assign t_3__32_ = t_2__32_ | t_2__36_;
  assign t_3__31_ = t_2__31_ | t_2__35_;
  assign t_3__30_ = t_2__30_ | t_2__34_;
  assign t_3__29_ = t_2__29_ | t_2__33_;
  assign t_3__28_ = t_2__28_ | t_2__32_;
  assign t_3__27_ = t_2__27_ | t_2__31_;
  assign t_3__26_ = t_2__26_ | t_2__30_;
  assign t_3__25_ = t_2__25_ | t_2__29_;
  assign t_3__24_ = t_2__24_ | t_2__28_;
  assign t_3__23_ = t_2__23_ | t_2__27_;
  assign t_3__22_ = t_2__22_ | t_2__26_;
  assign t_3__21_ = t_2__21_ | t_2__25_;
  assign t_3__20_ = t_2__20_ | t_2__24_;
  assign t_3__19_ = t_2__19_ | t_2__23_;
  assign t_3__18_ = t_2__18_ | t_2__22_;
  assign t_3__17_ = t_2__17_ | t_2__21_;
  assign t_3__16_ = t_2__16_ | t_2__20_;
  assign t_3__15_ = t_2__15_ | t_2__19_;
  assign t_3__14_ = t_2__14_ | t_2__18_;
  assign t_3__13_ = t_2__13_ | t_2__17_;
  assign t_3__12_ = t_2__12_ | t_2__16_;
  assign t_3__11_ = t_2__11_ | t_2__15_;
  assign t_3__10_ = t_2__10_ | t_2__14_;
  assign t_3__9_ = t_2__9_ | t_2__13_;
  assign t_3__8_ = t_2__8_ | t_2__12_;
  assign t_3__7_ = t_2__7_ | t_2__11_;
  assign t_3__6_ = t_2__6_ | t_2__10_;
  assign t_3__5_ = t_2__5_ | t_2__9_;
  assign t_3__4_ = t_2__4_ | t_2__8_;
  assign t_3__3_ = t_2__3_ | t_2__7_;
  assign t_3__2_ = t_2__2_ | t_2__6_;
  assign t_3__1_ = t_2__1_ | t_2__5_;
  assign t_3__0_ = t_2__0_ | t_2__4_;
  assign t_4__127_ = t_3__127_ | 1'b0;
  assign t_4__126_ = t_3__126_ | 1'b0;
  assign t_4__125_ = t_3__125_ | 1'b0;
  assign t_4__124_ = t_3__124_ | 1'b0;
  assign t_4__123_ = t_3__123_ | 1'b0;
  assign t_4__122_ = t_3__122_ | 1'b0;
  assign t_4__121_ = t_3__121_ | 1'b0;
  assign t_4__120_ = t_3__120_ | 1'b0;
  assign t_4__119_ = t_3__119_ | t_3__127_;
  assign t_4__118_ = t_3__118_ | t_3__126_;
  assign t_4__117_ = t_3__117_ | t_3__125_;
  assign t_4__116_ = t_3__116_ | t_3__124_;
  assign t_4__115_ = t_3__115_ | t_3__123_;
  assign t_4__114_ = t_3__114_ | t_3__122_;
  assign t_4__113_ = t_3__113_ | t_3__121_;
  assign t_4__112_ = t_3__112_ | t_3__120_;
  assign t_4__111_ = t_3__111_ | t_3__119_;
  assign t_4__110_ = t_3__110_ | t_3__118_;
  assign t_4__109_ = t_3__109_ | t_3__117_;
  assign t_4__108_ = t_3__108_ | t_3__116_;
  assign t_4__107_ = t_3__107_ | t_3__115_;
  assign t_4__106_ = t_3__106_ | t_3__114_;
  assign t_4__105_ = t_3__105_ | t_3__113_;
  assign t_4__104_ = t_3__104_ | t_3__112_;
  assign t_4__103_ = t_3__103_ | t_3__111_;
  assign t_4__102_ = t_3__102_ | t_3__110_;
  assign t_4__101_ = t_3__101_ | t_3__109_;
  assign t_4__100_ = t_3__100_ | t_3__108_;
  assign t_4__99_ = t_3__99_ | t_3__107_;
  assign t_4__98_ = t_3__98_ | t_3__106_;
  assign t_4__97_ = t_3__97_ | t_3__105_;
  assign t_4__96_ = t_3__96_ | t_3__104_;
  assign t_4__95_ = t_3__95_ | t_3__103_;
  assign t_4__94_ = t_3__94_ | t_3__102_;
  assign t_4__93_ = t_3__93_ | t_3__101_;
  assign t_4__92_ = t_3__92_ | t_3__100_;
  assign t_4__91_ = t_3__91_ | t_3__99_;
  assign t_4__90_ = t_3__90_ | t_3__98_;
  assign t_4__89_ = t_3__89_ | t_3__97_;
  assign t_4__88_ = t_3__88_ | t_3__96_;
  assign t_4__87_ = t_3__87_ | t_3__95_;
  assign t_4__86_ = t_3__86_ | t_3__94_;
  assign t_4__85_ = t_3__85_ | t_3__93_;
  assign t_4__84_ = t_3__84_ | t_3__92_;
  assign t_4__83_ = t_3__83_ | t_3__91_;
  assign t_4__82_ = t_3__82_ | t_3__90_;
  assign t_4__81_ = t_3__81_ | t_3__89_;
  assign t_4__80_ = t_3__80_ | t_3__88_;
  assign t_4__79_ = t_3__79_ | t_3__87_;
  assign t_4__78_ = t_3__78_ | t_3__86_;
  assign t_4__77_ = t_3__77_ | t_3__85_;
  assign t_4__76_ = t_3__76_ | t_3__84_;
  assign t_4__75_ = t_3__75_ | t_3__83_;
  assign t_4__74_ = t_3__74_ | t_3__82_;
  assign t_4__73_ = t_3__73_ | t_3__81_;
  assign t_4__72_ = t_3__72_ | t_3__80_;
  assign t_4__71_ = t_3__71_ | t_3__79_;
  assign t_4__70_ = t_3__70_ | t_3__78_;
  assign t_4__69_ = t_3__69_ | t_3__77_;
  assign t_4__68_ = t_3__68_ | t_3__76_;
  assign t_4__67_ = t_3__67_ | t_3__75_;
  assign t_4__66_ = t_3__66_ | t_3__74_;
  assign t_4__65_ = t_3__65_ | t_3__73_;
  assign t_4__64_ = t_3__64_ | t_3__72_;
  assign t_4__63_ = t_3__63_ | t_3__71_;
  assign t_4__62_ = t_3__62_ | t_3__70_;
  assign t_4__61_ = t_3__61_ | t_3__69_;
  assign t_4__60_ = t_3__60_ | t_3__68_;
  assign t_4__59_ = t_3__59_ | t_3__67_;
  assign t_4__58_ = t_3__58_ | t_3__66_;
  assign t_4__57_ = t_3__57_ | t_3__65_;
  assign t_4__56_ = t_3__56_ | t_3__64_;
  assign t_4__55_ = t_3__55_ | t_3__63_;
  assign t_4__54_ = t_3__54_ | t_3__62_;
  assign t_4__53_ = t_3__53_ | t_3__61_;
  assign t_4__52_ = t_3__52_ | t_3__60_;
  assign t_4__51_ = t_3__51_ | t_3__59_;
  assign t_4__50_ = t_3__50_ | t_3__58_;
  assign t_4__49_ = t_3__49_ | t_3__57_;
  assign t_4__48_ = t_3__48_ | t_3__56_;
  assign t_4__47_ = t_3__47_ | t_3__55_;
  assign t_4__46_ = t_3__46_ | t_3__54_;
  assign t_4__45_ = t_3__45_ | t_3__53_;
  assign t_4__44_ = t_3__44_ | t_3__52_;
  assign t_4__43_ = t_3__43_ | t_3__51_;
  assign t_4__42_ = t_3__42_ | t_3__50_;
  assign t_4__41_ = t_3__41_ | t_3__49_;
  assign t_4__40_ = t_3__40_ | t_3__48_;
  assign t_4__39_ = t_3__39_ | t_3__47_;
  assign t_4__38_ = t_3__38_ | t_3__46_;
  assign t_4__37_ = t_3__37_ | t_3__45_;
  assign t_4__36_ = t_3__36_ | t_3__44_;
  assign t_4__35_ = t_3__35_ | t_3__43_;
  assign t_4__34_ = t_3__34_ | t_3__42_;
  assign t_4__33_ = t_3__33_ | t_3__41_;
  assign t_4__32_ = t_3__32_ | t_3__40_;
  assign t_4__31_ = t_3__31_ | t_3__39_;
  assign t_4__30_ = t_3__30_ | t_3__38_;
  assign t_4__29_ = t_3__29_ | t_3__37_;
  assign t_4__28_ = t_3__28_ | t_3__36_;
  assign t_4__27_ = t_3__27_ | t_3__35_;
  assign t_4__26_ = t_3__26_ | t_3__34_;
  assign t_4__25_ = t_3__25_ | t_3__33_;
  assign t_4__24_ = t_3__24_ | t_3__32_;
  assign t_4__23_ = t_3__23_ | t_3__31_;
  assign t_4__22_ = t_3__22_ | t_3__30_;
  assign t_4__21_ = t_3__21_ | t_3__29_;
  assign t_4__20_ = t_3__20_ | t_3__28_;
  assign t_4__19_ = t_3__19_ | t_3__27_;
  assign t_4__18_ = t_3__18_ | t_3__26_;
  assign t_4__17_ = t_3__17_ | t_3__25_;
  assign t_4__16_ = t_3__16_ | t_3__24_;
  assign t_4__15_ = t_3__15_ | t_3__23_;
  assign t_4__14_ = t_3__14_ | t_3__22_;
  assign t_4__13_ = t_3__13_ | t_3__21_;
  assign t_4__12_ = t_3__12_ | t_3__20_;
  assign t_4__11_ = t_3__11_ | t_3__19_;
  assign t_4__10_ = t_3__10_ | t_3__18_;
  assign t_4__9_ = t_3__9_ | t_3__17_;
  assign t_4__8_ = t_3__8_ | t_3__16_;
  assign t_4__7_ = t_3__7_ | t_3__15_;
  assign t_4__6_ = t_3__6_ | t_3__14_;
  assign t_4__5_ = t_3__5_ | t_3__13_;
  assign t_4__4_ = t_3__4_ | t_3__12_;
  assign t_4__3_ = t_3__3_ | t_3__11_;
  assign t_4__2_ = t_3__2_ | t_3__10_;
  assign t_4__1_ = t_3__1_ | t_3__9_;
  assign t_4__0_ = t_3__0_ | t_3__8_;
  assign t_5__127_ = t_4__127_ | 1'b0;
  assign t_5__126_ = t_4__126_ | 1'b0;
  assign t_5__125_ = t_4__125_ | 1'b0;
  assign t_5__124_ = t_4__124_ | 1'b0;
  assign t_5__123_ = t_4__123_ | 1'b0;
  assign t_5__122_ = t_4__122_ | 1'b0;
  assign t_5__121_ = t_4__121_ | 1'b0;
  assign t_5__120_ = t_4__120_ | 1'b0;
  assign t_5__119_ = t_4__119_ | 1'b0;
  assign t_5__118_ = t_4__118_ | 1'b0;
  assign t_5__117_ = t_4__117_ | 1'b0;
  assign t_5__116_ = t_4__116_ | 1'b0;
  assign t_5__115_ = t_4__115_ | 1'b0;
  assign t_5__114_ = t_4__114_ | 1'b0;
  assign t_5__113_ = t_4__113_ | 1'b0;
  assign t_5__112_ = t_4__112_ | 1'b0;
  assign t_5__111_ = t_4__111_ | t_4__127_;
  assign t_5__110_ = t_4__110_ | t_4__126_;
  assign t_5__109_ = t_4__109_ | t_4__125_;
  assign t_5__108_ = t_4__108_ | t_4__124_;
  assign t_5__107_ = t_4__107_ | t_4__123_;
  assign t_5__106_ = t_4__106_ | t_4__122_;
  assign t_5__105_ = t_4__105_ | t_4__121_;
  assign t_5__104_ = t_4__104_ | t_4__120_;
  assign t_5__103_ = t_4__103_ | t_4__119_;
  assign t_5__102_ = t_4__102_ | t_4__118_;
  assign t_5__101_ = t_4__101_ | t_4__117_;
  assign t_5__100_ = t_4__100_ | t_4__116_;
  assign t_5__99_ = t_4__99_ | t_4__115_;
  assign t_5__98_ = t_4__98_ | t_4__114_;
  assign t_5__97_ = t_4__97_ | t_4__113_;
  assign t_5__96_ = t_4__96_ | t_4__112_;
  assign t_5__95_ = t_4__95_ | t_4__111_;
  assign t_5__94_ = t_4__94_ | t_4__110_;
  assign t_5__93_ = t_4__93_ | t_4__109_;
  assign t_5__92_ = t_4__92_ | t_4__108_;
  assign t_5__91_ = t_4__91_ | t_4__107_;
  assign t_5__90_ = t_4__90_ | t_4__106_;
  assign t_5__89_ = t_4__89_ | t_4__105_;
  assign t_5__88_ = t_4__88_ | t_4__104_;
  assign t_5__87_ = t_4__87_ | t_4__103_;
  assign t_5__86_ = t_4__86_ | t_4__102_;
  assign t_5__85_ = t_4__85_ | t_4__101_;
  assign t_5__84_ = t_4__84_ | t_4__100_;
  assign t_5__83_ = t_4__83_ | t_4__99_;
  assign t_5__82_ = t_4__82_ | t_4__98_;
  assign t_5__81_ = t_4__81_ | t_4__97_;
  assign t_5__80_ = t_4__80_ | t_4__96_;
  assign t_5__79_ = t_4__79_ | t_4__95_;
  assign t_5__78_ = t_4__78_ | t_4__94_;
  assign t_5__77_ = t_4__77_ | t_4__93_;
  assign t_5__76_ = t_4__76_ | t_4__92_;
  assign t_5__75_ = t_4__75_ | t_4__91_;
  assign t_5__74_ = t_4__74_ | t_4__90_;
  assign t_5__73_ = t_4__73_ | t_4__89_;
  assign t_5__72_ = t_4__72_ | t_4__88_;
  assign t_5__71_ = t_4__71_ | t_4__87_;
  assign t_5__70_ = t_4__70_ | t_4__86_;
  assign t_5__69_ = t_4__69_ | t_4__85_;
  assign t_5__68_ = t_4__68_ | t_4__84_;
  assign t_5__67_ = t_4__67_ | t_4__83_;
  assign t_5__66_ = t_4__66_ | t_4__82_;
  assign t_5__65_ = t_4__65_ | t_4__81_;
  assign t_5__64_ = t_4__64_ | t_4__80_;
  assign t_5__63_ = t_4__63_ | t_4__79_;
  assign t_5__62_ = t_4__62_ | t_4__78_;
  assign t_5__61_ = t_4__61_ | t_4__77_;
  assign t_5__60_ = t_4__60_ | t_4__76_;
  assign t_5__59_ = t_4__59_ | t_4__75_;
  assign t_5__58_ = t_4__58_ | t_4__74_;
  assign t_5__57_ = t_4__57_ | t_4__73_;
  assign t_5__56_ = t_4__56_ | t_4__72_;
  assign t_5__55_ = t_4__55_ | t_4__71_;
  assign t_5__54_ = t_4__54_ | t_4__70_;
  assign t_5__53_ = t_4__53_ | t_4__69_;
  assign t_5__52_ = t_4__52_ | t_4__68_;
  assign t_5__51_ = t_4__51_ | t_4__67_;
  assign t_5__50_ = t_4__50_ | t_4__66_;
  assign t_5__49_ = t_4__49_ | t_4__65_;
  assign t_5__48_ = t_4__48_ | t_4__64_;
  assign t_5__47_ = t_4__47_ | t_4__63_;
  assign t_5__46_ = t_4__46_ | t_4__62_;
  assign t_5__45_ = t_4__45_ | t_4__61_;
  assign t_5__44_ = t_4__44_ | t_4__60_;
  assign t_5__43_ = t_4__43_ | t_4__59_;
  assign t_5__42_ = t_4__42_ | t_4__58_;
  assign t_5__41_ = t_4__41_ | t_4__57_;
  assign t_5__40_ = t_4__40_ | t_4__56_;
  assign t_5__39_ = t_4__39_ | t_4__55_;
  assign t_5__38_ = t_4__38_ | t_4__54_;
  assign t_5__37_ = t_4__37_ | t_4__53_;
  assign t_5__36_ = t_4__36_ | t_4__52_;
  assign t_5__35_ = t_4__35_ | t_4__51_;
  assign t_5__34_ = t_4__34_ | t_4__50_;
  assign t_5__33_ = t_4__33_ | t_4__49_;
  assign t_5__32_ = t_4__32_ | t_4__48_;
  assign t_5__31_ = t_4__31_ | t_4__47_;
  assign t_5__30_ = t_4__30_ | t_4__46_;
  assign t_5__29_ = t_4__29_ | t_4__45_;
  assign t_5__28_ = t_4__28_ | t_4__44_;
  assign t_5__27_ = t_4__27_ | t_4__43_;
  assign t_5__26_ = t_4__26_ | t_4__42_;
  assign t_5__25_ = t_4__25_ | t_4__41_;
  assign t_5__24_ = t_4__24_ | t_4__40_;
  assign t_5__23_ = t_4__23_ | t_4__39_;
  assign t_5__22_ = t_4__22_ | t_4__38_;
  assign t_5__21_ = t_4__21_ | t_4__37_;
  assign t_5__20_ = t_4__20_ | t_4__36_;
  assign t_5__19_ = t_4__19_ | t_4__35_;
  assign t_5__18_ = t_4__18_ | t_4__34_;
  assign t_5__17_ = t_4__17_ | t_4__33_;
  assign t_5__16_ = t_4__16_ | t_4__32_;
  assign t_5__15_ = t_4__15_ | t_4__31_;
  assign t_5__14_ = t_4__14_ | t_4__30_;
  assign t_5__13_ = t_4__13_ | t_4__29_;
  assign t_5__12_ = t_4__12_ | t_4__28_;
  assign t_5__11_ = t_4__11_ | t_4__27_;
  assign t_5__10_ = t_4__10_ | t_4__26_;
  assign t_5__9_ = t_4__9_ | t_4__25_;
  assign t_5__8_ = t_4__8_ | t_4__24_;
  assign t_5__7_ = t_4__7_ | t_4__23_;
  assign t_5__6_ = t_4__6_ | t_4__22_;
  assign t_5__5_ = t_4__5_ | t_4__21_;
  assign t_5__4_ = t_4__4_ | t_4__20_;
  assign t_5__3_ = t_4__3_ | t_4__19_;
  assign t_5__2_ = t_4__2_ | t_4__18_;
  assign t_5__1_ = t_4__1_ | t_4__17_;
  assign t_5__0_ = t_4__0_ | t_4__16_;
  assign t_6__127_ = t_5__127_ | 1'b0;
  assign t_6__126_ = t_5__126_ | 1'b0;
  assign t_6__125_ = t_5__125_ | 1'b0;
  assign t_6__124_ = t_5__124_ | 1'b0;
  assign t_6__123_ = t_5__123_ | 1'b0;
  assign t_6__122_ = t_5__122_ | 1'b0;
  assign t_6__121_ = t_5__121_ | 1'b0;
  assign t_6__120_ = t_5__120_ | 1'b0;
  assign t_6__119_ = t_5__119_ | 1'b0;
  assign t_6__118_ = t_5__118_ | 1'b0;
  assign t_6__117_ = t_5__117_ | 1'b0;
  assign t_6__116_ = t_5__116_ | 1'b0;
  assign t_6__115_ = t_5__115_ | 1'b0;
  assign t_6__114_ = t_5__114_ | 1'b0;
  assign t_6__113_ = t_5__113_ | 1'b0;
  assign t_6__112_ = t_5__112_ | 1'b0;
  assign t_6__111_ = t_5__111_ | 1'b0;
  assign t_6__110_ = t_5__110_ | 1'b0;
  assign t_6__109_ = t_5__109_ | 1'b0;
  assign t_6__108_ = t_5__108_ | 1'b0;
  assign t_6__107_ = t_5__107_ | 1'b0;
  assign t_6__106_ = t_5__106_ | 1'b0;
  assign t_6__105_ = t_5__105_ | 1'b0;
  assign t_6__104_ = t_5__104_ | 1'b0;
  assign t_6__103_ = t_5__103_ | 1'b0;
  assign t_6__102_ = t_5__102_ | 1'b0;
  assign t_6__101_ = t_5__101_ | 1'b0;
  assign t_6__100_ = t_5__100_ | 1'b0;
  assign t_6__99_ = t_5__99_ | 1'b0;
  assign t_6__98_ = t_5__98_ | 1'b0;
  assign t_6__97_ = t_5__97_ | 1'b0;
  assign t_6__96_ = t_5__96_ | 1'b0;
  assign t_6__95_ = t_5__95_ | t_5__127_;
  assign t_6__94_ = t_5__94_ | t_5__126_;
  assign t_6__93_ = t_5__93_ | t_5__125_;
  assign t_6__92_ = t_5__92_ | t_5__124_;
  assign t_6__91_ = t_5__91_ | t_5__123_;
  assign t_6__90_ = t_5__90_ | t_5__122_;
  assign t_6__89_ = t_5__89_ | t_5__121_;
  assign t_6__88_ = t_5__88_ | t_5__120_;
  assign t_6__87_ = t_5__87_ | t_5__119_;
  assign t_6__86_ = t_5__86_ | t_5__118_;
  assign t_6__85_ = t_5__85_ | t_5__117_;
  assign t_6__84_ = t_5__84_ | t_5__116_;
  assign t_6__83_ = t_5__83_ | t_5__115_;
  assign t_6__82_ = t_5__82_ | t_5__114_;
  assign t_6__81_ = t_5__81_ | t_5__113_;
  assign t_6__80_ = t_5__80_ | t_5__112_;
  assign t_6__79_ = t_5__79_ | t_5__111_;
  assign t_6__78_ = t_5__78_ | t_5__110_;
  assign t_6__77_ = t_5__77_ | t_5__109_;
  assign t_6__76_ = t_5__76_ | t_5__108_;
  assign t_6__75_ = t_5__75_ | t_5__107_;
  assign t_6__74_ = t_5__74_ | t_5__106_;
  assign t_6__73_ = t_5__73_ | t_5__105_;
  assign t_6__72_ = t_5__72_ | t_5__104_;
  assign t_6__71_ = t_5__71_ | t_5__103_;
  assign t_6__70_ = t_5__70_ | t_5__102_;
  assign t_6__69_ = t_5__69_ | t_5__101_;
  assign t_6__68_ = t_5__68_ | t_5__100_;
  assign t_6__67_ = t_5__67_ | t_5__99_;
  assign t_6__66_ = t_5__66_ | t_5__98_;
  assign t_6__65_ = t_5__65_ | t_5__97_;
  assign t_6__64_ = t_5__64_ | t_5__96_;
  assign t_6__63_ = t_5__63_ | t_5__95_;
  assign t_6__62_ = t_5__62_ | t_5__94_;
  assign t_6__61_ = t_5__61_ | t_5__93_;
  assign t_6__60_ = t_5__60_ | t_5__92_;
  assign t_6__59_ = t_5__59_ | t_5__91_;
  assign t_6__58_ = t_5__58_ | t_5__90_;
  assign t_6__57_ = t_5__57_ | t_5__89_;
  assign t_6__56_ = t_5__56_ | t_5__88_;
  assign t_6__55_ = t_5__55_ | t_5__87_;
  assign t_6__54_ = t_5__54_ | t_5__86_;
  assign t_6__53_ = t_5__53_ | t_5__85_;
  assign t_6__52_ = t_5__52_ | t_5__84_;
  assign t_6__51_ = t_5__51_ | t_5__83_;
  assign t_6__50_ = t_5__50_ | t_5__82_;
  assign t_6__49_ = t_5__49_ | t_5__81_;
  assign t_6__48_ = t_5__48_ | t_5__80_;
  assign t_6__47_ = t_5__47_ | t_5__79_;
  assign t_6__46_ = t_5__46_ | t_5__78_;
  assign t_6__45_ = t_5__45_ | t_5__77_;
  assign t_6__44_ = t_5__44_ | t_5__76_;
  assign t_6__43_ = t_5__43_ | t_5__75_;
  assign t_6__42_ = t_5__42_ | t_5__74_;
  assign t_6__41_ = t_5__41_ | t_5__73_;
  assign t_6__40_ = t_5__40_ | t_5__72_;
  assign t_6__39_ = t_5__39_ | t_5__71_;
  assign t_6__38_ = t_5__38_ | t_5__70_;
  assign t_6__37_ = t_5__37_ | t_5__69_;
  assign t_6__36_ = t_5__36_ | t_5__68_;
  assign t_6__35_ = t_5__35_ | t_5__67_;
  assign t_6__34_ = t_5__34_ | t_5__66_;
  assign t_6__33_ = t_5__33_ | t_5__65_;
  assign t_6__32_ = t_5__32_ | t_5__64_;
  assign t_6__31_ = t_5__31_ | t_5__63_;
  assign t_6__30_ = t_5__30_ | t_5__62_;
  assign t_6__29_ = t_5__29_ | t_5__61_;
  assign t_6__28_ = t_5__28_ | t_5__60_;
  assign t_6__27_ = t_5__27_ | t_5__59_;
  assign t_6__26_ = t_5__26_ | t_5__58_;
  assign t_6__25_ = t_5__25_ | t_5__57_;
  assign t_6__24_ = t_5__24_ | t_5__56_;
  assign t_6__23_ = t_5__23_ | t_5__55_;
  assign t_6__22_ = t_5__22_ | t_5__54_;
  assign t_6__21_ = t_5__21_ | t_5__53_;
  assign t_6__20_ = t_5__20_ | t_5__52_;
  assign t_6__19_ = t_5__19_ | t_5__51_;
  assign t_6__18_ = t_5__18_ | t_5__50_;
  assign t_6__17_ = t_5__17_ | t_5__49_;
  assign t_6__16_ = t_5__16_ | t_5__48_;
  assign t_6__15_ = t_5__15_ | t_5__47_;
  assign t_6__14_ = t_5__14_ | t_5__46_;
  assign t_6__13_ = t_5__13_ | t_5__45_;
  assign t_6__12_ = t_5__12_ | t_5__44_;
  assign t_6__11_ = t_5__11_ | t_5__43_;
  assign t_6__10_ = t_5__10_ | t_5__42_;
  assign t_6__9_ = t_5__9_ | t_5__41_;
  assign t_6__8_ = t_5__8_ | t_5__40_;
  assign t_6__7_ = t_5__7_ | t_5__39_;
  assign t_6__6_ = t_5__6_ | t_5__38_;
  assign t_6__5_ = t_5__5_ | t_5__37_;
  assign t_6__4_ = t_5__4_ | t_5__36_;
  assign t_6__3_ = t_5__3_ | t_5__35_;
  assign t_6__2_ = t_5__2_ | t_5__34_;
  assign t_6__1_ = t_5__1_ | t_5__33_;
  assign t_6__0_ = t_5__0_ | t_5__32_;
  assign o[127] = t_6__127_ | 1'b0;
  assign o[126] = t_6__126_ | 1'b0;
  assign o[125] = t_6__125_ | 1'b0;
  assign o[124] = t_6__124_ | 1'b0;
  assign o[123] = t_6__123_ | 1'b0;
  assign o[122] = t_6__122_ | 1'b0;
  assign o[121] = t_6__121_ | 1'b0;
  assign o[120] = t_6__120_ | 1'b0;
  assign o[119] = t_6__119_ | 1'b0;
  assign o[118] = t_6__118_ | 1'b0;
  assign o[117] = t_6__117_ | 1'b0;
  assign o[116] = t_6__116_ | 1'b0;
  assign o[115] = t_6__115_ | 1'b0;
  assign o[114] = t_6__114_ | 1'b0;
  assign o[113] = t_6__113_ | 1'b0;
  assign o[112] = t_6__112_ | 1'b0;
  assign o[111] = t_6__111_ | 1'b0;
  assign o[110] = t_6__110_ | 1'b0;
  assign o[109] = t_6__109_ | 1'b0;
  assign o[108] = t_6__108_ | 1'b0;
  assign o[107] = t_6__107_ | 1'b0;
  assign o[106] = t_6__106_ | 1'b0;
  assign o[105] = t_6__105_ | 1'b0;
  assign o[104] = t_6__104_ | 1'b0;
  assign o[103] = t_6__103_ | 1'b0;
  assign o[102] = t_6__102_ | 1'b0;
  assign o[101] = t_6__101_ | 1'b0;
  assign o[100] = t_6__100_ | 1'b0;
  assign o[99] = t_6__99_ | 1'b0;
  assign o[98] = t_6__98_ | 1'b0;
  assign o[97] = t_6__97_ | 1'b0;
  assign o[96] = t_6__96_ | 1'b0;
  assign o[95] = t_6__95_ | 1'b0;
  assign o[94] = t_6__94_ | 1'b0;
  assign o[93] = t_6__93_ | 1'b0;
  assign o[92] = t_6__92_ | 1'b0;
  assign o[91] = t_6__91_ | 1'b0;
  assign o[90] = t_6__90_ | 1'b0;
  assign o[89] = t_6__89_ | 1'b0;
  assign o[88] = t_6__88_ | 1'b0;
  assign o[87] = t_6__87_ | 1'b0;
  assign o[86] = t_6__86_ | 1'b0;
  assign o[85] = t_6__85_ | 1'b0;
  assign o[84] = t_6__84_ | 1'b0;
  assign o[83] = t_6__83_ | 1'b0;
  assign o[82] = t_6__82_ | 1'b0;
  assign o[81] = t_6__81_ | 1'b0;
  assign o[80] = t_6__80_ | 1'b0;
  assign o[79] = t_6__79_ | 1'b0;
  assign o[78] = t_6__78_ | 1'b0;
  assign o[77] = t_6__77_ | 1'b0;
  assign o[76] = t_6__76_ | 1'b0;
  assign o[75] = t_6__75_ | 1'b0;
  assign o[74] = t_6__74_ | 1'b0;
  assign o[73] = t_6__73_ | 1'b0;
  assign o[72] = t_6__72_ | 1'b0;
  assign o[71] = t_6__71_ | 1'b0;
  assign o[70] = t_6__70_ | 1'b0;
  assign o[69] = t_6__69_ | 1'b0;
  assign o[68] = t_6__68_ | 1'b0;
  assign o[67] = t_6__67_ | 1'b0;
  assign o[66] = t_6__66_ | 1'b0;
  assign o[65] = t_6__65_ | 1'b0;
  assign o[64] = t_6__64_ | 1'b0;
  assign o[63] = t_6__63_ | t_6__127_;
  assign o[62] = t_6__62_ | t_6__126_;
  assign o[61] = t_6__61_ | t_6__125_;
  assign o[60] = t_6__60_ | t_6__124_;
  assign o[59] = t_6__59_ | t_6__123_;
  assign o[58] = t_6__58_ | t_6__122_;
  assign o[57] = t_6__57_ | t_6__121_;
  assign o[56] = t_6__56_ | t_6__120_;
  assign o[55] = t_6__55_ | t_6__119_;
  assign o[54] = t_6__54_ | t_6__118_;
  assign o[53] = t_6__53_ | t_6__117_;
  assign o[52] = t_6__52_ | t_6__116_;
  assign o[51] = t_6__51_ | t_6__115_;
  assign o[50] = t_6__50_ | t_6__114_;
  assign o[49] = t_6__49_ | t_6__113_;
  assign o[48] = t_6__48_ | t_6__112_;
  assign o[47] = t_6__47_ | t_6__111_;
  assign o[46] = t_6__46_ | t_6__110_;
  assign o[45] = t_6__45_ | t_6__109_;
  assign o[44] = t_6__44_ | t_6__108_;
  assign o[43] = t_6__43_ | t_6__107_;
  assign o[42] = t_6__42_ | t_6__106_;
  assign o[41] = t_6__41_ | t_6__105_;
  assign o[40] = t_6__40_ | t_6__104_;
  assign o[39] = t_6__39_ | t_6__103_;
  assign o[38] = t_6__38_ | t_6__102_;
  assign o[37] = t_6__37_ | t_6__101_;
  assign o[36] = t_6__36_ | t_6__100_;
  assign o[35] = t_6__35_ | t_6__99_;
  assign o[34] = t_6__34_ | t_6__98_;
  assign o[33] = t_6__33_ | t_6__97_;
  assign o[32] = t_6__32_ | t_6__96_;
  assign o[31] = t_6__31_ | t_6__95_;
  assign o[30] = t_6__30_ | t_6__94_;
  assign o[29] = t_6__29_ | t_6__93_;
  assign o[28] = t_6__28_ | t_6__92_;
  assign o[27] = t_6__27_ | t_6__91_;
  assign o[26] = t_6__26_ | t_6__90_;
  assign o[25] = t_6__25_ | t_6__89_;
  assign o[24] = t_6__24_ | t_6__88_;
  assign o[23] = t_6__23_ | t_6__87_;
  assign o[22] = t_6__22_ | t_6__86_;
  assign o[21] = t_6__21_ | t_6__85_;
  assign o[20] = t_6__20_ | t_6__84_;
  assign o[19] = t_6__19_ | t_6__83_;
  assign o[18] = t_6__18_ | t_6__82_;
  assign o[17] = t_6__17_ | t_6__81_;
  assign o[16] = t_6__16_ | t_6__80_;
  assign o[15] = t_6__15_ | t_6__79_;
  assign o[14] = t_6__14_ | t_6__78_;
  assign o[13] = t_6__13_ | t_6__77_;
  assign o[12] = t_6__12_ | t_6__76_;
  assign o[11] = t_6__11_ | t_6__75_;
  assign o[10] = t_6__10_ | t_6__74_;
  assign o[9] = t_6__9_ | t_6__73_;
  assign o[8] = t_6__8_ | t_6__72_;
  assign o[7] = t_6__7_ | t_6__71_;
  assign o[6] = t_6__6_ | t_6__70_;
  assign o[5] = t_6__5_ | t_6__69_;
  assign o[4] = t_6__4_ | t_6__68_;
  assign o[3] = t_6__3_ | t_6__67_;
  assign o[2] = t_6__2_ | t_6__66_;
  assign o[1] = t_6__1_ | t_6__65_;
  assign o[0] = t_6__0_ | t_6__64_;

endmodule



module bsg_priority_encode_one_hot_out_width_p128_lo_to_hi_p0
(
  i,
  o
);

  input [127:0] i;
  output [127:0] o;
  wire [127:0] o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126;
  wire [126:0] scan_lo;

  bsg_scan_width_p128_or_p1_lo_to_hi_p0
  genblk1_scan
  (
    .i(i),
    .o({ o[127:127], scan_lo })
  );

  assign o[126] = scan_lo[126] & N0;
  assign N0 = ~o[127];
  assign o[125] = scan_lo[125] & N1;
  assign N1 = ~scan_lo[126];
  assign o[124] = scan_lo[124] & N2;
  assign N2 = ~scan_lo[125];
  assign o[123] = scan_lo[123] & N3;
  assign N3 = ~scan_lo[124];
  assign o[122] = scan_lo[122] & N4;
  assign N4 = ~scan_lo[123];
  assign o[121] = scan_lo[121] & N5;
  assign N5 = ~scan_lo[122];
  assign o[120] = scan_lo[120] & N6;
  assign N6 = ~scan_lo[121];
  assign o[119] = scan_lo[119] & N7;
  assign N7 = ~scan_lo[120];
  assign o[118] = scan_lo[118] & N8;
  assign N8 = ~scan_lo[119];
  assign o[117] = scan_lo[117] & N9;
  assign N9 = ~scan_lo[118];
  assign o[116] = scan_lo[116] & N10;
  assign N10 = ~scan_lo[117];
  assign o[115] = scan_lo[115] & N11;
  assign N11 = ~scan_lo[116];
  assign o[114] = scan_lo[114] & N12;
  assign N12 = ~scan_lo[115];
  assign o[113] = scan_lo[113] & N13;
  assign N13 = ~scan_lo[114];
  assign o[112] = scan_lo[112] & N14;
  assign N14 = ~scan_lo[113];
  assign o[111] = scan_lo[111] & N15;
  assign N15 = ~scan_lo[112];
  assign o[110] = scan_lo[110] & N16;
  assign N16 = ~scan_lo[111];
  assign o[109] = scan_lo[109] & N17;
  assign N17 = ~scan_lo[110];
  assign o[108] = scan_lo[108] & N18;
  assign N18 = ~scan_lo[109];
  assign o[107] = scan_lo[107] & N19;
  assign N19 = ~scan_lo[108];
  assign o[106] = scan_lo[106] & N20;
  assign N20 = ~scan_lo[107];
  assign o[105] = scan_lo[105] & N21;
  assign N21 = ~scan_lo[106];
  assign o[104] = scan_lo[104] & N22;
  assign N22 = ~scan_lo[105];
  assign o[103] = scan_lo[103] & N23;
  assign N23 = ~scan_lo[104];
  assign o[102] = scan_lo[102] & N24;
  assign N24 = ~scan_lo[103];
  assign o[101] = scan_lo[101] & N25;
  assign N25 = ~scan_lo[102];
  assign o[100] = scan_lo[100] & N26;
  assign N26 = ~scan_lo[101];
  assign o[99] = scan_lo[99] & N27;
  assign N27 = ~scan_lo[100];
  assign o[98] = scan_lo[98] & N28;
  assign N28 = ~scan_lo[99];
  assign o[97] = scan_lo[97] & N29;
  assign N29 = ~scan_lo[98];
  assign o[96] = scan_lo[96] & N30;
  assign N30 = ~scan_lo[97];
  assign o[95] = scan_lo[95] & N31;
  assign N31 = ~scan_lo[96];
  assign o[94] = scan_lo[94] & N32;
  assign N32 = ~scan_lo[95];
  assign o[93] = scan_lo[93] & N33;
  assign N33 = ~scan_lo[94];
  assign o[92] = scan_lo[92] & N34;
  assign N34 = ~scan_lo[93];
  assign o[91] = scan_lo[91] & N35;
  assign N35 = ~scan_lo[92];
  assign o[90] = scan_lo[90] & N36;
  assign N36 = ~scan_lo[91];
  assign o[89] = scan_lo[89] & N37;
  assign N37 = ~scan_lo[90];
  assign o[88] = scan_lo[88] & N38;
  assign N38 = ~scan_lo[89];
  assign o[87] = scan_lo[87] & N39;
  assign N39 = ~scan_lo[88];
  assign o[86] = scan_lo[86] & N40;
  assign N40 = ~scan_lo[87];
  assign o[85] = scan_lo[85] & N41;
  assign N41 = ~scan_lo[86];
  assign o[84] = scan_lo[84] & N42;
  assign N42 = ~scan_lo[85];
  assign o[83] = scan_lo[83] & N43;
  assign N43 = ~scan_lo[84];
  assign o[82] = scan_lo[82] & N44;
  assign N44 = ~scan_lo[83];
  assign o[81] = scan_lo[81] & N45;
  assign N45 = ~scan_lo[82];
  assign o[80] = scan_lo[80] & N46;
  assign N46 = ~scan_lo[81];
  assign o[79] = scan_lo[79] & N47;
  assign N47 = ~scan_lo[80];
  assign o[78] = scan_lo[78] & N48;
  assign N48 = ~scan_lo[79];
  assign o[77] = scan_lo[77] & N49;
  assign N49 = ~scan_lo[78];
  assign o[76] = scan_lo[76] & N50;
  assign N50 = ~scan_lo[77];
  assign o[75] = scan_lo[75] & N51;
  assign N51 = ~scan_lo[76];
  assign o[74] = scan_lo[74] & N52;
  assign N52 = ~scan_lo[75];
  assign o[73] = scan_lo[73] & N53;
  assign N53 = ~scan_lo[74];
  assign o[72] = scan_lo[72] & N54;
  assign N54 = ~scan_lo[73];
  assign o[71] = scan_lo[71] & N55;
  assign N55 = ~scan_lo[72];
  assign o[70] = scan_lo[70] & N56;
  assign N56 = ~scan_lo[71];
  assign o[69] = scan_lo[69] & N57;
  assign N57 = ~scan_lo[70];
  assign o[68] = scan_lo[68] & N58;
  assign N58 = ~scan_lo[69];
  assign o[67] = scan_lo[67] & N59;
  assign N59 = ~scan_lo[68];
  assign o[66] = scan_lo[66] & N60;
  assign N60 = ~scan_lo[67];
  assign o[65] = scan_lo[65] & N61;
  assign N61 = ~scan_lo[66];
  assign o[64] = scan_lo[64] & N62;
  assign N62 = ~scan_lo[65];
  assign o[63] = scan_lo[63] & N63;
  assign N63 = ~scan_lo[64];
  assign o[62] = scan_lo[62] & N64;
  assign N64 = ~scan_lo[63];
  assign o[61] = scan_lo[61] & N65;
  assign N65 = ~scan_lo[62];
  assign o[60] = scan_lo[60] & N66;
  assign N66 = ~scan_lo[61];
  assign o[59] = scan_lo[59] & N67;
  assign N67 = ~scan_lo[60];
  assign o[58] = scan_lo[58] & N68;
  assign N68 = ~scan_lo[59];
  assign o[57] = scan_lo[57] & N69;
  assign N69 = ~scan_lo[58];
  assign o[56] = scan_lo[56] & N70;
  assign N70 = ~scan_lo[57];
  assign o[55] = scan_lo[55] & N71;
  assign N71 = ~scan_lo[56];
  assign o[54] = scan_lo[54] & N72;
  assign N72 = ~scan_lo[55];
  assign o[53] = scan_lo[53] & N73;
  assign N73 = ~scan_lo[54];
  assign o[52] = scan_lo[52] & N74;
  assign N74 = ~scan_lo[53];
  assign o[51] = scan_lo[51] & N75;
  assign N75 = ~scan_lo[52];
  assign o[50] = scan_lo[50] & N76;
  assign N76 = ~scan_lo[51];
  assign o[49] = scan_lo[49] & N77;
  assign N77 = ~scan_lo[50];
  assign o[48] = scan_lo[48] & N78;
  assign N78 = ~scan_lo[49];
  assign o[47] = scan_lo[47] & N79;
  assign N79 = ~scan_lo[48];
  assign o[46] = scan_lo[46] & N80;
  assign N80 = ~scan_lo[47];
  assign o[45] = scan_lo[45] & N81;
  assign N81 = ~scan_lo[46];
  assign o[44] = scan_lo[44] & N82;
  assign N82 = ~scan_lo[45];
  assign o[43] = scan_lo[43] & N83;
  assign N83 = ~scan_lo[44];
  assign o[42] = scan_lo[42] & N84;
  assign N84 = ~scan_lo[43];
  assign o[41] = scan_lo[41] & N85;
  assign N85 = ~scan_lo[42];
  assign o[40] = scan_lo[40] & N86;
  assign N86 = ~scan_lo[41];
  assign o[39] = scan_lo[39] & N87;
  assign N87 = ~scan_lo[40];
  assign o[38] = scan_lo[38] & N88;
  assign N88 = ~scan_lo[39];
  assign o[37] = scan_lo[37] & N89;
  assign N89 = ~scan_lo[38];
  assign o[36] = scan_lo[36] & N90;
  assign N90 = ~scan_lo[37];
  assign o[35] = scan_lo[35] & N91;
  assign N91 = ~scan_lo[36];
  assign o[34] = scan_lo[34] & N92;
  assign N92 = ~scan_lo[35];
  assign o[33] = scan_lo[33] & N93;
  assign N93 = ~scan_lo[34];
  assign o[32] = scan_lo[32] & N94;
  assign N94 = ~scan_lo[33];
  assign o[31] = scan_lo[31] & N95;
  assign N95 = ~scan_lo[32];
  assign o[30] = scan_lo[30] & N96;
  assign N96 = ~scan_lo[31];
  assign o[29] = scan_lo[29] & N97;
  assign N97 = ~scan_lo[30];
  assign o[28] = scan_lo[28] & N98;
  assign N98 = ~scan_lo[29];
  assign o[27] = scan_lo[27] & N99;
  assign N99 = ~scan_lo[28];
  assign o[26] = scan_lo[26] & N100;
  assign N100 = ~scan_lo[27];
  assign o[25] = scan_lo[25] & N101;
  assign N101 = ~scan_lo[26];
  assign o[24] = scan_lo[24] & N102;
  assign N102 = ~scan_lo[25];
  assign o[23] = scan_lo[23] & N103;
  assign N103 = ~scan_lo[24];
  assign o[22] = scan_lo[22] & N104;
  assign N104 = ~scan_lo[23];
  assign o[21] = scan_lo[21] & N105;
  assign N105 = ~scan_lo[22];
  assign o[20] = scan_lo[20] & N106;
  assign N106 = ~scan_lo[21];
  assign o[19] = scan_lo[19] & N107;
  assign N107 = ~scan_lo[20];
  assign o[18] = scan_lo[18] & N108;
  assign N108 = ~scan_lo[19];
  assign o[17] = scan_lo[17] & N109;
  assign N109 = ~scan_lo[18];
  assign o[16] = scan_lo[16] & N110;
  assign N110 = ~scan_lo[17];
  assign o[15] = scan_lo[15] & N111;
  assign N111 = ~scan_lo[16];
  assign o[14] = scan_lo[14] & N112;
  assign N112 = ~scan_lo[15];
  assign o[13] = scan_lo[13] & N113;
  assign N113 = ~scan_lo[14];
  assign o[12] = scan_lo[12] & N114;
  assign N114 = ~scan_lo[13];
  assign o[11] = scan_lo[11] & N115;
  assign N115 = ~scan_lo[12];
  assign o[10] = scan_lo[10] & N116;
  assign N116 = ~scan_lo[11];
  assign o[9] = scan_lo[9] & N117;
  assign N117 = ~scan_lo[10];
  assign o[8] = scan_lo[8] & N118;
  assign N118 = ~scan_lo[9];
  assign o[7] = scan_lo[7] & N119;
  assign N119 = ~scan_lo[8];
  assign o[6] = scan_lo[6] & N120;
  assign N120 = ~scan_lo[7];
  assign o[5] = scan_lo[5] & N121;
  assign N121 = ~scan_lo[6];
  assign o[4] = scan_lo[4] & N122;
  assign N122 = ~scan_lo[5];
  assign o[3] = scan_lo[3] & N123;
  assign N123 = ~scan_lo[4];
  assign o[2] = scan_lo[2] & N124;
  assign N124 = ~scan_lo[3];
  assign o[1] = scan_lo[1] & N125;
  assign N125 = ~scan_lo[2];
  assign o[0] = scan_lo[0] & N126;
  assign N126 = ~scan_lo[1];

endmodule



module bsg_arb_fixed_inputs_p128_lo_to_hi_p0
(
  ready_i,
  reqs_i,
  grants_o
);

  input [127:0] reqs_i;
  output [127:0] grants_o;
  input ready_i;
  wire [127:0] grants_o,grants_unmasked_lo;

  bsg_priority_encode_one_hot_out_width_p128_lo_to_hi_p0
  enc
  (
    .i(reqs_i),
    .o(grants_unmasked_lo)
  );

  assign grants_o[127] = grants_unmasked_lo[127] & ready_i;
  assign grants_o[126] = grants_unmasked_lo[126] & ready_i;
  assign grants_o[125] = grants_unmasked_lo[125] & ready_i;
  assign grants_o[124] = grants_unmasked_lo[124] & ready_i;
  assign grants_o[123] = grants_unmasked_lo[123] & ready_i;
  assign grants_o[122] = grants_unmasked_lo[122] & ready_i;
  assign grants_o[121] = grants_unmasked_lo[121] & ready_i;
  assign grants_o[120] = grants_unmasked_lo[120] & ready_i;
  assign grants_o[119] = grants_unmasked_lo[119] & ready_i;
  assign grants_o[118] = grants_unmasked_lo[118] & ready_i;
  assign grants_o[117] = grants_unmasked_lo[117] & ready_i;
  assign grants_o[116] = grants_unmasked_lo[116] & ready_i;
  assign grants_o[115] = grants_unmasked_lo[115] & ready_i;
  assign grants_o[114] = grants_unmasked_lo[114] & ready_i;
  assign grants_o[113] = grants_unmasked_lo[113] & ready_i;
  assign grants_o[112] = grants_unmasked_lo[112] & ready_i;
  assign grants_o[111] = grants_unmasked_lo[111] & ready_i;
  assign grants_o[110] = grants_unmasked_lo[110] & ready_i;
  assign grants_o[109] = grants_unmasked_lo[109] & ready_i;
  assign grants_o[108] = grants_unmasked_lo[108] & ready_i;
  assign grants_o[107] = grants_unmasked_lo[107] & ready_i;
  assign grants_o[106] = grants_unmasked_lo[106] & ready_i;
  assign grants_o[105] = grants_unmasked_lo[105] & ready_i;
  assign grants_o[104] = grants_unmasked_lo[104] & ready_i;
  assign grants_o[103] = grants_unmasked_lo[103] & ready_i;
  assign grants_o[102] = grants_unmasked_lo[102] & ready_i;
  assign grants_o[101] = grants_unmasked_lo[101] & ready_i;
  assign grants_o[100] = grants_unmasked_lo[100] & ready_i;
  assign grants_o[99] = grants_unmasked_lo[99] & ready_i;
  assign grants_o[98] = grants_unmasked_lo[98] & ready_i;
  assign grants_o[97] = grants_unmasked_lo[97] & ready_i;
  assign grants_o[96] = grants_unmasked_lo[96] & ready_i;
  assign grants_o[95] = grants_unmasked_lo[95] & ready_i;
  assign grants_o[94] = grants_unmasked_lo[94] & ready_i;
  assign grants_o[93] = grants_unmasked_lo[93] & ready_i;
  assign grants_o[92] = grants_unmasked_lo[92] & ready_i;
  assign grants_o[91] = grants_unmasked_lo[91] & ready_i;
  assign grants_o[90] = grants_unmasked_lo[90] & ready_i;
  assign grants_o[89] = grants_unmasked_lo[89] & ready_i;
  assign grants_o[88] = grants_unmasked_lo[88] & ready_i;
  assign grants_o[87] = grants_unmasked_lo[87] & ready_i;
  assign grants_o[86] = grants_unmasked_lo[86] & ready_i;
  assign grants_o[85] = grants_unmasked_lo[85] & ready_i;
  assign grants_o[84] = grants_unmasked_lo[84] & ready_i;
  assign grants_o[83] = grants_unmasked_lo[83] & ready_i;
  assign grants_o[82] = grants_unmasked_lo[82] & ready_i;
  assign grants_o[81] = grants_unmasked_lo[81] & ready_i;
  assign grants_o[80] = grants_unmasked_lo[80] & ready_i;
  assign grants_o[79] = grants_unmasked_lo[79] & ready_i;
  assign grants_o[78] = grants_unmasked_lo[78] & ready_i;
  assign grants_o[77] = grants_unmasked_lo[77] & ready_i;
  assign grants_o[76] = grants_unmasked_lo[76] & ready_i;
  assign grants_o[75] = grants_unmasked_lo[75] & ready_i;
  assign grants_o[74] = grants_unmasked_lo[74] & ready_i;
  assign grants_o[73] = grants_unmasked_lo[73] & ready_i;
  assign grants_o[72] = grants_unmasked_lo[72] & ready_i;
  assign grants_o[71] = grants_unmasked_lo[71] & ready_i;
  assign grants_o[70] = grants_unmasked_lo[70] & ready_i;
  assign grants_o[69] = grants_unmasked_lo[69] & ready_i;
  assign grants_o[68] = grants_unmasked_lo[68] & ready_i;
  assign grants_o[67] = grants_unmasked_lo[67] & ready_i;
  assign grants_o[66] = grants_unmasked_lo[66] & ready_i;
  assign grants_o[65] = grants_unmasked_lo[65] & ready_i;
  assign grants_o[64] = grants_unmasked_lo[64] & ready_i;
  assign grants_o[63] = grants_unmasked_lo[63] & ready_i;
  assign grants_o[62] = grants_unmasked_lo[62] & ready_i;
  assign grants_o[61] = grants_unmasked_lo[61] & ready_i;
  assign grants_o[60] = grants_unmasked_lo[60] & ready_i;
  assign grants_o[59] = grants_unmasked_lo[59] & ready_i;
  assign grants_o[58] = grants_unmasked_lo[58] & ready_i;
  assign grants_o[57] = grants_unmasked_lo[57] & ready_i;
  assign grants_o[56] = grants_unmasked_lo[56] & ready_i;
  assign grants_o[55] = grants_unmasked_lo[55] & ready_i;
  assign grants_o[54] = grants_unmasked_lo[54] & ready_i;
  assign grants_o[53] = grants_unmasked_lo[53] & ready_i;
  assign grants_o[52] = grants_unmasked_lo[52] & ready_i;
  assign grants_o[51] = grants_unmasked_lo[51] & ready_i;
  assign grants_o[50] = grants_unmasked_lo[50] & ready_i;
  assign grants_o[49] = grants_unmasked_lo[49] & ready_i;
  assign grants_o[48] = grants_unmasked_lo[48] & ready_i;
  assign grants_o[47] = grants_unmasked_lo[47] & ready_i;
  assign grants_o[46] = grants_unmasked_lo[46] & ready_i;
  assign grants_o[45] = grants_unmasked_lo[45] & ready_i;
  assign grants_o[44] = grants_unmasked_lo[44] & ready_i;
  assign grants_o[43] = grants_unmasked_lo[43] & ready_i;
  assign grants_o[42] = grants_unmasked_lo[42] & ready_i;
  assign grants_o[41] = grants_unmasked_lo[41] & ready_i;
  assign grants_o[40] = grants_unmasked_lo[40] & ready_i;
  assign grants_o[39] = grants_unmasked_lo[39] & ready_i;
  assign grants_o[38] = grants_unmasked_lo[38] & ready_i;
  assign grants_o[37] = grants_unmasked_lo[37] & ready_i;
  assign grants_o[36] = grants_unmasked_lo[36] & ready_i;
  assign grants_o[35] = grants_unmasked_lo[35] & ready_i;
  assign grants_o[34] = grants_unmasked_lo[34] & ready_i;
  assign grants_o[33] = grants_unmasked_lo[33] & ready_i;
  assign grants_o[32] = grants_unmasked_lo[32] & ready_i;
  assign grants_o[31] = grants_unmasked_lo[31] & ready_i;
  assign grants_o[30] = grants_unmasked_lo[30] & ready_i;
  assign grants_o[29] = grants_unmasked_lo[29] & ready_i;
  assign grants_o[28] = grants_unmasked_lo[28] & ready_i;
  assign grants_o[27] = grants_unmasked_lo[27] & ready_i;
  assign grants_o[26] = grants_unmasked_lo[26] & ready_i;
  assign grants_o[25] = grants_unmasked_lo[25] & ready_i;
  assign grants_o[24] = grants_unmasked_lo[24] & ready_i;
  assign grants_o[23] = grants_unmasked_lo[23] & ready_i;
  assign grants_o[22] = grants_unmasked_lo[22] & ready_i;
  assign grants_o[21] = grants_unmasked_lo[21] & ready_i;
  assign grants_o[20] = grants_unmasked_lo[20] & ready_i;
  assign grants_o[19] = grants_unmasked_lo[19] & ready_i;
  assign grants_o[18] = grants_unmasked_lo[18] & ready_i;
  assign grants_o[17] = grants_unmasked_lo[17] & ready_i;
  assign grants_o[16] = grants_unmasked_lo[16] & ready_i;
  assign grants_o[15] = grants_unmasked_lo[15] & ready_i;
  assign grants_o[14] = grants_unmasked_lo[14] & ready_i;
  assign grants_o[13] = grants_unmasked_lo[13] & ready_i;
  assign grants_o[12] = grants_unmasked_lo[12] & ready_i;
  assign grants_o[11] = grants_unmasked_lo[11] & ready_i;
  assign grants_o[10] = grants_unmasked_lo[10] & ready_i;
  assign grants_o[9] = grants_unmasked_lo[9] & ready_i;
  assign grants_o[8] = grants_unmasked_lo[8] & ready_i;
  assign grants_o[7] = grants_unmasked_lo[7] & ready_i;
  assign grants_o[6] = grants_unmasked_lo[6] & ready_i;
  assign grants_o[5] = grants_unmasked_lo[5] & ready_i;
  assign grants_o[4] = grants_unmasked_lo[4] & ready_i;
  assign grants_o[3] = grants_unmasked_lo[3] & ready_i;
  assign grants_o[2] = grants_unmasked_lo[2] & ready_i;
  assign grants_o[1] = grants_unmasked_lo[1] & ready_i;
  assign grants_o[0] = grants_unmasked_lo[0] & ready_i;

endmodule



module bsg_locking_arb_fixed
(
  clk_i,
  ready_i,
  unlock_i,
  reqs_i,
  grants_o
);

  input [127:0] reqs_i;
  output [127:0] grants_o;
  input clk_i;
  input ready_i;
  input unlock_i;
  wire [127:0] grants_o,not_req_mask_r,req_mask_r;
  wire n_0_net_,n_1_net__127_,n_1_net__126_,n_1_net__125_,n_1_net__124_,n_1_net__123_,
  n_1_net__122_,n_1_net__121_,n_1_net__120_,n_1_net__119_,n_1_net__118_,
  n_1_net__117_,n_1_net__116_,n_1_net__115_,n_1_net__114_,n_1_net__113_,n_1_net__112_,
  n_1_net__111_,n_1_net__110_,n_1_net__109_,n_1_net__108_,n_1_net__107_,n_1_net__106_,
  n_1_net__105_,n_1_net__104_,n_1_net__103_,n_1_net__102_,n_1_net__101_,
  n_1_net__100_,n_1_net__99_,n_1_net__98_,n_1_net__97_,n_1_net__96_,n_1_net__95_,n_1_net__94_,
  n_1_net__93_,n_1_net__92_,n_1_net__91_,n_1_net__90_,n_1_net__89_,n_1_net__88_,
  n_1_net__87_,n_1_net__86_,n_1_net__85_,n_1_net__84_,n_1_net__83_,n_1_net__82_,
  n_1_net__81_,n_1_net__80_,n_1_net__79_,n_1_net__78_,n_1_net__77_,n_1_net__76_,
  n_1_net__75_,n_1_net__74_,n_1_net__73_,n_1_net__72_,n_1_net__71_,n_1_net__70_,
  n_1_net__69_,n_1_net__68_,n_1_net__67_,n_1_net__66_,n_1_net__65_,n_1_net__64_,
  n_1_net__63_,n_1_net__62_,n_1_net__61_,n_1_net__60_,n_1_net__59_,n_1_net__58_,n_1_net__57_,
  n_1_net__56_,n_1_net__55_,n_1_net__54_,n_1_net__53_,n_1_net__52_,n_1_net__51_,
  n_1_net__50_,n_1_net__49_,n_1_net__48_,n_1_net__47_,n_1_net__46_,n_1_net__45_,
  n_1_net__44_,n_1_net__43_,n_1_net__42_,n_1_net__41_,n_1_net__40_,n_1_net__39_,
  n_1_net__38_,n_1_net__37_,n_1_net__36_,n_1_net__35_,n_1_net__34_,n_1_net__33_,
  n_1_net__32_,n_1_net__31_,n_1_net__30_,n_1_net__29_,n_1_net__28_,n_1_net__27_,
  n_1_net__26_,n_1_net__25_,n_1_net__24_,n_1_net__23_,n_1_net__22_,n_1_net__21_,
  n_1_net__20_,n_1_net__19_,n_1_net__18_,n_1_net__17_,n_1_net__16_,n_1_net__15_,n_1_net__14_,
  n_1_net__13_,n_1_net__12_,n_1_net__11_,n_1_net__10_,n_1_net__9_,n_1_net__8_,
  n_1_net__7_,n_1_net__6_,n_1_net__5_,n_1_net__4_,n_1_net__3_,n_1_net__2_,n_1_net__1_,
  n_1_net__0_,n_2_net__127_,n_2_net__126_,n_2_net__125_,n_2_net__124_,
  n_2_net__123_,n_2_net__122_,n_2_net__121_,n_2_net__120_,n_2_net__119_,n_2_net__118_,
  n_2_net__117_,n_2_net__116_,n_2_net__115_,n_2_net__114_,n_2_net__113_,n_2_net__112_,
  n_2_net__111_,n_2_net__110_,n_2_net__109_,n_2_net__108_,n_2_net__107_,n_2_net__106_,
  n_2_net__105_,n_2_net__104_,n_2_net__103_,n_2_net__102_,n_2_net__101_,
  n_2_net__100_,n_2_net__99_,n_2_net__98_,n_2_net__97_,n_2_net__96_,n_2_net__95_,
  n_2_net__94_,n_2_net__93_,n_2_net__92_,n_2_net__91_,n_2_net__90_,n_2_net__89_,n_2_net__88_,
  n_2_net__87_,n_2_net__86_,n_2_net__85_,n_2_net__84_,n_2_net__83_,n_2_net__82_,
  n_2_net__81_,n_2_net__80_,n_2_net__79_,n_2_net__78_,n_2_net__77_,n_2_net__76_,
  n_2_net__75_,n_2_net__74_,n_2_net__73_,n_2_net__72_,n_2_net__71_,n_2_net__70_,
  n_2_net__69_,n_2_net__68_,n_2_net__67_,n_2_net__66_,n_2_net__65_,n_2_net__64_,
  n_2_net__63_,n_2_net__62_,n_2_net__61_,n_2_net__60_,n_2_net__59_,n_2_net__58_,
  n_2_net__57_,n_2_net__56_,n_2_net__55_,n_2_net__54_,n_2_net__53_,n_2_net__52_,n_2_net__51_,
  n_2_net__50_,n_2_net__49_,n_2_net__48_,n_2_net__47_,n_2_net__46_,n_2_net__45_,
  n_2_net__44_,n_2_net__43_,n_2_net__42_,n_2_net__41_,n_2_net__40_,n_2_net__39_,
  n_2_net__38_,n_2_net__37_,n_2_net__36_,n_2_net__35_,n_2_net__34_,n_2_net__33_,
  n_2_net__32_,n_2_net__31_,n_2_net__30_,n_2_net__29_,n_2_net__28_,n_2_net__27_,
  n_2_net__26_,n_2_net__25_,n_2_net__24_,n_2_net__23_,n_2_net__22_,n_2_net__21_,
  n_2_net__20_,n_2_net__19_,n_2_net__18_,n_2_net__17_,n_2_net__16_,n_2_net__15_,
  n_2_net__14_,n_2_net__13_,n_2_net__12_,n_2_net__11_,n_2_net__10_,n_2_net__9_,n_2_net__8_,
  n_2_net__7_,n_2_net__6_,n_2_net__5_,n_2_net__4_,n_2_net__3_,n_2_net__2_,
  n_2_net__1_,n_2_net__0_,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,
  N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,
  N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,
  N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,
  N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,
  N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,
  N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
  N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,
  N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253;

  bsg_dff_reset_en_width_p128
  req_words_reg
  (
    .clk_i(clk_i),
    .reset_i(unlock_i),
    .en_i(n_0_net_),
    .data_i({ n_1_net__127_, n_1_net__126_, n_1_net__125_, n_1_net__124_, n_1_net__123_, n_1_net__122_, n_1_net__121_, n_1_net__120_, n_1_net__119_, n_1_net__118_, n_1_net__117_, n_1_net__116_, n_1_net__115_, n_1_net__114_, n_1_net__113_, n_1_net__112_, n_1_net__111_, n_1_net__110_, n_1_net__109_, n_1_net__108_, n_1_net__107_, n_1_net__106_, n_1_net__105_, n_1_net__104_, n_1_net__103_, n_1_net__102_, n_1_net__101_, n_1_net__100_, n_1_net__99_, n_1_net__98_, n_1_net__97_, n_1_net__96_, n_1_net__95_, n_1_net__94_, n_1_net__93_, n_1_net__92_, n_1_net__91_, n_1_net__90_, n_1_net__89_, n_1_net__88_, n_1_net__87_, n_1_net__86_, n_1_net__85_, n_1_net__84_, n_1_net__83_, n_1_net__82_, n_1_net__81_, n_1_net__80_, n_1_net__79_, n_1_net__78_, n_1_net__77_, n_1_net__76_, n_1_net__75_, n_1_net__74_, n_1_net__73_, n_1_net__72_, n_1_net__71_, n_1_net__70_, n_1_net__69_, n_1_net__68_, n_1_net__67_, n_1_net__66_, n_1_net__65_, n_1_net__64_, n_1_net__63_, n_1_net__62_, n_1_net__61_, n_1_net__60_, n_1_net__59_, n_1_net__58_, n_1_net__57_, n_1_net__56_, n_1_net__55_, n_1_net__54_, n_1_net__53_, n_1_net__52_, n_1_net__51_, n_1_net__50_, n_1_net__49_, n_1_net__48_, n_1_net__47_, n_1_net__46_, n_1_net__45_, n_1_net__44_, n_1_net__43_, n_1_net__42_, n_1_net__41_, n_1_net__40_, n_1_net__39_, n_1_net__38_, n_1_net__37_, n_1_net__36_, n_1_net__35_, n_1_net__34_, n_1_net__33_, n_1_net__32_, n_1_net__31_, n_1_net__30_, n_1_net__29_, n_1_net__28_, n_1_net__27_, n_1_net__26_, n_1_net__25_, n_1_net__24_, n_1_net__23_, n_1_net__22_, n_1_net__21_, n_1_net__20_, n_1_net__19_, n_1_net__18_, n_1_net__17_, n_1_net__16_, n_1_net__15_, n_1_net__14_, n_1_net__13_, n_1_net__12_, n_1_net__11_, n_1_net__10_, n_1_net__9_, n_1_net__8_, n_1_net__7_, n_1_net__6_, n_1_net__5_, n_1_net__4_, n_1_net__3_, n_1_net__2_, n_1_net__1_, n_1_net__0_ }),
    .data_o(not_req_mask_r)
  );


  bsg_arb_fixed_inputs_p128_lo_to_hi_p0
  fixed_arb
  (
    .ready_i(ready_i),
    .reqs_i({ n_2_net__127_, n_2_net__126_, n_2_net__125_, n_2_net__124_, n_2_net__123_, n_2_net__122_, n_2_net__121_, n_2_net__120_, n_2_net__119_, n_2_net__118_, n_2_net__117_, n_2_net__116_, n_2_net__115_, n_2_net__114_, n_2_net__113_, n_2_net__112_, n_2_net__111_, n_2_net__110_, n_2_net__109_, n_2_net__108_, n_2_net__107_, n_2_net__106_, n_2_net__105_, n_2_net__104_, n_2_net__103_, n_2_net__102_, n_2_net__101_, n_2_net__100_, n_2_net__99_, n_2_net__98_, n_2_net__97_, n_2_net__96_, n_2_net__95_, n_2_net__94_, n_2_net__93_, n_2_net__92_, n_2_net__91_, n_2_net__90_, n_2_net__89_, n_2_net__88_, n_2_net__87_, n_2_net__86_, n_2_net__85_, n_2_net__84_, n_2_net__83_, n_2_net__82_, n_2_net__81_, n_2_net__80_, n_2_net__79_, n_2_net__78_, n_2_net__77_, n_2_net__76_, n_2_net__75_, n_2_net__74_, n_2_net__73_, n_2_net__72_, n_2_net__71_, n_2_net__70_, n_2_net__69_, n_2_net__68_, n_2_net__67_, n_2_net__66_, n_2_net__65_, n_2_net__64_, n_2_net__63_, n_2_net__62_, n_2_net__61_, n_2_net__60_, n_2_net__59_, n_2_net__58_, n_2_net__57_, n_2_net__56_, n_2_net__55_, n_2_net__54_, n_2_net__53_, n_2_net__52_, n_2_net__51_, n_2_net__50_, n_2_net__49_, n_2_net__48_, n_2_net__47_, n_2_net__46_, n_2_net__45_, n_2_net__44_, n_2_net__43_, n_2_net__42_, n_2_net__41_, n_2_net__40_, n_2_net__39_, n_2_net__38_, n_2_net__37_, n_2_net__36_, n_2_net__35_, n_2_net__34_, n_2_net__33_, n_2_net__32_, n_2_net__31_, n_2_net__30_, n_2_net__29_, n_2_net__28_, n_2_net__27_, n_2_net__26_, n_2_net__25_, n_2_net__24_, n_2_net__23_, n_2_net__22_, n_2_net__21_, n_2_net__20_, n_2_net__19_, n_2_net__18_, n_2_net__17_, n_2_net__16_, n_2_net__15_, n_2_net__14_, n_2_net__13_, n_2_net__12_, n_2_net__11_, n_2_net__10_, n_2_net__9_, n_2_net__8_, n_2_net__7_, n_2_net__6_, n_2_net__5_, n_2_net__4_, n_2_net__3_, n_2_net__2_, n_2_net__1_, n_2_net__0_ }),
    .grants_o(grants_o)
  );

  assign n_1_net__127_ = ~grants_o[127];
  assign n_1_net__126_ = ~grants_o[126];
  assign n_1_net__125_ = ~grants_o[125];
  assign n_1_net__124_ = ~grants_o[124];
  assign n_1_net__123_ = ~grants_o[123];
  assign n_1_net__122_ = ~grants_o[122];
  assign n_1_net__121_ = ~grants_o[121];
  assign n_1_net__120_ = ~grants_o[120];
  assign n_1_net__119_ = ~grants_o[119];
  assign n_1_net__118_ = ~grants_o[118];
  assign n_1_net__117_ = ~grants_o[117];
  assign n_1_net__116_ = ~grants_o[116];
  assign n_1_net__115_ = ~grants_o[115];
  assign n_1_net__114_ = ~grants_o[114];
  assign n_1_net__113_ = ~grants_o[113];
  assign n_1_net__112_ = ~grants_o[112];
  assign n_1_net__111_ = ~grants_o[111];
  assign n_1_net__110_ = ~grants_o[110];
  assign n_1_net__109_ = ~grants_o[109];
  assign n_1_net__108_ = ~grants_o[108];
  assign n_1_net__107_ = ~grants_o[107];
  assign n_1_net__106_ = ~grants_o[106];
  assign n_1_net__105_ = ~grants_o[105];
  assign n_1_net__104_ = ~grants_o[104];
  assign n_1_net__103_ = ~grants_o[103];
  assign n_1_net__102_ = ~grants_o[102];
  assign n_1_net__101_ = ~grants_o[101];
  assign n_1_net__100_ = ~grants_o[100];
  assign n_1_net__99_ = ~grants_o[99];
  assign n_1_net__98_ = ~grants_o[98];
  assign n_1_net__97_ = ~grants_o[97];
  assign n_1_net__96_ = ~grants_o[96];
  assign n_1_net__95_ = ~grants_o[95];
  assign n_1_net__94_ = ~grants_o[94];
  assign n_1_net__93_ = ~grants_o[93];
  assign n_1_net__92_ = ~grants_o[92];
  assign n_1_net__91_ = ~grants_o[91];
  assign n_1_net__90_ = ~grants_o[90];
  assign n_1_net__89_ = ~grants_o[89];
  assign n_1_net__88_ = ~grants_o[88];
  assign n_1_net__87_ = ~grants_o[87];
  assign n_1_net__86_ = ~grants_o[86];
  assign n_1_net__85_ = ~grants_o[85];
  assign n_1_net__84_ = ~grants_o[84];
  assign n_1_net__83_ = ~grants_o[83];
  assign n_1_net__82_ = ~grants_o[82];
  assign n_1_net__81_ = ~grants_o[81];
  assign n_1_net__80_ = ~grants_o[80];
  assign n_1_net__79_ = ~grants_o[79];
  assign n_1_net__78_ = ~grants_o[78];
  assign n_1_net__77_ = ~grants_o[77];
  assign n_1_net__76_ = ~grants_o[76];
  assign n_1_net__75_ = ~grants_o[75];
  assign n_1_net__74_ = ~grants_o[74];
  assign n_1_net__73_ = ~grants_o[73];
  assign n_1_net__72_ = ~grants_o[72];
  assign n_1_net__71_ = ~grants_o[71];
  assign n_1_net__70_ = ~grants_o[70];
  assign n_1_net__69_ = ~grants_o[69];
  assign n_1_net__68_ = ~grants_o[68];
  assign n_1_net__67_ = ~grants_o[67];
  assign n_1_net__66_ = ~grants_o[66];
  assign n_1_net__65_ = ~grants_o[65];
  assign n_1_net__64_ = ~grants_o[64];
  assign n_1_net__63_ = ~grants_o[63];
  assign n_1_net__62_ = ~grants_o[62];
  assign n_1_net__61_ = ~grants_o[61];
  assign n_1_net__60_ = ~grants_o[60];
  assign n_1_net__59_ = ~grants_o[59];
  assign n_1_net__58_ = ~grants_o[58];
  assign n_1_net__57_ = ~grants_o[57];
  assign n_1_net__56_ = ~grants_o[56];
  assign n_1_net__55_ = ~grants_o[55];
  assign n_1_net__54_ = ~grants_o[54];
  assign n_1_net__53_ = ~grants_o[53];
  assign n_1_net__52_ = ~grants_o[52];
  assign n_1_net__51_ = ~grants_o[51];
  assign n_1_net__50_ = ~grants_o[50];
  assign n_1_net__49_ = ~grants_o[49];
  assign n_1_net__48_ = ~grants_o[48];
  assign n_1_net__47_ = ~grants_o[47];
  assign n_1_net__46_ = ~grants_o[46];
  assign n_1_net__45_ = ~grants_o[45];
  assign n_1_net__44_ = ~grants_o[44];
  assign n_1_net__43_ = ~grants_o[43];
  assign n_1_net__42_ = ~grants_o[42];
  assign n_1_net__41_ = ~grants_o[41];
  assign n_1_net__40_ = ~grants_o[40];
  assign n_1_net__39_ = ~grants_o[39];
  assign n_1_net__38_ = ~grants_o[38];
  assign n_1_net__37_ = ~grants_o[37];
  assign n_1_net__36_ = ~grants_o[36];
  assign n_1_net__35_ = ~grants_o[35];
  assign n_1_net__34_ = ~grants_o[34];
  assign n_1_net__33_ = ~grants_o[33];
  assign n_1_net__32_ = ~grants_o[32];
  assign n_1_net__31_ = ~grants_o[31];
  assign n_1_net__30_ = ~grants_o[30];
  assign n_1_net__29_ = ~grants_o[29];
  assign n_1_net__28_ = ~grants_o[28];
  assign n_1_net__27_ = ~grants_o[27];
  assign n_1_net__26_ = ~grants_o[26];
  assign n_1_net__25_ = ~grants_o[25];
  assign n_1_net__24_ = ~grants_o[24];
  assign n_1_net__23_ = ~grants_o[23];
  assign n_1_net__22_ = ~grants_o[22];
  assign n_1_net__21_ = ~grants_o[21];
  assign n_1_net__20_ = ~grants_o[20];
  assign n_1_net__19_ = ~grants_o[19];
  assign n_1_net__18_ = ~grants_o[18];
  assign n_1_net__17_ = ~grants_o[17];
  assign n_1_net__16_ = ~grants_o[16];
  assign n_1_net__15_ = ~grants_o[15];
  assign n_1_net__14_ = ~grants_o[14];
  assign n_1_net__13_ = ~grants_o[13];
  assign n_1_net__12_ = ~grants_o[12];
  assign n_1_net__11_ = ~grants_o[11];
  assign n_1_net__10_ = ~grants_o[10];
  assign n_1_net__9_ = ~grants_o[9];
  assign n_1_net__8_ = ~grants_o[8];
  assign n_1_net__7_ = ~grants_o[7];
  assign n_1_net__6_ = ~grants_o[6];
  assign n_1_net__5_ = ~grants_o[5];
  assign n_1_net__4_ = ~grants_o[4];
  assign n_1_net__3_ = ~grants_o[3];
  assign n_1_net__2_ = ~grants_o[2];
  assign n_1_net__1_ = ~grants_o[1];
  assign n_1_net__0_ = ~grants_o[0];
  assign n_0_net_ = N126 & N253;
  assign N126 = N125 & req_mask_r[0];
  assign N125 = N124 & req_mask_r[1];
  assign N124 = N123 & req_mask_r[2];
  assign N123 = N122 & req_mask_r[3];
  assign N122 = N121 & req_mask_r[4];
  assign N121 = N120 & req_mask_r[5];
  assign N120 = N119 & req_mask_r[6];
  assign N119 = N118 & req_mask_r[7];
  assign N118 = N117 & req_mask_r[8];
  assign N117 = N116 & req_mask_r[9];
  assign N116 = N115 & req_mask_r[10];
  assign N115 = N114 & req_mask_r[11];
  assign N114 = N113 & req_mask_r[12];
  assign N113 = N112 & req_mask_r[13];
  assign N112 = N111 & req_mask_r[14];
  assign N111 = N110 & req_mask_r[15];
  assign N110 = N109 & req_mask_r[16];
  assign N109 = N108 & req_mask_r[17];
  assign N108 = N107 & req_mask_r[18];
  assign N107 = N106 & req_mask_r[19];
  assign N106 = N105 & req_mask_r[20];
  assign N105 = N104 & req_mask_r[21];
  assign N104 = N103 & req_mask_r[22];
  assign N103 = N102 & req_mask_r[23];
  assign N102 = N101 & req_mask_r[24];
  assign N101 = N100 & req_mask_r[25];
  assign N100 = N99 & req_mask_r[26];
  assign N99 = N98 & req_mask_r[27];
  assign N98 = N97 & req_mask_r[28];
  assign N97 = N96 & req_mask_r[29];
  assign N96 = N95 & req_mask_r[30];
  assign N95 = N94 & req_mask_r[31];
  assign N94 = N93 & req_mask_r[32];
  assign N93 = N92 & req_mask_r[33];
  assign N92 = N91 & req_mask_r[34];
  assign N91 = N90 & req_mask_r[35];
  assign N90 = N89 & req_mask_r[36];
  assign N89 = N88 & req_mask_r[37];
  assign N88 = N87 & req_mask_r[38];
  assign N87 = N86 & req_mask_r[39];
  assign N86 = N85 & req_mask_r[40];
  assign N85 = N84 & req_mask_r[41];
  assign N84 = N83 & req_mask_r[42];
  assign N83 = N82 & req_mask_r[43];
  assign N82 = N81 & req_mask_r[44];
  assign N81 = N80 & req_mask_r[45];
  assign N80 = N79 & req_mask_r[46];
  assign N79 = N78 & req_mask_r[47];
  assign N78 = N77 & req_mask_r[48];
  assign N77 = N76 & req_mask_r[49];
  assign N76 = N75 & req_mask_r[50];
  assign N75 = N74 & req_mask_r[51];
  assign N74 = N73 & req_mask_r[52];
  assign N73 = N72 & req_mask_r[53];
  assign N72 = N71 & req_mask_r[54];
  assign N71 = N70 & req_mask_r[55];
  assign N70 = N69 & req_mask_r[56];
  assign N69 = N68 & req_mask_r[57];
  assign N68 = N67 & req_mask_r[58];
  assign N67 = N66 & req_mask_r[59];
  assign N66 = N65 & req_mask_r[60];
  assign N65 = N64 & req_mask_r[61];
  assign N64 = N63 & req_mask_r[62];
  assign N63 = N62 & req_mask_r[63];
  assign N62 = N61 & req_mask_r[64];
  assign N61 = N60 & req_mask_r[65];
  assign N60 = N59 & req_mask_r[66];
  assign N59 = N58 & req_mask_r[67];
  assign N58 = N57 & req_mask_r[68];
  assign N57 = N56 & req_mask_r[69];
  assign N56 = N55 & req_mask_r[70];
  assign N55 = N54 & req_mask_r[71];
  assign N54 = N53 & req_mask_r[72];
  assign N53 = N52 & req_mask_r[73];
  assign N52 = N51 & req_mask_r[74];
  assign N51 = N50 & req_mask_r[75];
  assign N50 = N49 & req_mask_r[76];
  assign N49 = N48 & req_mask_r[77];
  assign N48 = N47 & req_mask_r[78];
  assign N47 = N46 & req_mask_r[79];
  assign N46 = N45 & req_mask_r[80];
  assign N45 = N44 & req_mask_r[81];
  assign N44 = N43 & req_mask_r[82];
  assign N43 = N42 & req_mask_r[83];
  assign N42 = N41 & req_mask_r[84];
  assign N41 = N40 & req_mask_r[85];
  assign N40 = N39 & req_mask_r[86];
  assign N39 = N38 & req_mask_r[87];
  assign N38 = N37 & req_mask_r[88];
  assign N37 = N36 & req_mask_r[89];
  assign N36 = N35 & req_mask_r[90];
  assign N35 = N34 & req_mask_r[91];
  assign N34 = N33 & req_mask_r[92];
  assign N33 = N32 & req_mask_r[93];
  assign N32 = N31 & req_mask_r[94];
  assign N31 = N30 & req_mask_r[95];
  assign N30 = N29 & req_mask_r[96];
  assign N29 = N28 & req_mask_r[97];
  assign N28 = N27 & req_mask_r[98];
  assign N27 = N26 & req_mask_r[99];
  assign N26 = N25 & req_mask_r[100];
  assign N25 = N24 & req_mask_r[101];
  assign N24 = N23 & req_mask_r[102];
  assign N23 = N22 & req_mask_r[103];
  assign N22 = N21 & req_mask_r[104];
  assign N21 = N20 & req_mask_r[105];
  assign N20 = N19 & req_mask_r[106];
  assign N19 = N18 & req_mask_r[107];
  assign N18 = N17 & req_mask_r[108];
  assign N17 = N16 & req_mask_r[109];
  assign N16 = N15 & req_mask_r[110];
  assign N15 = N14 & req_mask_r[111];
  assign N14 = N13 & req_mask_r[112];
  assign N13 = N12 & req_mask_r[113];
  assign N12 = N11 & req_mask_r[114];
  assign N11 = N10 & req_mask_r[115];
  assign N10 = N9 & req_mask_r[116];
  assign N9 = N8 & req_mask_r[117];
  assign N8 = N7 & req_mask_r[118];
  assign N7 = N6 & req_mask_r[119];
  assign N6 = N5 & req_mask_r[120];
  assign N5 = N4 & req_mask_r[121];
  assign N4 = N3 & req_mask_r[122];
  assign N3 = N2 & req_mask_r[123];
  assign N2 = N1 & req_mask_r[124];
  assign N1 = N0 & req_mask_r[125];
  assign N0 = req_mask_r[127] & req_mask_r[126];
  assign N253 = N252 | grants_o[0];
  assign N252 = N251 | grants_o[1];
  assign N251 = N250 | grants_o[2];
  assign N250 = N249 | grants_o[3];
  assign N249 = N248 | grants_o[4];
  assign N248 = N247 | grants_o[5];
  assign N247 = N246 | grants_o[6];
  assign N246 = N245 | grants_o[7];
  assign N245 = N244 | grants_o[8];
  assign N244 = N243 | grants_o[9];
  assign N243 = N242 | grants_o[10];
  assign N242 = N241 | grants_o[11];
  assign N241 = N240 | grants_o[12];
  assign N240 = N239 | grants_o[13];
  assign N239 = N238 | grants_o[14];
  assign N238 = N237 | grants_o[15];
  assign N237 = N236 | grants_o[16];
  assign N236 = N235 | grants_o[17];
  assign N235 = N234 | grants_o[18];
  assign N234 = N233 | grants_o[19];
  assign N233 = N232 | grants_o[20];
  assign N232 = N231 | grants_o[21];
  assign N231 = N230 | grants_o[22];
  assign N230 = N229 | grants_o[23];
  assign N229 = N228 | grants_o[24];
  assign N228 = N227 | grants_o[25];
  assign N227 = N226 | grants_o[26];
  assign N226 = N225 | grants_o[27];
  assign N225 = N224 | grants_o[28];
  assign N224 = N223 | grants_o[29];
  assign N223 = N222 | grants_o[30];
  assign N222 = N221 | grants_o[31];
  assign N221 = N220 | grants_o[32];
  assign N220 = N219 | grants_o[33];
  assign N219 = N218 | grants_o[34];
  assign N218 = N217 | grants_o[35];
  assign N217 = N216 | grants_o[36];
  assign N216 = N215 | grants_o[37];
  assign N215 = N214 | grants_o[38];
  assign N214 = N213 | grants_o[39];
  assign N213 = N212 | grants_o[40];
  assign N212 = N211 | grants_o[41];
  assign N211 = N210 | grants_o[42];
  assign N210 = N209 | grants_o[43];
  assign N209 = N208 | grants_o[44];
  assign N208 = N207 | grants_o[45];
  assign N207 = N206 | grants_o[46];
  assign N206 = N205 | grants_o[47];
  assign N205 = N204 | grants_o[48];
  assign N204 = N203 | grants_o[49];
  assign N203 = N202 | grants_o[50];
  assign N202 = N201 | grants_o[51];
  assign N201 = N200 | grants_o[52];
  assign N200 = N199 | grants_o[53];
  assign N199 = N198 | grants_o[54];
  assign N198 = N197 | grants_o[55];
  assign N197 = N196 | grants_o[56];
  assign N196 = N195 | grants_o[57];
  assign N195 = N194 | grants_o[58];
  assign N194 = N193 | grants_o[59];
  assign N193 = N192 | grants_o[60];
  assign N192 = N191 | grants_o[61];
  assign N191 = N190 | grants_o[62];
  assign N190 = N189 | grants_o[63];
  assign N189 = N188 | grants_o[64];
  assign N188 = N187 | grants_o[65];
  assign N187 = N186 | grants_o[66];
  assign N186 = N185 | grants_o[67];
  assign N185 = N184 | grants_o[68];
  assign N184 = N183 | grants_o[69];
  assign N183 = N182 | grants_o[70];
  assign N182 = N181 | grants_o[71];
  assign N181 = N180 | grants_o[72];
  assign N180 = N179 | grants_o[73];
  assign N179 = N178 | grants_o[74];
  assign N178 = N177 | grants_o[75];
  assign N177 = N176 | grants_o[76];
  assign N176 = N175 | grants_o[77];
  assign N175 = N174 | grants_o[78];
  assign N174 = N173 | grants_o[79];
  assign N173 = N172 | grants_o[80];
  assign N172 = N171 | grants_o[81];
  assign N171 = N170 | grants_o[82];
  assign N170 = N169 | grants_o[83];
  assign N169 = N168 | grants_o[84];
  assign N168 = N167 | grants_o[85];
  assign N167 = N166 | grants_o[86];
  assign N166 = N165 | grants_o[87];
  assign N165 = N164 | grants_o[88];
  assign N164 = N163 | grants_o[89];
  assign N163 = N162 | grants_o[90];
  assign N162 = N161 | grants_o[91];
  assign N161 = N160 | grants_o[92];
  assign N160 = N159 | grants_o[93];
  assign N159 = N158 | grants_o[94];
  assign N158 = N157 | grants_o[95];
  assign N157 = N156 | grants_o[96];
  assign N156 = N155 | grants_o[97];
  assign N155 = N154 | grants_o[98];
  assign N154 = N153 | grants_o[99];
  assign N153 = N152 | grants_o[100];
  assign N152 = N151 | grants_o[101];
  assign N151 = N150 | grants_o[102];
  assign N150 = N149 | grants_o[103];
  assign N149 = N148 | grants_o[104];
  assign N148 = N147 | grants_o[105];
  assign N147 = N146 | grants_o[106];
  assign N146 = N145 | grants_o[107];
  assign N145 = N144 | grants_o[108];
  assign N144 = N143 | grants_o[109];
  assign N143 = N142 | grants_o[110];
  assign N142 = N141 | grants_o[111];
  assign N141 = N140 | grants_o[112];
  assign N140 = N139 | grants_o[113];
  assign N139 = N138 | grants_o[114];
  assign N138 = N137 | grants_o[115];
  assign N137 = N136 | grants_o[116];
  assign N136 = N135 | grants_o[117];
  assign N135 = N134 | grants_o[118];
  assign N134 = N133 | grants_o[119];
  assign N133 = N132 | grants_o[120];
  assign N132 = N131 | grants_o[121];
  assign N131 = N130 | grants_o[122];
  assign N130 = N129 | grants_o[123];
  assign N129 = N128 | grants_o[124];
  assign N128 = N127 | grants_o[125];
  assign N127 = grants_o[127] | grants_o[126];
  assign req_mask_r[127] = ~not_req_mask_r[127];
  assign req_mask_r[126] = ~not_req_mask_r[126];
  assign req_mask_r[125] = ~not_req_mask_r[125];
  assign req_mask_r[124] = ~not_req_mask_r[124];
  assign req_mask_r[123] = ~not_req_mask_r[123];
  assign req_mask_r[122] = ~not_req_mask_r[122];
  assign req_mask_r[121] = ~not_req_mask_r[121];
  assign req_mask_r[120] = ~not_req_mask_r[120];
  assign req_mask_r[119] = ~not_req_mask_r[119];
  assign req_mask_r[118] = ~not_req_mask_r[118];
  assign req_mask_r[117] = ~not_req_mask_r[117];
  assign req_mask_r[116] = ~not_req_mask_r[116];
  assign req_mask_r[115] = ~not_req_mask_r[115];
  assign req_mask_r[114] = ~not_req_mask_r[114];
  assign req_mask_r[113] = ~not_req_mask_r[113];
  assign req_mask_r[112] = ~not_req_mask_r[112];
  assign req_mask_r[111] = ~not_req_mask_r[111];
  assign req_mask_r[110] = ~not_req_mask_r[110];
  assign req_mask_r[109] = ~not_req_mask_r[109];
  assign req_mask_r[108] = ~not_req_mask_r[108];
  assign req_mask_r[107] = ~not_req_mask_r[107];
  assign req_mask_r[106] = ~not_req_mask_r[106];
  assign req_mask_r[105] = ~not_req_mask_r[105];
  assign req_mask_r[104] = ~not_req_mask_r[104];
  assign req_mask_r[103] = ~not_req_mask_r[103];
  assign req_mask_r[102] = ~not_req_mask_r[102];
  assign req_mask_r[101] = ~not_req_mask_r[101];
  assign req_mask_r[100] = ~not_req_mask_r[100];
  assign req_mask_r[99] = ~not_req_mask_r[99];
  assign req_mask_r[98] = ~not_req_mask_r[98];
  assign req_mask_r[97] = ~not_req_mask_r[97];
  assign req_mask_r[96] = ~not_req_mask_r[96];
  assign req_mask_r[95] = ~not_req_mask_r[95];
  assign req_mask_r[94] = ~not_req_mask_r[94];
  assign req_mask_r[93] = ~not_req_mask_r[93];
  assign req_mask_r[92] = ~not_req_mask_r[92];
  assign req_mask_r[91] = ~not_req_mask_r[91];
  assign req_mask_r[90] = ~not_req_mask_r[90];
  assign req_mask_r[89] = ~not_req_mask_r[89];
  assign req_mask_r[88] = ~not_req_mask_r[88];
  assign req_mask_r[87] = ~not_req_mask_r[87];
  assign req_mask_r[86] = ~not_req_mask_r[86];
  assign req_mask_r[85] = ~not_req_mask_r[85];
  assign req_mask_r[84] = ~not_req_mask_r[84];
  assign req_mask_r[83] = ~not_req_mask_r[83];
  assign req_mask_r[82] = ~not_req_mask_r[82];
  assign req_mask_r[81] = ~not_req_mask_r[81];
  assign req_mask_r[80] = ~not_req_mask_r[80];
  assign req_mask_r[79] = ~not_req_mask_r[79];
  assign req_mask_r[78] = ~not_req_mask_r[78];
  assign req_mask_r[77] = ~not_req_mask_r[77];
  assign req_mask_r[76] = ~not_req_mask_r[76];
  assign req_mask_r[75] = ~not_req_mask_r[75];
  assign req_mask_r[74] = ~not_req_mask_r[74];
  assign req_mask_r[73] = ~not_req_mask_r[73];
  assign req_mask_r[72] = ~not_req_mask_r[72];
  assign req_mask_r[71] = ~not_req_mask_r[71];
  assign req_mask_r[70] = ~not_req_mask_r[70];
  assign req_mask_r[69] = ~not_req_mask_r[69];
  assign req_mask_r[68] = ~not_req_mask_r[68];
  assign req_mask_r[67] = ~not_req_mask_r[67];
  assign req_mask_r[66] = ~not_req_mask_r[66];
  assign req_mask_r[65] = ~not_req_mask_r[65];
  assign req_mask_r[64] = ~not_req_mask_r[64];
  assign req_mask_r[63] = ~not_req_mask_r[63];
  assign req_mask_r[62] = ~not_req_mask_r[62];
  assign req_mask_r[61] = ~not_req_mask_r[61];
  assign req_mask_r[60] = ~not_req_mask_r[60];
  assign req_mask_r[59] = ~not_req_mask_r[59];
  assign req_mask_r[58] = ~not_req_mask_r[58];
  assign req_mask_r[57] = ~not_req_mask_r[57];
  assign req_mask_r[56] = ~not_req_mask_r[56];
  assign req_mask_r[55] = ~not_req_mask_r[55];
  assign req_mask_r[54] = ~not_req_mask_r[54];
  assign req_mask_r[53] = ~not_req_mask_r[53];
  assign req_mask_r[52] = ~not_req_mask_r[52];
  assign req_mask_r[51] = ~not_req_mask_r[51];
  assign req_mask_r[50] = ~not_req_mask_r[50];
  assign req_mask_r[49] = ~not_req_mask_r[49];
  assign req_mask_r[48] = ~not_req_mask_r[48];
  assign req_mask_r[47] = ~not_req_mask_r[47];
  assign req_mask_r[46] = ~not_req_mask_r[46];
  assign req_mask_r[45] = ~not_req_mask_r[45];
  assign req_mask_r[44] = ~not_req_mask_r[44];
  assign req_mask_r[43] = ~not_req_mask_r[43];
  assign req_mask_r[42] = ~not_req_mask_r[42];
  assign req_mask_r[41] = ~not_req_mask_r[41];
  assign req_mask_r[40] = ~not_req_mask_r[40];
  assign req_mask_r[39] = ~not_req_mask_r[39];
  assign req_mask_r[38] = ~not_req_mask_r[38];
  assign req_mask_r[37] = ~not_req_mask_r[37];
  assign req_mask_r[36] = ~not_req_mask_r[36];
  assign req_mask_r[35] = ~not_req_mask_r[35];
  assign req_mask_r[34] = ~not_req_mask_r[34];
  assign req_mask_r[33] = ~not_req_mask_r[33];
  assign req_mask_r[32] = ~not_req_mask_r[32];
  assign req_mask_r[31] = ~not_req_mask_r[31];
  assign req_mask_r[30] = ~not_req_mask_r[30];
  assign req_mask_r[29] = ~not_req_mask_r[29];
  assign req_mask_r[28] = ~not_req_mask_r[28];
  assign req_mask_r[27] = ~not_req_mask_r[27];
  assign req_mask_r[26] = ~not_req_mask_r[26];
  assign req_mask_r[25] = ~not_req_mask_r[25];
  assign req_mask_r[24] = ~not_req_mask_r[24];
  assign req_mask_r[23] = ~not_req_mask_r[23];
  assign req_mask_r[22] = ~not_req_mask_r[22];
  assign req_mask_r[21] = ~not_req_mask_r[21];
  assign req_mask_r[20] = ~not_req_mask_r[20];
  assign req_mask_r[19] = ~not_req_mask_r[19];
  assign req_mask_r[18] = ~not_req_mask_r[18];
  assign req_mask_r[17] = ~not_req_mask_r[17];
  assign req_mask_r[16] = ~not_req_mask_r[16];
  assign req_mask_r[15] = ~not_req_mask_r[15];
  assign req_mask_r[14] = ~not_req_mask_r[14];
  assign req_mask_r[13] = ~not_req_mask_r[13];
  assign req_mask_r[12] = ~not_req_mask_r[12];
  assign req_mask_r[11] = ~not_req_mask_r[11];
  assign req_mask_r[10] = ~not_req_mask_r[10];
  assign req_mask_r[9] = ~not_req_mask_r[9];
  assign req_mask_r[8] = ~not_req_mask_r[8];
  assign req_mask_r[7] = ~not_req_mask_r[7];
  assign req_mask_r[6] = ~not_req_mask_r[6];
  assign req_mask_r[5] = ~not_req_mask_r[5];
  assign req_mask_r[4] = ~not_req_mask_r[4];
  assign req_mask_r[3] = ~not_req_mask_r[3];
  assign req_mask_r[2] = ~not_req_mask_r[2];
  assign req_mask_r[1] = ~not_req_mask_r[1];
  assign req_mask_r[0] = ~not_req_mask_r[0];
  assign n_2_net__127_ = reqs_i[127] & req_mask_r[127];
  assign n_2_net__126_ = reqs_i[126] & req_mask_r[126];
  assign n_2_net__125_ = reqs_i[125] & req_mask_r[125];
  assign n_2_net__124_ = reqs_i[124] & req_mask_r[124];
  assign n_2_net__123_ = reqs_i[123] & req_mask_r[123];
  assign n_2_net__122_ = reqs_i[122] & req_mask_r[122];
  assign n_2_net__121_ = reqs_i[121] & req_mask_r[121];
  assign n_2_net__120_ = reqs_i[120] & req_mask_r[120];
  assign n_2_net__119_ = reqs_i[119] & req_mask_r[119];
  assign n_2_net__118_ = reqs_i[118] & req_mask_r[118];
  assign n_2_net__117_ = reqs_i[117] & req_mask_r[117];
  assign n_2_net__116_ = reqs_i[116] & req_mask_r[116];
  assign n_2_net__115_ = reqs_i[115] & req_mask_r[115];
  assign n_2_net__114_ = reqs_i[114] & req_mask_r[114];
  assign n_2_net__113_ = reqs_i[113] & req_mask_r[113];
  assign n_2_net__112_ = reqs_i[112] & req_mask_r[112];
  assign n_2_net__111_ = reqs_i[111] & req_mask_r[111];
  assign n_2_net__110_ = reqs_i[110] & req_mask_r[110];
  assign n_2_net__109_ = reqs_i[109] & req_mask_r[109];
  assign n_2_net__108_ = reqs_i[108] & req_mask_r[108];
  assign n_2_net__107_ = reqs_i[107] & req_mask_r[107];
  assign n_2_net__106_ = reqs_i[106] & req_mask_r[106];
  assign n_2_net__105_ = reqs_i[105] & req_mask_r[105];
  assign n_2_net__104_ = reqs_i[104] & req_mask_r[104];
  assign n_2_net__103_ = reqs_i[103] & req_mask_r[103];
  assign n_2_net__102_ = reqs_i[102] & req_mask_r[102];
  assign n_2_net__101_ = reqs_i[101] & req_mask_r[101];
  assign n_2_net__100_ = reqs_i[100] & req_mask_r[100];
  assign n_2_net__99_ = reqs_i[99] & req_mask_r[99];
  assign n_2_net__98_ = reqs_i[98] & req_mask_r[98];
  assign n_2_net__97_ = reqs_i[97] & req_mask_r[97];
  assign n_2_net__96_ = reqs_i[96] & req_mask_r[96];
  assign n_2_net__95_ = reqs_i[95] & req_mask_r[95];
  assign n_2_net__94_ = reqs_i[94] & req_mask_r[94];
  assign n_2_net__93_ = reqs_i[93] & req_mask_r[93];
  assign n_2_net__92_ = reqs_i[92] & req_mask_r[92];
  assign n_2_net__91_ = reqs_i[91] & req_mask_r[91];
  assign n_2_net__90_ = reqs_i[90] & req_mask_r[90];
  assign n_2_net__89_ = reqs_i[89] & req_mask_r[89];
  assign n_2_net__88_ = reqs_i[88] & req_mask_r[88];
  assign n_2_net__87_ = reqs_i[87] & req_mask_r[87];
  assign n_2_net__86_ = reqs_i[86] & req_mask_r[86];
  assign n_2_net__85_ = reqs_i[85] & req_mask_r[85];
  assign n_2_net__84_ = reqs_i[84] & req_mask_r[84];
  assign n_2_net__83_ = reqs_i[83] & req_mask_r[83];
  assign n_2_net__82_ = reqs_i[82] & req_mask_r[82];
  assign n_2_net__81_ = reqs_i[81] & req_mask_r[81];
  assign n_2_net__80_ = reqs_i[80] & req_mask_r[80];
  assign n_2_net__79_ = reqs_i[79] & req_mask_r[79];
  assign n_2_net__78_ = reqs_i[78] & req_mask_r[78];
  assign n_2_net__77_ = reqs_i[77] & req_mask_r[77];
  assign n_2_net__76_ = reqs_i[76] & req_mask_r[76];
  assign n_2_net__75_ = reqs_i[75] & req_mask_r[75];
  assign n_2_net__74_ = reqs_i[74] & req_mask_r[74];
  assign n_2_net__73_ = reqs_i[73] & req_mask_r[73];
  assign n_2_net__72_ = reqs_i[72] & req_mask_r[72];
  assign n_2_net__71_ = reqs_i[71] & req_mask_r[71];
  assign n_2_net__70_ = reqs_i[70] & req_mask_r[70];
  assign n_2_net__69_ = reqs_i[69] & req_mask_r[69];
  assign n_2_net__68_ = reqs_i[68] & req_mask_r[68];
  assign n_2_net__67_ = reqs_i[67] & req_mask_r[67];
  assign n_2_net__66_ = reqs_i[66] & req_mask_r[66];
  assign n_2_net__65_ = reqs_i[65] & req_mask_r[65];
  assign n_2_net__64_ = reqs_i[64] & req_mask_r[64];
  assign n_2_net__63_ = reqs_i[63] & req_mask_r[63];
  assign n_2_net__62_ = reqs_i[62] & req_mask_r[62];
  assign n_2_net__61_ = reqs_i[61] & req_mask_r[61];
  assign n_2_net__60_ = reqs_i[60] & req_mask_r[60];
  assign n_2_net__59_ = reqs_i[59] & req_mask_r[59];
  assign n_2_net__58_ = reqs_i[58] & req_mask_r[58];
  assign n_2_net__57_ = reqs_i[57] & req_mask_r[57];
  assign n_2_net__56_ = reqs_i[56] & req_mask_r[56];
  assign n_2_net__55_ = reqs_i[55] & req_mask_r[55];
  assign n_2_net__54_ = reqs_i[54] & req_mask_r[54];
  assign n_2_net__53_ = reqs_i[53] & req_mask_r[53];
  assign n_2_net__52_ = reqs_i[52] & req_mask_r[52];
  assign n_2_net__51_ = reqs_i[51] & req_mask_r[51];
  assign n_2_net__50_ = reqs_i[50] & req_mask_r[50];
  assign n_2_net__49_ = reqs_i[49] & req_mask_r[49];
  assign n_2_net__48_ = reqs_i[48] & req_mask_r[48];
  assign n_2_net__47_ = reqs_i[47] & req_mask_r[47];
  assign n_2_net__46_ = reqs_i[46] & req_mask_r[46];
  assign n_2_net__45_ = reqs_i[45] & req_mask_r[45];
  assign n_2_net__44_ = reqs_i[44] & req_mask_r[44];
  assign n_2_net__43_ = reqs_i[43] & req_mask_r[43];
  assign n_2_net__42_ = reqs_i[42] & req_mask_r[42];
  assign n_2_net__41_ = reqs_i[41] & req_mask_r[41];
  assign n_2_net__40_ = reqs_i[40] & req_mask_r[40];
  assign n_2_net__39_ = reqs_i[39] & req_mask_r[39];
  assign n_2_net__38_ = reqs_i[38] & req_mask_r[38];
  assign n_2_net__37_ = reqs_i[37] & req_mask_r[37];
  assign n_2_net__36_ = reqs_i[36] & req_mask_r[36];
  assign n_2_net__35_ = reqs_i[35] & req_mask_r[35];
  assign n_2_net__34_ = reqs_i[34] & req_mask_r[34];
  assign n_2_net__33_ = reqs_i[33] & req_mask_r[33];
  assign n_2_net__32_ = reqs_i[32] & req_mask_r[32];
  assign n_2_net__31_ = reqs_i[31] & req_mask_r[31];
  assign n_2_net__30_ = reqs_i[30] & req_mask_r[30];
  assign n_2_net__29_ = reqs_i[29] & req_mask_r[29];
  assign n_2_net__28_ = reqs_i[28] & req_mask_r[28];
  assign n_2_net__27_ = reqs_i[27] & req_mask_r[27];
  assign n_2_net__26_ = reqs_i[26] & req_mask_r[26];
  assign n_2_net__25_ = reqs_i[25] & req_mask_r[25];
  assign n_2_net__24_ = reqs_i[24] & req_mask_r[24];
  assign n_2_net__23_ = reqs_i[23] & req_mask_r[23];
  assign n_2_net__22_ = reqs_i[22] & req_mask_r[22];
  assign n_2_net__21_ = reqs_i[21] & req_mask_r[21];
  assign n_2_net__20_ = reqs_i[20] & req_mask_r[20];
  assign n_2_net__19_ = reqs_i[19] & req_mask_r[19];
  assign n_2_net__18_ = reqs_i[18] & req_mask_r[18];
  assign n_2_net__17_ = reqs_i[17] & req_mask_r[17];
  assign n_2_net__16_ = reqs_i[16] & req_mask_r[16];
  assign n_2_net__15_ = reqs_i[15] & req_mask_r[15];
  assign n_2_net__14_ = reqs_i[14] & req_mask_r[14];
  assign n_2_net__13_ = reqs_i[13] & req_mask_r[13];
  assign n_2_net__12_ = reqs_i[12] & req_mask_r[12];
  assign n_2_net__11_ = reqs_i[11] & req_mask_r[11];
  assign n_2_net__10_ = reqs_i[10] & req_mask_r[10];
  assign n_2_net__9_ = reqs_i[9] & req_mask_r[9];
  assign n_2_net__8_ = reqs_i[8] & req_mask_r[8];
  assign n_2_net__7_ = reqs_i[7] & req_mask_r[7];
  assign n_2_net__6_ = reqs_i[6] & req_mask_r[6];
  assign n_2_net__5_ = reqs_i[5] & req_mask_r[5];
  assign n_2_net__4_ = reqs_i[4] & req_mask_r[4];
  assign n_2_net__3_ = reqs_i[3] & req_mask_r[3];
  assign n_2_net__2_ = reqs_i[2] & req_mask_r[2];
  assign n_2_net__1_ = reqs_i[1] & req_mask_r[1];
  assign n_2_net__0_ = reqs_i[0] & req_mask_r[0];

endmodule

