

module top
(
  clk,
  reset,
  valid_i,
  data_i,
  yumi_o,
  in_top_channel_i,
  out_top_channel_i,
  valid_o,
  data_o,
  ready_i
);

  input [15:0] valid_i;
  input [1023:0] data_i;
  output [15:0] yumi_o;
  input [3:0] in_top_channel_i;
  input [2:0] out_top_channel_i;
  output [7:0] valid_o;
  output [511:0] data_o;
  input [7:0] ready_i;
  input clk;
  input reset;

  bsg_round_robin_fifo_to_fifo
  wrapper
  (
    .valid_i(valid_i),
    .data_i(data_i),
    .yumi_o(yumi_o),
    .in_top_channel_i(in_top_channel_i),
    .out_top_channel_i(out_top_channel_i),
    .valid_o(valid_o),
    .data_o(data_o),
    .ready_i(ready_i),
    .clk(clk),
    .reset(reset)
  );


endmodule



module bsg_make_2D_array_width_p64_items_p8
(
  i,
  o
);

  input [511:0] i;
  output [511:0] o;
  wire [511:0] o;
  assign o[511] = i[511];
  assign o[510] = i[510];
  assign o[509] = i[509];
  assign o[508] = i[508];
  assign o[507] = i[507];
  assign o[506] = i[506];
  assign o[505] = i[505];
  assign o[504] = i[504];
  assign o[503] = i[503];
  assign o[502] = i[502];
  assign o[501] = i[501];
  assign o[500] = i[500];
  assign o[499] = i[499];
  assign o[498] = i[498];
  assign o[497] = i[497];
  assign o[496] = i[496];
  assign o[495] = i[495];
  assign o[494] = i[494];
  assign o[493] = i[493];
  assign o[492] = i[492];
  assign o[491] = i[491];
  assign o[490] = i[490];
  assign o[489] = i[489];
  assign o[488] = i[488];
  assign o[487] = i[487];
  assign o[486] = i[486];
  assign o[485] = i[485];
  assign o[484] = i[484];
  assign o[483] = i[483];
  assign o[482] = i[482];
  assign o[481] = i[481];
  assign o[480] = i[480];
  assign o[479] = i[479];
  assign o[478] = i[478];
  assign o[477] = i[477];
  assign o[476] = i[476];
  assign o[475] = i[475];
  assign o[474] = i[474];
  assign o[473] = i[473];
  assign o[472] = i[472];
  assign o[471] = i[471];
  assign o[470] = i[470];
  assign o[469] = i[469];
  assign o[468] = i[468];
  assign o[467] = i[467];
  assign o[466] = i[466];
  assign o[465] = i[465];
  assign o[464] = i[464];
  assign o[463] = i[463];
  assign o[462] = i[462];
  assign o[461] = i[461];
  assign o[460] = i[460];
  assign o[459] = i[459];
  assign o[458] = i[458];
  assign o[457] = i[457];
  assign o[456] = i[456];
  assign o[455] = i[455];
  assign o[454] = i[454];
  assign o[453] = i[453];
  assign o[452] = i[452];
  assign o[451] = i[451];
  assign o[450] = i[450];
  assign o[449] = i[449];
  assign o[448] = i[448];
  assign o[447] = i[447];
  assign o[446] = i[446];
  assign o[445] = i[445];
  assign o[444] = i[444];
  assign o[443] = i[443];
  assign o[442] = i[442];
  assign o[441] = i[441];
  assign o[440] = i[440];
  assign o[439] = i[439];
  assign o[438] = i[438];
  assign o[437] = i[437];
  assign o[436] = i[436];
  assign o[435] = i[435];
  assign o[434] = i[434];
  assign o[433] = i[433];
  assign o[432] = i[432];
  assign o[431] = i[431];
  assign o[430] = i[430];
  assign o[429] = i[429];
  assign o[428] = i[428];
  assign o[427] = i[427];
  assign o[426] = i[426];
  assign o[425] = i[425];
  assign o[424] = i[424];
  assign o[423] = i[423];
  assign o[422] = i[422];
  assign o[421] = i[421];
  assign o[420] = i[420];
  assign o[419] = i[419];
  assign o[418] = i[418];
  assign o[417] = i[417];
  assign o[416] = i[416];
  assign o[415] = i[415];
  assign o[414] = i[414];
  assign o[413] = i[413];
  assign o[412] = i[412];
  assign o[411] = i[411];
  assign o[410] = i[410];
  assign o[409] = i[409];
  assign o[408] = i[408];
  assign o[407] = i[407];
  assign o[406] = i[406];
  assign o[405] = i[405];
  assign o[404] = i[404];
  assign o[403] = i[403];
  assign o[402] = i[402];
  assign o[401] = i[401];
  assign o[400] = i[400];
  assign o[399] = i[399];
  assign o[398] = i[398];
  assign o[397] = i[397];
  assign o[396] = i[396];
  assign o[395] = i[395];
  assign o[394] = i[394];
  assign o[393] = i[393];
  assign o[392] = i[392];
  assign o[391] = i[391];
  assign o[390] = i[390];
  assign o[389] = i[389];
  assign o[388] = i[388];
  assign o[387] = i[387];
  assign o[386] = i[386];
  assign o[385] = i[385];
  assign o[384] = i[384];
  assign o[383] = i[383];
  assign o[382] = i[382];
  assign o[381] = i[381];
  assign o[380] = i[380];
  assign o[379] = i[379];
  assign o[378] = i[378];
  assign o[377] = i[377];
  assign o[376] = i[376];
  assign o[375] = i[375];
  assign o[374] = i[374];
  assign o[373] = i[373];
  assign o[372] = i[372];
  assign o[371] = i[371];
  assign o[370] = i[370];
  assign o[369] = i[369];
  assign o[368] = i[368];
  assign o[367] = i[367];
  assign o[366] = i[366];
  assign o[365] = i[365];
  assign o[364] = i[364];
  assign o[363] = i[363];
  assign o[362] = i[362];
  assign o[361] = i[361];
  assign o[360] = i[360];
  assign o[359] = i[359];
  assign o[358] = i[358];
  assign o[357] = i[357];
  assign o[356] = i[356];
  assign o[355] = i[355];
  assign o[354] = i[354];
  assign o[353] = i[353];
  assign o[352] = i[352];
  assign o[351] = i[351];
  assign o[350] = i[350];
  assign o[349] = i[349];
  assign o[348] = i[348];
  assign o[347] = i[347];
  assign o[346] = i[346];
  assign o[345] = i[345];
  assign o[344] = i[344];
  assign o[343] = i[343];
  assign o[342] = i[342];
  assign o[341] = i[341];
  assign o[340] = i[340];
  assign o[339] = i[339];
  assign o[338] = i[338];
  assign o[337] = i[337];
  assign o[336] = i[336];
  assign o[335] = i[335];
  assign o[334] = i[334];
  assign o[333] = i[333];
  assign o[332] = i[332];
  assign o[331] = i[331];
  assign o[330] = i[330];
  assign o[329] = i[329];
  assign o[328] = i[328];
  assign o[327] = i[327];
  assign o[326] = i[326];
  assign o[325] = i[325];
  assign o[324] = i[324];
  assign o[323] = i[323];
  assign o[322] = i[322];
  assign o[321] = i[321];
  assign o[320] = i[320];
  assign o[319] = i[319];
  assign o[318] = i[318];
  assign o[317] = i[317];
  assign o[316] = i[316];
  assign o[315] = i[315];
  assign o[314] = i[314];
  assign o[313] = i[313];
  assign o[312] = i[312];
  assign o[311] = i[311];
  assign o[310] = i[310];
  assign o[309] = i[309];
  assign o[308] = i[308];
  assign o[307] = i[307];
  assign o[306] = i[306];
  assign o[305] = i[305];
  assign o[304] = i[304];
  assign o[303] = i[303];
  assign o[302] = i[302];
  assign o[301] = i[301];
  assign o[300] = i[300];
  assign o[299] = i[299];
  assign o[298] = i[298];
  assign o[297] = i[297];
  assign o[296] = i[296];
  assign o[295] = i[295];
  assign o[294] = i[294];
  assign o[293] = i[293];
  assign o[292] = i[292];
  assign o[291] = i[291];
  assign o[290] = i[290];
  assign o[289] = i[289];
  assign o[288] = i[288];
  assign o[287] = i[287];
  assign o[286] = i[286];
  assign o[285] = i[285];
  assign o[284] = i[284];
  assign o[283] = i[283];
  assign o[282] = i[282];
  assign o[281] = i[281];
  assign o[280] = i[280];
  assign o[279] = i[279];
  assign o[278] = i[278];
  assign o[277] = i[277];
  assign o[276] = i[276];
  assign o[275] = i[275];
  assign o[274] = i[274];
  assign o[273] = i[273];
  assign o[272] = i[272];
  assign o[271] = i[271];
  assign o[270] = i[270];
  assign o[269] = i[269];
  assign o[268] = i[268];
  assign o[267] = i[267];
  assign o[266] = i[266];
  assign o[265] = i[265];
  assign o[264] = i[264];
  assign o[263] = i[263];
  assign o[262] = i[262];
  assign o[261] = i[261];
  assign o[260] = i[260];
  assign o[259] = i[259];
  assign o[258] = i[258];
  assign o[257] = i[257];
  assign o[256] = i[256];
  assign o[255] = i[255];
  assign o[254] = i[254];
  assign o[253] = i[253];
  assign o[252] = i[252];
  assign o[251] = i[251];
  assign o[250] = i[250];
  assign o[249] = i[249];
  assign o[248] = i[248];
  assign o[247] = i[247];
  assign o[246] = i[246];
  assign o[245] = i[245];
  assign o[244] = i[244];
  assign o[243] = i[243];
  assign o[242] = i[242];
  assign o[241] = i[241];
  assign o[240] = i[240];
  assign o[239] = i[239];
  assign o[238] = i[238];
  assign o[237] = i[237];
  assign o[236] = i[236];
  assign o[235] = i[235];
  assign o[234] = i[234];
  assign o[233] = i[233];
  assign o[232] = i[232];
  assign o[231] = i[231];
  assign o[230] = i[230];
  assign o[229] = i[229];
  assign o[228] = i[228];
  assign o[227] = i[227];
  assign o[226] = i[226];
  assign o[225] = i[225];
  assign o[224] = i[224];
  assign o[223] = i[223];
  assign o[222] = i[222];
  assign o[221] = i[221];
  assign o[220] = i[220];
  assign o[219] = i[219];
  assign o[218] = i[218];
  assign o[217] = i[217];
  assign o[216] = i[216];
  assign o[215] = i[215];
  assign o[214] = i[214];
  assign o[213] = i[213];
  assign o[212] = i[212];
  assign o[211] = i[211];
  assign o[210] = i[210];
  assign o[209] = i[209];
  assign o[208] = i[208];
  assign o[207] = i[207];
  assign o[206] = i[206];
  assign o[205] = i[205];
  assign o[204] = i[204];
  assign o[203] = i[203];
  assign o[202] = i[202];
  assign o[201] = i[201];
  assign o[200] = i[200];
  assign o[199] = i[199];
  assign o[198] = i[198];
  assign o[197] = i[197];
  assign o[196] = i[196];
  assign o[195] = i[195];
  assign o[194] = i[194];
  assign o[193] = i[193];
  assign o[192] = i[192];
  assign o[191] = i[191];
  assign o[190] = i[190];
  assign o[189] = i[189];
  assign o[188] = i[188];
  assign o[187] = i[187];
  assign o[186] = i[186];
  assign o[185] = i[185];
  assign o[184] = i[184];
  assign o[183] = i[183];
  assign o[182] = i[182];
  assign o[181] = i[181];
  assign o[180] = i[180];
  assign o[179] = i[179];
  assign o[178] = i[178];
  assign o[177] = i[177];
  assign o[176] = i[176];
  assign o[175] = i[175];
  assign o[174] = i[174];
  assign o[173] = i[173];
  assign o[172] = i[172];
  assign o[171] = i[171];
  assign o[170] = i[170];
  assign o[169] = i[169];
  assign o[168] = i[168];
  assign o[167] = i[167];
  assign o[166] = i[166];
  assign o[165] = i[165];
  assign o[164] = i[164];
  assign o[163] = i[163];
  assign o[162] = i[162];
  assign o[161] = i[161];
  assign o[160] = i[160];
  assign o[159] = i[159];
  assign o[158] = i[158];
  assign o[157] = i[157];
  assign o[156] = i[156];
  assign o[155] = i[155];
  assign o[154] = i[154];
  assign o[153] = i[153];
  assign o[152] = i[152];
  assign o[151] = i[151];
  assign o[150] = i[150];
  assign o[149] = i[149];
  assign o[148] = i[148];
  assign o[147] = i[147];
  assign o[146] = i[146];
  assign o[145] = i[145];
  assign o[144] = i[144];
  assign o[143] = i[143];
  assign o[142] = i[142];
  assign o[141] = i[141];
  assign o[140] = i[140];
  assign o[139] = i[139];
  assign o[138] = i[138];
  assign o[137] = i[137];
  assign o[136] = i[136];
  assign o[135] = i[135];
  assign o[134] = i[134];
  assign o[133] = i[133];
  assign o[132] = i[132];
  assign o[131] = i[131];
  assign o[130] = i[130];
  assign o[129] = i[129];
  assign o[128] = i[128];
  assign o[127] = i[127];
  assign o[126] = i[126];
  assign o[125] = i[125];
  assign o[124] = i[124];
  assign o[123] = i[123];
  assign o[122] = i[122];
  assign o[121] = i[121];
  assign o[120] = i[120];
  assign o[119] = i[119];
  assign o[118] = i[118];
  assign o[117] = i[117];
  assign o[116] = i[116];
  assign o[115] = i[115];
  assign o[114] = i[114];
  assign o[113] = i[113];
  assign o[112] = i[112];
  assign o[111] = i[111];
  assign o[110] = i[110];
  assign o[109] = i[109];
  assign o[108] = i[108];
  assign o[107] = i[107];
  assign o[106] = i[106];
  assign o[105] = i[105];
  assign o[104] = i[104];
  assign o[103] = i[103];
  assign o[102] = i[102];
  assign o[101] = i[101];
  assign o[100] = i[100];
  assign o[99] = i[99];
  assign o[98] = i[98];
  assign o[97] = i[97];
  assign o[96] = i[96];
  assign o[95] = i[95];
  assign o[94] = i[94];
  assign o[93] = i[93];
  assign o[92] = i[92];
  assign o[91] = i[91];
  assign o[90] = i[90];
  assign o[89] = i[89];
  assign o[88] = i[88];
  assign o[87] = i[87];
  assign o[86] = i[86];
  assign o[85] = i[85];
  assign o[84] = i[84];
  assign o[83] = i[83];
  assign o[82] = i[82];
  assign o[81] = i[81];
  assign o[80] = i[80];
  assign o[79] = i[79];
  assign o[78] = i[78];
  assign o[77] = i[77];
  assign o[76] = i[76];
  assign o[75] = i[75];
  assign o[74] = i[74];
  assign o[73] = i[73];
  assign o[72] = i[72];
  assign o[71] = i[71];
  assign o[70] = i[70];
  assign o[69] = i[69];
  assign o[68] = i[68];
  assign o[67] = i[67];
  assign o[66] = i[66];
  assign o[65] = i[65];
  assign o[64] = i[64];
  assign o[63] = i[63];
  assign o[62] = i[62];
  assign o[61] = i[61];
  assign o[60] = i[60];
  assign o[59] = i[59];
  assign o[58] = i[58];
  assign o[57] = i[57];
  assign o[56] = i[56];
  assign o[55] = i[55];
  assign o[54] = i[54];
  assign o[53] = i[53];
  assign o[52] = i[52];
  assign o[51] = i[51];
  assign o[50] = i[50];
  assign o[49] = i[49];
  assign o[48] = i[48];
  assign o[47] = i[47];
  assign o[46] = i[46];
  assign o[45] = i[45];
  assign o[44] = i[44];
  assign o[43] = i[43];
  assign o[42] = i[42];
  assign o[41] = i[41];
  assign o[40] = i[40];
  assign o[39] = i[39];
  assign o[38] = i[38];
  assign o[37] = i[37];
  assign o[36] = i[36];
  assign o[35] = i[35];
  assign o[34] = i[34];
  assign o[33] = i[33];
  assign o[32] = i[32];
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_rotate_right_width_p16
(
  data_i,
  rot_i,
  o
);

  input [15:0] data_i;
  input [3:0] rot_i;
  output [15:0] o;
  wire [15:0] o;
  wire SYNOPSYS_UNCONNECTED_1,SYNOPSYS_UNCONNECTED_2,SYNOPSYS_UNCONNECTED_3,
  SYNOPSYS_UNCONNECTED_4,SYNOPSYS_UNCONNECTED_5,SYNOPSYS_UNCONNECTED_6,
  SYNOPSYS_UNCONNECTED_7,SYNOPSYS_UNCONNECTED_8,SYNOPSYS_UNCONNECTED_9,SYNOPSYS_UNCONNECTED_10,
  SYNOPSYS_UNCONNECTED_11,SYNOPSYS_UNCONNECTED_12,SYNOPSYS_UNCONNECTED_13,
  SYNOPSYS_UNCONNECTED_14,SYNOPSYS_UNCONNECTED_15;
  assign { SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, o } = { data_i[14:0], data_i } >> rot_i;

endmodule



module bsg_circular_ptr_slots_p16_max_add_p8
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [3:0] add_i;
  output [3:0] o;
  output [3:0] n_o;
  input clk;
  input reset_i;
  wire [3:0] n_o;
  wire N0,N1,N2,N3,N4,N5,N6;
  reg [3:0] o;
  assign n_o = o + add_i;
  assign { N6, N5, N4, N3 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N1)? n_o : 1'b0;
  assign N0 = reset_i;
  assign N1 = N2;
  assign N2 = ~reset_i;

  always @(posedge clk) begin
    if(1'b1) begin
      { o[3:0] } <= { N6, N5, N4, N3 };
    end 
  end


endmodule



module bsg_rr_f2f_input_width_p64_num_in_p16_middle_meet_p8
(
  clk,
  reset,
  valid_i,
  data_i,
  data_head_o,
  valid_head_o,
  go_channels_i,
  go_cnt_i,
  yumi_o
);

  input [15:0] valid_i;
  input [1023:0] data_i;
  output [511:0] data_head_o;
  output [7:0] valid_head_o;
  input [7:0] go_channels_i;
  input [3:0] go_cnt_i;
  output [15:0] yumi_o;
  input clk;
  input reset;
  wire [511:0] data_head_o,data_head_o_flat_pretrunc;
  wire [7:0] valid_head_o;
  wire [15:0] yumi_o;
  wire SYNOPSYS_UNCONNECTED_1,SYNOPSYS_UNCONNECTED_2,SYNOPSYS_UNCONNECTED_3,
  SYNOPSYS_UNCONNECTED_4,SYNOPSYS_UNCONNECTED_5,SYNOPSYS_UNCONNECTED_6,
  SYNOPSYS_UNCONNECTED_7,SYNOPSYS_UNCONNECTED_8,SYNOPSYS_UNCONNECTED_9,SYNOPSYS_UNCONNECTED_10,
  SYNOPSYS_UNCONNECTED_11,SYNOPSYS_UNCONNECTED_12,SYNOPSYS_UNCONNECTED_13,
  SYNOPSYS_UNCONNECTED_14,SYNOPSYS_UNCONNECTED_15,SYNOPSYS_UNCONNECTED_16,SYNOPSYS_UNCONNECTED_17,
  SYNOPSYS_UNCONNECTED_18,SYNOPSYS_UNCONNECTED_19,SYNOPSYS_UNCONNECTED_20,
  SYNOPSYS_UNCONNECTED_21,SYNOPSYS_UNCONNECTED_22,SYNOPSYS_UNCONNECTED_23,
  SYNOPSYS_UNCONNECTED_24,SYNOPSYS_UNCONNECTED_25,SYNOPSYS_UNCONNECTED_26,SYNOPSYS_UNCONNECTED_27,
  SYNOPSYS_UNCONNECTED_28,SYNOPSYS_UNCONNECTED_29,SYNOPSYS_UNCONNECTED_30,
  SYNOPSYS_UNCONNECTED_31,SYNOPSYS_UNCONNECTED_32,SYNOPSYS_UNCONNECTED_33,
  SYNOPSYS_UNCONNECTED_34,SYNOPSYS_UNCONNECTED_35,SYNOPSYS_UNCONNECTED_36,SYNOPSYS_UNCONNECTED_37,
  SYNOPSYS_UNCONNECTED_38,SYNOPSYS_UNCONNECTED_39,SYNOPSYS_UNCONNECTED_40,
  SYNOPSYS_UNCONNECTED_41,SYNOPSYS_UNCONNECTED_42,SYNOPSYS_UNCONNECTED_43,
  SYNOPSYS_UNCONNECTED_44,SYNOPSYS_UNCONNECTED_45,SYNOPSYS_UNCONNECTED_46,SYNOPSYS_UNCONNECTED_47,
  SYNOPSYS_UNCONNECTED_48,SYNOPSYS_UNCONNECTED_49,SYNOPSYS_UNCONNECTED_50,
  SYNOPSYS_UNCONNECTED_51,SYNOPSYS_UNCONNECTED_52,SYNOPSYS_UNCONNECTED_53,
  SYNOPSYS_UNCONNECTED_54,SYNOPSYS_UNCONNECTED_55,SYNOPSYS_UNCONNECTED_56,SYNOPSYS_UNCONNECTED_57,
  SYNOPSYS_UNCONNECTED_58,SYNOPSYS_UNCONNECTED_59,SYNOPSYS_UNCONNECTED_60,
  SYNOPSYS_UNCONNECTED_61,SYNOPSYS_UNCONNECTED_62,SYNOPSYS_UNCONNECTED_63,
  SYNOPSYS_UNCONNECTED_64,SYNOPSYS_UNCONNECTED_65,SYNOPSYS_UNCONNECTED_66,SYNOPSYS_UNCONNECTED_67,
  SYNOPSYS_UNCONNECTED_68,SYNOPSYS_UNCONNECTED_69,SYNOPSYS_UNCONNECTED_70,
  SYNOPSYS_UNCONNECTED_71,SYNOPSYS_UNCONNECTED_72,SYNOPSYS_UNCONNECTED_73,
  SYNOPSYS_UNCONNECTED_74,SYNOPSYS_UNCONNECTED_75,SYNOPSYS_UNCONNECTED_76,SYNOPSYS_UNCONNECTED_77,
  SYNOPSYS_UNCONNECTED_78,SYNOPSYS_UNCONNECTED_79,SYNOPSYS_UNCONNECTED_80,
  SYNOPSYS_UNCONNECTED_81,SYNOPSYS_UNCONNECTED_82,SYNOPSYS_UNCONNECTED_83,
  SYNOPSYS_UNCONNECTED_84,SYNOPSYS_UNCONNECTED_85,SYNOPSYS_UNCONNECTED_86,SYNOPSYS_UNCONNECTED_87,
  SYNOPSYS_UNCONNECTED_88,SYNOPSYS_UNCONNECTED_89,SYNOPSYS_UNCONNECTED_90,
  SYNOPSYS_UNCONNECTED_91,SYNOPSYS_UNCONNECTED_92,SYNOPSYS_UNCONNECTED_93,
  SYNOPSYS_UNCONNECTED_94,SYNOPSYS_UNCONNECTED_95,SYNOPSYS_UNCONNECTED_96,SYNOPSYS_UNCONNECTED_97,
  SYNOPSYS_UNCONNECTED_98,SYNOPSYS_UNCONNECTED_99,SYNOPSYS_UNCONNECTED_100,
  SYNOPSYS_UNCONNECTED_101,SYNOPSYS_UNCONNECTED_102,SYNOPSYS_UNCONNECTED_103,
  SYNOPSYS_UNCONNECTED_104,SYNOPSYS_UNCONNECTED_105,SYNOPSYS_UNCONNECTED_106,
  SYNOPSYS_UNCONNECTED_107,SYNOPSYS_UNCONNECTED_108,SYNOPSYS_UNCONNECTED_109,
  SYNOPSYS_UNCONNECTED_110,SYNOPSYS_UNCONNECTED_111,SYNOPSYS_UNCONNECTED_112,SYNOPSYS_UNCONNECTED_113,
  SYNOPSYS_UNCONNECTED_114,SYNOPSYS_UNCONNECTED_115,SYNOPSYS_UNCONNECTED_116,
  SYNOPSYS_UNCONNECTED_117,SYNOPSYS_UNCONNECTED_118,SYNOPSYS_UNCONNECTED_119,
  SYNOPSYS_UNCONNECTED_120,SYNOPSYS_UNCONNECTED_121,SYNOPSYS_UNCONNECTED_122,
  SYNOPSYS_UNCONNECTED_123,SYNOPSYS_UNCONNECTED_124,SYNOPSYS_UNCONNECTED_125,
  SYNOPSYS_UNCONNECTED_126,SYNOPSYS_UNCONNECTED_127,SYNOPSYS_UNCONNECTED_128,SYNOPSYS_UNCONNECTED_129,
  SYNOPSYS_UNCONNECTED_130,SYNOPSYS_UNCONNECTED_131,SYNOPSYS_UNCONNECTED_132,
  SYNOPSYS_UNCONNECTED_133,SYNOPSYS_UNCONNECTED_134,SYNOPSYS_UNCONNECTED_135,
  SYNOPSYS_UNCONNECTED_136,SYNOPSYS_UNCONNECTED_137,SYNOPSYS_UNCONNECTED_138,
  SYNOPSYS_UNCONNECTED_139,SYNOPSYS_UNCONNECTED_140,SYNOPSYS_UNCONNECTED_141,
  SYNOPSYS_UNCONNECTED_142,SYNOPSYS_UNCONNECTED_143,SYNOPSYS_UNCONNECTED_144,SYNOPSYS_UNCONNECTED_145,
  SYNOPSYS_UNCONNECTED_146,SYNOPSYS_UNCONNECTED_147,SYNOPSYS_UNCONNECTED_148,
  SYNOPSYS_UNCONNECTED_149,SYNOPSYS_UNCONNECTED_150,SYNOPSYS_UNCONNECTED_151,
  SYNOPSYS_UNCONNECTED_152,SYNOPSYS_UNCONNECTED_153,SYNOPSYS_UNCONNECTED_154,
  SYNOPSYS_UNCONNECTED_155,SYNOPSYS_UNCONNECTED_156,SYNOPSYS_UNCONNECTED_157,
  SYNOPSYS_UNCONNECTED_158,SYNOPSYS_UNCONNECTED_159,SYNOPSYS_UNCONNECTED_160,SYNOPSYS_UNCONNECTED_161,
  SYNOPSYS_UNCONNECTED_162,SYNOPSYS_UNCONNECTED_163,SYNOPSYS_UNCONNECTED_164,
  SYNOPSYS_UNCONNECTED_165,SYNOPSYS_UNCONNECTED_166,SYNOPSYS_UNCONNECTED_167,
  SYNOPSYS_UNCONNECTED_168,SYNOPSYS_UNCONNECTED_169,SYNOPSYS_UNCONNECTED_170,
  SYNOPSYS_UNCONNECTED_171,SYNOPSYS_UNCONNECTED_172,SYNOPSYS_UNCONNECTED_173,
  SYNOPSYS_UNCONNECTED_174,SYNOPSYS_UNCONNECTED_175,SYNOPSYS_UNCONNECTED_176,SYNOPSYS_UNCONNECTED_177,
  SYNOPSYS_UNCONNECTED_178,SYNOPSYS_UNCONNECTED_179,SYNOPSYS_UNCONNECTED_180,
  SYNOPSYS_UNCONNECTED_181,SYNOPSYS_UNCONNECTED_182,SYNOPSYS_UNCONNECTED_183,
  SYNOPSYS_UNCONNECTED_184,SYNOPSYS_UNCONNECTED_185,SYNOPSYS_UNCONNECTED_186,
  SYNOPSYS_UNCONNECTED_187,SYNOPSYS_UNCONNECTED_188,SYNOPSYS_UNCONNECTED_189,
  SYNOPSYS_UNCONNECTED_190,SYNOPSYS_UNCONNECTED_191,SYNOPSYS_UNCONNECTED_192,SYNOPSYS_UNCONNECTED_193,
  SYNOPSYS_UNCONNECTED_194,SYNOPSYS_UNCONNECTED_195,SYNOPSYS_UNCONNECTED_196,
  SYNOPSYS_UNCONNECTED_197,SYNOPSYS_UNCONNECTED_198,SYNOPSYS_UNCONNECTED_199,
  SYNOPSYS_UNCONNECTED_200,SYNOPSYS_UNCONNECTED_201,SYNOPSYS_UNCONNECTED_202,
  SYNOPSYS_UNCONNECTED_203,SYNOPSYS_UNCONNECTED_204,SYNOPSYS_UNCONNECTED_205,
  SYNOPSYS_UNCONNECTED_206,SYNOPSYS_UNCONNECTED_207,SYNOPSYS_UNCONNECTED_208,SYNOPSYS_UNCONNECTED_209,
  SYNOPSYS_UNCONNECTED_210,SYNOPSYS_UNCONNECTED_211,SYNOPSYS_UNCONNECTED_212,
  SYNOPSYS_UNCONNECTED_213,SYNOPSYS_UNCONNECTED_214,SYNOPSYS_UNCONNECTED_215,
  SYNOPSYS_UNCONNECTED_216,SYNOPSYS_UNCONNECTED_217,SYNOPSYS_UNCONNECTED_218,
  SYNOPSYS_UNCONNECTED_219,SYNOPSYS_UNCONNECTED_220,SYNOPSYS_UNCONNECTED_221,
  SYNOPSYS_UNCONNECTED_222,SYNOPSYS_UNCONNECTED_223,SYNOPSYS_UNCONNECTED_224,SYNOPSYS_UNCONNECTED_225,
  SYNOPSYS_UNCONNECTED_226,SYNOPSYS_UNCONNECTED_227,SYNOPSYS_UNCONNECTED_228,
  SYNOPSYS_UNCONNECTED_229,SYNOPSYS_UNCONNECTED_230,SYNOPSYS_UNCONNECTED_231,
  SYNOPSYS_UNCONNECTED_232,SYNOPSYS_UNCONNECTED_233,SYNOPSYS_UNCONNECTED_234,
  SYNOPSYS_UNCONNECTED_235,SYNOPSYS_UNCONNECTED_236,SYNOPSYS_UNCONNECTED_237,
  SYNOPSYS_UNCONNECTED_238,SYNOPSYS_UNCONNECTED_239,SYNOPSYS_UNCONNECTED_240,SYNOPSYS_UNCONNECTED_241,
  SYNOPSYS_UNCONNECTED_242,SYNOPSYS_UNCONNECTED_243,SYNOPSYS_UNCONNECTED_244,
  SYNOPSYS_UNCONNECTED_245,SYNOPSYS_UNCONNECTED_246,SYNOPSYS_UNCONNECTED_247,
  SYNOPSYS_UNCONNECTED_248,SYNOPSYS_UNCONNECTED_249,SYNOPSYS_UNCONNECTED_250,
  SYNOPSYS_UNCONNECTED_251,SYNOPSYS_UNCONNECTED_252,SYNOPSYS_UNCONNECTED_253,
  SYNOPSYS_UNCONNECTED_254,SYNOPSYS_UNCONNECTED_255,SYNOPSYS_UNCONNECTED_256,SYNOPSYS_UNCONNECTED_257,
  SYNOPSYS_UNCONNECTED_258,SYNOPSYS_UNCONNECTED_259,SYNOPSYS_UNCONNECTED_260,
  SYNOPSYS_UNCONNECTED_261,SYNOPSYS_UNCONNECTED_262,SYNOPSYS_UNCONNECTED_263,
  SYNOPSYS_UNCONNECTED_264,SYNOPSYS_UNCONNECTED_265,SYNOPSYS_UNCONNECTED_266,
  SYNOPSYS_UNCONNECTED_267,SYNOPSYS_UNCONNECTED_268,SYNOPSYS_UNCONNECTED_269,
  SYNOPSYS_UNCONNECTED_270,SYNOPSYS_UNCONNECTED_271,SYNOPSYS_UNCONNECTED_272,SYNOPSYS_UNCONNECTED_273,
  SYNOPSYS_UNCONNECTED_274,SYNOPSYS_UNCONNECTED_275,SYNOPSYS_UNCONNECTED_276,
  SYNOPSYS_UNCONNECTED_277,SYNOPSYS_UNCONNECTED_278,SYNOPSYS_UNCONNECTED_279,
  SYNOPSYS_UNCONNECTED_280,SYNOPSYS_UNCONNECTED_281,SYNOPSYS_UNCONNECTED_282,
  SYNOPSYS_UNCONNECTED_283,SYNOPSYS_UNCONNECTED_284,SYNOPSYS_UNCONNECTED_285,
  SYNOPSYS_UNCONNECTED_286,SYNOPSYS_UNCONNECTED_287,SYNOPSYS_UNCONNECTED_288,SYNOPSYS_UNCONNECTED_289,
  SYNOPSYS_UNCONNECTED_290,SYNOPSYS_UNCONNECTED_291,SYNOPSYS_UNCONNECTED_292,
  SYNOPSYS_UNCONNECTED_293,SYNOPSYS_UNCONNECTED_294,SYNOPSYS_UNCONNECTED_295,
  SYNOPSYS_UNCONNECTED_296,SYNOPSYS_UNCONNECTED_297,SYNOPSYS_UNCONNECTED_298,
  SYNOPSYS_UNCONNECTED_299,SYNOPSYS_UNCONNECTED_300,SYNOPSYS_UNCONNECTED_301,
  SYNOPSYS_UNCONNECTED_302,SYNOPSYS_UNCONNECTED_303,SYNOPSYS_UNCONNECTED_304,SYNOPSYS_UNCONNECTED_305,
  SYNOPSYS_UNCONNECTED_306,SYNOPSYS_UNCONNECTED_307,SYNOPSYS_UNCONNECTED_308,
  SYNOPSYS_UNCONNECTED_309,SYNOPSYS_UNCONNECTED_310,SYNOPSYS_UNCONNECTED_311,
  SYNOPSYS_UNCONNECTED_312,SYNOPSYS_UNCONNECTED_313,SYNOPSYS_UNCONNECTED_314,
  SYNOPSYS_UNCONNECTED_315,SYNOPSYS_UNCONNECTED_316,SYNOPSYS_UNCONNECTED_317,
  SYNOPSYS_UNCONNECTED_318,SYNOPSYS_UNCONNECTED_319,SYNOPSYS_UNCONNECTED_320,SYNOPSYS_UNCONNECTED_321,
  SYNOPSYS_UNCONNECTED_322,SYNOPSYS_UNCONNECTED_323,SYNOPSYS_UNCONNECTED_324,
  SYNOPSYS_UNCONNECTED_325,SYNOPSYS_UNCONNECTED_326,SYNOPSYS_UNCONNECTED_327,
  SYNOPSYS_UNCONNECTED_328,SYNOPSYS_UNCONNECTED_329,SYNOPSYS_UNCONNECTED_330,
  SYNOPSYS_UNCONNECTED_331,SYNOPSYS_UNCONNECTED_332,SYNOPSYS_UNCONNECTED_333,
  SYNOPSYS_UNCONNECTED_334,SYNOPSYS_UNCONNECTED_335,SYNOPSYS_UNCONNECTED_336,SYNOPSYS_UNCONNECTED_337,
  SYNOPSYS_UNCONNECTED_338,SYNOPSYS_UNCONNECTED_339,SYNOPSYS_UNCONNECTED_340,
  SYNOPSYS_UNCONNECTED_341,SYNOPSYS_UNCONNECTED_342,SYNOPSYS_UNCONNECTED_343,
  SYNOPSYS_UNCONNECTED_344,SYNOPSYS_UNCONNECTED_345,SYNOPSYS_UNCONNECTED_346,
  SYNOPSYS_UNCONNECTED_347,SYNOPSYS_UNCONNECTED_348,SYNOPSYS_UNCONNECTED_349,
  SYNOPSYS_UNCONNECTED_350,SYNOPSYS_UNCONNECTED_351,SYNOPSYS_UNCONNECTED_352,SYNOPSYS_UNCONNECTED_353,
  SYNOPSYS_UNCONNECTED_354,SYNOPSYS_UNCONNECTED_355,SYNOPSYS_UNCONNECTED_356,
  SYNOPSYS_UNCONNECTED_357,SYNOPSYS_UNCONNECTED_358,SYNOPSYS_UNCONNECTED_359,
  SYNOPSYS_UNCONNECTED_360,SYNOPSYS_UNCONNECTED_361,SYNOPSYS_UNCONNECTED_362,
  SYNOPSYS_UNCONNECTED_363,SYNOPSYS_UNCONNECTED_364,SYNOPSYS_UNCONNECTED_365,
  SYNOPSYS_UNCONNECTED_366,SYNOPSYS_UNCONNECTED_367,SYNOPSYS_UNCONNECTED_368,SYNOPSYS_UNCONNECTED_369,
  SYNOPSYS_UNCONNECTED_370,SYNOPSYS_UNCONNECTED_371,SYNOPSYS_UNCONNECTED_372,
  SYNOPSYS_UNCONNECTED_373,SYNOPSYS_UNCONNECTED_374,SYNOPSYS_UNCONNECTED_375,
  SYNOPSYS_UNCONNECTED_376,SYNOPSYS_UNCONNECTED_377,SYNOPSYS_UNCONNECTED_378,
  SYNOPSYS_UNCONNECTED_379,SYNOPSYS_UNCONNECTED_380,SYNOPSYS_UNCONNECTED_381,
  SYNOPSYS_UNCONNECTED_382,SYNOPSYS_UNCONNECTED_383,SYNOPSYS_UNCONNECTED_384,SYNOPSYS_UNCONNECTED_385,
  SYNOPSYS_UNCONNECTED_386,SYNOPSYS_UNCONNECTED_387,SYNOPSYS_UNCONNECTED_388,
  SYNOPSYS_UNCONNECTED_389,SYNOPSYS_UNCONNECTED_390,SYNOPSYS_UNCONNECTED_391,
  SYNOPSYS_UNCONNECTED_392,SYNOPSYS_UNCONNECTED_393,SYNOPSYS_UNCONNECTED_394,
  SYNOPSYS_UNCONNECTED_395,SYNOPSYS_UNCONNECTED_396,SYNOPSYS_UNCONNECTED_397,
  SYNOPSYS_UNCONNECTED_398,SYNOPSYS_UNCONNECTED_399,SYNOPSYS_UNCONNECTED_400,SYNOPSYS_UNCONNECTED_401,
  SYNOPSYS_UNCONNECTED_402,SYNOPSYS_UNCONNECTED_403,SYNOPSYS_UNCONNECTED_404,
  SYNOPSYS_UNCONNECTED_405,SYNOPSYS_UNCONNECTED_406,SYNOPSYS_UNCONNECTED_407,
  SYNOPSYS_UNCONNECTED_408,SYNOPSYS_UNCONNECTED_409,SYNOPSYS_UNCONNECTED_410,
  SYNOPSYS_UNCONNECTED_411,SYNOPSYS_UNCONNECTED_412,SYNOPSYS_UNCONNECTED_413,
  SYNOPSYS_UNCONNECTED_414,SYNOPSYS_UNCONNECTED_415,SYNOPSYS_UNCONNECTED_416,SYNOPSYS_UNCONNECTED_417,
  SYNOPSYS_UNCONNECTED_418,SYNOPSYS_UNCONNECTED_419,SYNOPSYS_UNCONNECTED_420,
  SYNOPSYS_UNCONNECTED_421,SYNOPSYS_UNCONNECTED_422,SYNOPSYS_UNCONNECTED_423,
  SYNOPSYS_UNCONNECTED_424,SYNOPSYS_UNCONNECTED_425,SYNOPSYS_UNCONNECTED_426,
  SYNOPSYS_UNCONNECTED_427,SYNOPSYS_UNCONNECTED_428,SYNOPSYS_UNCONNECTED_429,
  SYNOPSYS_UNCONNECTED_430,SYNOPSYS_UNCONNECTED_431,SYNOPSYS_UNCONNECTED_432,SYNOPSYS_UNCONNECTED_433,
  SYNOPSYS_UNCONNECTED_434,SYNOPSYS_UNCONNECTED_435,SYNOPSYS_UNCONNECTED_436,
  SYNOPSYS_UNCONNECTED_437,SYNOPSYS_UNCONNECTED_438,SYNOPSYS_UNCONNECTED_439,
  SYNOPSYS_UNCONNECTED_440,SYNOPSYS_UNCONNECTED_441,SYNOPSYS_UNCONNECTED_442,
  SYNOPSYS_UNCONNECTED_443,SYNOPSYS_UNCONNECTED_444,SYNOPSYS_UNCONNECTED_445,
  SYNOPSYS_UNCONNECTED_446,SYNOPSYS_UNCONNECTED_447,SYNOPSYS_UNCONNECTED_448,SYNOPSYS_UNCONNECTED_449,
  SYNOPSYS_UNCONNECTED_450,SYNOPSYS_UNCONNECTED_451,SYNOPSYS_UNCONNECTED_452,
  SYNOPSYS_UNCONNECTED_453,SYNOPSYS_UNCONNECTED_454,SYNOPSYS_UNCONNECTED_455,
  SYNOPSYS_UNCONNECTED_456,SYNOPSYS_UNCONNECTED_457,SYNOPSYS_UNCONNECTED_458,
  SYNOPSYS_UNCONNECTED_459,SYNOPSYS_UNCONNECTED_460,SYNOPSYS_UNCONNECTED_461,
  SYNOPSYS_UNCONNECTED_462,SYNOPSYS_UNCONNECTED_463,SYNOPSYS_UNCONNECTED_464,SYNOPSYS_UNCONNECTED_465,
  SYNOPSYS_UNCONNECTED_466,SYNOPSYS_UNCONNECTED_467,SYNOPSYS_UNCONNECTED_468,
  SYNOPSYS_UNCONNECTED_469,SYNOPSYS_UNCONNECTED_470,SYNOPSYS_UNCONNECTED_471,
  SYNOPSYS_UNCONNECTED_472,SYNOPSYS_UNCONNECTED_473,SYNOPSYS_UNCONNECTED_474,
  SYNOPSYS_UNCONNECTED_475,SYNOPSYS_UNCONNECTED_476,SYNOPSYS_UNCONNECTED_477,
  SYNOPSYS_UNCONNECTED_478,SYNOPSYS_UNCONNECTED_479,SYNOPSYS_UNCONNECTED_480,SYNOPSYS_UNCONNECTED_481,
  SYNOPSYS_UNCONNECTED_482,SYNOPSYS_UNCONNECTED_483,SYNOPSYS_UNCONNECTED_484,
  SYNOPSYS_UNCONNECTED_485,SYNOPSYS_UNCONNECTED_486,SYNOPSYS_UNCONNECTED_487,
  SYNOPSYS_UNCONNECTED_488,SYNOPSYS_UNCONNECTED_489,SYNOPSYS_UNCONNECTED_490,
  SYNOPSYS_UNCONNECTED_491,SYNOPSYS_UNCONNECTED_492,SYNOPSYS_UNCONNECTED_493,
  SYNOPSYS_UNCONNECTED_494,SYNOPSYS_UNCONNECTED_495,SYNOPSYS_UNCONNECTED_496,SYNOPSYS_UNCONNECTED_497,
  SYNOPSYS_UNCONNECTED_498,SYNOPSYS_UNCONNECTED_499,SYNOPSYS_UNCONNECTED_500,
  SYNOPSYS_UNCONNECTED_501,SYNOPSYS_UNCONNECTED_502,SYNOPSYS_UNCONNECTED_503,
  SYNOPSYS_UNCONNECTED_504,SYNOPSYS_UNCONNECTED_505,SYNOPSYS_UNCONNECTED_506,
  SYNOPSYS_UNCONNECTED_507,SYNOPSYS_UNCONNECTED_508,SYNOPSYS_UNCONNECTED_509,
  SYNOPSYS_UNCONNECTED_510,SYNOPSYS_UNCONNECTED_511,SYNOPSYS_UNCONNECTED_512,SYNOPSYS_UNCONNECTED_513,
  SYNOPSYS_UNCONNECTED_514,SYNOPSYS_UNCONNECTED_515,SYNOPSYS_UNCONNECTED_516,
  SYNOPSYS_UNCONNECTED_517,SYNOPSYS_UNCONNECTED_518,SYNOPSYS_UNCONNECTED_519,
  SYNOPSYS_UNCONNECTED_520,SYNOPSYS_UNCONNECTED_521,SYNOPSYS_UNCONNECTED_522,
  SYNOPSYS_UNCONNECTED_523,SYNOPSYS_UNCONNECTED_524,SYNOPSYS_UNCONNECTED_525,
  SYNOPSYS_UNCONNECTED_526,SYNOPSYS_UNCONNECTED_527,SYNOPSYS_UNCONNECTED_528,SYNOPSYS_UNCONNECTED_529,
  SYNOPSYS_UNCONNECTED_530,SYNOPSYS_UNCONNECTED_531,SYNOPSYS_UNCONNECTED_532,
  SYNOPSYS_UNCONNECTED_533,SYNOPSYS_UNCONNECTED_534,SYNOPSYS_UNCONNECTED_535,
  SYNOPSYS_UNCONNECTED_536,SYNOPSYS_UNCONNECTED_537,SYNOPSYS_UNCONNECTED_538,
  SYNOPSYS_UNCONNECTED_539,SYNOPSYS_UNCONNECTED_540,SYNOPSYS_UNCONNECTED_541,
  SYNOPSYS_UNCONNECTED_542,SYNOPSYS_UNCONNECTED_543,SYNOPSYS_UNCONNECTED_544,SYNOPSYS_UNCONNECTED_545,
  SYNOPSYS_UNCONNECTED_546,SYNOPSYS_UNCONNECTED_547,SYNOPSYS_UNCONNECTED_548,
  SYNOPSYS_UNCONNECTED_549,SYNOPSYS_UNCONNECTED_550,SYNOPSYS_UNCONNECTED_551,
  SYNOPSYS_UNCONNECTED_552,SYNOPSYS_UNCONNECTED_553,SYNOPSYS_UNCONNECTED_554,
  SYNOPSYS_UNCONNECTED_555,SYNOPSYS_UNCONNECTED_556,SYNOPSYS_UNCONNECTED_557,
  SYNOPSYS_UNCONNECTED_558,SYNOPSYS_UNCONNECTED_559,SYNOPSYS_UNCONNECTED_560,SYNOPSYS_UNCONNECTED_561,
  SYNOPSYS_UNCONNECTED_562,SYNOPSYS_UNCONNECTED_563,SYNOPSYS_UNCONNECTED_564,
  SYNOPSYS_UNCONNECTED_565,SYNOPSYS_UNCONNECTED_566,SYNOPSYS_UNCONNECTED_567,
  SYNOPSYS_UNCONNECTED_568,SYNOPSYS_UNCONNECTED_569,SYNOPSYS_UNCONNECTED_570,
  SYNOPSYS_UNCONNECTED_571,SYNOPSYS_UNCONNECTED_572,SYNOPSYS_UNCONNECTED_573,
  SYNOPSYS_UNCONNECTED_574,SYNOPSYS_UNCONNECTED_575,SYNOPSYS_UNCONNECTED_576,SYNOPSYS_UNCONNECTED_577,
  SYNOPSYS_UNCONNECTED_578,SYNOPSYS_UNCONNECTED_579,SYNOPSYS_UNCONNECTED_580,
  SYNOPSYS_UNCONNECTED_581,SYNOPSYS_UNCONNECTED_582,SYNOPSYS_UNCONNECTED_583,
  SYNOPSYS_UNCONNECTED_584,SYNOPSYS_UNCONNECTED_585,SYNOPSYS_UNCONNECTED_586,
  SYNOPSYS_UNCONNECTED_587,SYNOPSYS_UNCONNECTED_588,SYNOPSYS_UNCONNECTED_589,
  SYNOPSYS_UNCONNECTED_590,SYNOPSYS_UNCONNECTED_591,SYNOPSYS_UNCONNECTED_592,SYNOPSYS_UNCONNECTED_593,
  SYNOPSYS_UNCONNECTED_594,SYNOPSYS_UNCONNECTED_595,SYNOPSYS_UNCONNECTED_596,
  SYNOPSYS_UNCONNECTED_597,SYNOPSYS_UNCONNECTED_598,SYNOPSYS_UNCONNECTED_599,
  SYNOPSYS_UNCONNECTED_600,SYNOPSYS_UNCONNECTED_601,SYNOPSYS_UNCONNECTED_602,
  SYNOPSYS_UNCONNECTED_603,SYNOPSYS_UNCONNECTED_604,SYNOPSYS_UNCONNECTED_605,
  SYNOPSYS_UNCONNECTED_606,SYNOPSYS_UNCONNECTED_607,SYNOPSYS_UNCONNECTED_608,SYNOPSYS_UNCONNECTED_609,
  SYNOPSYS_UNCONNECTED_610,SYNOPSYS_UNCONNECTED_611,SYNOPSYS_UNCONNECTED_612,
  SYNOPSYS_UNCONNECTED_613,SYNOPSYS_UNCONNECTED_614,SYNOPSYS_UNCONNECTED_615,
  SYNOPSYS_UNCONNECTED_616,SYNOPSYS_UNCONNECTED_617,SYNOPSYS_UNCONNECTED_618,
  SYNOPSYS_UNCONNECTED_619,SYNOPSYS_UNCONNECTED_620,SYNOPSYS_UNCONNECTED_621,
  SYNOPSYS_UNCONNECTED_622,SYNOPSYS_UNCONNECTED_623,SYNOPSYS_UNCONNECTED_624,SYNOPSYS_UNCONNECTED_625,
  SYNOPSYS_UNCONNECTED_626,SYNOPSYS_UNCONNECTED_627,SYNOPSYS_UNCONNECTED_628,
  SYNOPSYS_UNCONNECTED_629,SYNOPSYS_UNCONNECTED_630,SYNOPSYS_UNCONNECTED_631,
  SYNOPSYS_UNCONNECTED_632,SYNOPSYS_UNCONNECTED_633,SYNOPSYS_UNCONNECTED_634,
  SYNOPSYS_UNCONNECTED_635,SYNOPSYS_UNCONNECTED_636,SYNOPSYS_UNCONNECTED_637,
  SYNOPSYS_UNCONNECTED_638,SYNOPSYS_UNCONNECTED_639,SYNOPSYS_UNCONNECTED_640,SYNOPSYS_UNCONNECTED_641,
  SYNOPSYS_UNCONNECTED_642,SYNOPSYS_UNCONNECTED_643,SYNOPSYS_UNCONNECTED_644,
  SYNOPSYS_UNCONNECTED_645,SYNOPSYS_UNCONNECTED_646,SYNOPSYS_UNCONNECTED_647,
  SYNOPSYS_UNCONNECTED_648,SYNOPSYS_UNCONNECTED_649,SYNOPSYS_UNCONNECTED_650,
  SYNOPSYS_UNCONNECTED_651,SYNOPSYS_UNCONNECTED_652,SYNOPSYS_UNCONNECTED_653,
  SYNOPSYS_UNCONNECTED_654,SYNOPSYS_UNCONNECTED_655,SYNOPSYS_UNCONNECTED_656,SYNOPSYS_UNCONNECTED_657,
  SYNOPSYS_UNCONNECTED_658,SYNOPSYS_UNCONNECTED_659,SYNOPSYS_UNCONNECTED_660,
  SYNOPSYS_UNCONNECTED_661,SYNOPSYS_UNCONNECTED_662,SYNOPSYS_UNCONNECTED_663,
  SYNOPSYS_UNCONNECTED_664,SYNOPSYS_UNCONNECTED_665,SYNOPSYS_UNCONNECTED_666,
  SYNOPSYS_UNCONNECTED_667,SYNOPSYS_UNCONNECTED_668,SYNOPSYS_UNCONNECTED_669,
  SYNOPSYS_UNCONNECTED_670,SYNOPSYS_UNCONNECTED_671,SYNOPSYS_UNCONNECTED_672,SYNOPSYS_UNCONNECTED_673,
  SYNOPSYS_UNCONNECTED_674,SYNOPSYS_UNCONNECTED_675,SYNOPSYS_UNCONNECTED_676,
  SYNOPSYS_UNCONNECTED_677,SYNOPSYS_UNCONNECTED_678,SYNOPSYS_UNCONNECTED_679,
  SYNOPSYS_UNCONNECTED_680,SYNOPSYS_UNCONNECTED_681,SYNOPSYS_UNCONNECTED_682,
  SYNOPSYS_UNCONNECTED_683,SYNOPSYS_UNCONNECTED_684,SYNOPSYS_UNCONNECTED_685,
  SYNOPSYS_UNCONNECTED_686,SYNOPSYS_UNCONNECTED_687,SYNOPSYS_UNCONNECTED_688,SYNOPSYS_UNCONNECTED_689,
  SYNOPSYS_UNCONNECTED_690,SYNOPSYS_UNCONNECTED_691,SYNOPSYS_UNCONNECTED_692,
  SYNOPSYS_UNCONNECTED_693,SYNOPSYS_UNCONNECTED_694,SYNOPSYS_UNCONNECTED_695,
  SYNOPSYS_UNCONNECTED_696,SYNOPSYS_UNCONNECTED_697,SYNOPSYS_UNCONNECTED_698,
  SYNOPSYS_UNCONNECTED_699,SYNOPSYS_UNCONNECTED_700,SYNOPSYS_UNCONNECTED_701,
  SYNOPSYS_UNCONNECTED_702,SYNOPSYS_UNCONNECTED_703,SYNOPSYS_UNCONNECTED_704,SYNOPSYS_UNCONNECTED_705,
  SYNOPSYS_UNCONNECTED_706,SYNOPSYS_UNCONNECTED_707,SYNOPSYS_UNCONNECTED_708,
  SYNOPSYS_UNCONNECTED_709,SYNOPSYS_UNCONNECTED_710,SYNOPSYS_UNCONNECTED_711,
  SYNOPSYS_UNCONNECTED_712,SYNOPSYS_UNCONNECTED_713,SYNOPSYS_UNCONNECTED_714,
  SYNOPSYS_UNCONNECTED_715,SYNOPSYS_UNCONNECTED_716,SYNOPSYS_UNCONNECTED_717,
  SYNOPSYS_UNCONNECTED_718,SYNOPSYS_UNCONNECTED_719,SYNOPSYS_UNCONNECTED_720,SYNOPSYS_UNCONNECTED_721,
  SYNOPSYS_UNCONNECTED_722,SYNOPSYS_UNCONNECTED_723,SYNOPSYS_UNCONNECTED_724,
  SYNOPSYS_UNCONNECTED_725,SYNOPSYS_UNCONNECTED_726,SYNOPSYS_UNCONNECTED_727,
  SYNOPSYS_UNCONNECTED_728,SYNOPSYS_UNCONNECTED_729,SYNOPSYS_UNCONNECTED_730,
  SYNOPSYS_UNCONNECTED_731,SYNOPSYS_UNCONNECTED_732,SYNOPSYS_UNCONNECTED_733,
  SYNOPSYS_UNCONNECTED_734,SYNOPSYS_UNCONNECTED_735,SYNOPSYS_UNCONNECTED_736,SYNOPSYS_UNCONNECTED_737,
  SYNOPSYS_UNCONNECTED_738,SYNOPSYS_UNCONNECTED_739,SYNOPSYS_UNCONNECTED_740,
  SYNOPSYS_UNCONNECTED_741,SYNOPSYS_UNCONNECTED_742,SYNOPSYS_UNCONNECTED_743,
  SYNOPSYS_UNCONNECTED_744,SYNOPSYS_UNCONNECTED_745,SYNOPSYS_UNCONNECTED_746,
  SYNOPSYS_UNCONNECTED_747,SYNOPSYS_UNCONNECTED_748,SYNOPSYS_UNCONNECTED_749,
  SYNOPSYS_UNCONNECTED_750,SYNOPSYS_UNCONNECTED_751,SYNOPSYS_UNCONNECTED_752,SYNOPSYS_UNCONNECTED_753,
  SYNOPSYS_UNCONNECTED_754,SYNOPSYS_UNCONNECTED_755,SYNOPSYS_UNCONNECTED_756,
  SYNOPSYS_UNCONNECTED_757,SYNOPSYS_UNCONNECTED_758,SYNOPSYS_UNCONNECTED_759,
  SYNOPSYS_UNCONNECTED_760,SYNOPSYS_UNCONNECTED_761,SYNOPSYS_UNCONNECTED_762,
  SYNOPSYS_UNCONNECTED_763,SYNOPSYS_UNCONNECTED_764,SYNOPSYS_UNCONNECTED_765,
  SYNOPSYS_UNCONNECTED_766,SYNOPSYS_UNCONNECTED_767,SYNOPSYS_UNCONNECTED_768,SYNOPSYS_UNCONNECTED_769,
  SYNOPSYS_UNCONNECTED_770,SYNOPSYS_UNCONNECTED_771,SYNOPSYS_UNCONNECTED_772,
  SYNOPSYS_UNCONNECTED_773,SYNOPSYS_UNCONNECTED_774,SYNOPSYS_UNCONNECTED_775,
  SYNOPSYS_UNCONNECTED_776,SYNOPSYS_UNCONNECTED_777,SYNOPSYS_UNCONNECTED_778,
  SYNOPSYS_UNCONNECTED_779,SYNOPSYS_UNCONNECTED_780,SYNOPSYS_UNCONNECTED_781,
  SYNOPSYS_UNCONNECTED_782,SYNOPSYS_UNCONNECTED_783,SYNOPSYS_UNCONNECTED_784,SYNOPSYS_UNCONNECTED_785,
  SYNOPSYS_UNCONNECTED_786,SYNOPSYS_UNCONNECTED_787,SYNOPSYS_UNCONNECTED_788,
  SYNOPSYS_UNCONNECTED_789,SYNOPSYS_UNCONNECTED_790,SYNOPSYS_UNCONNECTED_791,
  SYNOPSYS_UNCONNECTED_792,SYNOPSYS_UNCONNECTED_793,SYNOPSYS_UNCONNECTED_794,
  SYNOPSYS_UNCONNECTED_795,SYNOPSYS_UNCONNECTED_796,SYNOPSYS_UNCONNECTED_797,
  SYNOPSYS_UNCONNECTED_798,SYNOPSYS_UNCONNECTED_799,SYNOPSYS_UNCONNECTED_800,SYNOPSYS_UNCONNECTED_801,
  SYNOPSYS_UNCONNECTED_802,SYNOPSYS_UNCONNECTED_803,SYNOPSYS_UNCONNECTED_804,
  SYNOPSYS_UNCONNECTED_805,SYNOPSYS_UNCONNECTED_806,SYNOPSYS_UNCONNECTED_807,
  SYNOPSYS_UNCONNECTED_808,SYNOPSYS_UNCONNECTED_809,SYNOPSYS_UNCONNECTED_810,
  SYNOPSYS_UNCONNECTED_811,SYNOPSYS_UNCONNECTED_812,SYNOPSYS_UNCONNECTED_813,
  SYNOPSYS_UNCONNECTED_814,SYNOPSYS_UNCONNECTED_815,SYNOPSYS_UNCONNECTED_816,SYNOPSYS_UNCONNECTED_817,
  SYNOPSYS_UNCONNECTED_818,SYNOPSYS_UNCONNECTED_819,SYNOPSYS_UNCONNECTED_820,
  SYNOPSYS_UNCONNECTED_821,SYNOPSYS_UNCONNECTED_822,SYNOPSYS_UNCONNECTED_823,
  SYNOPSYS_UNCONNECTED_824,SYNOPSYS_UNCONNECTED_825,SYNOPSYS_UNCONNECTED_826,
  SYNOPSYS_UNCONNECTED_827,SYNOPSYS_UNCONNECTED_828,SYNOPSYS_UNCONNECTED_829,
  SYNOPSYS_UNCONNECTED_830,SYNOPSYS_UNCONNECTED_831,SYNOPSYS_UNCONNECTED_832,SYNOPSYS_UNCONNECTED_833,
  SYNOPSYS_UNCONNECTED_834,SYNOPSYS_UNCONNECTED_835,SYNOPSYS_UNCONNECTED_836,
  SYNOPSYS_UNCONNECTED_837,SYNOPSYS_UNCONNECTED_838,SYNOPSYS_UNCONNECTED_839,
  SYNOPSYS_UNCONNECTED_840,SYNOPSYS_UNCONNECTED_841,SYNOPSYS_UNCONNECTED_842,
  SYNOPSYS_UNCONNECTED_843,SYNOPSYS_UNCONNECTED_844,SYNOPSYS_UNCONNECTED_845,
  SYNOPSYS_UNCONNECTED_846,SYNOPSYS_UNCONNECTED_847,SYNOPSYS_UNCONNECTED_848,SYNOPSYS_UNCONNECTED_849,
  SYNOPSYS_UNCONNECTED_850,SYNOPSYS_UNCONNECTED_851,SYNOPSYS_UNCONNECTED_852,
  SYNOPSYS_UNCONNECTED_853,SYNOPSYS_UNCONNECTED_854,SYNOPSYS_UNCONNECTED_855,
  SYNOPSYS_UNCONNECTED_856,SYNOPSYS_UNCONNECTED_857,SYNOPSYS_UNCONNECTED_858,
  SYNOPSYS_UNCONNECTED_859,SYNOPSYS_UNCONNECTED_860,SYNOPSYS_UNCONNECTED_861,
  SYNOPSYS_UNCONNECTED_862,SYNOPSYS_UNCONNECTED_863,SYNOPSYS_UNCONNECTED_864,SYNOPSYS_UNCONNECTED_865,
  SYNOPSYS_UNCONNECTED_866,SYNOPSYS_UNCONNECTED_867,SYNOPSYS_UNCONNECTED_868,
  SYNOPSYS_UNCONNECTED_869,SYNOPSYS_UNCONNECTED_870,SYNOPSYS_UNCONNECTED_871,
  SYNOPSYS_UNCONNECTED_872,SYNOPSYS_UNCONNECTED_873,SYNOPSYS_UNCONNECTED_874,
  SYNOPSYS_UNCONNECTED_875,SYNOPSYS_UNCONNECTED_876,SYNOPSYS_UNCONNECTED_877,
  SYNOPSYS_UNCONNECTED_878,SYNOPSYS_UNCONNECTED_879,SYNOPSYS_UNCONNECTED_880,SYNOPSYS_UNCONNECTED_881,
  SYNOPSYS_UNCONNECTED_882,SYNOPSYS_UNCONNECTED_883,SYNOPSYS_UNCONNECTED_884,
  SYNOPSYS_UNCONNECTED_885,SYNOPSYS_UNCONNECTED_886,SYNOPSYS_UNCONNECTED_887,
  SYNOPSYS_UNCONNECTED_888,SYNOPSYS_UNCONNECTED_889,SYNOPSYS_UNCONNECTED_890,
  SYNOPSYS_UNCONNECTED_891,SYNOPSYS_UNCONNECTED_892,SYNOPSYS_UNCONNECTED_893,
  SYNOPSYS_UNCONNECTED_894,SYNOPSYS_UNCONNECTED_895,SYNOPSYS_UNCONNECTED_896,SYNOPSYS_UNCONNECTED_897,
  SYNOPSYS_UNCONNECTED_898,SYNOPSYS_UNCONNECTED_899,SYNOPSYS_UNCONNECTED_900,
  SYNOPSYS_UNCONNECTED_901,SYNOPSYS_UNCONNECTED_902,SYNOPSYS_UNCONNECTED_903,
  SYNOPSYS_UNCONNECTED_904,SYNOPSYS_UNCONNECTED_905,SYNOPSYS_UNCONNECTED_906,
  SYNOPSYS_UNCONNECTED_907,SYNOPSYS_UNCONNECTED_908,SYNOPSYS_UNCONNECTED_909,
  SYNOPSYS_UNCONNECTED_910,SYNOPSYS_UNCONNECTED_911,SYNOPSYS_UNCONNECTED_912,SYNOPSYS_UNCONNECTED_913,
  SYNOPSYS_UNCONNECTED_914,SYNOPSYS_UNCONNECTED_915,SYNOPSYS_UNCONNECTED_916,
  SYNOPSYS_UNCONNECTED_917,SYNOPSYS_UNCONNECTED_918,SYNOPSYS_UNCONNECTED_919,
  SYNOPSYS_UNCONNECTED_920,SYNOPSYS_UNCONNECTED_921,SYNOPSYS_UNCONNECTED_922,
  SYNOPSYS_UNCONNECTED_923,SYNOPSYS_UNCONNECTED_924,SYNOPSYS_UNCONNECTED_925,
  SYNOPSYS_UNCONNECTED_926,SYNOPSYS_UNCONNECTED_927,SYNOPSYS_UNCONNECTED_928,SYNOPSYS_UNCONNECTED_929,
  SYNOPSYS_UNCONNECTED_930,SYNOPSYS_UNCONNECTED_931,SYNOPSYS_UNCONNECTED_932,
  SYNOPSYS_UNCONNECTED_933,SYNOPSYS_UNCONNECTED_934,SYNOPSYS_UNCONNECTED_935,
  SYNOPSYS_UNCONNECTED_936,SYNOPSYS_UNCONNECTED_937,SYNOPSYS_UNCONNECTED_938,
  SYNOPSYS_UNCONNECTED_939,SYNOPSYS_UNCONNECTED_940,SYNOPSYS_UNCONNECTED_941,
  SYNOPSYS_UNCONNECTED_942,SYNOPSYS_UNCONNECTED_943,SYNOPSYS_UNCONNECTED_944,SYNOPSYS_UNCONNECTED_945,
  SYNOPSYS_UNCONNECTED_946,SYNOPSYS_UNCONNECTED_947,SYNOPSYS_UNCONNECTED_948,
  SYNOPSYS_UNCONNECTED_949,SYNOPSYS_UNCONNECTED_950,SYNOPSYS_UNCONNECTED_951,
  SYNOPSYS_UNCONNECTED_952,SYNOPSYS_UNCONNECTED_953,SYNOPSYS_UNCONNECTED_954,
  SYNOPSYS_UNCONNECTED_955,SYNOPSYS_UNCONNECTED_956,SYNOPSYS_UNCONNECTED_957,
  SYNOPSYS_UNCONNECTED_958,SYNOPSYS_UNCONNECTED_959,SYNOPSYS_UNCONNECTED_960,SYNOPSYS_UNCONNECTED_961,
  SYNOPSYS_UNCONNECTED_962,SYNOPSYS_UNCONNECTED_963,SYNOPSYS_UNCONNECTED_964,
  SYNOPSYS_UNCONNECTED_965,SYNOPSYS_UNCONNECTED_966,SYNOPSYS_UNCONNECTED_967,
  SYNOPSYS_UNCONNECTED_968,SYNOPSYS_UNCONNECTED_969,SYNOPSYS_UNCONNECTED_970,
  SYNOPSYS_UNCONNECTED_971,SYNOPSYS_UNCONNECTED_972,SYNOPSYS_UNCONNECTED_973,
  SYNOPSYS_UNCONNECTED_974,SYNOPSYS_UNCONNECTED_975,SYNOPSYS_UNCONNECTED_976,SYNOPSYS_UNCONNECTED_977,
  SYNOPSYS_UNCONNECTED_978,SYNOPSYS_UNCONNECTED_979,SYNOPSYS_UNCONNECTED_980,
  SYNOPSYS_UNCONNECTED_981,SYNOPSYS_UNCONNECTED_982,SYNOPSYS_UNCONNECTED_983,
  SYNOPSYS_UNCONNECTED_984,SYNOPSYS_UNCONNECTED_985,SYNOPSYS_UNCONNECTED_986,
  SYNOPSYS_UNCONNECTED_987,SYNOPSYS_UNCONNECTED_988,SYNOPSYS_UNCONNECTED_989,
  SYNOPSYS_UNCONNECTED_990,SYNOPSYS_UNCONNECTED_991,SYNOPSYS_UNCONNECTED_992,SYNOPSYS_UNCONNECTED_993,
  SYNOPSYS_UNCONNECTED_994,SYNOPSYS_UNCONNECTED_995,SYNOPSYS_UNCONNECTED_996,
  SYNOPSYS_UNCONNECTED_997,SYNOPSYS_UNCONNECTED_998,SYNOPSYS_UNCONNECTED_999,
  SYNOPSYS_UNCONNECTED_1000,SYNOPSYS_UNCONNECTED_1001,SYNOPSYS_UNCONNECTED_1002,
  SYNOPSYS_UNCONNECTED_1003,SYNOPSYS_UNCONNECTED_1004,SYNOPSYS_UNCONNECTED_1005,
  SYNOPSYS_UNCONNECTED_1006,SYNOPSYS_UNCONNECTED_1007,SYNOPSYS_UNCONNECTED_1008,
  SYNOPSYS_UNCONNECTED_1009,SYNOPSYS_UNCONNECTED_1010,SYNOPSYS_UNCONNECTED_1011,
  SYNOPSYS_UNCONNECTED_1012,SYNOPSYS_UNCONNECTED_1013,SYNOPSYS_UNCONNECTED_1014,
  SYNOPSYS_UNCONNECTED_1015,SYNOPSYS_UNCONNECTED_1016,SYNOPSYS_UNCONNECTED_1017,
  SYNOPSYS_UNCONNECTED_1018,SYNOPSYS_UNCONNECTED_1019,SYNOPSYS_UNCONNECTED_1020,SYNOPSYS_UNCONNECTED_1021,
  SYNOPSYS_UNCONNECTED_1022,SYNOPSYS_UNCONNECTED_1023,SYNOPSYS_UNCONNECTED_1024,
  SYNOPSYS_UNCONNECTED_1025,SYNOPSYS_UNCONNECTED_1026,SYNOPSYS_UNCONNECTED_1027,
  SYNOPSYS_UNCONNECTED_1028,SYNOPSYS_UNCONNECTED_1029,SYNOPSYS_UNCONNECTED_1030,
  SYNOPSYS_UNCONNECTED_1031,SYNOPSYS_UNCONNECTED_1032,SYNOPSYS_UNCONNECTED_1033,
  SYNOPSYS_UNCONNECTED_1034,SYNOPSYS_UNCONNECTED_1035,SYNOPSYS_UNCONNECTED_1036,
  SYNOPSYS_UNCONNECTED_1037,SYNOPSYS_UNCONNECTED_1038,SYNOPSYS_UNCONNECTED_1039,
  SYNOPSYS_UNCONNECTED_1040,SYNOPSYS_UNCONNECTED_1041,SYNOPSYS_UNCONNECTED_1042,
  SYNOPSYS_UNCONNECTED_1043,SYNOPSYS_UNCONNECTED_1044,SYNOPSYS_UNCONNECTED_1045,
  SYNOPSYS_UNCONNECTED_1046;
  wire [3:0] iptr_r,iptr_r_data;
  wire [15:8] valid_head_o_pretrunc;

  bsg_make_2D_array_width_p64_items_p8
  bm2Da
  (
    .i(data_head_o_flat_pretrunc),
    .o(data_head_o)
  );


  bsg_rotate_right_width_p16
  valid_rr
  (
    .data_i(valid_i),
    .rot_i(iptr_r),
    .o({ valid_head_o_pretrunc, valid_head_o })
  );


  bsg_circular_ptr_slots_p16_max_add_p8
  c_ptr
  (
    .clk(clk),
    .reset_i(reset),
    .add_i(go_cnt_i),
    .o(iptr_r),
    .n_o({ SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4 })
  );


  bsg_circular_ptr_slots_p16_max_add_p8
  c_ptr_data
  (
    .clk(clk),
    .reset_i(reset),
    .add_i(go_cnt_i),
    .o(iptr_r_data),
    .n_o({ SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8 })
  );

  assign { yumi_o, SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, go_channels_i, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, go_channels_i[7:1] } << iptr_r;
  assign { SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_415, SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_417, SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_419, SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_421, SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_423, SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_425, SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_427, SYNOPSYS_UNCONNECTED_428, SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_430, SYNOPSYS_UNCONNECTED_431, SYNOPSYS_UNCONNECTED_432, SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_434, SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_436, SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_438, SYNOPSYS_UNCONNECTED_439, SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441, SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443, SYNOPSYS_UNCONNECTED_444, SYNOPSYS_UNCONNECTED_445, SYNOPSYS_UNCONNECTED_446, SYNOPSYS_UNCONNECTED_447, SYNOPSYS_UNCONNECTED_448, SYNOPSYS_UNCONNECTED_449, SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_451, SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_453, SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_455, SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457, SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_459, SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461, SYNOPSYS_UNCONNECTED_462, SYNOPSYS_UNCONNECTED_463, SYNOPSYS_UNCONNECTED_464, SYNOPSYS_UNCONNECTED_465, SYNOPSYS_UNCONNECTED_466, SYNOPSYS_UNCONNECTED_467, SYNOPSYS_UNCONNECTED_468, SYNOPSYS_UNCONNECTED_469, SYNOPSYS_UNCONNECTED_470, SYNOPSYS_UNCONNECTED_471, SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_473, SYNOPSYS_UNCONNECTED_474, SYNOPSYS_UNCONNECTED_475, SYNOPSYS_UNCONNECTED_476, SYNOPSYS_UNCONNECTED_477, SYNOPSYS_UNCONNECTED_478, SYNOPSYS_UNCONNECTED_479, SYNOPSYS_UNCONNECTED_480, SYNOPSYS_UNCONNECTED_481, SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_483, SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_485, SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_487, SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_489, SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_491, SYNOPSYS_UNCONNECTED_492, SYNOPSYS_UNCONNECTED_493, SYNOPSYS_UNCONNECTED_494, SYNOPSYS_UNCONNECTED_495, SYNOPSYS_UNCONNECTED_496, SYNOPSYS_UNCONNECTED_497, SYNOPSYS_UNCONNECTED_498, SYNOPSYS_UNCONNECTED_499, SYNOPSYS_UNCONNECTED_500, SYNOPSYS_UNCONNECTED_501, SYNOPSYS_UNCONNECTED_502, SYNOPSYS_UNCONNECTED_503, SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_505, SYNOPSYS_UNCONNECTED_506, SYNOPSYS_UNCONNECTED_507, SYNOPSYS_UNCONNECTED_508, SYNOPSYS_UNCONNECTED_509, SYNOPSYS_UNCONNECTED_510, SYNOPSYS_UNCONNECTED_511, SYNOPSYS_UNCONNECTED_512, SYNOPSYS_UNCONNECTED_513, SYNOPSYS_UNCONNECTED_514, SYNOPSYS_UNCONNECTED_515, SYNOPSYS_UNCONNECTED_516, SYNOPSYS_UNCONNECTED_517, SYNOPSYS_UNCONNECTED_518, SYNOPSYS_UNCONNECTED_519, SYNOPSYS_UNCONNECTED_520, SYNOPSYS_UNCONNECTED_521, SYNOPSYS_UNCONNECTED_522, SYNOPSYS_UNCONNECTED_523, SYNOPSYS_UNCONNECTED_524, SYNOPSYS_UNCONNECTED_525, SYNOPSYS_UNCONNECTED_526, SYNOPSYS_UNCONNECTED_527, SYNOPSYS_UNCONNECTED_528, SYNOPSYS_UNCONNECTED_529, SYNOPSYS_UNCONNECTED_530, SYNOPSYS_UNCONNECTED_531, SYNOPSYS_UNCONNECTED_532, SYNOPSYS_UNCONNECTED_533, SYNOPSYS_UNCONNECTED_534, SYNOPSYS_UNCONNECTED_535, SYNOPSYS_UNCONNECTED_536, SYNOPSYS_UNCONNECTED_537, SYNOPSYS_UNCONNECTED_538, SYNOPSYS_UNCONNECTED_539, SYNOPSYS_UNCONNECTED_540, SYNOPSYS_UNCONNECTED_541, SYNOPSYS_UNCONNECTED_542, SYNOPSYS_UNCONNECTED_543, SYNOPSYS_UNCONNECTED_544, SYNOPSYS_UNCONNECTED_545, SYNOPSYS_UNCONNECTED_546, SYNOPSYS_UNCONNECTED_547, SYNOPSYS_UNCONNECTED_548, SYNOPSYS_UNCONNECTED_549, SYNOPSYS_UNCONNECTED_550, SYNOPSYS_UNCONNECTED_551, SYNOPSYS_UNCONNECTED_552, SYNOPSYS_UNCONNECTED_553, SYNOPSYS_UNCONNECTED_554, SYNOPSYS_UNCONNECTED_555, SYNOPSYS_UNCONNECTED_556, SYNOPSYS_UNCONNECTED_557, SYNOPSYS_UNCONNECTED_558, SYNOPSYS_UNCONNECTED_559, SYNOPSYS_UNCONNECTED_560, SYNOPSYS_UNCONNECTED_561, SYNOPSYS_UNCONNECTED_562, SYNOPSYS_UNCONNECTED_563, SYNOPSYS_UNCONNECTED_564, SYNOPSYS_UNCONNECTED_565, SYNOPSYS_UNCONNECTED_566, SYNOPSYS_UNCONNECTED_567, SYNOPSYS_UNCONNECTED_568, SYNOPSYS_UNCONNECTED_569, SYNOPSYS_UNCONNECTED_570, SYNOPSYS_UNCONNECTED_571, SYNOPSYS_UNCONNECTED_572, SYNOPSYS_UNCONNECTED_573, SYNOPSYS_UNCONNECTED_574, SYNOPSYS_UNCONNECTED_575, SYNOPSYS_UNCONNECTED_576, SYNOPSYS_UNCONNECTED_577, SYNOPSYS_UNCONNECTED_578, SYNOPSYS_UNCONNECTED_579, SYNOPSYS_UNCONNECTED_580, SYNOPSYS_UNCONNECTED_581, SYNOPSYS_UNCONNECTED_582, SYNOPSYS_UNCONNECTED_583, SYNOPSYS_UNCONNECTED_584, SYNOPSYS_UNCONNECTED_585, SYNOPSYS_UNCONNECTED_586, SYNOPSYS_UNCONNECTED_587, SYNOPSYS_UNCONNECTED_588, SYNOPSYS_UNCONNECTED_589, SYNOPSYS_UNCONNECTED_590, SYNOPSYS_UNCONNECTED_591, SYNOPSYS_UNCONNECTED_592, SYNOPSYS_UNCONNECTED_593, SYNOPSYS_UNCONNECTED_594, SYNOPSYS_UNCONNECTED_595, SYNOPSYS_UNCONNECTED_596, SYNOPSYS_UNCONNECTED_597, SYNOPSYS_UNCONNECTED_598, SYNOPSYS_UNCONNECTED_599, SYNOPSYS_UNCONNECTED_600, SYNOPSYS_UNCONNECTED_601, SYNOPSYS_UNCONNECTED_602, SYNOPSYS_UNCONNECTED_603, SYNOPSYS_UNCONNECTED_604, SYNOPSYS_UNCONNECTED_605, SYNOPSYS_UNCONNECTED_606, SYNOPSYS_UNCONNECTED_607, SYNOPSYS_UNCONNECTED_608, SYNOPSYS_UNCONNECTED_609, SYNOPSYS_UNCONNECTED_610, SYNOPSYS_UNCONNECTED_611, SYNOPSYS_UNCONNECTED_612, SYNOPSYS_UNCONNECTED_613, SYNOPSYS_UNCONNECTED_614, SYNOPSYS_UNCONNECTED_615, SYNOPSYS_UNCONNECTED_616, SYNOPSYS_UNCONNECTED_617, SYNOPSYS_UNCONNECTED_618, SYNOPSYS_UNCONNECTED_619, SYNOPSYS_UNCONNECTED_620, SYNOPSYS_UNCONNECTED_621, SYNOPSYS_UNCONNECTED_622, SYNOPSYS_UNCONNECTED_623, SYNOPSYS_UNCONNECTED_624, SYNOPSYS_UNCONNECTED_625, SYNOPSYS_UNCONNECTED_626, SYNOPSYS_UNCONNECTED_627, SYNOPSYS_UNCONNECTED_628, SYNOPSYS_UNCONNECTED_629, SYNOPSYS_UNCONNECTED_630, SYNOPSYS_UNCONNECTED_631, SYNOPSYS_UNCONNECTED_632, SYNOPSYS_UNCONNECTED_633, SYNOPSYS_UNCONNECTED_634, SYNOPSYS_UNCONNECTED_635, SYNOPSYS_UNCONNECTED_636, SYNOPSYS_UNCONNECTED_637, SYNOPSYS_UNCONNECTED_638, SYNOPSYS_UNCONNECTED_639, SYNOPSYS_UNCONNECTED_640, SYNOPSYS_UNCONNECTED_641, SYNOPSYS_UNCONNECTED_642, SYNOPSYS_UNCONNECTED_643, SYNOPSYS_UNCONNECTED_644, SYNOPSYS_UNCONNECTED_645, SYNOPSYS_UNCONNECTED_646, SYNOPSYS_UNCONNECTED_647, SYNOPSYS_UNCONNECTED_648, SYNOPSYS_UNCONNECTED_649, SYNOPSYS_UNCONNECTED_650, SYNOPSYS_UNCONNECTED_651, SYNOPSYS_UNCONNECTED_652, SYNOPSYS_UNCONNECTED_653, SYNOPSYS_UNCONNECTED_654, SYNOPSYS_UNCONNECTED_655, SYNOPSYS_UNCONNECTED_656, SYNOPSYS_UNCONNECTED_657, SYNOPSYS_UNCONNECTED_658, SYNOPSYS_UNCONNECTED_659, SYNOPSYS_UNCONNECTED_660, SYNOPSYS_UNCONNECTED_661, SYNOPSYS_UNCONNECTED_662, SYNOPSYS_UNCONNECTED_663, SYNOPSYS_UNCONNECTED_664, SYNOPSYS_UNCONNECTED_665, SYNOPSYS_UNCONNECTED_666, SYNOPSYS_UNCONNECTED_667, SYNOPSYS_UNCONNECTED_668, SYNOPSYS_UNCONNECTED_669, SYNOPSYS_UNCONNECTED_670, SYNOPSYS_UNCONNECTED_671, SYNOPSYS_UNCONNECTED_672, SYNOPSYS_UNCONNECTED_673, SYNOPSYS_UNCONNECTED_674, SYNOPSYS_UNCONNECTED_675, SYNOPSYS_UNCONNECTED_676, SYNOPSYS_UNCONNECTED_677, SYNOPSYS_UNCONNECTED_678, SYNOPSYS_UNCONNECTED_679, SYNOPSYS_UNCONNECTED_680, SYNOPSYS_UNCONNECTED_681, SYNOPSYS_UNCONNECTED_682, SYNOPSYS_UNCONNECTED_683, SYNOPSYS_UNCONNECTED_684, SYNOPSYS_UNCONNECTED_685, SYNOPSYS_UNCONNECTED_686, SYNOPSYS_UNCONNECTED_687, SYNOPSYS_UNCONNECTED_688, SYNOPSYS_UNCONNECTED_689, SYNOPSYS_UNCONNECTED_690, SYNOPSYS_UNCONNECTED_691, SYNOPSYS_UNCONNECTED_692, SYNOPSYS_UNCONNECTED_693, SYNOPSYS_UNCONNECTED_694, SYNOPSYS_UNCONNECTED_695, SYNOPSYS_UNCONNECTED_696, SYNOPSYS_UNCONNECTED_697, SYNOPSYS_UNCONNECTED_698, SYNOPSYS_UNCONNECTED_699, SYNOPSYS_UNCONNECTED_700, SYNOPSYS_UNCONNECTED_701, SYNOPSYS_UNCONNECTED_702, SYNOPSYS_UNCONNECTED_703, SYNOPSYS_UNCONNECTED_704, SYNOPSYS_UNCONNECTED_705, SYNOPSYS_UNCONNECTED_706, SYNOPSYS_UNCONNECTED_707, SYNOPSYS_UNCONNECTED_708, SYNOPSYS_UNCONNECTED_709, SYNOPSYS_UNCONNECTED_710, SYNOPSYS_UNCONNECTED_711, SYNOPSYS_UNCONNECTED_712, SYNOPSYS_UNCONNECTED_713, SYNOPSYS_UNCONNECTED_714, SYNOPSYS_UNCONNECTED_715, SYNOPSYS_UNCONNECTED_716, SYNOPSYS_UNCONNECTED_717, SYNOPSYS_UNCONNECTED_718, SYNOPSYS_UNCONNECTED_719, SYNOPSYS_UNCONNECTED_720, SYNOPSYS_UNCONNECTED_721, SYNOPSYS_UNCONNECTED_722, SYNOPSYS_UNCONNECTED_723, SYNOPSYS_UNCONNECTED_724, SYNOPSYS_UNCONNECTED_725, SYNOPSYS_UNCONNECTED_726, SYNOPSYS_UNCONNECTED_727, SYNOPSYS_UNCONNECTED_728, SYNOPSYS_UNCONNECTED_729, SYNOPSYS_UNCONNECTED_730, SYNOPSYS_UNCONNECTED_731, SYNOPSYS_UNCONNECTED_732, SYNOPSYS_UNCONNECTED_733, SYNOPSYS_UNCONNECTED_734, SYNOPSYS_UNCONNECTED_735, SYNOPSYS_UNCONNECTED_736, SYNOPSYS_UNCONNECTED_737, SYNOPSYS_UNCONNECTED_738, SYNOPSYS_UNCONNECTED_739, SYNOPSYS_UNCONNECTED_740, SYNOPSYS_UNCONNECTED_741, SYNOPSYS_UNCONNECTED_742, SYNOPSYS_UNCONNECTED_743, SYNOPSYS_UNCONNECTED_744, SYNOPSYS_UNCONNECTED_745, SYNOPSYS_UNCONNECTED_746, SYNOPSYS_UNCONNECTED_747, SYNOPSYS_UNCONNECTED_748, SYNOPSYS_UNCONNECTED_749, SYNOPSYS_UNCONNECTED_750, SYNOPSYS_UNCONNECTED_751, SYNOPSYS_UNCONNECTED_752, SYNOPSYS_UNCONNECTED_753, SYNOPSYS_UNCONNECTED_754, SYNOPSYS_UNCONNECTED_755, SYNOPSYS_UNCONNECTED_756, SYNOPSYS_UNCONNECTED_757, SYNOPSYS_UNCONNECTED_758, SYNOPSYS_UNCONNECTED_759, SYNOPSYS_UNCONNECTED_760, SYNOPSYS_UNCONNECTED_761, SYNOPSYS_UNCONNECTED_762, SYNOPSYS_UNCONNECTED_763, SYNOPSYS_UNCONNECTED_764, SYNOPSYS_UNCONNECTED_765, SYNOPSYS_UNCONNECTED_766, SYNOPSYS_UNCONNECTED_767, SYNOPSYS_UNCONNECTED_768, SYNOPSYS_UNCONNECTED_769, SYNOPSYS_UNCONNECTED_770, SYNOPSYS_UNCONNECTED_771, SYNOPSYS_UNCONNECTED_772, SYNOPSYS_UNCONNECTED_773, SYNOPSYS_UNCONNECTED_774, SYNOPSYS_UNCONNECTED_775, SYNOPSYS_UNCONNECTED_776, SYNOPSYS_UNCONNECTED_777, SYNOPSYS_UNCONNECTED_778, SYNOPSYS_UNCONNECTED_779, SYNOPSYS_UNCONNECTED_780, SYNOPSYS_UNCONNECTED_781, SYNOPSYS_UNCONNECTED_782, SYNOPSYS_UNCONNECTED_783, SYNOPSYS_UNCONNECTED_784, SYNOPSYS_UNCONNECTED_785, SYNOPSYS_UNCONNECTED_786, SYNOPSYS_UNCONNECTED_787, SYNOPSYS_UNCONNECTED_788, SYNOPSYS_UNCONNECTED_789, SYNOPSYS_UNCONNECTED_790, SYNOPSYS_UNCONNECTED_791, SYNOPSYS_UNCONNECTED_792, SYNOPSYS_UNCONNECTED_793, SYNOPSYS_UNCONNECTED_794, SYNOPSYS_UNCONNECTED_795, SYNOPSYS_UNCONNECTED_796, SYNOPSYS_UNCONNECTED_797, SYNOPSYS_UNCONNECTED_798, SYNOPSYS_UNCONNECTED_799, SYNOPSYS_UNCONNECTED_800, SYNOPSYS_UNCONNECTED_801, SYNOPSYS_UNCONNECTED_802, SYNOPSYS_UNCONNECTED_803, SYNOPSYS_UNCONNECTED_804, SYNOPSYS_UNCONNECTED_805, SYNOPSYS_UNCONNECTED_806, SYNOPSYS_UNCONNECTED_807, SYNOPSYS_UNCONNECTED_808, SYNOPSYS_UNCONNECTED_809, SYNOPSYS_UNCONNECTED_810, SYNOPSYS_UNCONNECTED_811, SYNOPSYS_UNCONNECTED_812, SYNOPSYS_UNCONNECTED_813, SYNOPSYS_UNCONNECTED_814, SYNOPSYS_UNCONNECTED_815, SYNOPSYS_UNCONNECTED_816, SYNOPSYS_UNCONNECTED_817, SYNOPSYS_UNCONNECTED_818, SYNOPSYS_UNCONNECTED_819, SYNOPSYS_UNCONNECTED_820, SYNOPSYS_UNCONNECTED_821, SYNOPSYS_UNCONNECTED_822, SYNOPSYS_UNCONNECTED_823, SYNOPSYS_UNCONNECTED_824, SYNOPSYS_UNCONNECTED_825, SYNOPSYS_UNCONNECTED_826, SYNOPSYS_UNCONNECTED_827, SYNOPSYS_UNCONNECTED_828, SYNOPSYS_UNCONNECTED_829, SYNOPSYS_UNCONNECTED_830, SYNOPSYS_UNCONNECTED_831, SYNOPSYS_UNCONNECTED_832, SYNOPSYS_UNCONNECTED_833, SYNOPSYS_UNCONNECTED_834, SYNOPSYS_UNCONNECTED_835, SYNOPSYS_UNCONNECTED_836, SYNOPSYS_UNCONNECTED_837, SYNOPSYS_UNCONNECTED_838, SYNOPSYS_UNCONNECTED_839, SYNOPSYS_UNCONNECTED_840, SYNOPSYS_UNCONNECTED_841, SYNOPSYS_UNCONNECTED_842, SYNOPSYS_UNCONNECTED_843, SYNOPSYS_UNCONNECTED_844, SYNOPSYS_UNCONNECTED_845, SYNOPSYS_UNCONNECTED_846, SYNOPSYS_UNCONNECTED_847, SYNOPSYS_UNCONNECTED_848, SYNOPSYS_UNCONNECTED_849, SYNOPSYS_UNCONNECTED_850, SYNOPSYS_UNCONNECTED_851, SYNOPSYS_UNCONNECTED_852, SYNOPSYS_UNCONNECTED_853, SYNOPSYS_UNCONNECTED_854, SYNOPSYS_UNCONNECTED_855, SYNOPSYS_UNCONNECTED_856, SYNOPSYS_UNCONNECTED_857, SYNOPSYS_UNCONNECTED_858, SYNOPSYS_UNCONNECTED_859, SYNOPSYS_UNCONNECTED_860, SYNOPSYS_UNCONNECTED_861, SYNOPSYS_UNCONNECTED_862, SYNOPSYS_UNCONNECTED_863, SYNOPSYS_UNCONNECTED_864, SYNOPSYS_UNCONNECTED_865, SYNOPSYS_UNCONNECTED_866, SYNOPSYS_UNCONNECTED_867, SYNOPSYS_UNCONNECTED_868, SYNOPSYS_UNCONNECTED_869, SYNOPSYS_UNCONNECTED_870, SYNOPSYS_UNCONNECTED_871, SYNOPSYS_UNCONNECTED_872, SYNOPSYS_UNCONNECTED_873, SYNOPSYS_UNCONNECTED_874, SYNOPSYS_UNCONNECTED_875, SYNOPSYS_UNCONNECTED_876, SYNOPSYS_UNCONNECTED_877, SYNOPSYS_UNCONNECTED_878, SYNOPSYS_UNCONNECTED_879, SYNOPSYS_UNCONNECTED_880, SYNOPSYS_UNCONNECTED_881, SYNOPSYS_UNCONNECTED_882, SYNOPSYS_UNCONNECTED_883, SYNOPSYS_UNCONNECTED_884, SYNOPSYS_UNCONNECTED_885, SYNOPSYS_UNCONNECTED_886, SYNOPSYS_UNCONNECTED_887, SYNOPSYS_UNCONNECTED_888, SYNOPSYS_UNCONNECTED_889, SYNOPSYS_UNCONNECTED_890, SYNOPSYS_UNCONNECTED_891, SYNOPSYS_UNCONNECTED_892, SYNOPSYS_UNCONNECTED_893, SYNOPSYS_UNCONNECTED_894, SYNOPSYS_UNCONNECTED_895, SYNOPSYS_UNCONNECTED_896, SYNOPSYS_UNCONNECTED_897, SYNOPSYS_UNCONNECTED_898, SYNOPSYS_UNCONNECTED_899, SYNOPSYS_UNCONNECTED_900, SYNOPSYS_UNCONNECTED_901, SYNOPSYS_UNCONNECTED_902, SYNOPSYS_UNCONNECTED_903, SYNOPSYS_UNCONNECTED_904, SYNOPSYS_UNCONNECTED_905, SYNOPSYS_UNCONNECTED_906, SYNOPSYS_UNCONNECTED_907, SYNOPSYS_UNCONNECTED_908, SYNOPSYS_UNCONNECTED_909, SYNOPSYS_UNCONNECTED_910, SYNOPSYS_UNCONNECTED_911, SYNOPSYS_UNCONNECTED_912, SYNOPSYS_UNCONNECTED_913, SYNOPSYS_UNCONNECTED_914, SYNOPSYS_UNCONNECTED_915, SYNOPSYS_UNCONNECTED_916, SYNOPSYS_UNCONNECTED_917, SYNOPSYS_UNCONNECTED_918, SYNOPSYS_UNCONNECTED_919, SYNOPSYS_UNCONNECTED_920, SYNOPSYS_UNCONNECTED_921, SYNOPSYS_UNCONNECTED_922, SYNOPSYS_UNCONNECTED_923, SYNOPSYS_UNCONNECTED_924, SYNOPSYS_UNCONNECTED_925, SYNOPSYS_UNCONNECTED_926, SYNOPSYS_UNCONNECTED_927, SYNOPSYS_UNCONNECTED_928, SYNOPSYS_UNCONNECTED_929, SYNOPSYS_UNCONNECTED_930, SYNOPSYS_UNCONNECTED_931, SYNOPSYS_UNCONNECTED_932, SYNOPSYS_UNCONNECTED_933, SYNOPSYS_UNCONNECTED_934, SYNOPSYS_UNCONNECTED_935, SYNOPSYS_UNCONNECTED_936, SYNOPSYS_UNCONNECTED_937, SYNOPSYS_UNCONNECTED_938, SYNOPSYS_UNCONNECTED_939, SYNOPSYS_UNCONNECTED_940, SYNOPSYS_UNCONNECTED_941, SYNOPSYS_UNCONNECTED_942, SYNOPSYS_UNCONNECTED_943, SYNOPSYS_UNCONNECTED_944, SYNOPSYS_UNCONNECTED_945, SYNOPSYS_UNCONNECTED_946, SYNOPSYS_UNCONNECTED_947, SYNOPSYS_UNCONNECTED_948, SYNOPSYS_UNCONNECTED_949, SYNOPSYS_UNCONNECTED_950, SYNOPSYS_UNCONNECTED_951, SYNOPSYS_UNCONNECTED_952, SYNOPSYS_UNCONNECTED_953, SYNOPSYS_UNCONNECTED_954, SYNOPSYS_UNCONNECTED_955, SYNOPSYS_UNCONNECTED_956, SYNOPSYS_UNCONNECTED_957, SYNOPSYS_UNCONNECTED_958, SYNOPSYS_UNCONNECTED_959, SYNOPSYS_UNCONNECTED_960, SYNOPSYS_UNCONNECTED_961, SYNOPSYS_UNCONNECTED_962, SYNOPSYS_UNCONNECTED_963, SYNOPSYS_UNCONNECTED_964, SYNOPSYS_UNCONNECTED_965, SYNOPSYS_UNCONNECTED_966, SYNOPSYS_UNCONNECTED_967, SYNOPSYS_UNCONNECTED_968, SYNOPSYS_UNCONNECTED_969, SYNOPSYS_UNCONNECTED_970, SYNOPSYS_UNCONNECTED_971, SYNOPSYS_UNCONNECTED_972, SYNOPSYS_UNCONNECTED_973, SYNOPSYS_UNCONNECTED_974, SYNOPSYS_UNCONNECTED_975, SYNOPSYS_UNCONNECTED_976, SYNOPSYS_UNCONNECTED_977, SYNOPSYS_UNCONNECTED_978, SYNOPSYS_UNCONNECTED_979, SYNOPSYS_UNCONNECTED_980, SYNOPSYS_UNCONNECTED_981, SYNOPSYS_UNCONNECTED_982, SYNOPSYS_UNCONNECTED_983, SYNOPSYS_UNCONNECTED_984, SYNOPSYS_UNCONNECTED_985, SYNOPSYS_UNCONNECTED_986, SYNOPSYS_UNCONNECTED_987, SYNOPSYS_UNCONNECTED_988, SYNOPSYS_UNCONNECTED_989, SYNOPSYS_UNCONNECTED_990, SYNOPSYS_UNCONNECTED_991, SYNOPSYS_UNCONNECTED_992, SYNOPSYS_UNCONNECTED_993, SYNOPSYS_UNCONNECTED_994, SYNOPSYS_UNCONNECTED_995, SYNOPSYS_UNCONNECTED_996, SYNOPSYS_UNCONNECTED_997, SYNOPSYS_UNCONNECTED_998, SYNOPSYS_UNCONNECTED_999, SYNOPSYS_UNCONNECTED_1000, SYNOPSYS_UNCONNECTED_1001, SYNOPSYS_UNCONNECTED_1002, SYNOPSYS_UNCONNECTED_1003, SYNOPSYS_UNCONNECTED_1004, SYNOPSYS_UNCONNECTED_1005, SYNOPSYS_UNCONNECTED_1006, SYNOPSYS_UNCONNECTED_1007, SYNOPSYS_UNCONNECTED_1008, SYNOPSYS_UNCONNECTED_1009, SYNOPSYS_UNCONNECTED_1010, SYNOPSYS_UNCONNECTED_1011, SYNOPSYS_UNCONNECTED_1012, SYNOPSYS_UNCONNECTED_1013, SYNOPSYS_UNCONNECTED_1014, SYNOPSYS_UNCONNECTED_1015, SYNOPSYS_UNCONNECTED_1016, SYNOPSYS_UNCONNECTED_1017, SYNOPSYS_UNCONNECTED_1018, SYNOPSYS_UNCONNECTED_1019, SYNOPSYS_UNCONNECTED_1020, SYNOPSYS_UNCONNECTED_1021, SYNOPSYS_UNCONNECTED_1022, SYNOPSYS_UNCONNECTED_1023, SYNOPSYS_UNCONNECTED_1024, SYNOPSYS_UNCONNECTED_1025, SYNOPSYS_UNCONNECTED_1026, SYNOPSYS_UNCONNECTED_1027, SYNOPSYS_UNCONNECTED_1028, SYNOPSYS_UNCONNECTED_1029, SYNOPSYS_UNCONNECTED_1030, SYNOPSYS_UNCONNECTED_1031, SYNOPSYS_UNCONNECTED_1032, SYNOPSYS_UNCONNECTED_1033, SYNOPSYS_UNCONNECTED_1034, SYNOPSYS_UNCONNECTED_1035, SYNOPSYS_UNCONNECTED_1036, SYNOPSYS_UNCONNECTED_1037, SYNOPSYS_UNCONNECTED_1038, SYNOPSYS_UNCONNECTED_1039, SYNOPSYS_UNCONNECTED_1040, SYNOPSYS_UNCONNECTED_1041, SYNOPSYS_UNCONNECTED_1042, SYNOPSYS_UNCONNECTED_1043, SYNOPSYS_UNCONNECTED_1044, SYNOPSYS_UNCONNECTED_1045, SYNOPSYS_UNCONNECTED_1046, data_head_o_flat_pretrunc } = { data_i[510:0], data_i } >> { iptr_r_data, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };

endmodule



module bsg_scan_width_p8_and_p1_lo_to_hi_p1
(
  i,
  o
);

  input [7:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__7_,t_1__6_,
  t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__7_ = i[0] & 1'b1;
  assign t_1__6_ = i[1] & i[0];
  assign t_1__5_ = i[2] & i[1];
  assign t_1__4_ = i[3] & i[2];
  assign t_1__3_ = i[4] & i[3];
  assign t_1__2_ = i[5] & i[4];
  assign t_1__1_ = i[6] & i[5];
  assign t_1__0_ = i[7] & i[6];
  assign t_2__7_ = t_1__7_ & 1'b1;
  assign t_2__6_ = t_1__6_ & 1'b1;
  assign t_2__5_ = t_1__5_ & t_1__7_;
  assign t_2__4_ = t_1__4_ & t_1__6_;
  assign t_2__3_ = t_1__3_ & t_1__5_;
  assign t_2__2_ = t_1__2_ & t_1__4_;
  assign t_2__1_ = t_1__1_ & t_1__3_;
  assign t_2__0_ = t_1__0_ & t_1__2_;
  assign o[0] = t_2__7_ & 1'b1;
  assign o[1] = t_2__6_ & 1'b1;
  assign o[2] = t_2__5_ & 1'b1;
  assign o[3] = t_2__4_ & 1'b1;
  assign o[4] = t_2__3_ & t_2__7_;
  assign o[5] = t_2__2_ & t_2__6_;
  assign o[6] = t_2__1_ & t_2__5_;
  assign o[7] = t_2__0_ & t_2__4_;

endmodule



module bsg_encode_one_hot_width_p1
(
  i,
  addr_o,
  v_o
);

  input [0:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  assign v_o = i[0];
  assign addr_o[0] = 1'b0;

endmodule



module bsg_encode_one_hot_width_p2
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o,aligned_vs;
  wire v_o;
  wire [1:0] aligned_addrs;

  bsg_encode_one_hot_width_p1
  aligned_left
  (
    .i(i[0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p1
  aligned_right
  (
    .i(i[1]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[0])
  );

  assign v_o = addr_o[0] | aligned_vs[0];

endmodule



module bsg_encode_one_hot_width_p4
(
  i,
  addr_o,
  v_o
);

  input [3:0] i;
  output [1:0] addr_o;
  output v_o;
  wire [1:0] addr_o,aligned_addrs;
  wire v_o;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p2
  aligned_left
  (
    .i(i[1:0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p2
  aligned_right
  (
    .i(i[3:2]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[1])
  );

  assign v_o = addr_o[1] | aligned_vs[0];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[1];

endmodule



module bsg_encode_one_hot_width_p8
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [3:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p4
  aligned_left
  (
    .i(i[3:0]),
    .addr_o(aligned_addrs[1:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p4
  aligned_right
  (
    .i(i[7:4]),
    .addr_o(aligned_addrs[3:2]),
    .v_o(addr_o[2])
  );

  assign v_o = addr_o[2] | aligned_vs[0];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[3];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[2];

endmodule



module bsg_encode_one_hot_width_p16
(
  i,
  addr_o,
  v_o
);

  input [15:0] i;
  output [3:0] addr_o;
  output v_o;
  wire [3:0] addr_o;
  wire v_o;
  wire [5:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p8
  aligned_left
  (
    .i(i[7:0]),
    .addr_o(aligned_addrs[2:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p8
  aligned_right
  (
    .i(i[15:8]),
    .addr_o(aligned_addrs[5:3]),
    .v_o(addr_o[3])
  );

  assign v_o = addr_o[3] | aligned_vs[0];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[5];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[4];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[3];

endmodule



module bsg_encode_one_hot_width_p9
(
  i,
  addr_o,
  v_o
);

  input [8:0] i;
  output [3:0] addr_o;
  output v_o;
  wire [3:0] addr_o;
  wire v_o;

  bsg_encode_one_hot_width_p16
  unaligned_align
  (
    .i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, i }),
    .addr_o(addr_o),
    .v_o(v_o)
  );


endmodule



module bsg_thermometer_count_width_p8
(
  i,
  o
);

  input [7:0] i;
  output [3:0] o;
  wire [3:0] o;
  wire N0,N1,N2,N3,N4,N5,N6;
  wire [7:0] big_one_hot;

  bsg_encode_one_hot_width_p9
  big_encode_one_hot
  (
    .i({ i[7:7], big_one_hot }),
    .addr_o(o)
  );

  assign big_one_hot[7] = N0 & i[6];
  assign N0 = ~i[7];
  assign big_one_hot[6] = N1 & i[5];
  assign N1 = ~i[6];
  assign big_one_hot[5] = N2 & i[4];
  assign N2 = ~i[5];
  assign big_one_hot[4] = N3 & i[3];
  assign N3 = ~i[4];
  assign big_one_hot[3] = N4 & i[2];
  assign N4 = ~i[3];
  assign big_one_hot[2] = N5 & i[1];
  assign N5 = ~i[2];
  assign big_one_hot[1] = N6 & i[0];
  assign N6 = ~i[1];
  assign big_one_hot[0] = ~i[0];

endmodule



module bsg_rr_f2f_middle_width_p64_middle_meet_p8
(
  valid_head_i,
  ready_head_i,
  go_channels_o,
  go_cnt_o
);

  input [7:0] valid_head_i;
  input [7:0] ready_head_i;
  output [7:0] go_channels_o;
  output [3:0] go_cnt_o;
  wire [7:0] go_channels_o,happy_channels;
  wire [3:0] go_cnt_o;

  bsg_scan_width_p8_and_p1_lo_to_hi_p1
  and_scan
  (
    .i(happy_channels),
    .o(go_channels_o)
  );


  bsg_thermometer_count_width_p8
  genblk1_genblk1_thermo
  (
    .i(go_channels_o),
    .o(go_cnt_o)
  );

  assign happy_channels[7] = valid_head_i[7] & ready_head_i[7];
  assign happy_channels[6] = valid_head_i[6] & ready_head_i[6];
  assign happy_channels[5] = valid_head_i[5] & ready_head_i[5];
  assign happy_channels[4] = valid_head_i[4] & ready_head_i[4];
  assign happy_channels[3] = valid_head_i[3] & ready_head_i[3];
  assign happy_channels[2] = valid_head_i[2] & ready_head_i[2];
  assign happy_channels[1] = valid_head_i[1] & ready_head_i[1];
  assign happy_channels[0] = valid_head_i[0] & ready_head_i[0];

endmodule



module bsg_rotate_right_width_p8
(
  data_i,
  rot_i,
  o
);

  input [7:0] data_i;
  input [2:0] rot_i;
  output [7:0] o;
  wire [7:0] o;
  wire SYNOPSYS_UNCONNECTED_1,SYNOPSYS_UNCONNECTED_2,SYNOPSYS_UNCONNECTED_3,
  SYNOPSYS_UNCONNECTED_4,SYNOPSYS_UNCONNECTED_5,SYNOPSYS_UNCONNECTED_6,
  SYNOPSYS_UNCONNECTED_7;
  assign { SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, o } = { data_i[6:0], data_i } >> rot_i;

endmodule



module bsg_circular_ptr_slots_p8_max_add_p8
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [3:0] add_i;
  output [2:0] o;
  output [2:0] n_o;
  input clk;
  input reset_i;
  wire [2:0] n_o;
  wire N0,N1,N2,N3,N4,N5;
  reg [2:0] o;
  assign n_o = o + add_i[2:0];
  assign { N5, N4, N3 } = (N0)? { 1'b0, 1'b0, 1'b0 } : 
                          (N1)? n_o : 1'b0;
  assign N0 = reset_i;
  assign N1 = N2;
  assign N2 = ~reset_i;

  always @(posedge clk) begin
    if(1'b1) begin
      { o[2:0] } <= { N5, N4, N3 };
    end 
  end


endmodule



module bsg_rr_f2f_output_width_p64_num_out_p8_middle_meet_p8
(
  clk,
  reset,
  ready_i,
  ready_head_o,
  go_channels_i,
  go_cnt_i,
  data_head_i,
  valid_o,
  data_o
);

  input [7:0] ready_i;
  output [7:0] ready_head_o;
  input [7:0] go_channels_i;
  input [3:0] go_cnt_i;
  input [511:0] data_head_i;
  output [7:0] valid_o;
  output [511:0] data_o;
  input clk;
  input reset;
  wire [7:0] ready_head_o,valid_o;
  wire [511:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,SYNOPSYS_UNCONNECTED_1,
  SYNOPSYS_UNCONNECTED_2,SYNOPSYS_UNCONNECTED_3,SYNOPSYS_UNCONNECTED_4,
  SYNOPSYS_UNCONNECTED_5,SYNOPSYS_UNCONNECTED_6,SYNOPSYS_UNCONNECTED_7,SYNOPSYS_UNCONNECTED_8,
  SYNOPSYS_UNCONNECTED_9,SYNOPSYS_UNCONNECTED_10,SYNOPSYS_UNCONNECTED_11,
  SYNOPSYS_UNCONNECTED_12,SYNOPSYS_UNCONNECTED_13;
  wire [2:0] optr_r,optr_r_data;

  bsg_rotate_right_width_p8
  ready_rr
  (
    .data_i(ready_i),
    .rot_i(optr_r),
    .o(ready_head_o)
  );


  bsg_circular_ptr_slots_p8_max_add_p8
  c_ptr
  (
    .clk(clk),
    .reset_i(reset),
    .add_i(go_cnt_i),
    .o(optr_r),
    .n_o({ SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3 })
  );


  bsg_circular_ptr_slots_p8_max_add_p8
  c_ptr_data
  (
    .clk(clk),
    .reset_i(reset),
    .add_i(go_cnt_i),
    .o(optr_r_data),
    .n_o({ SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6 })
  );

  assign { valid_o, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13 } = { go_channels_i, go_channels_i[7:1] } << optr_r;
  assign N224 = optr_r_data[0] & optr_r_data[1];
  assign N167 = N224 & optr_r_data[2];
  assign N225 = N0 & optr_r_data[1];
  assign N0 = ~optr_r_data[0];
  assign N166 = N225 & optr_r_data[2];
  assign N226 = optr_r_data[0] & N1;
  assign N1 = ~optr_r_data[1];
  assign N165 = N226 & optr_r_data[2];
  assign N227 = N2 & N3;
  assign N2 = ~optr_r_data[0];
  assign N3 = ~optr_r_data[1];
  assign N164 = N227 & optr_r_data[2];
  assign N228 = optr_r_data[0] & optr_r_data[1];
  assign N163 = N228 & N4;
  assign N4 = ~optr_r_data[2];
  assign N229 = N5 & optr_r_data[1];
  assign N5 = ~optr_r_data[0];
  assign N162 = N229 & N6;
  assign N6 = ~optr_r_data[2];
  assign N230 = optr_r_data[0] & N7;
  assign N7 = ~optr_r_data[1];
  assign N161 = N230 & N8;
  assign N8 = ~optr_r_data[2];
  assign N231 = N9 & N10;
  assign N9 = ~optr_r_data[0];
  assign N10 = ~optr_r_data[1];
  assign N160 = N231 & N11;
  assign N11 = ~optr_r_data[2];
  assign N232 = optr_r_data[0] & optr_r_data[1];
  assign N175 = N232 & optr_r_data[2];
  assign N233 = N12 & optr_r_data[1];
  assign N12 = ~optr_r_data[0];
  assign N174 = N233 & optr_r_data[2];
  assign N234 = optr_r_data[0] & N13;
  assign N13 = ~optr_r_data[1];
  assign N173 = N234 & optr_r_data[2];
  assign N235 = N14 & N15;
  assign N14 = ~optr_r_data[0];
  assign N15 = ~optr_r_data[1];
  assign N172 = N235 & optr_r_data[2];
  assign N236 = optr_r_data[0] & optr_r_data[1];
  assign N171 = N236 & N16;
  assign N16 = ~optr_r_data[2];
  assign N237 = N17 & optr_r_data[1];
  assign N17 = ~optr_r_data[0];
  assign N170 = N237 & N18;
  assign N18 = ~optr_r_data[2];
  assign N238 = optr_r_data[0] & N19;
  assign N19 = ~optr_r_data[1];
  assign N169 = N238 & N20;
  assign N20 = ~optr_r_data[2];
  assign N239 = N21 & N22;
  assign N21 = ~optr_r_data[0];
  assign N22 = ~optr_r_data[1];
  assign N168 = N239 & N23;
  assign N23 = ~optr_r_data[2];
  assign N240 = optr_r_data[0] & optr_r_data[1];
  assign N183 = N240 & optr_r_data[2];
  assign N241 = N24 & optr_r_data[1];
  assign N24 = ~optr_r_data[0];
  assign N182 = N241 & optr_r_data[2];
  assign N242 = optr_r_data[0] & N25;
  assign N25 = ~optr_r_data[1];
  assign N181 = N242 & optr_r_data[2];
  assign N243 = N26 & N27;
  assign N26 = ~optr_r_data[0];
  assign N27 = ~optr_r_data[1];
  assign N180 = N243 & optr_r_data[2];
  assign N244 = optr_r_data[0] & optr_r_data[1];
  assign N179 = N244 & N28;
  assign N28 = ~optr_r_data[2];
  assign N245 = N29 & optr_r_data[1];
  assign N29 = ~optr_r_data[0];
  assign N178 = N245 & N30;
  assign N30 = ~optr_r_data[2];
  assign N246 = optr_r_data[0] & N31;
  assign N31 = ~optr_r_data[1];
  assign N177 = N246 & N32;
  assign N32 = ~optr_r_data[2];
  assign N247 = N33 & N34;
  assign N33 = ~optr_r_data[0];
  assign N34 = ~optr_r_data[1];
  assign N176 = N247 & N35;
  assign N35 = ~optr_r_data[2];
  assign N248 = optr_r_data[0] & optr_r_data[1];
  assign N191 = N248 & optr_r_data[2];
  assign N249 = N36 & optr_r_data[1];
  assign N36 = ~optr_r_data[0];
  assign N190 = N249 & optr_r_data[2];
  assign N250 = optr_r_data[0] & N37;
  assign N37 = ~optr_r_data[1];
  assign N189 = N250 & optr_r_data[2];
  assign N251 = N38 & N39;
  assign N38 = ~optr_r_data[0];
  assign N39 = ~optr_r_data[1];
  assign N188 = N251 & optr_r_data[2];
  assign N252 = optr_r_data[0] & optr_r_data[1];
  assign N187 = N252 & N40;
  assign N40 = ~optr_r_data[2];
  assign N253 = N41 & optr_r_data[1];
  assign N41 = ~optr_r_data[0];
  assign N186 = N253 & N42;
  assign N42 = ~optr_r_data[2];
  assign N254 = optr_r_data[0] & N43;
  assign N43 = ~optr_r_data[1];
  assign N185 = N254 & N44;
  assign N44 = ~optr_r_data[2];
  assign N255 = N45 & N46;
  assign N45 = ~optr_r_data[0];
  assign N46 = ~optr_r_data[1];
  assign N184 = N255 & N47;
  assign N47 = ~optr_r_data[2];
  assign N256 = optr_r_data[0] & optr_r_data[1];
  assign N199 = N256 & optr_r_data[2];
  assign N257 = N48 & optr_r_data[1];
  assign N48 = ~optr_r_data[0];
  assign N198 = N257 & optr_r_data[2];
  assign N258 = optr_r_data[0] & N49;
  assign N49 = ~optr_r_data[1];
  assign N197 = N258 & optr_r_data[2];
  assign N259 = N50 & N51;
  assign N50 = ~optr_r_data[0];
  assign N51 = ~optr_r_data[1];
  assign N196 = N259 & optr_r_data[2];
  assign N260 = optr_r_data[0] & optr_r_data[1];
  assign N195 = N260 & N52;
  assign N52 = ~optr_r_data[2];
  assign N261 = N53 & optr_r_data[1];
  assign N53 = ~optr_r_data[0];
  assign N194 = N261 & N54;
  assign N54 = ~optr_r_data[2];
  assign N262 = optr_r_data[0] & N55;
  assign N55 = ~optr_r_data[1];
  assign N193 = N262 & N56;
  assign N56 = ~optr_r_data[2];
  assign N263 = N57 & N58;
  assign N57 = ~optr_r_data[0];
  assign N58 = ~optr_r_data[1];
  assign N192 = N263 & N59;
  assign N59 = ~optr_r_data[2];
  assign N264 = optr_r_data[0] & optr_r_data[1];
  assign N207 = N264 & optr_r_data[2];
  assign N265 = N60 & optr_r_data[1];
  assign N60 = ~optr_r_data[0];
  assign N206 = N265 & optr_r_data[2];
  assign N266 = optr_r_data[0] & N61;
  assign N61 = ~optr_r_data[1];
  assign N205 = N266 & optr_r_data[2];
  assign N267 = N62 & N63;
  assign N62 = ~optr_r_data[0];
  assign N63 = ~optr_r_data[1];
  assign N204 = N267 & optr_r_data[2];
  assign N268 = optr_r_data[0] & optr_r_data[1];
  assign N203 = N268 & N64;
  assign N64 = ~optr_r_data[2];
  assign N269 = N65 & optr_r_data[1];
  assign N65 = ~optr_r_data[0];
  assign N202 = N269 & N66;
  assign N66 = ~optr_r_data[2];
  assign N270 = optr_r_data[0] & N67;
  assign N67 = ~optr_r_data[1];
  assign N201 = N270 & N68;
  assign N68 = ~optr_r_data[2];
  assign N271 = N69 & N70;
  assign N69 = ~optr_r_data[0];
  assign N70 = ~optr_r_data[1];
  assign N200 = N271 & N71;
  assign N71 = ~optr_r_data[2];
  assign N272 = optr_r_data[0] & optr_r_data[1];
  assign N215 = N272 & optr_r_data[2];
  assign N273 = N72 & optr_r_data[1];
  assign N72 = ~optr_r_data[0];
  assign N214 = N273 & optr_r_data[2];
  assign N274 = optr_r_data[0] & N73;
  assign N73 = ~optr_r_data[1];
  assign N213 = N274 & optr_r_data[2];
  assign N275 = N74 & N75;
  assign N74 = ~optr_r_data[0];
  assign N75 = ~optr_r_data[1];
  assign N212 = N275 & optr_r_data[2];
  assign N276 = optr_r_data[0] & optr_r_data[1];
  assign N211 = N276 & N76;
  assign N76 = ~optr_r_data[2];
  assign N277 = N77 & optr_r_data[1];
  assign N77 = ~optr_r_data[0];
  assign N210 = N277 & N78;
  assign N78 = ~optr_r_data[2];
  assign N278 = optr_r_data[0] & N79;
  assign N79 = ~optr_r_data[1];
  assign N209 = N278 & N80;
  assign N80 = ~optr_r_data[2];
  assign N279 = N81 & N82;
  assign N81 = ~optr_r_data[0];
  assign N82 = ~optr_r_data[1];
  assign N208 = N279 & N83;
  assign N83 = ~optr_r_data[2];
  assign N280 = optr_r_data[0] & optr_r_data[1];
  assign N223 = N280 & optr_r_data[2];
  assign N281 = N84 & optr_r_data[1];
  assign N84 = ~optr_r_data[0];
  assign N222 = N281 & optr_r_data[2];
  assign N282 = optr_r_data[0] & N85;
  assign N85 = ~optr_r_data[1];
  assign N221 = N282 & optr_r_data[2];
  assign N283 = N86 & N87;
  assign N86 = ~optr_r_data[0];
  assign N87 = ~optr_r_data[1];
  assign N220 = N283 & optr_r_data[2];
  assign N284 = optr_r_data[0] & optr_r_data[1];
  assign N219 = N284 & N88;
  assign N88 = ~optr_r_data[2];
  assign N285 = N89 & optr_r_data[1];
  assign N89 = ~optr_r_data[0];
  assign N218 = N285 & N90;
  assign N90 = ~optr_r_data[2];
  assign N286 = optr_r_data[0] & N91;
  assign N91 = ~optr_r_data[1];
  assign N217 = N286 & N92;
  assign N92 = ~optr_r_data[2];
  assign N287 = N93 & N94;
  assign N93 = ~optr_r_data[0];
  assign N94 = ~optr_r_data[1];
  assign N216 = N287 & N95;
  assign N95 = ~optr_r_data[2];
  assign data_o[63:0] = (N96)? data_head_i[127:64] : 
                        (N97)? data_head_i[191:128] : 
                        (N98)? data_head_i[255:192] : 
                        (N99)? data_head_i[319:256] : 
                        (N100)? data_head_i[383:320] : 
                        (N101)? data_head_i[447:384] : 
                        (N102)? data_head_i[511:448] : 
                        (N103)? data_head_i[63:0] : 1'b0;
  assign N96 = N167;
  assign N97 = N166;
  assign N98 = N165;
  assign N99 = N164;
  assign N100 = N163;
  assign N101 = N162;
  assign N102 = N161;
  assign N103 = N160;
  assign data_o[127:64] = (N104)? data_head_i[191:128] : 
                          (N105)? data_head_i[255:192] : 
                          (N106)? data_head_i[319:256] : 
                          (N107)? data_head_i[383:320] : 
                          (N108)? data_head_i[447:384] : 
                          (N109)? data_head_i[511:448] : 
                          (N110)? data_head_i[63:0] : 
                          (N111)? data_head_i[127:64] : 1'b0;
  assign N104 = N175;
  assign N105 = N174;
  assign N106 = N173;
  assign N107 = N172;
  assign N108 = N171;
  assign N109 = N170;
  assign N110 = N169;
  assign N111 = N168;
  assign data_o[191:128] = (N112)? data_head_i[255:192] : 
                           (N113)? data_head_i[319:256] : 
                           (N114)? data_head_i[383:320] : 
                           (N115)? data_head_i[447:384] : 
                           (N116)? data_head_i[511:448] : 
                           (N117)? data_head_i[63:0] : 
                           (N118)? data_head_i[127:64] : 
                           (N119)? data_head_i[191:128] : 1'b0;
  assign N112 = N183;
  assign N113 = N182;
  assign N114 = N181;
  assign N115 = N180;
  assign N116 = N179;
  assign N117 = N178;
  assign N118 = N177;
  assign N119 = N176;
  assign data_o[255:192] = (N120)? data_head_i[319:256] : 
                           (N121)? data_head_i[383:320] : 
                           (N122)? data_head_i[447:384] : 
                           (N123)? data_head_i[511:448] : 
                           (N124)? data_head_i[63:0] : 
                           (N125)? data_head_i[127:64] : 
                           (N126)? data_head_i[191:128] : 
                           (N127)? data_head_i[255:192] : 1'b0;
  assign N120 = N191;
  assign N121 = N190;
  assign N122 = N189;
  assign N123 = N188;
  assign N124 = N187;
  assign N125 = N186;
  assign N126 = N185;
  assign N127 = N184;
  assign data_o[319:256] = (N128)? data_head_i[383:320] : 
                           (N129)? data_head_i[447:384] : 
                           (N130)? data_head_i[511:448] : 
                           (N131)? data_head_i[63:0] : 
                           (N132)? data_head_i[127:64] : 
                           (N133)? data_head_i[191:128] : 
                           (N134)? data_head_i[255:192] : 
                           (N135)? data_head_i[319:256] : 1'b0;
  assign N128 = N199;
  assign N129 = N198;
  assign N130 = N197;
  assign N131 = N196;
  assign N132 = N195;
  assign N133 = N194;
  assign N134 = N193;
  assign N135 = N192;
  assign data_o[383:320] = (N136)? data_head_i[447:384] : 
                           (N137)? data_head_i[511:448] : 
                           (N138)? data_head_i[63:0] : 
                           (N139)? data_head_i[127:64] : 
                           (N140)? data_head_i[191:128] : 
                           (N141)? data_head_i[255:192] : 
                           (N142)? data_head_i[319:256] : 
                           (N143)? data_head_i[383:320] : 1'b0;
  assign N136 = N207;
  assign N137 = N206;
  assign N138 = N205;
  assign N139 = N204;
  assign N140 = N203;
  assign N141 = N202;
  assign N142 = N201;
  assign N143 = N200;
  assign data_o[447:384] = (N144)? data_head_i[511:448] : 
                           (N145)? data_head_i[63:0] : 
                           (N146)? data_head_i[127:64] : 
                           (N147)? data_head_i[191:128] : 
                           (N148)? data_head_i[255:192] : 
                           (N149)? data_head_i[319:256] : 
                           (N150)? data_head_i[383:320] : 
                           (N151)? data_head_i[447:384] : 1'b0;
  assign N144 = N215;
  assign N145 = N214;
  assign N146 = N213;
  assign N147 = N212;
  assign N148 = N211;
  assign N149 = N210;
  assign N150 = N209;
  assign N151 = N208;
  assign data_o[511:448] = (N152)? data_head_i[63:0] : 
                           (N153)? data_head_i[127:64] : 
                           (N154)? data_head_i[191:128] : 
                           (N155)? data_head_i[255:192] : 
                           (N156)? data_head_i[319:256] : 
                           (N157)? data_head_i[383:320] : 
                           (N158)? data_head_i[447:384] : 
                           (N159)? data_head_i[511:448] : 1'b0;
  assign N152 = N223;
  assign N153 = N222;
  assign N154 = N221;
  assign N155 = N220;
  assign N156 = N219;
  assign N157 = N218;
  assign N158 = N217;
  assign N159 = N216;

endmodule



module bsg_round_robin_fifo_to_fifo
(
  clk,
  reset,
  valid_i,
  data_i,
  yumi_o,
  in_top_channel_i,
  out_top_channel_i,
  valid_o,
  data_o,
  ready_i
);

  input [15:0] valid_i;
  input [1023:0] data_i;
  output [15:0] yumi_o;
  input [3:0] in_top_channel_i;
  input [2:0] out_top_channel_i;
  output [7:0] valid_o;
  output [511:0] data_o;
  input [7:0] ready_i;
  input clk;
  input reset;
  wire [15:0] yumi_o;
  wire [7:0] valid_o,go_channels;
  wire [511:0] data_o,data_o_flat,oc_7__out_chan_data_head_array;
  wire yumi_int_o_15__15_,yumi_int_o_15__14_,yumi_int_o_15__13_,yumi_int_o_15__12_,
  yumi_int_o_15__11_,yumi_int_o_15__10_,yumi_int_o_15__9_,yumi_int_o_15__8_,
  yumi_int_o_15__7_,yumi_int_o_15__6_,yumi_int_o_15__5_,yumi_int_o_15__4_,yumi_int_o_15__3_,
  yumi_int_o_15__2_,yumi_int_o_15__1_,yumi_int_o_15__0_,N0,N1,N2,N3,N4,N5,N6,N7,
  N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,
  N29,N30,N31,valid_int_o_7__7_,valid_int_o_7__6_,valid_int_o_7__5_,
  valid_int_o_7__4_,valid_int_o_7__3_,valid_int_o_7__2_,valid_int_o_7__1_,valid_int_o_7__0_,N32,
  N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,data_int_o_7__511_,
  data_int_o_7__510_,data_int_o_7__509_,data_int_o_7__508_,data_int_o_7__507_,
  data_int_o_7__506_,data_int_o_7__505_,data_int_o_7__504_,data_int_o_7__503_,
  data_int_o_7__502_,data_int_o_7__501_,data_int_o_7__500_,data_int_o_7__499_,
  data_int_o_7__498_,data_int_o_7__497_,data_int_o_7__496_,data_int_o_7__495_,data_int_o_7__494_,
  data_int_o_7__493_,data_int_o_7__492_,data_int_o_7__491_,data_int_o_7__490_,
  data_int_o_7__489_,data_int_o_7__488_,data_int_o_7__487_,data_int_o_7__486_,
  data_int_o_7__485_,data_int_o_7__484_,data_int_o_7__483_,data_int_o_7__482_,
  data_int_o_7__481_,data_int_o_7__480_,data_int_o_7__479_,data_int_o_7__478_,
  data_int_o_7__477_,data_int_o_7__476_,data_int_o_7__475_,data_int_o_7__474_,data_int_o_7__473_,
  data_int_o_7__472_,data_int_o_7__471_,data_int_o_7__470_,data_int_o_7__469_,
  data_int_o_7__468_,data_int_o_7__467_,data_int_o_7__466_,data_int_o_7__465_,
  data_int_o_7__464_,data_int_o_7__463_,data_int_o_7__462_,data_int_o_7__461_,
  data_int_o_7__460_,data_int_o_7__459_,data_int_o_7__458_,data_int_o_7__457_,data_int_o_7__456_,
  data_int_o_7__455_,data_int_o_7__454_,data_int_o_7__453_,data_int_o_7__452_,
  data_int_o_7__451_,data_int_o_7__450_,data_int_o_7__449_,data_int_o_7__448_,
  data_int_o_7__447_,data_int_o_7__446_,data_int_o_7__445_,data_int_o_7__444_,
  data_int_o_7__443_,data_int_o_7__442_,data_int_o_7__441_,data_int_o_7__440_,
  data_int_o_7__439_,data_int_o_7__438_,data_int_o_7__437_,data_int_o_7__436_,data_int_o_7__435_,
  data_int_o_7__434_,data_int_o_7__433_,data_int_o_7__432_,data_int_o_7__431_,
  data_int_o_7__430_,data_int_o_7__429_,data_int_o_7__428_,data_int_o_7__427_,
  data_int_o_7__426_,data_int_o_7__425_,data_int_o_7__424_,data_int_o_7__423_,
  data_int_o_7__422_,data_int_o_7__421_,data_int_o_7__420_,data_int_o_7__419_,
  data_int_o_7__418_,data_int_o_7__417_,data_int_o_7__416_,data_int_o_7__415_,data_int_o_7__414_,
  data_int_o_7__413_,data_int_o_7__412_,data_int_o_7__411_,data_int_o_7__410_,
  data_int_o_7__409_,data_int_o_7__408_,data_int_o_7__407_,data_int_o_7__406_,
  data_int_o_7__405_,data_int_o_7__404_,data_int_o_7__403_,data_int_o_7__402_,
  data_int_o_7__401_,data_int_o_7__400_,data_int_o_7__399_,data_int_o_7__398_,
  data_int_o_7__397_,data_int_o_7__396_,data_int_o_7__395_,data_int_o_7__394_,data_int_o_7__393_,
  data_int_o_7__392_,data_int_o_7__391_,data_int_o_7__390_,data_int_o_7__389_,
  data_int_o_7__388_,data_int_o_7__387_,data_int_o_7__386_,data_int_o_7__385_,
  data_int_o_7__384_,data_int_o_7__383_,data_int_o_7__382_,data_int_o_7__381_,
  data_int_o_7__380_,data_int_o_7__379_,data_int_o_7__378_,data_int_o_7__377_,data_int_o_7__376_,
  data_int_o_7__375_,data_int_o_7__374_,data_int_o_7__373_,data_int_o_7__372_,
  data_int_o_7__371_,data_int_o_7__370_,data_int_o_7__369_,data_int_o_7__368_,
  data_int_o_7__367_,data_int_o_7__366_,data_int_o_7__365_,data_int_o_7__364_,
  data_int_o_7__363_,data_int_o_7__362_,data_int_o_7__361_,data_int_o_7__360_,
  data_int_o_7__359_,data_int_o_7__358_,data_int_o_7__357_,data_int_o_7__356_,data_int_o_7__355_,
  data_int_o_7__354_,data_int_o_7__353_,data_int_o_7__352_,data_int_o_7__351_,
  data_int_o_7__350_,data_int_o_7__349_,data_int_o_7__348_,data_int_o_7__347_,
  data_int_o_7__346_,data_int_o_7__345_,data_int_o_7__344_,data_int_o_7__343_,
  data_int_o_7__342_,data_int_o_7__341_,data_int_o_7__340_,data_int_o_7__339_,
  data_int_o_7__338_,data_int_o_7__337_,data_int_o_7__336_,data_int_o_7__335_,data_int_o_7__334_,
  data_int_o_7__333_,data_int_o_7__332_,data_int_o_7__331_,data_int_o_7__330_,
  data_int_o_7__329_,data_int_o_7__328_,data_int_o_7__327_,data_int_o_7__326_,
  data_int_o_7__325_,data_int_o_7__324_,data_int_o_7__323_,data_int_o_7__322_,
  data_int_o_7__321_,data_int_o_7__320_,data_int_o_7__319_,data_int_o_7__318_,
  data_int_o_7__317_,data_int_o_7__316_,data_int_o_7__315_,data_int_o_7__314_,data_int_o_7__313_,
  data_int_o_7__312_,data_int_o_7__311_,data_int_o_7__310_,data_int_o_7__309_,
  data_int_o_7__308_,data_int_o_7__307_,data_int_o_7__306_,data_int_o_7__305_,
  data_int_o_7__304_,data_int_o_7__303_,data_int_o_7__302_,data_int_o_7__301_,
  data_int_o_7__300_,data_int_o_7__299_,data_int_o_7__298_,data_int_o_7__297_,data_int_o_7__296_,
  data_int_o_7__295_,data_int_o_7__294_,data_int_o_7__293_,data_int_o_7__292_,
  data_int_o_7__291_,data_int_o_7__290_,data_int_o_7__289_,data_int_o_7__288_,
  data_int_o_7__287_,data_int_o_7__286_,data_int_o_7__285_,data_int_o_7__284_,
  data_int_o_7__283_,data_int_o_7__282_,data_int_o_7__281_,data_int_o_7__280_,
  data_int_o_7__279_,data_int_o_7__278_,data_int_o_7__277_,data_int_o_7__276_,data_int_o_7__275_,
  data_int_o_7__274_,data_int_o_7__273_,data_int_o_7__272_,data_int_o_7__271_,
  data_int_o_7__270_,data_int_o_7__269_,data_int_o_7__268_,data_int_o_7__267_,
  data_int_o_7__266_,data_int_o_7__265_,data_int_o_7__264_,data_int_o_7__263_,
  data_int_o_7__262_,data_int_o_7__261_,data_int_o_7__260_,data_int_o_7__259_,
  data_int_o_7__258_,data_int_o_7__257_,data_int_o_7__256_,data_int_o_7__255_,data_int_o_7__254_,
  data_int_o_7__253_,data_int_o_7__252_,data_int_o_7__251_,data_int_o_7__250_,
  data_int_o_7__249_,data_int_o_7__248_,data_int_o_7__247_,data_int_o_7__246_,
  data_int_o_7__245_,data_int_o_7__244_,data_int_o_7__243_,data_int_o_7__242_,
  data_int_o_7__241_,data_int_o_7__240_,data_int_o_7__239_,data_int_o_7__238_,
  data_int_o_7__237_,data_int_o_7__236_,data_int_o_7__235_,data_int_o_7__234_,data_int_o_7__233_,
  data_int_o_7__232_,data_int_o_7__231_,data_int_o_7__230_,data_int_o_7__229_,
  data_int_o_7__228_,data_int_o_7__227_,data_int_o_7__226_,data_int_o_7__225_,
  data_int_o_7__224_,data_int_o_7__223_,data_int_o_7__222_,data_int_o_7__221_,
  data_int_o_7__220_,data_int_o_7__219_,data_int_o_7__218_,data_int_o_7__217_,data_int_o_7__216_,
  data_int_o_7__215_,data_int_o_7__214_,data_int_o_7__213_,data_int_o_7__212_,
  data_int_o_7__211_,data_int_o_7__210_,data_int_o_7__209_,data_int_o_7__208_,
  data_int_o_7__207_,data_int_o_7__206_,data_int_o_7__205_,data_int_o_7__204_,
  data_int_o_7__203_,data_int_o_7__202_,data_int_o_7__201_,data_int_o_7__200_,
  data_int_o_7__199_,data_int_o_7__198_,data_int_o_7__197_,data_int_o_7__196_,data_int_o_7__195_,
  data_int_o_7__194_,data_int_o_7__193_,data_int_o_7__192_,data_int_o_7__191_,
  data_int_o_7__190_,data_int_o_7__189_,data_int_o_7__188_,data_int_o_7__187_,
  data_int_o_7__186_,data_int_o_7__185_,data_int_o_7__184_,data_int_o_7__183_,
  data_int_o_7__182_,data_int_o_7__181_,data_int_o_7__180_,data_int_o_7__179_,
  data_int_o_7__178_,data_int_o_7__177_,data_int_o_7__176_,data_int_o_7__175_,data_int_o_7__174_,
  data_int_o_7__173_,data_int_o_7__172_,data_int_o_7__171_,data_int_o_7__170_,
  data_int_o_7__169_,data_int_o_7__168_,data_int_o_7__167_,data_int_o_7__166_,
  data_int_o_7__165_,data_int_o_7__164_,data_int_o_7__163_,data_int_o_7__162_,
  data_int_o_7__161_,data_int_o_7__160_,data_int_o_7__159_,data_int_o_7__158_,
  data_int_o_7__157_,data_int_o_7__156_,data_int_o_7__155_,data_int_o_7__154_,data_int_o_7__153_,
  data_int_o_7__152_,data_int_o_7__151_,data_int_o_7__150_,data_int_o_7__149_,
  data_int_o_7__148_,data_int_o_7__147_,data_int_o_7__146_,data_int_o_7__145_,
  data_int_o_7__144_,data_int_o_7__143_,data_int_o_7__142_,data_int_o_7__141_,
  data_int_o_7__140_,data_int_o_7__139_,data_int_o_7__138_,data_int_o_7__137_,data_int_o_7__136_,
  data_int_o_7__135_,data_int_o_7__134_,data_int_o_7__133_,data_int_o_7__132_,
  data_int_o_7__131_,data_int_o_7__130_,data_int_o_7__129_,data_int_o_7__128_,
  data_int_o_7__127_,data_int_o_7__126_,data_int_o_7__125_,data_int_o_7__124_,
  data_int_o_7__123_,data_int_o_7__122_,data_int_o_7__121_,data_int_o_7__120_,
  data_int_o_7__119_,data_int_o_7__118_,data_int_o_7__117_,data_int_o_7__116_,data_int_o_7__115_,
  data_int_o_7__114_,data_int_o_7__113_,data_int_o_7__112_,data_int_o_7__111_,
  data_int_o_7__110_,data_int_o_7__109_,data_int_o_7__108_,data_int_o_7__107_,
  data_int_o_7__106_,data_int_o_7__105_,data_int_o_7__104_,data_int_o_7__103_,
  data_int_o_7__102_,data_int_o_7__101_,data_int_o_7__100_,data_int_o_7__99_,data_int_o_7__98_,
  data_int_o_7__97_,data_int_o_7__96_,data_int_o_7__95_,data_int_o_7__94_,
  data_int_o_7__93_,data_int_o_7__92_,data_int_o_7__91_,data_int_o_7__90_,
  data_int_o_7__89_,data_int_o_7__88_,data_int_o_7__87_,data_int_o_7__86_,data_int_o_7__85_,
  data_int_o_7__84_,data_int_o_7__83_,data_int_o_7__82_,data_int_o_7__81_,
  data_int_o_7__80_,data_int_o_7__79_,data_int_o_7__78_,data_int_o_7__77_,data_int_o_7__76_,
  data_int_o_7__75_,data_int_o_7__74_,data_int_o_7__73_,data_int_o_7__72_,
  data_int_o_7__71_,data_int_o_7__70_,data_int_o_7__69_,data_int_o_7__68_,data_int_o_7__67_,
  data_int_o_7__66_,data_int_o_7__65_,data_int_o_7__64_,data_int_o_7__63_,
  data_int_o_7__62_,data_int_o_7__61_,data_int_o_7__60_,data_int_o_7__59_,data_int_o_7__58_,
  data_int_o_7__57_,data_int_o_7__56_,data_int_o_7__55_,data_int_o_7__54_,
  data_int_o_7__53_,data_int_o_7__52_,data_int_o_7__51_,data_int_o_7__50_,
  data_int_o_7__49_,data_int_o_7__48_,data_int_o_7__47_,data_int_o_7__46_,data_int_o_7__45_,
  data_int_o_7__44_,data_int_o_7__43_,data_int_o_7__42_,data_int_o_7__41_,
  data_int_o_7__40_,data_int_o_7__39_,data_int_o_7__38_,data_int_o_7__37_,data_int_o_7__36_,
  data_int_o_7__35_,data_int_o_7__34_,data_int_o_7__33_,data_int_o_7__32_,
  data_int_o_7__31_,data_int_o_7__30_,data_int_o_7__29_,data_int_o_7__28_,data_int_o_7__27_,
  data_int_o_7__26_,data_int_o_7__25_,data_int_o_7__24_,data_int_o_7__23_,
  data_int_o_7__22_,data_int_o_7__21_,data_int_o_7__20_,data_int_o_7__19_,data_int_o_7__18_,
  data_int_o_7__17_,data_int_o_7__16_,data_int_o_7__15_,data_int_o_7__14_,
  data_int_o_7__13_,data_int_o_7__12_,data_int_o_7__11_,data_int_o_7__10_,
  data_int_o_7__9_,data_int_o_7__8_,data_int_o_7__7_,data_int_o_7__6_,data_int_o_7__5_,
  data_int_o_7__4_,data_int_o_7__3_,data_int_o_7__2_,data_int_o_7__1_,data_int_o_7__0_,N47,
  N48,N49,N50,N51,N52,N53,N54,data_head_15__511_,data_head_15__510_,
  data_head_15__509_,data_head_15__508_,data_head_15__507_,data_head_15__506_,data_head_15__505_,
  data_head_15__504_,data_head_15__503_,data_head_15__502_,data_head_15__501_,
  data_head_15__500_,data_head_15__499_,data_head_15__498_,data_head_15__497_,
  data_head_15__496_,data_head_15__495_,data_head_15__494_,data_head_15__493_,
  data_head_15__492_,data_head_15__491_,data_head_15__490_,data_head_15__489_,
  data_head_15__488_,data_head_15__487_,data_head_15__486_,data_head_15__485_,data_head_15__484_,
  data_head_15__483_,data_head_15__482_,data_head_15__481_,data_head_15__480_,
  data_head_15__479_,data_head_15__478_,data_head_15__477_,data_head_15__476_,
  data_head_15__475_,data_head_15__474_,data_head_15__473_,data_head_15__472_,
  data_head_15__471_,data_head_15__470_,data_head_15__469_,data_head_15__468_,
  data_head_15__467_,data_head_15__466_,data_head_15__465_,data_head_15__464_,data_head_15__463_,
  data_head_15__462_,data_head_15__461_,data_head_15__460_,data_head_15__459_,
  data_head_15__458_,data_head_15__457_,data_head_15__456_,data_head_15__455_,
  data_head_15__454_,data_head_15__453_,data_head_15__452_,data_head_15__451_,
  data_head_15__450_,data_head_15__449_,data_head_15__448_,data_head_15__447_,data_head_15__446_,
  data_head_15__445_,data_head_15__444_,data_head_15__443_,data_head_15__442_,
  data_head_15__441_,data_head_15__440_,data_head_15__439_,data_head_15__438_,
  data_head_15__437_,data_head_15__436_,data_head_15__435_,data_head_15__434_,
  data_head_15__433_,data_head_15__432_,data_head_15__431_,data_head_15__430_,
  data_head_15__429_,data_head_15__428_,data_head_15__427_,data_head_15__426_,data_head_15__425_,
  data_head_15__424_,data_head_15__423_,data_head_15__422_,data_head_15__421_,
  data_head_15__420_,data_head_15__419_,data_head_15__418_,data_head_15__417_,
  data_head_15__416_,data_head_15__415_,data_head_15__414_,data_head_15__413_,
  data_head_15__412_,data_head_15__411_,data_head_15__410_,data_head_15__409_,
  data_head_15__408_,data_head_15__407_,data_head_15__406_,data_head_15__405_,data_head_15__404_,
  data_head_15__403_,data_head_15__402_,data_head_15__401_,data_head_15__400_,
  data_head_15__399_,data_head_15__398_,data_head_15__397_,data_head_15__396_,
  data_head_15__395_,data_head_15__394_,data_head_15__393_,data_head_15__392_,
  data_head_15__391_,data_head_15__390_,data_head_15__389_,data_head_15__388_,
  data_head_15__387_,data_head_15__386_,data_head_15__385_,data_head_15__384_,data_head_15__383_,
  data_head_15__382_,data_head_15__381_,data_head_15__380_,data_head_15__379_,
  data_head_15__378_,data_head_15__377_,data_head_15__376_,data_head_15__375_,
  data_head_15__374_,data_head_15__373_,data_head_15__372_,data_head_15__371_,
  data_head_15__370_,data_head_15__369_,data_head_15__368_,data_head_15__367_,data_head_15__366_,
  data_head_15__365_,data_head_15__364_,data_head_15__363_,data_head_15__362_,
  data_head_15__361_,data_head_15__360_,data_head_15__359_,data_head_15__358_,
  data_head_15__357_,data_head_15__356_,data_head_15__355_,data_head_15__354_,
  data_head_15__353_,data_head_15__352_,data_head_15__351_,data_head_15__350_,
  data_head_15__349_,data_head_15__348_,data_head_15__347_,data_head_15__346_,data_head_15__345_,
  data_head_15__344_,data_head_15__343_,data_head_15__342_,data_head_15__341_,
  data_head_15__340_,data_head_15__339_,data_head_15__338_,data_head_15__337_,
  data_head_15__336_,data_head_15__335_,data_head_15__334_,data_head_15__333_,
  data_head_15__332_,data_head_15__331_,data_head_15__330_,data_head_15__329_,
  data_head_15__328_,data_head_15__327_,data_head_15__326_,data_head_15__325_,data_head_15__324_,
  data_head_15__323_,data_head_15__322_,data_head_15__321_,data_head_15__320_,
  data_head_15__319_,data_head_15__318_,data_head_15__317_,data_head_15__316_,
  data_head_15__315_,data_head_15__314_,data_head_15__313_,data_head_15__312_,
  data_head_15__311_,data_head_15__310_,data_head_15__309_,data_head_15__308_,
  data_head_15__307_,data_head_15__306_,data_head_15__305_,data_head_15__304_,data_head_15__303_,
  data_head_15__302_,data_head_15__301_,data_head_15__300_,data_head_15__299_,
  data_head_15__298_,data_head_15__297_,data_head_15__296_,data_head_15__295_,
  data_head_15__294_,data_head_15__293_,data_head_15__292_,data_head_15__291_,
  data_head_15__290_,data_head_15__289_,data_head_15__288_,data_head_15__287_,data_head_15__286_,
  data_head_15__285_,data_head_15__284_,data_head_15__283_,data_head_15__282_,
  data_head_15__281_,data_head_15__280_,data_head_15__279_,data_head_15__278_,
  data_head_15__277_,data_head_15__276_,data_head_15__275_,data_head_15__274_,
  data_head_15__273_,data_head_15__272_,data_head_15__271_,data_head_15__270_,
  data_head_15__269_,data_head_15__268_,data_head_15__267_,data_head_15__266_,data_head_15__265_,
  data_head_15__264_,data_head_15__263_,data_head_15__262_,data_head_15__261_,
  data_head_15__260_,data_head_15__259_,data_head_15__258_,data_head_15__257_,
  data_head_15__256_,data_head_15__255_,data_head_15__254_,data_head_15__253_,
  data_head_15__252_,data_head_15__251_,data_head_15__250_,data_head_15__249_,
  data_head_15__248_,data_head_15__247_,data_head_15__246_,data_head_15__245_,data_head_15__244_,
  data_head_15__243_,data_head_15__242_,data_head_15__241_,data_head_15__240_,
  data_head_15__239_,data_head_15__238_,data_head_15__237_,data_head_15__236_,
  data_head_15__235_,data_head_15__234_,data_head_15__233_,data_head_15__232_,
  data_head_15__231_,data_head_15__230_,data_head_15__229_,data_head_15__228_,
  data_head_15__227_,data_head_15__226_,data_head_15__225_,data_head_15__224_,data_head_15__223_,
  data_head_15__222_,data_head_15__221_,data_head_15__220_,data_head_15__219_,
  data_head_15__218_,data_head_15__217_,data_head_15__216_,data_head_15__215_,
  data_head_15__214_,data_head_15__213_,data_head_15__212_,data_head_15__211_,
  data_head_15__210_,data_head_15__209_,data_head_15__208_,data_head_15__207_,data_head_15__206_,
  data_head_15__205_,data_head_15__204_,data_head_15__203_,data_head_15__202_,
  data_head_15__201_,data_head_15__200_,data_head_15__199_,data_head_15__198_,
  data_head_15__197_,data_head_15__196_,data_head_15__195_,data_head_15__194_,
  data_head_15__193_,data_head_15__192_,data_head_15__191_,data_head_15__190_,
  data_head_15__189_,data_head_15__188_,data_head_15__187_,data_head_15__186_,data_head_15__185_,
  data_head_15__184_,data_head_15__183_,data_head_15__182_,data_head_15__181_,
  data_head_15__180_,data_head_15__179_,data_head_15__178_,data_head_15__177_,
  data_head_15__176_,data_head_15__175_,data_head_15__174_,data_head_15__173_,
  data_head_15__172_,data_head_15__171_,data_head_15__170_,data_head_15__169_,
  data_head_15__168_,data_head_15__167_,data_head_15__166_,data_head_15__165_,data_head_15__164_,
  data_head_15__163_,data_head_15__162_,data_head_15__161_,data_head_15__160_,
  data_head_15__159_,data_head_15__158_,data_head_15__157_,data_head_15__156_,
  data_head_15__155_,data_head_15__154_,data_head_15__153_,data_head_15__152_,
  data_head_15__151_,data_head_15__150_,data_head_15__149_,data_head_15__148_,
  data_head_15__147_,data_head_15__146_,data_head_15__145_,data_head_15__144_,data_head_15__143_,
  data_head_15__142_,data_head_15__141_,data_head_15__140_,data_head_15__139_,
  data_head_15__138_,data_head_15__137_,data_head_15__136_,data_head_15__135_,
  data_head_15__134_,data_head_15__133_,data_head_15__132_,data_head_15__131_,
  data_head_15__130_,data_head_15__129_,data_head_15__128_,data_head_15__127_,data_head_15__126_,
  data_head_15__125_,data_head_15__124_,data_head_15__123_,data_head_15__122_,
  data_head_15__121_,data_head_15__120_,data_head_15__119_,data_head_15__118_,
  data_head_15__117_,data_head_15__116_,data_head_15__115_,data_head_15__114_,
  data_head_15__113_,data_head_15__112_,data_head_15__111_,data_head_15__110_,
  data_head_15__109_,data_head_15__108_,data_head_15__107_,data_head_15__106_,data_head_15__105_,
  data_head_15__104_,data_head_15__103_,data_head_15__102_,data_head_15__101_,
  data_head_15__100_,data_head_15__99_,data_head_15__98_,data_head_15__97_,
  data_head_15__96_,data_head_15__95_,data_head_15__94_,data_head_15__93_,data_head_15__92_,
  data_head_15__91_,data_head_15__90_,data_head_15__89_,data_head_15__88_,
  data_head_15__87_,data_head_15__86_,data_head_15__85_,data_head_15__84_,data_head_15__83_,
  data_head_15__82_,data_head_15__81_,data_head_15__80_,data_head_15__79_,
  data_head_15__78_,data_head_15__77_,data_head_15__76_,data_head_15__75_,
  data_head_15__74_,data_head_15__73_,data_head_15__72_,data_head_15__71_,data_head_15__70_,
  data_head_15__69_,data_head_15__68_,data_head_15__67_,data_head_15__66_,
  data_head_15__65_,data_head_15__64_,data_head_15__63_,data_head_15__62_,data_head_15__61_,
  data_head_15__60_,data_head_15__59_,data_head_15__58_,data_head_15__57_,
  data_head_15__56_,data_head_15__55_,data_head_15__54_,data_head_15__53_,data_head_15__52_,
  data_head_15__51_,data_head_15__50_,data_head_15__49_,data_head_15__48_,
  data_head_15__47_,data_head_15__46_,data_head_15__45_,data_head_15__44_,data_head_15__43_,
  data_head_15__42_,data_head_15__41_,data_head_15__40_,data_head_15__39_,
  data_head_15__38_,data_head_15__37_,data_head_15__36_,data_head_15__35_,
  data_head_15__34_,data_head_15__33_,data_head_15__32_,data_head_15__31_,data_head_15__30_,
  data_head_15__29_,data_head_15__28_,data_head_15__27_,data_head_15__26_,
  data_head_15__25_,data_head_15__24_,data_head_15__23_,data_head_15__22_,data_head_15__21_,
  data_head_15__20_,data_head_15__19_,data_head_15__18_,data_head_15__17_,
  data_head_15__16_,data_head_15__15_,data_head_15__14_,data_head_15__13_,data_head_15__12_,
  data_head_15__11_,data_head_15__10_,data_head_15__9_,data_head_15__8_,
  data_head_15__7_,data_head_15__6_,data_head_15__5_,data_head_15__4_,data_head_15__3_,
  data_head_15__2_,data_head_15__1_,data_head_15__0_,n_0_net_,valid_head_15__7_,
  valid_head_15__6_,valid_head_15__5_,valid_head_15__4_,valid_head_15__3_,
  valid_head_15__2_,valid_head_15__1_,valid_head_15__0_,n_2_net__7_,n_2_net__6_,n_2_net__5_,
  n_2_net__4_,n_2_net__3_,n_2_net__2_,n_2_net__1_,n_2_net__0_,n_3_net__7_,n_3_net__6_,
  n_3_net__5_,n_3_net__4_,n_3_net__3_,n_3_net__2_,n_3_net__1_,n_3_net__0_,
  ready_head_7__7_,ready_head_7__6_,ready_head_7__5_,ready_head_7__4_,ready_head_7__3_,
  ready_head_7__2_,ready_head_7__1_,ready_head_7__0_,N55,N56,N57,N58,N59,n_4_net__511_,
  n_4_net__510_,n_4_net__509_,n_4_net__508_,n_4_net__507_,n_4_net__506_,
  n_4_net__505_,n_4_net__504_,n_4_net__503_,n_4_net__502_,n_4_net__501_,n_4_net__500_,
  n_4_net__499_,n_4_net__498_,n_4_net__497_,n_4_net__496_,n_4_net__495_,n_4_net__494_,
  n_4_net__493_,n_4_net__492_,n_4_net__491_,n_4_net__490_,n_4_net__489_,
  n_4_net__488_,n_4_net__487_,n_4_net__486_,n_4_net__485_,n_4_net__484_,n_4_net__483_,
  n_4_net__482_,n_4_net__481_,n_4_net__480_,n_4_net__479_,n_4_net__478_,n_4_net__477_,
  n_4_net__476_,n_4_net__475_,n_4_net__474_,n_4_net__473_,n_4_net__472_,n_4_net__471_,
  n_4_net__470_,n_4_net__469_,n_4_net__468_,n_4_net__467_,n_4_net__466_,
  n_4_net__465_,n_4_net__464_,n_4_net__463_,n_4_net__462_,n_4_net__461_,n_4_net__460_,
  n_4_net__459_,n_4_net__458_,n_4_net__457_,n_4_net__456_,n_4_net__455_,n_4_net__454_,
  n_4_net__453_,n_4_net__452_,n_4_net__451_,n_4_net__450_,n_4_net__449_,
  n_4_net__448_,n_4_net__447_,n_4_net__446_,n_4_net__445_,n_4_net__444_,n_4_net__443_,
  n_4_net__442_,n_4_net__441_,n_4_net__440_,n_4_net__439_,n_4_net__438_,n_4_net__437_,
  n_4_net__436_,n_4_net__435_,n_4_net__434_,n_4_net__433_,n_4_net__432_,n_4_net__431_,
  n_4_net__430_,n_4_net__429_,n_4_net__428_,n_4_net__427_,n_4_net__426_,
  n_4_net__425_,n_4_net__424_,n_4_net__423_,n_4_net__422_,n_4_net__421_,n_4_net__420_,
  n_4_net__419_,n_4_net__418_,n_4_net__417_,n_4_net__416_,n_4_net__415_,n_4_net__414_,
  n_4_net__413_,n_4_net__412_,n_4_net__411_,n_4_net__410_,n_4_net__409_,
  n_4_net__408_,n_4_net__407_,n_4_net__406_,n_4_net__405_,n_4_net__404_,n_4_net__403_,
  n_4_net__402_,n_4_net__401_,n_4_net__400_,n_4_net__399_,n_4_net__398_,n_4_net__397_,
  n_4_net__396_,n_4_net__395_,n_4_net__394_,n_4_net__393_,n_4_net__392_,n_4_net__391_,
  n_4_net__390_,n_4_net__389_,n_4_net__388_,n_4_net__387_,n_4_net__386_,
  n_4_net__385_,n_4_net__384_,n_4_net__383_,n_4_net__382_,n_4_net__381_,n_4_net__380_,
  n_4_net__379_,n_4_net__378_,n_4_net__377_,n_4_net__376_,n_4_net__375_,n_4_net__374_,
  n_4_net__373_,n_4_net__372_,n_4_net__371_,n_4_net__370_,n_4_net__369_,
  n_4_net__368_,n_4_net__367_,n_4_net__366_,n_4_net__365_,n_4_net__364_,n_4_net__363_,
  n_4_net__362_,n_4_net__361_,n_4_net__360_,n_4_net__359_,n_4_net__358_,n_4_net__357_,
  n_4_net__356_,n_4_net__355_,n_4_net__354_,n_4_net__353_,n_4_net__352_,n_4_net__351_,
  n_4_net__350_,n_4_net__349_,n_4_net__348_,n_4_net__347_,n_4_net__346_,
  n_4_net__345_,n_4_net__344_,n_4_net__343_,n_4_net__342_,n_4_net__341_,n_4_net__340_,
  n_4_net__339_,n_4_net__338_,n_4_net__337_,n_4_net__336_,n_4_net__335_,n_4_net__334_,
  n_4_net__333_,n_4_net__332_,n_4_net__331_,n_4_net__330_,n_4_net__329_,
  n_4_net__328_,n_4_net__327_,n_4_net__326_,n_4_net__325_,n_4_net__324_,n_4_net__323_,
  n_4_net__322_,n_4_net__321_,n_4_net__320_,n_4_net__319_,n_4_net__318_,n_4_net__317_,
  n_4_net__316_,n_4_net__315_,n_4_net__314_,n_4_net__313_,n_4_net__312_,n_4_net__311_,
  n_4_net__310_,n_4_net__309_,n_4_net__308_,n_4_net__307_,n_4_net__306_,
  n_4_net__305_,n_4_net__304_,n_4_net__303_,n_4_net__302_,n_4_net__301_,n_4_net__300_,
  n_4_net__299_,n_4_net__298_,n_4_net__297_,n_4_net__296_,n_4_net__295_,n_4_net__294_,
  n_4_net__293_,n_4_net__292_,n_4_net__291_,n_4_net__290_,n_4_net__289_,
  n_4_net__288_,n_4_net__287_,n_4_net__286_,n_4_net__285_,n_4_net__284_,n_4_net__283_,
  n_4_net__282_,n_4_net__281_,n_4_net__280_,n_4_net__279_,n_4_net__278_,n_4_net__277_,
  n_4_net__276_,n_4_net__275_,n_4_net__274_,n_4_net__273_,n_4_net__272_,n_4_net__271_,
  n_4_net__270_,n_4_net__269_,n_4_net__268_,n_4_net__267_,n_4_net__266_,
  n_4_net__265_,n_4_net__264_,n_4_net__263_,n_4_net__262_,n_4_net__261_,n_4_net__260_,
  n_4_net__259_,n_4_net__258_,n_4_net__257_,n_4_net__256_,n_4_net__255_,n_4_net__254_,
  n_4_net__253_,n_4_net__252_,n_4_net__251_,n_4_net__250_,n_4_net__249_,
  n_4_net__248_,n_4_net__247_,n_4_net__246_,n_4_net__245_,n_4_net__244_,n_4_net__243_,
  n_4_net__242_,n_4_net__241_,n_4_net__240_,n_4_net__239_,n_4_net__238_,n_4_net__237_,
  n_4_net__236_,n_4_net__235_,n_4_net__234_,n_4_net__233_,n_4_net__232_,n_4_net__231_,
  n_4_net__230_,n_4_net__229_,n_4_net__228_,n_4_net__227_,n_4_net__226_,
  n_4_net__225_,n_4_net__224_,n_4_net__223_,n_4_net__222_,n_4_net__221_,n_4_net__220_,
  n_4_net__219_,n_4_net__218_,n_4_net__217_,n_4_net__216_,n_4_net__215_,n_4_net__214_,
  n_4_net__213_,n_4_net__212_,n_4_net__211_,n_4_net__210_,n_4_net__209_,
  n_4_net__208_,n_4_net__207_,n_4_net__206_,n_4_net__205_,n_4_net__204_,n_4_net__203_,
  n_4_net__202_,n_4_net__201_,n_4_net__200_,n_4_net__199_,n_4_net__198_,n_4_net__197_,
  n_4_net__196_,n_4_net__195_,n_4_net__194_,n_4_net__193_,n_4_net__192_,n_4_net__191_,
  n_4_net__190_,n_4_net__189_,n_4_net__188_,n_4_net__187_,n_4_net__186_,
  n_4_net__185_,n_4_net__184_,n_4_net__183_,n_4_net__182_,n_4_net__181_,n_4_net__180_,
  n_4_net__179_,n_4_net__178_,n_4_net__177_,n_4_net__176_,n_4_net__175_,n_4_net__174_,
  n_4_net__173_,n_4_net__172_,n_4_net__171_,n_4_net__170_,n_4_net__169_,
  n_4_net__168_,n_4_net__167_,n_4_net__166_,n_4_net__165_,n_4_net__164_,n_4_net__163_,
  n_4_net__162_,n_4_net__161_,n_4_net__160_,n_4_net__159_,n_4_net__158_,n_4_net__157_,
  n_4_net__156_,n_4_net__155_,n_4_net__154_,n_4_net__153_,n_4_net__152_,n_4_net__151_,
  n_4_net__150_,n_4_net__149_,n_4_net__148_,n_4_net__147_,n_4_net__146_,
  n_4_net__145_,n_4_net__144_,n_4_net__143_,n_4_net__142_,n_4_net__141_,n_4_net__140_,
  n_4_net__139_,n_4_net__138_,n_4_net__137_,n_4_net__136_,n_4_net__135_,n_4_net__134_,
  n_4_net__133_,n_4_net__132_,n_4_net__131_,n_4_net__130_,n_4_net__129_,
  n_4_net__128_,n_4_net__127_,n_4_net__126_,n_4_net__125_,n_4_net__124_,n_4_net__123_,
  n_4_net__122_,n_4_net__121_,n_4_net__120_,n_4_net__119_,n_4_net__118_,n_4_net__117_,
  n_4_net__116_,n_4_net__115_,n_4_net__114_,n_4_net__113_,n_4_net__112_,n_4_net__111_,
  n_4_net__110_,n_4_net__109_,n_4_net__108_,n_4_net__107_,n_4_net__106_,
  n_4_net__105_,n_4_net__104_,n_4_net__103_,n_4_net__102_,n_4_net__101_,n_4_net__100_,
  n_4_net__99_,n_4_net__98_,n_4_net__97_,n_4_net__96_,n_4_net__95_,n_4_net__94_,
  n_4_net__93_,n_4_net__92_,n_4_net__91_,n_4_net__90_,n_4_net__89_,n_4_net__88_,
  n_4_net__87_,n_4_net__86_,n_4_net__85_,n_4_net__84_,n_4_net__83_,n_4_net__82_,n_4_net__81_,
  n_4_net__80_,n_4_net__79_,n_4_net__78_,n_4_net__77_,n_4_net__76_,n_4_net__75_,
  n_4_net__74_,n_4_net__73_,n_4_net__72_,n_4_net__71_,n_4_net__70_,n_4_net__69_,
  n_4_net__68_,n_4_net__67_,n_4_net__66_,n_4_net__65_,n_4_net__64_,n_4_net__63_,
  n_4_net__62_,n_4_net__61_,n_4_net__60_,n_4_net__59_,n_4_net__58_,n_4_net__57_,
  n_4_net__56_,n_4_net__55_,n_4_net__54_,n_4_net__53_,n_4_net__52_,n_4_net__51_,
  n_4_net__50_,n_4_net__49_,n_4_net__48_,n_4_net__47_,n_4_net__46_,n_4_net__45_,
  n_4_net__44_,n_4_net__43_,n_4_net__42_,n_4_net__41_,n_4_net__40_,n_4_net__39_,n_4_net__38_,
  n_4_net__37_,n_4_net__36_,n_4_net__35_,n_4_net__34_,n_4_net__33_,n_4_net__32_,
  n_4_net__31_,n_4_net__30_,n_4_net__29_,n_4_net__28_,n_4_net__27_,n_4_net__26_,
  n_4_net__25_,n_4_net__24_,n_4_net__23_,n_4_net__22_,n_4_net__21_,n_4_net__20_,
  n_4_net__19_,n_4_net__18_,n_4_net__17_,n_4_net__16_,n_4_net__15_,n_4_net__14_,
  n_4_net__13_,n_4_net__12_,n_4_net__11_,n_4_net__10_,n_4_net__9_,n_4_net__8_,n_4_net__7_,
  n_4_net__6_,n_4_net__5_,n_4_net__4_,n_4_net__3_,n_4_net__2_,n_4_net__1_,
  n_4_net__0_,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,n_5_net_,N76,
  N77,N78,N79,N80,N81,N82;
  wire [3:0] go_cnt;
  assign yumi_o[15] = (N16)? 1'b0 : 
                      (N18)? 1'b0 : 
                      (N20)? 1'b0 : 
                      (N22)? 1'b0 : 
                      (N24)? 1'b0 : 
                      (N26)? 1'b0 : 
                      (N28)? 1'b0 : 
                      (N30)? 1'b0 : 
                      (N17)? 1'b0 : 
                      (N19)? 1'b0 : 
                      (N21)? 1'b0 : 
                      (N23)? 1'b0 : 
                      (N25)? 1'b0 : 
                      (N27)? 1'b0 : 
                      (N29)? 1'b0 : 
                      (N31)? yumi_int_o_15__15_ : 1'b0;
  assign yumi_o[14] = (N16)? 1'b0 : 
                      (N18)? 1'b0 : 
                      (N20)? 1'b0 : 
                      (N22)? 1'b0 : 
                      (N24)? 1'b0 : 
                      (N26)? 1'b0 : 
                      (N28)? 1'b0 : 
                      (N30)? 1'b0 : 
                      (N17)? 1'b0 : 
                      (N19)? 1'b0 : 
                      (N21)? 1'b0 : 
                      (N23)? 1'b0 : 
                      (N25)? 1'b0 : 
                      (N27)? 1'b0 : 
                      (N29)? 1'b0 : 
                      (N31)? yumi_int_o_15__14_ : 1'b0;
  assign yumi_o[13] = (N16)? 1'b0 : 
                      (N18)? 1'b0 : 
                      (N20)? 1'b0 : 
                      (N22)? 1'b0 : 
                      (N24)? 1'b0 : 
                      (N26)? 1'b0 : 
                      (N28)? 1'b0 : 
                      (N30)? 1'b0 : 
                      (N17)? 1'b0 : 
                      (N19)? 1'b0 : 
                      (N21)? 1'b0 : 
                      (N23)? 1'b0 : 
                      (N25)? 1'b0 : 
                      (N27)? 1'b0 : 
                      (N29)? 1'b0 : 
                      (N31)? yumi_int_o_15__13_ : 1'b0;
  assign yumi_o[12] = (N16)? 1'b0 : 
                      (N18)? 1'b0 : 
                      (N20)? 1'b0 : 
                      (N22)? 1'b0 : 
                      (N24)? 1'b0 : 
                      (N26)? 1'b0 : 
                      (N28)? 1'b0 : 
                      (N30)? 1'b0 : 
                      (N17)? 1'b0 : 
                      (N19)? 1'b0 : 
                      (N21)? 1'b0 : 
                      (N23)? 1'b0 : 
                      (N25)? 1'b0 : 
                      (N27)? 1'b0 : 
                      (N29)? 1'b0 : 
                      (N31)? yumi_int_o_15__12_ : 1'b0;
  assign yumi_o[11] = (N16)? 1'b0 : 
                      (N18)? 1'b0 : 
                      (N20)? 1'b0 : 
                      (N22)? 1'b0 : 
                      (N24)? 1'b0 : 
                      (N26)? 1'b0 : 
                      (N28)? 1'b0 : 
                      (N30)? 1'b0 : 
                      (N17)? 1'b0 : 
                      (N19)? 1'b0 : 
                      (N21)? 1'b0 : 
                      (N23)? 1'b0 : 
                      (N25)? 1'b0 : 
                      (N27)? 1'b0 : 
                      (N29)? 1'b0 : 
                      (N31)? yumi_int_o_15__11_ : 1'b0;
  assign yumi_o[10] = (N16)? 1'b0 : 
                      (N18)? 1'b0 : 
                      (N20)? 1'b0 : 
                      (N22)? 1'b0 : 
                      (N24)? 1'b0 : 
                      (N26)? 1'b0 : 
                      (N28)? 1'b0 : 
                      (N30)? 1'b0 : 
                      (N17)? 1'b0 : 
                      (N19)? 1'b0 : 
                      (N21)? 1'b0 : 
                      (N23)? 1'b0 : 
                      (N25)? 1'b0 : 
                      (N27)? 1'b0 : 
                      (N29)? 1'b0 : 
                      (N31)? yumi_int_o_15__10_ : 1'b0;
  assign yumi_o[9] = (N16)? 1'b0 : 
                     (N18)? 1'b0 : 
                     (N20)? 1'b0 : 
                     (N22)? 1'b0 : 
                     (N24)? 1'b0 : 
                     (N26)? 1'b0 : 
                     (N28)? 1'b0 : 
                     (N30)? 1'b0 : 
                     (N17)? 1'b0 : 
                     (N19)? 1'b0 : 
                     (N21)? 1'b0 : 
                     (N23)? 1'b0 : 
                     (N25)? 1'b0 : 
                     (N27)? 1'b0 : 
                     (N29)? 1'b0 : 
                     (N31)? yumi_int_o_15__9_ : 1'b0;
  assign yumi_o[8] = (N16)? 1'b0 : 
                     (N18)? 1'b0 : 
                     (N20)? 1'b0 : 
                     (N22)? 1'b0 : 
                     (N24)? 1'b0 : 
                     (N26)? 1'b0 : 
                     (N28)? 1'b0 : 
                     (N30)? 1'b0 : 
                     (N17)? 1'b0 : 
                     (N19)? 1'b0 : 
                     (N21)? 1'b0 : 
                     (N23)? 1'b0 : 
                     (N25)? 1'b0 : 
                     (N27)? 1'b0 : 
                     (N29)? 1'b0 : 
                     (N31)? yumi_int_o_15__8_ : 1'b0;
  assign yumi_o[7] = (N16)? 1'b0 : 
                     (N18)? 1'b0 : 
                     (N20)? 1'b0 : 
                     (N22)? 1'b0 : 
                     (N24)? 1'b0 : 
                     (N26)? 1'b0 : 
                     (N28)? 1'b0 : 
                     (N30)? 1'b0 : 
                     (N17)? 1'b0 : 
                     (N19)? 1'b0 : 
                     (N21)? 1'b0 : 
                     (N23)? 1'b0 : 
                     (N25)? 1'b0 : 
                     (N27)? 1'b0 : 
                     (N29)? 1'b0 : 
                     (N31)? yumi_int_o_15__7_ : 1'b0;
  assign yumi_o[6] = (N16)? 1'b0 : 
                     (N18)? 1'b0 : 
                     (N20)? 1'b0 : 
                     (N22)? 1'b0 : 
                     (N24)? 1'b0 : 
                     (N26)? 1'b0 : 
                     (N28)? 1'b0 : 
                     (N30)? 1'b0 : 
                     (N17)? 1'b0 : 
                     (N19)? 1'b0 : 
                     (N21)? 1'b0 : 
                     (N23)? 1'b0 : 
                     (N25)? 1'b0 : 
                     (N27)? 1'b0 : 
                     (N29)? 1'b0 : 
                     (N31)? yumi_int_o_15__6_ : 1'b0;
  assign yumi_o[5] = (N16)? 1'b0 : 
                     (N18)? 1'b0 : 
                     (N20)? 1'b0 : 
                     (N22)? 1'b0 : 
                     (N24)? 1'b0 : 
                     (N26)? 1'b0 : 
                     (N28)? 1'b0 : 
                     (N30)? 1'b0 : 
                     (N17)? 1'b0 : 
                     (N19)? 1'b0 : 
                     (N21)? 1'b0 : 
                     (N23)? 1'b0 : 
                     (N25)? 1'b0 : 
                     (N27)? 1'b0 : 
                     (N29)? 1'b0 : 
                     (N31)? yumi_int_o_15__5_ : 1'b0;
  assign yumi_o[4] = (N16)? 1'b0 : 
                     (N18)? 1'b0 : 
                     (N20)? 1'b0 : 
                     (N22)? 1'b0 : 
                     (N24)? 1'b0 : 
                     (N26)? 1'b0 : 
                     (N28)? 1'b0 : 
                     (N30)? 1'b0 : 
                     (N17)? 1'b0 : 
                     (N19)? 1'b0 : 
                     (N21)? 1'b0 : 
                     (N23)? 1'b0 : 
                     (N25)? 1'b0 : 
                     (N27)? 1'b0 : 
                     (N29)? 1'b0 : 
                     (N31)? yumi_int_o_15__4_ : 1'b0;
  assign yumi_o[3] = (N16)? 1'b0 : 
                     (N18)? 1'b0 : 
                     (N20)? 1'b0 : 
                     (N22)? 1'b0 : 
                     (N24)? 1'b0 : 
                     (N26)? 1'b0 : 
                     (N28)? 1'b0 : 
                     (N30)? 1'b0 : 
                     (N17)? 1'b0 : 
                     (N19)? 1'b0 : 
                     (N21)? 1'b0 : 
                     (N23)? 1'b0 : 
                     (N25)? 1'b0 : 
                     (N27)? 1'b0 : 
                     (N29)? 1'b0 : 
                     (N31)? yumi_int_o_15__3_ : 1'b0;
  assign yumi_o[2] = (N16)? 1'b0 : 
                     (N18)? 1'b0 : 
                     (N20)? 1'b0 : 
                     (N22)? 1'b0 : 
                     (N24)? 1'b0 : 
                     (N26)? 1'b0 : 
                     (N28)? 1'b0 : 
                     (N30)? 1'b0 : 
                     (N17)? 1'b0 : 
                     (N19)? 1'b0 : 
                     (N21)? 1'b0 : 
                     (N23)? 1'b0 : 
                     (N25)? 1'b0 : 
                     (N27)? 1'b0 : 
                     (N29)? 1'b0 : 
                     (N31)? yumi_int_o_15__2_ : 1'b0;
  assign yumi_o[1] = (N16)? 1'b0 : 
                     (N18)? 1'b0 : 
                     (N20)? 1'b0 : 
                     (N22)? 1'b0 : 
                     (N24)? 1'b0 : 
                     (N26)? 1'b0 : 
                     (N28)? 1'b0 : 
                     (N30)? 1'b0 : 
                     (N17)? 1'b0 : 
                     (N19)? 1'b0 : 
                     (N21)? 1'b0 : 
                     (N23)? 1'b0 : 
                     (N25)? 1'b0 : 
                     (N27)? 1'b0 : 
                     (N29)? 1'b0 : 
                     (N31)? yumi_int_o_15__1_ : 1'b0;
  assign yumi_o[0] = (N16)? 1'b0 : 
                     (N18)? 1'b0 : 
                     (N20)? 1'b0 : 
                     (N22)? 1'b0 : 
                     (N24)? 1'b0 : 
                     (N26)? 1'b0 : 
                     (N28)? 1'b0 : 
                     (N30)? 1'b0 : 
                     (N17)? 1'b0 : 
                     (N19)? 1'b0 : 
                     (N21)? 1'b0 : 
                     (N23)? 1'b0 : 
                     (N25)? 1'b0 : 
                     (N27)? 1'b0 : 
                     (N29)? 1'b0 : 
                     (N31)? yumi_int_o_15__0_ : 1'b0;
  assign valid_o[7] = (N39)? 1'b0 : 
                      (N41)? 1'b0 : 
                      (N43)? 1'b0 : 
                      (N45)? 1'b0 : 
                      (N40)? 1'b0 : 
                      (N42)? 1'b0 : 
                      (N44)? 1'b0 : 
                      (N46)? valid_int_o_7__7_ : 1'b0;
  assign valid_o[6] = (N39)? 1'b0 : 
                      (N41)? 1'b0 : 
                      (N43)? 1'b0 : 
                      (N45)? 1'b0 : 
                      (N40)? 1'b0 : 
                      (N42)? 1'b0 : 
                      (N44)? 1'b0 : 
                      (N46)? valid_int_o_7__6_ : 1'b0;
  assign valid_o[5] = (N39)? 1'b0 : 
                      (N41)? 1'b0 : 
                      (N43)? 1'b0 : 
                      (N45)? 1'b0 : 
                      (N40)? 1'b0 : 
                      (N42)? 1'b0 : 
                      (N44)? 1'b0 : 
                      (N46)? valid_int_o_7__5_ : 1'b0;
  assign valid_o[4] = (N39)? 1'b0 : 
                      (N41)? 1'b0 : 
                      (N43)? 1'b0 : 
                      (N45)? 1'b0 : 
                      (N40)? 1'b0 : 
                      (N42)? 1'b0 : 
                      (N44)? 1'b0 : 
                      (N46)? valid_int_o_7__4_ : 1'b0;
  assign valid_o[3] = (N39)? 1'b0 : 
                      (N41)? 1'b0 : 
                      (N43)? 1'b0 : 
                      (N45)? 1'b0 : 
                      (N40)? 1'b0 : 
                      (N42)? 1'b0 : 
                      (N44)? 1'b0 : 
                      (N46)? valid_int_o_7__3_ : 1'b0;
  assign valid_o[2] = (N39)? 1'b0 : 
                      (N41)? 1'b0 : 
                      (N43)? 1'b0 : 
                      (N45)? 1'b0 : 
                      (N40)? 1'b0 : 
                      (N42)? 1'b0 : 
                      (N44)? 1'b0 : 
                      (N46)? valid_int_o_7__2_ : 1'b0;
  assign valid_o[1] = (N39)? 1'b0 : 
                      (N41)? 1'b0 : 
                      (N43)? 1'b0 : 
                      (N45)? 1'b0 : 
                      (N40)? 1'b0 : 
                      (N42)? 1'b0 : 
                      (N44)? 1'b0 : 
                      (N46)? valid_int_o_7__1_ : 1'b0;
  assign valid_o[0] = (N39)? 1'b0 : 
                      (N41)? 1'b0 : 
                      (N43)? 1'b0 : 
                      (N45)? 1'b0 : 
                      (N40)? 1'b0 : 
                      (N42)? 1'b0 : 
                      (N44)? 1'b0 : 
                      (N46)? valid_int_o_7__0_ : 1'b0;
  assign data_o_flat[511] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__511_ : 1'b0;
  assign data_o_flat[510] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__510_ : 1'b0;
  assign data_o_flat[509] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__509_ : 1'b0;
  assign data_o_flat[508] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__508_ : 1'b0;
  assign data_o_flat[507] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__507_ : 1'b0;
  assign data_o_flat[506] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__506_ : 1'b0;
  assign data_o_flat[505] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__505_ : 1'b0;
  assign data_o_flat[504] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__504_ : 1'b0;
  assign data_o_flat[503] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__503_ : 1'b0;
  assign data_o_flat[502] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__502_ : 1'b0;
  assign data_o_flat[501] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__501_ : 1'b0;
  assign data_o_flat[500] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__500_ : 1'b0;
  assign data_o_flat[499] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__499_ : 1'b0;
  assign data_o_flat[498] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__498_ : 1'b0;
  assign data_o_flat[497] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__497_ : 1'b0;
  assign data_o_flat[496] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__496_ : 1'b0;
  assign data_o_flat[495] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__495_ : 1'b0;
  assign data_o_flat[494] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__494_ : 1'b0;
  assign data_o_flat[493] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__493_ : 1'b0;
  assign data_o_flat[492] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__492_ : 1'b0;
  assign data_o_flat[491] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__491_ : 1'b0;
  assign data_o_flat[490] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__490_ : 1'b0;
  assign data_o_flat[489] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__489_ : 1'b0;
  assign data_o_flat[488] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__488_ : 1'b0;
  assign data_o_flat[487] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__487_ : 1'b0;
  assign data_o_flat[486] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__486_ : 1'b0;
  assign data_o_flat[485] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__485_ : 1'b0;
  assign data_o_flat[484] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__484_ : 1'b0;
  assign data_o_flat[483] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__483_ : 1'b0;
  assign data_o_flat[482] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__482_ : 1'b0;
  assign data_o_flat[481] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__481_ : 1'b0;
  assign data_o_flat[480] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__480_ : 1'b0;
  assign data_o_flat[479] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__479_ : 1'b0;
  assign data_o_flat[478] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__478_ : 1'b0;
  assign data_o_flat[477] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__477_ : 1'b0;
  assign data_o_flat[476] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__476_ : 1'b0;
  assign data_o_flat[475] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__475_ : 1'b0;
  assign data_o_flat[474] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__474_ : 1'b0;
  assign data_o_flat[473] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__473_ : 1'b0;
  assign data_o_flat[472] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__472_ : 1'b0;
  assign data_o_flat[471] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__471_ : 1'b0;
  assign data_o_flat[470] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__470_ : 1'b0;
  assign data_o_flat[469] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__469_ : 1'b0;
  assign data_o_flat[468] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__468_ : 1'b0;
  assign data_o_flat[467] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__467_ : 1'b0;
  assign data_o_flat[466] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__466_ : 1'b0;
  assign data_o_flat[465] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__465_ : 1'b0;
  assign data_o_flat[464] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__464_ : 1'b0;
  assign data_o_flat[463] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__463_ : 1'b0;
  assign data_o_flat[462] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__462_ : 1'b0;
  assign data_o_flat[461] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__461_ : 1'b0;
  assign data_o_flat[460] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__460_ : 1'b0;
  assign data_o_flat[459] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__459_ : 1'b0;
  assign data_o_flat[458] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__458_ : 1'b0;
  assign data_o_flat[457] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__457_ : 1'b0;
  assign data_o_flat[456] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__456_ : 1'b0;
  assign data_o_flat[455] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__455_ : 1'b0;
  assign data_o_flat[454] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__454_ : 1'b0;
  assign data_o_flat[453] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__453_ : 1'b0;
  assign data_o_flat[452] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__452_ : 1'b0;
  assign data_o_flat[451] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__451_ : 1'b0;
  assign data_o_flat[450] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__450_ : 1'b0;
  assign data_o_flat[449] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__449_ : 1'b0;
  assign data_o_flat[448] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__448_ : 1'b0;
  assign data_o_flat[447] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__447_ : 1'b0;
  assign data_o_flat[446] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__446_ : 1'b0;
  assign data_o_flat[445] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__445_ : 1'b0;
  assign data_o_flat[444] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__444_ : 1'b0;
  assign data_o_flat[443] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__443_ : 1'b0;
  assign data_o_flat[442] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__442_ : 1'b0;
  assign data_o_flat[441] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__441_ : 1'b0;
  assign data_o_flat[440] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__440_ : 1'b0;
  assign data_o_flat[439] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__439_ : 1'b0;
  assign data_o_flat[438] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__438_ : 1'b0;
  assign data_o_flat[437] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__437_ : 1'b0;
  assign data_o_flat[436] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__436_ : 1'b0;
  assign data_o_flat[435] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__435_ : 1'b0;
  assign data_o_flat[434] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__434_ : 1'b0;
  assign data_o_flat[433] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__433_ : 1'b0;
  assign data_o_flat[432] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__432_ : 1'b0;
  assign data_o_flat[431] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__431_ : 1'b0;
  assign data_o_flat[430] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__430_ : 1'b0;
  assign data_o_flat[429] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__429_ : 1'b0;
  assign data_o_flat[428] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__428_ : 1'b0;
  assign data_o_flat[427] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__427_ : 1'b0;
  assign data_o_flat[426] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__426_ : 1'b0;
  assign data_o_flat[425] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__425_ : 1'b0;
  assign data_o_flat[424] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__424_ : 1'b0;
  assign data_o_flat[423] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__423_ : 1'b0;
  assign data_o_flat[422] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__422_ : 1'b0;
  assign data_o_flat[421] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__421_ : 1'b0;
  assign data_o_flat[420] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__420_ : 1'b0;
  assign data_o_flat[419] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__419_ : 1'b0;
  assign data_o_flat[418] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__418_ : 1'b0;
  assign data_o_flat[417] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__417_ : 1'b0;
  assign data_o_flat[416] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__416_ : 1'b0;
  assign data_o_flat[415] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__415_ : 1'b0;
  assign data_o_flat[414] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__414_ : 1'b0;
  assign data_o_flat[413] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__413_ : 1'b0;
  assign data_o_flat[412] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__412_ : 1'b0;
  assign data_o_flat[411] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__411_ : 1'b0;
  assign data_o_flat[410] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__410_ : 1'b0;
  assign data_o_flat[409] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__409_ : 1'b0;
  assign data_o_flat[408] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__408_ : 1'b0;
  assign data_o_flat[407] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__407_ : 1'b0;
  assign data_o_flat[406] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__406_ : 1'b0;
  assign data_o_flat[405] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__405_ : 1'b0;
  assign data_o_flat[404] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__404_ : 1'b0;
  assign data_o_flat[403] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__403_ : 1'b0;
  assign data_o_flat[402] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__402_ : 1'b0;
  assign data_o_flat[401] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__401_ : 1'b0;
  assign data_o_flat[400] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__400_ : 1'b0;
  assign data_o_flat[399] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__399_ : 1'b0;
  assign data_o_flat[398] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__398_ : 1'b0;
  assign data_o_flat[397] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__397_ : 1'b0;
  assign data_o_flat[396] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__396_ : 1'b0;
  assign data_o_flat[395] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__395_ : 1'b0;
  assign data_o_flat[394] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__394_ : 1'b0;
  assign data_o_flat[393] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__393_ : 1'b0;
  assign data_o_flat[392] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__392_ : 1'b0;
  assign data_o_flat[391] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__391_ : 1'b0;
  assign data_o_flat[390] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__390_ : 1'b0;
  assign data_o_flat[389] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__389_ : 1'b0;
  assign data_o_flat[388] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__388_ : 1'b0;
  assign data_o_flat[387] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__387_ : 1'b0;
  assign data_o_flat[386] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__386_ : 1'b0;
  assign data_o_flat[385] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__385_ : 1'b0;
  assign data_o_flat[384] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__384_ : 1'b0;
  assign data_o_flat[383] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__383_ : 1'b0;
  assign data_o_flat[382] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__382_ : 1'b0;
  assign data_o_flat[381] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__381_ : 1'b0;
  assign data_o_flat[380] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__380_ : 1'b0;
  assign data_o_flat[379] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__379_ : 1'b0;
  assign data_o_flat[378] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__378_ : 1'b0;
  assign data_o_flat[377] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__377_ : 1'b0;
  assign data_o_flat[376] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__376_ : 1'b0;
  assign data_o_flat[375] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__375_ : 1'b0;
  assign data_o_flat[374] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__374_ : 1'b0;
  assign data_o_flat[373] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__373_ : 1'b0;
  assign data_o_flat[372] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__372_ : 1'b0;
  assign data_o_flat[371] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__371_ : 1'b0;
  assign data_o_flat[370] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__370_ : 1'b0;
  assign data_o_flat[369] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__369_ : 1'b0;
  assign data_o_flat[368] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__368_ : 1'b0;
  assign data_o_flat[367] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__367_ : 1'b0;
  assign data_o_flat[366] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__366_ : 1'b0;
  assign data_o_flat[365] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__365_ : 1'b0;
  assign data_o_flat[364] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__364_ : 1'b0;
  assign data_o_flat[363] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__363_ : 1'b0;
  assign data_o_flat[362] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__362_ : 1'b0;
  assign data_o_flat[361] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__361_ : 1'b0;
  assign data_o_flat[360] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__360_ : 1'b0;
  assign data_o_flat[359] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__359_ : 1'b0;
  assign data_o_flat[358] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__358_ : 1'b0;
  assign data_o_flat[357] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__357_ : 1'b0;
  assign data_o_flat[356] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__356_ : 1'b0;
  assign data_o_flat[355] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__355_ : 1'b0;
  assign data_o_flat[354] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__354_ : 1'b0;
  assign data_o_flat[353] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__353_ : 1'b0;
  assign data_o_flat[352] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__352_ : 1'b0;
  assign data_o_flat[351] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__351_ : 1'b0;
  assign data_o_flat[350] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__350_ : 1'b0;
  assign data_o_flat[349] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__349_ : 1'b0;
  assign data_o_flat[348] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__348_ : 1'b0;
  assign data_o_flat[347] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__347_ : 1'b0;
  assign data_o_flat[346] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__346_ : 1'b0;
  assign data_o_flat[345] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__345_ : 1'b0;
  assign data_o_flat[344] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__344_ : 1'b0;
  assign data_o_flat[343] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__343_ : 1'b0;
  assign data_o_flat[342] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__342_ : 1'b0;
  assign data_o_flat[341] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__341_ : 1'b0;
  assign data_o_flat[340] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__340_ : 1'b0;
  assign data_o_flat[339] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__339_ : 1'b0;
  assign data_o_flat[338] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__338_ : 1'b0;
  assign data_o_flat[337] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__337_ : 1'b0;
  assign data_o_flat[336] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__336_ : 1'b0;
  assign data_o_flat[335] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__335_ : 1'b0;
  assign data_o_flat[334] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__334_ : 1'b0;
  assign data_o_flat[333] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__333_ : 1'b0;
  assign data_o_flat[332] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__332_ : 1'b0;
  assign data_o_flat[331] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__331_ : 1'b0;
  assign data_o_flat[330] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__330_ : 1'b0;
  assign data_o_flat[329] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__329_ : 1'b0;
  assign data_o_flat[328] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__328_ : 1'b0;
  assign data_o_flat[327] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__327_ : 1'b0;
  assign data_o_flat[326] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__326_ : 1'b0;
  assign data_o_flat[325] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__325_ : 1'b0;
  assign data_o_flat[324] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__324_ : 1'b0;
  assign data_o_flat[323] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__323_ : 1'b0;
  assign data_o_flat[322] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__322_ : 1'b0;
  assign data_o_flat[321] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__321_ : 1'b0;
  assign data_o_flat[320] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__320_ : 1'b0;
  assign data_o_flat[319] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__319_ : 1'b0;
  assign data_o_flat[318] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__318_ : 1'b0;
  assign data_o_flat[317] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__317_ : 1'b0;
  assign data_o_flat[316] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__316_ : 1'b0;
  assign data_o_flat[315] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__315_ : 1'b0;
  assign data_o_flat[314] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__314_ : 1'b0;
  assign data_o_flat[313] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__313_ : 1'b0;
  assign data_o_flat[312] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__312_ : 1'b0;
  assign data_o_flat[311] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__311_ : 1'b0;
  assign data_o_flat[310] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__310_ : 1'b0;
  assign data_o_flat[309] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__309_ : 1'b0;
  assign data_o_flat[308] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__308_ : 1'b0;
  assign data_o_flat[307] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__307_ : 1'b0;
  assign data_o_flat[306] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__306_ : 1'b0;
  assign data_o_flat[305] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__305_ : 1'b0;
  assign data_o_flat[304] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__304_ : 1'b0;
  assign data_o_flat[303] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__303_ : 1'b0;
  assign data_o_flat[302] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__302_ : 1'b0;
  assign data_o_flat[301] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__301_ : 1'b0;
  assign data_o_flat[300] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__300_ : 1'b0;
  assign data_o_flat[299] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__299_ : 1'b0;
  assign data_o_flat[298] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__298_ : 1'b0;
  assign data_o_flat[297] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__297_ : 1'b0;
  assign data_o_flat[296] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__296_ : 1'b0;
  assign data_o_flat[295] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__295_ : 1'b0;
  assign data_o_flat[294] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__294_ : 1'b0;
  assign data_o_flat[293] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__293_ : 1'b0;
  assign data_o_flat[292] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__292_ : 1'b0;
  assign data_o_flat[291] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__291_ : 1'b0;
  assign data_o_flat[290] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__290_ : 1'b0;
  assign data_o_flat[289] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__289_ : 1'b0;
  assign data_o_flat[288] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__288_ : 1'b0;
  assign data_o_flat[287] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__287_ : 1'b0;
  assign data_o_flat[286] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__286_ : 1'b0;
  assign data_o_flat[285] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__285_ : 1'b0;
  assign data_o_flat[284] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__284_ : 1'b0;
  assign data_o_flat[283] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__283_ : 1'b0;
  assign data_o_flat[282] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__282_ : 1'b0;
  assign data_o_flat[281] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__281_ : 1'b0;
  assign data_o_flat[280] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__280_ : 1'b0;
  assign data_o_flat[279] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__279_ : 1'b0;
  assign data_o_flat[278] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__278_ : 1'b0;
  assign data_o_flat[277] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__277_ : 1'b0;
  assign data_o_flat[276] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__276_ : 1'b0;
  assign data_o_flat[275] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__275_ : 1'b0;
  assign data_o_flat[274] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__274_ : 1'b0;
  assign data_o_flat[273] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__273_ : 1'b0;
  assign data_o_flat[272] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__272_ : 1'b0;
  assign data_o_flat[271] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__271_ : 1'b0;
  assign data_o_flat[270] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__270_ : 1'b0;
  assign data_o_flat[269] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__269_ : 1'b0;
  assign data_o_flat[268] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__268_ : 1'b0;
  assign data_o_flat[267] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__267_ : 1'b0;
  assign data_o_flat[266] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__266_ : 1'b0;
  assign data_o_flat[265] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__265_ : 1'b0;
  assign data_o_flat[264] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__264_ : 1'b0;
  assign data_o_flat[263] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__263_ : 1'b0;
  assign data_o_flat[262] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__262_ : 1'b0;
  assign data_o_flat[261] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__261_ : 1'b0;
  assign data_o_flat[260] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__260_ : 1'b0;
  assign data_o_flat[259] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__259_ : 1'b0;
  assign data_o_flat[258] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__258_ : 1'b0;
  assign data_o_flat[257] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__257_ : 1'b0;
  assign data_o_flat[256] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__256_ : 1'b0;
  assign data_o_flat[255] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__255_ : 1'b0;
  assign data_o_flat[254] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__254_ : 1'b0;
  assign data_o_flat[253] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__253_ : 1'b0;
  assign data_o_flat[252] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__252_ : 1'b0;
  assign data_o_flat[251] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__251_ : 1'b0;
  assign data_o_flat[250] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__250_ : 1'b0;
  assign data_o_flat[249] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__249_ : 1'b0;
  assign data_o_flat[248] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__248_ : 1'b0;
  assign data_o_flat[247] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__247_ : 1'b0;
  assign data_o_flat[246] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__246_ : 1'b0;
  assign data_o_flat[245] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__245_ : 1'b0;
  assign data_o_flat[244] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__244_ : 1'b0;
  assign data_o_flat[243] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__243_ : 1'b0;
  assign data_o_flat[242] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__242_ : 1'b0;
  assign data_o_flat[241] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__241_ : 1'b0;
  assign data_o_flat[240] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__240_ : 1'b0;
  assign data_o_flat[239] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__239_ : 1'b0;
  assign data_o_flat[238] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__238_ : 1'b0;
  assign data_o_flat[237] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__237_ : 1'b0;
  assign data_o_flat[236] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__236_ : 1'b0;
  assign data_o_flat[235] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__235_ : 1'b0;
  assign data_o_flat[234] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__234_ : 1'b0;
  assign data_o_flat[233] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__233_ : 1'b0;
  assign data_o_flat[232] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__232_ : 1'b0;
  assign data_o_flat[231] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__231_ : 1'b0;
  assign data_o_flat[230] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__230_ : 1'b0;
  assign data_o_flat[229] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__229_ : 1'b0;
  assign data_o_flat[228] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__228_ : 1'b0;
  assign data_o_flat[227] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__227_ : 1'b0;
  assign data_o_flat[226] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__226_ : 1'b0;
  assign data_o_flat[225] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__225_ : 1'b0;
  assign data_o_flat[224] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__224_ : 1'b0;
  assign data_o_flat[223] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__223_ : 1'b0;
  assign data_o_flat[222] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__222_ : 1'b0;
  assign data_o_flat[221] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__221_ : 1'b0;
  assign data_o_flat[220] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__220_ : 1'b0;
  assign data_o_flat[219] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__219_ : 1'b0;
  assign data_o_flat[218] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__218_ : 1'b0;
  assign data_o_flat[217] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__217_ : 1'b0;
  assign data_o_flat[216] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__216_ : 1'b0;
  assign data_o_flat[215] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__215_ : 1'b0;
  assign data_o_flat[214] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__214_ : 1'b0;
  assign data_o_flat[213] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__213_ : 1'b0;
  assign data_o_flat[212] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__212_ : 1'b0;
  assign data_o_flat[211] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__211_ : 1'b0;
  assign data_o_flat[210] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__210_ : 1'b0;
  assign data_o_flat[209] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__209_ : 1'b0;
  assign data_o_flat[208] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__208_ : 1'b0;
  assign data_o_flat[207] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__207_ : 1'b0;
  assign data_o_flat[206] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__206_ : 1'b0;
  assign data_o_flat[205] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__205_ : 1'b0;
  assign data_o_flat[204] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__204_ : 1'b0;
  assign data_o_flat[203] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__203_ : 1'b0;
  assign data_o_flat[202] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__202_ : 1'b0;
  assign data_o_flat[201] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__201_ : 1'b0;
  assign data_o_flat[200] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__200_ : 1'b0;
  assign data_o_flat[199] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__199_ : 1'b0;
  assign data_o_flat[198] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__198_ : 1'b0;
  assign data_o_flat[197] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__197_ : 1'b0;
  assign data_o_flat[196] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__196_ : 1'b0;
  assign data_o_flat[195] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__195_ : 1'b0;
  assign data_o_flat[194] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__194_ : 1'b0;
  assign data_o_flat[193] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__193_ : 1'b0;
  assign data_o_flat[192] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__192_ : 1'b0;
  assign data_o_flat[191] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__191_ : 1'b0;
  assign data_o_flat[190] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__190_ : 1'b0;
  assign data_o_flat[189] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__189_ : 1'b0;
  assign data_o_flat[188] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__188_ : 1'b0;
  assign data_o_flat[187] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__187_ : 1'b0;
  assign data_o_flat[186] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__186_ : 1'b0;
  assign data_o_flat[185] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__185_ : 1'b0;
  assign data_o_flat[184] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__184_ : 1'b0;
  assign data_o_flat[183] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__183_ : 1'b0;
  assign data_o_flat[182] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__182_ : 1'b0;
  assign data_o_flat[181] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__181_ : 1'b0;
  assign data_o_flat[180] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__180_ : 1'b0;
  assign data_o_flat[179] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__179_ : 1'b0;
  assign data_o_flat[178] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__178_ : 1'b0;
  assign data_o_flat[177] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__177_ : 1'b0;
  assign data_o_flat[176] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__176_ : 1'b0;
  assign data_o_flat[175] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__175_ : 1'b0;
  assign data_o_flat[174] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__174_ : 1'b0;
  assign data_o_flat[173] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__173_ : 1'b0;
  assign data_o_flat[172] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__172_ : 1'b0;
  assign data_o_flat[171] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__171_ : 1'b0;
  assign data_o_flat[170] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__170_ : 1'b0;
  assign data_o_flat[169] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__169_ : 1'b0;
  assign data_o_flat[168] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__168_ : 1'b0;
  assign data_o_flat[167] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__167_ : 1'b0;
  assign data_o_flat[166] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__166_ : 1'b0;
  assign data_o_flat[165] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__165_ : 1'b0;
  assign data_o_flat[164] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__164_ : 1'b0;
  assign data_o_flat[163] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__163_ : 1'b0;
  assign data_o_flat[162] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__162_ : 1'b0;
  assign data_o_flat[161] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__161_ : 1'b0;
  assign data_o_flat[160] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__160_ : 1'b0;
  assign data_o_flat[159] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__159_ : 1'b0;
  assign data_o_flat[158] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__158_ : 1'b0;
  assign data_o_flat[157] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__157_ : 1'b0;
  assign data_o_flat[156] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__156_ : 1'b0;
  assign data_o_flat[155] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__155_ : 1'b0;
  assign data_o_flat[154] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__154_ : 1'b0;
  assign data_o_flat[153] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__153_ : 1'b0;
  assign data_o_flat[152] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__152_ : 1'b0;
  assign data_o_flat[151] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__151_ : 1'b0;
  assign data_o_flat[150] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__150_ : 1'b0;
  assign data_o_flat[149] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__149_ : 1'b0;
  assign data_o_flat[148] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__148_ : 1'b0;
  assign data_o_flat[147] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__147_ : 1'b0;
  assign data_o_flat[146] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__146_ : 1'b0;
  assign data_o_flat[145] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__145_ : 1'b0;
  assign data_o_flat[144] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__144_ : 1'b0;
  assign data_o_flat[143] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__143_ : 1'b0;
  assign data_o_flat[142] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__142_ : 1'b0;
  assign data_o_flat[141] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__141_ : 1'b0;
  assign data_o_flat[140] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__140_ : 1'b0;
  assign data_o_flat[139] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__139_ : 1'b0;
  assign data_o_flat[138] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__138_ : 1'b0;
  assign data_o_flat[137] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__137_ : 1'b0;
  assign data_o_flat[136] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__136_ : 1'b0;
  assign data_o_flat[135] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__135_ : 1'b0;
  assign data_o_flat[134] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__134_ : 1'b0;
  assign data_o_flat[133] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__133_ : 1'b0;
  assign data_o_flat[132] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__132_ : 1'b0;
  assign data_o_flat[131] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__131_ : 1'b0;
  assign data_o_flat[130] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__130_ : 1'b0;
  assign data_o_flat[129] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__129_ : 1'b0;
  assign data_o_flat[128] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__128_ : 1'b0;
  assign data_o_flat[127] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__127_ : 1'b0;
  assign data_o_flat[126] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__126_ : 1'b0;
  assign data_o_flat[125] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__125_ : 1'b0;
  assign data_o_flat[124] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__124_ : 1'b0;
  assign data_o_flat[123] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__123_ : 1'b0;
  assign data_o_flat[122] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__122_ : 1'b0;
  assign data_o_flat[121] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__121_ : 1'b0;
  assign data_o_flat[120] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__120_ : 1'b0;
  assign data_o_flat[119] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__119_ : 1'b0;
  assign data_o_flat[118] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__118_ : 1'b0;
  assign data_o_flat[117] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__117_ : 1'b0;
  assign data_o_flat[116] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__116_ : 1'b0;
  assign data_o_flat[115] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__115_ : 1'b0;
  assign data_o_flat[114] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__114_ : 1'b0;
  assign data_o_flat[113] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__113_ : 1'b0;
  assign data_o_flat[112] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__112_ : 1'b0;
  assign data_o_flat[111] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__111_ : 1'b0;
  assign data_o_flat[110] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__110_ : 1'b0;
  assign data_o_flat[109] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__109_ : 1'b0;
  assign data_o_flat[108] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__108_ : 1'b0;
  assign data_o_flat[107] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__107_ : 1'b0;
  assign data_o_flat[106] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__106_ : 1'b0;
  assign data_o_flat[105] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__105_ : 1'b0;
  assign data_o_flat[104] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__104_ : 1'b0;
  assign data_o_flat[103] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__103_ : 1'b0;
  assign data_o_flat[102] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__102_ : 1'b0;
  assign data_o_flat[101] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__101_ : 1'b0;
  assign data_o_flat[100] = (N47)? 1'b0 : 
                            (N49)? 1'b0 : 
                            (N51)? 1'b0 : 
                            (N53)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N50)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N54)? data_int_o_7__100_ : 1'b0;
  assign data_o_flat[99] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__99_ : 1'b0;
  assign data_o_flat[98] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__98_ : 1'b0;
  assign data_o_flat[97] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__97_ : 1'b0;
  assign data_o_flat[96] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__96_ : 1'b0;
  assign data_o_flat[95] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__95_ : 1'b0;
  assign data_o_flat[94] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__94_ : 1'b0;
  assign data_o_flat[93] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__93_ : 1'b0;
  assign data_o_flat[92] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__92_ : 1'b0;
  assign data_o_flat[91] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__91_ : 1'b0;
  assign data_o_flat[90] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__90_ : 1'b0;
  assign data_o_flat[89] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__89_ : 1'b0;
  assign data_o_flat[88] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__88_ : 1'b0;
  assign data_o_flat[87] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__87_ : 1'b0;
  assign data_o_flat[86] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__86_ : 1'b0;
  assign data_o_flat[85] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__85_ : 1'b0;
  assign data_o_flat[84] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__84_ : 1'b0;
  assign data_o_flat[83] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__83_ : 1'b0;
  assign data_o_flat[82] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__82_ : 1'b0;
  assign data_o_flat[81] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__81_ : 1'b0;
  assign data_o_flat[80] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__80_ : 1'b0;
  assign data_o_flat[79] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__79_ : 1'b0;
  assign data_o_flat[78] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__78_ : 1'b0;
  assign data_o_flat[77] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__77_ : 1'b0;
  assign data_o_flat[76] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__76_ : 1'b0;
  assign data_o_flat[75] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__75_ : 1'b0;
  assign data_o_flat[74] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__74_ : 1'b0;
  assign data_o_flat[73] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__73_ : 1'b0;
  assign data_o_flat[72] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__72_ : 1'b0;
  assign data_o_flat[71] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__71_ : 1'b0;
  assign data_o_flat[70] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__70_ : 1'b0;
  assign data_o_flat[69] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__69_ : 1'b0;
  assign data_o_flat[68] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__68_ : 1'b0;
  assign data_o_flat[67] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__67_ : 1'b0;
  assign data_o_flat[66] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__66_ : 1'b0;
  assign data_o_flat[65] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__65_ : 1'b0;
  assign data_o_flat[64] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__64_ : 1'b0;
  assign data_o_flat[63] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__63_ : 1'b0;
  assign data_o_flat[62] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__62_ : 1'b0;
  assign data_o_flat[61] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__61_ : 1'b0;
  assign data_o_flat[60] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__60_ : 1'b0;
  assign data_o_flat[59] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__59_ : 1'b0;
  assign data_o_flat[58] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__58_ : 1'b0;
  assign data_o_flat[57] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__57_ : 1'b0;
  assign data_o_flat[56] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__56_ : 1'b0;
  assign data_o_flat[55] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__55_ : 1'b0;
  assign data_o_flat[54] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__54_ : 1'b0;
  assign data_o_flat[53] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__53_ : 1'b0;
  assign data_o_flat[52] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__52_ : 1'b0;
  assign data_o_flat[51] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__51_ : 1'b0;
  assign data_o_flat[50] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__50_ : 1'b0;
  assign data_o_flat[49] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__49_ : 1'b0;
  assign data_o_flat[48] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__48_ : 1'b0;
  assign data_o_flat[47] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__47_ : 1'b0;
  assign data_o_flat[46] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__46_ : 1'b0;
  assign data_o_flat[45] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__45_ : 1'b0;
  assign data_o_flat[44] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__44_ : 1'b0;
  assign data_o_flat[43] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__43_ : 1'b0;
  assign data_o_flat[42] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__42_ : 1'b0;
  assign data_o_flat[41] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__41_ : 1'b0;
  assign data_o_flat[40] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__40_ : 1'b0;
  assign data_o_flat[39] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__39_ : 1'b0;
  assign data_o_flat[38] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__38_ : 1'b0;
  assign data_o_flat[37] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__37_ : 1'b0;
  assign data_o_flat[36] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__36_ : 1'b0;
  assign data_o_flat[35] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__35_ : 1'b0;
  assign data_o_flat[34] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__34_ : 1'b0;
  assign data_o_flat[33] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__33_ : 1'b0;
  assign data_o_flat[32] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__32_ : 1'b0;
  assign data_o_flat[31] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__31_ : 1'b0;
  assign data_o_flat[30] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__30_ : 1'b0;
  assign data_o_flat[29] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__29_ : 1'b0;
  assign data_o_flat[28] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__28_ : 1'b0;
  assign data_o_flat[27] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__27_ : 1'b0;
  assign data_o_flat[26] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__26_ : 1'b0;
  assign data_o_flat[25] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__25_ : 1'b0;
  assign data_o_flat[24] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__24_ : 1'b0;
  assign data_o_flat[23] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__23_ : 1'b0;
  assign data_o_flat[22] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__22_ : 1'b0;
  assign data_o_flat[21] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__21_ : 1'b0;
  assign data_o_flat[20] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__20_ : 1'b0;
  assign data_o_flat[19] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__19_ : 1'b0;
  assign data_o_flat[18] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__18_ : 1'b0;
  assign data_o_flat[17] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__17_ : 1'b0;
  assign data_o_flat[16] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__16_ : 1'b0;
  assign data_o_flat[15] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__15_ : 1'b0;
  assign data_o_flat[14] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__14_ : 1'b0;
  assign data_o_flat[13] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__13_ : 1'b0;
  assign data_o_flat[12] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__12_ : 1'b0;
  assign data_o_flat[11] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__11_ : 1'b0;
  assign data_o_flat[10] = (N47)? 1'b0 : 
                           (N49)? 1'b0 : 
                           (N51)? 1'b0 : 
                           (N53)? 1'b0 : 
                           (N48)? 1'b0 : 
                           (N50)? 1'b0 : 
                           (N52)? 1'b0 : 
                           (N54)? data_int_o_7__10_ : 1'b0;
  assign data_o_flat[9] = (N47)? 1'b0 : 
                          (N49)? 1'b0 : 
                          (N51)? 1'b0 : 
                          (N53)? 1'b0 : 
                          (N48)? 1'b0 : 
                          (N50)? 1'b0 : 
                          (N52)? 1'b0 : 
                          (N54)? data_int_o_7__9_ : 1'b0;
  assign data_o_flat[8] = (N47)? 1'b0 : 
                          (N49)? 1'b0 : 
                          (N51)? 1'b0 : 
                          (N53)? 1'b0 : 
                          (N48)? 1'b0 : 
                          (N50)? 1'b0 : 
                          (N52)? 1'b0 : 
                          (N54)? data_int_o_7__8_ : 1'b0;
  assign data_o_flat[7] = (N47)? 1'b0 : 
                          (N49)? 1'b0 : 
                          (N51)? 1'b0 : 
                          (N53)? 1'b0 : 
                          (N48)? 1'b0 : 
                          (N50)? 1'b0 : 
                          (N52)? 1'b0 : 
                          (N54)? data_int_o_7__7_ : 1'b0;
  assign data_o_flat[6] = (N47)? 1'b0 : 
                          (N49)? 1'b0 : 
                          (N51)? 1'b0 : 
                          (N53)? 1'b0 : 
                          (N48)? 1'b0 : 
                          (N50)? 1'b0 : 
                          (N52)? 1'b0 : 
                          (N54)? data_int_o_7__6_ : 1'b0;
  assign data_o_flat[5] = (N47)? 1'b0 : 
                          (N49)? 1'b0 : 
                          (N51)? 1'b0 : 
                          (N53)? 1'b0 : 
                          (N48)? 1'b0 : 
                          (N50)? 1'b0 : 
                          (N52)? 1'b0 : 
                          (N54)? data_int_o_7__5_ : 1'b0;
  assign data_o_flat[4] = (N47)? 1'b0 : 
                          (N49)? 1'b0 : 
                          (N51)? 1'b0 : 
                          (N53)? 1'b0 : 
                          (N48)? 1'b0 : 
                          (N50)? 1'b0 : 
                          (N52)? 1'b0 : 
                          (N54)? data_int_o_7__4_ : 1'b0;
  assign data_o_flat[3] = (N47)? 1'b0 : 
                          (N49)? 1'b0 : 
                          (N51)? 1'b0 : 
                          (N53)? 1'b0 : 
                          (N48)? 1'b0 : 
                          (N50)? 1'b0 : 
                          (N52)? 1'b0 : 
                          (N54)? data_int_o_7__3_ : 1'b0;
  assign data_o_flat[2] = (N47)? 1'b0 : 
                          (N49)? 1'b0 : 
                          (N51)? 1'b0 : 
                          (N53)? 1'b0 : 
                          (N48)? 1'b0 : 
                          (N50)? 1'b0 : 
                          (N52)? 1'b0 : 
                          (N54)? data_int_o_7__2_ : 1'b0;
  assign data_o_flat[1] = (N47)? 1'b0 : 
                          (N49)? 1'b0 : 
                          (N51)? 1'b0 : 
                          (N53)? 1'b0 : 
                          (N48)? 1'b0 : 
                          (N50)? 1'b0 : 
                          (N52)? 1'b0 : 
                          (N54)? data_int_o_7__1_ : 1'b0;
  assign data_o_flat[0] = (N47)? 1'b0 : 
                          (N49)? 1'b0 : 
                          (N51)? 1'b0 : 
                          (N53)? 1'b0 : 
                          (N48)? 1'b0 : 
                          (N50)? 1'b0 : 
                          (N52)? 1'b0 : 
                          (N54)? data_int_o_7__0_ : 1'b0;

  bsg_make_2D_array_width_p64_items_p8
  bm2Da
  (
    .i(data_o_flat),
    .o(data_o)
  );


  bsg_rr_f2f_input_width_p64_num_in_p16_middle_meet_p8
  ic_15__in_chan_bsg_rr_ff_in
  (
    .clk(clk),
    .reset(n_0_net_),
    .valid_i(valid_i),
    .data_i(data_i),
    .data_head_o({ data_head_15__511_, data_head_15__510_, data_head_15__509_, data_head_15__508_, data_head_15__507_, data_head_15__506_, data_head_15__505_, data_head_15__504_, data_head_15__503_, data_head_15__502_, data_head_15__501_, data_head_15__500_, data_head_15__499_, data_head_15__498_, data_head_15__497_, data_head_15__496_, data_head_15__495_, data_head_15__494_, data_head_15__493_, data_head_15__492_, data_head_15__491_, data_head_15__490_, data_head_15__489_, data_head_15__488_, data_head_15__487_, data_head_15__486_, data_head_15__485_, data_head_15__484_, data_head_15__483_, data_head_15__482_, data_head_15__481_, data_head_15__480_, data_head_15__479_, data_head_15__478_, data_head_15__477_, data_head_15__476_, data_head_15__475_, data_head_15__474_, data_head_15__473_, data_head_15__472_, data_head_15__471_, data_head_15__470_, data_head_15__469_, data_head_15__468_, data_head_15__467_, data_head_15__466_, data_head_15__465_, data_head_15__464_, data_head_15__463_, data_head_15__462_, data_head_15__461_, data_head_15__460_, data_head_15__459_, data_head_15__458_, data_head_15__457_, data_head_15__456_, data_head_15__455_, data_head_15__454_, data_head_15__453_, data_head_15__452_, data_head_15__451_, data_head_15__450_, data_head_15__449_, data_head_15__448_, data_head_15__447_, data_head_15__446_, data_head_15__445_, data_head_15__444_, data_head_15__443_, data_head_15__442_, data_head_15__441_, data_head_15__440_, data_head_15__439_, data_head_15__438_, data_head_15__437_, data_head_15__436_, data_head_15__435_, data_head_15__434_, data_head_15__433_, data_head_15__432_, data_head_15__431_, data_head_15__430_, data_head_15__429_, data_head_15__428_, data_head_15__427_, data_head_15__426_, data_head_15__425_, data_head_15__424_, data_head_15__423_, data_head_15__422_, data_head_15__421_, data_head_15__420_, data_head_15__419_, data_head_15__418_, data_head_15__417_, data_head_15__416_, data_head_15__415_, data_head_15__414_, data_head_15__413_, data_head_15__412_, data_head_15__411_, data_head_15__410_, data_head_15__409_, data_head_15__408_, data_head_15__407_, data_head_15__406_, data_head_15__405_, data_head_15__404_, data_head_15__403_, data_head_15__402_, data_head_15__401_, data_head_15__400_, data_head_15__399_, data_head_15__398_, data_head_15__397_, data_head_15__396_, data_head_15__395_, data_head_15__394_, data_head_15__393_, data_head_15__392_, data_head_15__391_, data_head_15__390_, data_head_15__389_, data_head_15__388_, data_head_15__387_, data_head_15__386_, data_head_15__385_, data_head_15__384_, data_head_15__383_, data_head_15__382_, data_head_15__381_, data_head_15__380_, data_head_15__379_, data_head_15__378_, data_head_15__377_, data_head_15__376_, data_head_15__375_, data_head_15__374_, data_head_15__373_, data_head_15__372_, data_head_15__371_, data_head_15__370_, data_head_15__369_, data_head_15__368_, data_head_15__367_, data_head_15__366_, data_head_15__365_, data_head_15__364_, data_head_15__363_, data_head_15__362_, data_head_15__361_, data_head_15__360_, data_head_15__359_, data_head_15__358_, data_head_15__357_, data_head_15__356_, data_head_15__355_, data_head_15__354_, data_head_15__353_, data_head_15__352_, data_head_15__351_, data_head_15__350_, data_head_15__349_, data_head_15__348_, data_head_15__347_, data_head_15__346_, data_head_15__345_, data_head_15__344_, data_head_15__343_, data_head_15__342_, data_head_15__341_, data_head_15__340_, data_head_15__339_, data_head_15__338_, data_head_15__337_, data_head_15__336_, data_head_15__335_, data_head_15__334_, data_head_15__333_, data_head_15__332_, data_head_15__331_, data_head_15__330_, data_head_15__329_, data_head_15__328_, data_head_15__327_, data_head_15__326_, data_head_15__325_, data_head_15__324_, data_head_15__323_, data_head_15__322_, data_head_15__321_, data_head_15__320_, data_head_15__319_, data_head_15__318_, data_head_15__317_, data_head_15__316_, data_head_15__315_, data_head_15__314_, data_head_15__313_, data_head_15__312_, data_head_15__311_, data_head_15__310_, data_head_15__309_, data_head_15__308_, data_head_15__307_, data_head_15__306_, data_head_15__305_, data_head_15__304_, data_head_15__303_, data_head_15__302_, data_head_15__301_, data_head_15__300_, data_head_15__299_, data_head_15__298_, data_head_15__297_, data_head_15__296_, data_head_15__295_, data_head_15__294_, data_head_15__293_, data_head_15__292_, data_head_15__291_, data_head_15__290_, data_head_15__289_, data_head_15__288_, data_head_15__287_, data_head_15__286_, data_head_15__285_, data_head_15__284_, data_head_15__283_, data_head_15__282_, data_head_15__281_, data_head_15__280_, data_head_15__279_, data_head_15__278_, data_head_15__277_, data_head_15__276_, data_head_15__275_, data_head_15__274_, data_head_15__273_, data_head_15__272_, data_head_15__271_, data_head_15__270_, data_head_15__269_, data_head_15__268_, data_head_15__267_, data_head_15__266_, data_head_15__265_, data_head_15__264_, data_head_15__263_, data_head_15__262_, data_head_15__261_, data_head_15__260_, data_head_15__259_, data_head_15__258_, data_head_15__257_, data_head_15__256_, data_head_15__255_, data_head_15__254_, data_head_15__253_, data_head_15__252_, data_head_15__251_, data_head_15__250_, data_head_15__249_, data_head_15__248_, data_head_15__247_, data_head_15__246_, data_head_15__245_, data_head_15__244_, data_head_15__243_, data_head_15__242_, data_head_15__241_, data_head_15__240_, data_head_15__239_, data_head_15__238_, data_head_15__237_, data_head_15__236_, data_head_15__235_, data_head_15__234_, data_head_15__233_, data_head_15__232_, data_head_15__231_, data_head_15__230_, data_head_15__229_, data_head_15__228_, data_head_15__227_, data_head_15__226_, data_head_15__225_, data_head_15__224_, data_head_15__223_, data_head_15__222_, data_head_15__221_, data_head_15__220_, data_head_15__219_, data_head_15__218_, data_head_15__217_, data_head_15__216_, data_head_15__215_, data_head_15__214_, data_head_15__213_, data_head_15__212_, data_head_15__211_, data_head_15__210_, data_head_15__209_, data_head_15__208_, data_head_15__207_, data_head_15__206_, data_head_15__205_, data_head_15__204_, data_head_15__203_, data_head_15__202_, data_head_15__201_, data_head_15__200_, data_head_15__199_, data_head_15__198_, data_head_15__197_, data_head_15__196_, data_head_15__195_, data_head_15__194_, data_head_15__193_, data_head_15__192_, data_head_15__191_, data_head_15__190_, data_head_15__189_, data_head_15__188_, data_head_15__187_, data_head_15__186_, data_head_15__185_, data_head_15__184_, data_head_15__183_, data_head_15__182_, data_head_15__181_, data_head_15__180_, data_head_15__179_, data_head_15__178_, data_head_15__177_, data_head_15__176_, data_head_15__175_, data_head_15__174_, data_head_15__173_, data_head_15__172_, data_head_15__171_, data_head_15__170_, data_head_15__169_, data_head_15__168_, data_head_15__167_, data_head_15__166_, data_head_15__165_, data_head_15__164_, data_head_15__163_, data_head_15__162_, data_head_15__161_, data_head_15__160_, data_head_15__159_, data_head_15__158_, data_head_15__157_, data_head_15__156_, data_head_15__155_, data_head_15__154_, data_head_15__153_, data_head_15__152_, data_head_15__151_, data_head_15__150_, data_head_15__149_, data_head_15__148_, data_head_15__147_, data_head_15__146_, data_head_15__145_, data_head_15__144_, data_head_15__143_, data_head_15__142_, data_head_15__141_, data_head_15__140_, data_head_15__139_, data_head_15__138_, data_head_15__137_, data_head_15__136_, data_head_15__135_, data_head_15__134_, data_head_15__133_, data_head_15__132_, data_head_15__131_, data_head_15__130_, data_head_15__129_, data_head_15__128_, data_head_15__127_, data_head_15__126_, data_head_15__125_, data_head_15__124_, data_head_15__123_, data_head_15__122_, data_head_15__121_, data_head_15__120_, data_head_15__119_, data_head_15__118_, data_head_15__117_, data_head_15__116_, data_head_15__115_, data_head_15__114_, data_head_15__113_, data_head_15__112_, data_head_15__111_, data_head_15__110_, data_head_15__109_, data_head_15__108_, data_head_15__107_, data_head_15__106_, data_head_15__105_, data_head_15__104_, data_head_15__103_, data_head_15__102_, data_head_15__101_, data_head_15__100_, data_head_15__99_, data_head_15__98_, data_head_15__97_, data_head_15__96_, data_head_15__95_, data_head_15__94_, data_head_15__93_, data_head_15__92_, data_head_15__91_, data_head_15__90_, data_head_15__89_, data_head_15__88_, data_head_15__87_, data_head_15__86_, data_head_15__85_, data_head_15__84_, data_head_15__83_, data_head_15__82_, data_head_15__81_, data_head_15__80_, data_head_15__79_, data_head_15__78_, data_head_15__77_, data_head_15__76_, data_head_15__75_, data_head_15__74_, data_head_15__73_, data_head_15__72_, data_head_15__71_, data_head_15__70_, data_head_15__69_, data_head_15__68_, data_head_15__67_, data_head_15__66_, data_head_15__65_, data_head_15__64_, data_head_15__63_, data_head_15__62_, data_head_15__61_, data_head_15__60_, data_head_15__59_, data_head_15__58_, data_head_15__57_, data_head_15__56_, data_head_15__55_, data_head_15__54_, data_head_15__53_, data_head_15__52_, data_head_15__51_, data_head_15__50_, data_head_15__49_, data_head_15__48_, data_head_15__47_, data_head_15__46_, data_head_15__45_, data_head_15__44_, data_head_15__43_, data_head_15__42_, data_head_15__41_, data_head_15__40_, data_head_15__39_, data_head_15__38_, data_head_15__37_, data_head_15__36_, data_head_15__35_, data_head_15__34_, data_head_15__33_, data_head_15__32_, data_head_15__31_, data_head_15__30_, data_head_15__29_, data_head_15__28_, data_head_15__27_, data_head_15__26_, data_head_15__25_, data_head_15__24_, data_head_15__23_, data_head_15__22_, data_head_15__21_, data_head_15__20_, data_head_15__19_, data_head_15__18_, data_head_15__17_, data_head_15__16_, data_head_15__15_, data_head_15__14_, data_head_15__13_, data_head_15__12_, data_head_15__11_, data_head_15__10_, data_head_15__9_, data_head_15__8_, data_head_15__7_, data_head_15__6_, data_head_15__5_, data_head_15__4_, data_head_15__3_, data_head_15__2_, data_head_15__1_, data_head_15__0_ }),
    .valid_head_o({ valid_head_15__7_, valid_head_15__6_, valid_head_15__5_, valid_head_15__4_, valid_head_15__3_, valid_head_15__2_, valid_head_15__1_, valid_head_15__0_ }),
    .go_channels_i(go_channels),
    .go_cnt_i(go_cnt),
    .yumi_o({ yumi_int_o_15__15_, yumi_int_o_15__14_, yumi_int_o_15__13_, yumi_int_o_15__12_, yumi_int_o_15__11_, yumi_int_o_15__10_, yumi_int_o_15__9_, yumi_int_o_15__8_, yumi_int_o_15__7_, yumi_int_o_15__6_, yumi_int_o_15__5_, yumi_int_o_15__4_, yumi_int_o_15__3_, yumi_int_o_15__2_, yumi_int_o_15__1_, yumi_int_o_15__0_ })
  );


  bsg_rr_f2f_middle_width_p64_middle_meet_p8
  brrf2fm
  (
    .valid_head_i({ n_2_net__7_, n_2_net__6_, n_2_net__5_, n_2_net__4_, n_2_net__3_, n_2_net__2_, n_2_net__1_, n_2_net__0_ }),
    .ready_head_i({ n_3_net__7_, n_3_net__6_, n_3_net__5_, n_3_net__4_, n_3_net__3_, n_3_net__2_, n_3_net__1_, n_3_net__0_ }),
    .go_channels_o(go_channels),
    .go_cnt_o(go_cnt)
  );

  assign n_3_net__7_ = (N39)? 1'b0 : 
                       (N41)? 1'b0 : 
                       (N43)? 1'b0 : 
                       (N55)? 1'b0 : 
                       (N40)? 1'b0 : 
                       (N42)? 1'b0 : 
                       (N44)? 1'b0 : 
                       (N56)? ready_head_7__7_ : 1'b0;
  assign n_3_net__6_ = (N39)? 1'b0 : 
                       (N41)? 1'b0 : 
                       (N43)? 1'b0 : 
                       (N55)? 1'b0 : 
                       (N40)? 1'b0 : 
                       (N42)? 1'b0 : 
                       (N44)? 1'b0 : 
                       (N56)? ready_head_7__6_ : 1'b0;
  assign n_3_net__5_ = (N39)? 1'b0 : 
                       (N41)? 1'b0 : 
                       (N43)? 1'b0 : 
                       (N55)? 1'b0 : 
                       (N40)? 1'b0 : 
                       (N42)? 1'b0 : 
                       (N44)? 1'b0 : 
                       (N56)? ready_head_7__5_ : 1'b0;
  assign n_3_net__4_ = (N39)? 1'b0 : 
                       (N41)? 1'b0 : 
                       (N43)? 1'b0 : 
                       (N55)? 1'b0 : 
                       (N40)? 1'b0 : 
                       (N42)? 1'b0 : 
                       (N44)? 1'b0 : 
                       (N56)? ready_head_7__4_ : 1'b0;
  assign n_3_net__3_ = (N39)? 1'b0 : 
                       (N41)? 1'b0 : 
                       (N43)? 1'b0 : 
                       (N55)? 1'b0 : 
                       (N40)? 1'b0 : 
                       (N42)? 1'b0 : 
                       (N44)? 1'b0 : 
                       (N56)? ready_head_7__3_ : 1'b0;
  assign n_3_net__2_ = (N39)? 1'b0 : 
                       (N41)? 1'b0 : 
                       (N43)? 1'b0 : 
                       (N55)? 1'b0 : 
                       (N40)? 1'b0 : 
                       (N42)? 1'b0 : 
                       (N44)? 1'b0 : 
                       (N56)? ready_head_7__2_ : 1'b0;
  assign n_3_net__1_ = (N39)? 1'b0 : 
                       (N41)? 1'b0 : 
                       (N43)? 1'b0 : 
                       (N55)? 1'b0 : 
                       (N40)? 1'b0 : 
                       (N42)? 1'b0 : 
                       (N44)? 1'b0 : 
                       (N56)? ready_head_7__1_ : 1'b0;
  assign n_3_net__0_ = (N39)? 1'b0 : 
                       (N41)? 1'b0 : 
                       (N43)? 1'b0 : 
                       (N55)? 1'b0 : 
                       (N40)? 1'b0 : 
                       (N42)? 1'b0 : 
                       (N44)? 1'b0 : 
                       (N56)? ready_head_7__0_ : 1'b0;
  assign n_2_net__7_ = (N16)? 1'b0 : 
                       (N18)? 1'b0 : 
                       (N20)? 1'b0 : 
                       (N57)? 1'b0 : 
                       (N24)? 1'b0 : 
                       (N26)? 1'b0 : 
                       (N28)? 1'b0 : 
                       (N30)? 1'b0 : 
                       (N17)? 1'b0 : 
                       (N19)? 1'b0 : 
                       (N21)? 1'b0 : 
                       (N58)? 1'b0 : 
                       (N25)? 1'b0 : 
                       (N27)? 1'b0 : 
                       (N29)? 1'b0 : 
                       (N59)? valid_head_15__7_ : 1'b0;
  assign n_2_net__6_ = (N16)? 1'b0 : 
                       (N18)? 1'b0 : 
                       (N20)? 1'b0 : 
                       (N57)? 1'b0 : 
                       (N24)? 1'b0 : 
                       (N26)? 1'b0 : 
                       (N28)? 1'b0 : 
                       (N30)? 1'b0 : 
                       (N17)? 1'b0 : 
                       (N19)? 1'b0 : 
                       (N21)? 1'b0 : 
                       (N58)? 1'b0 : 
                       (N25)? 1'b0 : 
                       (N27)? 1'b0 : 
                       (N29)? 1'b0 : 
                       (N59)? valid_head_15__6_ : 1'b0;
  assign n_2_net__5_ = (N16)? 1'b0 : 
                       (N18)? 1'b0 : 
                       (N20)? 1'b0 : 
                       (N57)? 1'b0 : 
                       (N24)? 1'b0 : 
                       (N26)? 1'b0 : 
                       (N28)? 1'b0 : 
                       (N30)? 1'b0 : 
                       (N17)? 1'b0 : 
                       (N19)? 1'b0 : 
                       (N21)? 1'b0 : 
                       (N58)? 1'b0 : 
                       (N25)? 1'b0 : 
                       (N27)? 1'b0 : 
                       (N29)? 1'b0 : 
                       (N59)? valid_head_15__5_ : 1'b0;
  assign n_2_net__4_ = (N16)? 1'b0 : 
                       (N18)? 1'b0 : 
                       (N20)? 1'b0 : 
                       (N57)? 1'b0 : 
                       (N24)? 1'b0 : 
                       (N26)? 1'b0 : 
                       (N28)? 1'b0 : 
                       (N30)? 1'b0 : 
                       (N17)? 1'b0 : 
                       (N19)? 1'b0 : 
                       (N21)? 1'b0 : 
                       (N58)? 1'b0 : 
                       (N25)? 1'b0 : 
                       (N27)? 1'b0 : 
                       (N29)? 1'b0 : 
                       (N59)? valid_head_15__4_ : 1'b0;
  assign n_2_net__3_ = (N16)? 1'b0 : 
                       (N18)? 1'b0 : 
                       (N20)? 1'b0 : 
                       (N57)? 1'b0 : 
                       (N24)? 1'b0 : 
                       (N26)? 1'b0 : 
                       (N28)? 1'b0 : 
                       (N30)? 1'b0 : 
                       (N17)? 1'b0 : 
                       (N19)? 1'b0 : 
                       (N21)? 1'b0 : 
                       (N58)? 1'b0 : 
                       (N25)? 1'b0 : 
                       (N27)? 1'b0 : 
                       (N29)? 1'b0 : 
                       (N59)? valid_head_15__3_ : 1'b0;
  assign n_2_net__2_ = (N16)? 1'b0 : 
                       (N18)? 1'b0 : 
                       (N20)? 1'b0 : 
                       (N57)? 1'b0 : 
                       (N24)? 1'b0 : 
                       (N26)? 1'b0 : 
                       (N28)? 1'b0 : 
                       (N30)? 1'b0 : 
                       (N17)? 1'b0 : 
                       (N19)? 1'b0 : 
                       (N21)? 1'b0 : 
                       (N58)? 1'b0 : 
                       (N25)? 1'b0 : 
                       (N27)? 1'b0 : 
                       (N29)? 1'b0 : 
                       (N59)? valid_head_15__2_ : 1'b0;
  assign n_2_net__1_ = (N16)? 1'b0 : 
                       (N18)? 1'b0 : 
                       (N20)? 1'b0 : 
                       (N57)? 1'b0 : 
                       (N24)? 1'b0 : 
                       (N26)? 1'b0 : 
                       (N28)? 1'b0 : 
                       (N30)? 1'b0 : 
                       (N17)? 1'b0 : 
                       (N19)? 1'b0 : 
                       (N21)? 1'b0 : 
                       (N58)? 1'b0 : 
                       (N25)? 1'b0 : 
                       (N27)? 1'b0 : 
                       (N29)? 1'b0 : 
                       (N59)? valid_head_15__1_ : 1'b0;
  assign n_2_net__0_ = (N16)? 1'b0 : 
                       (N18)? 1'b0 : 
                       (N20)? 1'b0 : 
                       (N57)? 1'b0 : 
                       (N24)? 1'b0 : 
                       (N26)? 1'b0 : 
                       (N28)? 1'b0 : 
                       (N30)? 1'b0 : 
                       (N17)? 1'b0 : 
                       (N19)? 1'b0 : 
                       (N21)? 1'b0 : 
                       (N58)? 1'b0 : 
                       (N25)? 1'b0 : 
                       (N27)? 1'b0 : 
                       (N29)? 1'b0 : 
                       (N59)? valid_head_15__0_ : 1'b0;

  bsg_make_2D_array_width_p64_items_p8
  oc_7__out_chan_bm2Da
  (
    .i({ n_4_net__511_, n_4_net__510_, n_4_net__509_, n_4_net__508_, n_4_net__507_, n_4_net__506_, n_4_net__505_, n_4_net__504_, n_4_net__503_, n_4_net__502_, n_4_net__501_, n_4_net__500_, n_4_net__499_, n_4_net__498_, n_4_net__497_, n_4_net__496_, n_4_net__495_, n_4_net__494_, n_4_net__493_, n_4_net__492_, n_4_net__491_, n_4_net__490_, n_4_net__489_, n_4_net__488_, n_4_net__487_, n_4_net__486_, n_4_net__485_, n_4_net__484_, n_4_net__483_, n_4_net__482_, n_4_net__481_, n_4_net__480_, n_4_net__479_, n_4_net__478_, n_4_net__477_, n_4_net__476_, n_4_net__475_, n_4_net__474_, n_4_net__473_, n_4_net__472_, n_4_net__471_, n_4_net__470_, n_4_net__469_, n_4_net__468_, n_4_net__467_, n_4_net__466_, n_4_net__465_, n_4_net__464_, n_4_net__463_, n_4_net__462_, n_4_net__461_, n_4_net__460_, n_4_net__459_, n_4_net__458_, n_4_net__457_, n_4_net__456_, n_4_net__455_, n_4_net__454_, n_4_net__453_, n_4_net__452_, n_4_net__451_, n_4_net__450_, n_4_net__449_, n_4_net__448_, n_4_net__447_, n_4_net__446_, n_4_net__445_, n_4_net__444_, n_4_net__443_, n_4_net__442_, n_4_net__441_, n_4_net__440_, n_4_net__439_, n_4_net__438_, n_4_net__437_, n_4_net__436_, n_4_net__435_, n_4_net__434_, n_4_net__433_, n_4_net__432_, n_4_net__431_, n_4_net__430_, n_4_net__429_, n_4_net__428_, n_4_net__427_, n_4_net__426_, n_4_net__425_, n_4_net__424_, n_4_net__423_, n_4_net__422_, n_4_net__421_, n_4_net__420_, n_4_net__419_, n_4_net__418_, n_4_net__417_, n_4_net__416_, n_4_net__415_, n_4_net__414_, n_4_net__413_, n_4_net__412_, n_4_net__411_, n_4_net__410_, n_4_net__409_, n_4_net__408_, n_4_net__407_, n_4_net__406_, n_4_net__405_, n_4_net__404_, n_4_net__403_, n_4_net__402_, n_4_net__401_, n_4_net__400_, n_4_net__399_, n_4_net__398_, n_4_net__397_, n_4_net__396_, n_4_net__395_, n_4_net__394_, n_4_net__393_, n_4_net__392_, n_4_net__391_, n_4_net__390_, n_4_net__389_, n_4_net__388_, n_4_net__387_, n_4_net__386_, n_4_net__385_, n_4_net__384_, n_4_net__383_, n_4_net__382_, n_4_net__381_, n_4_net__380_, n_4_net__379_, n_4_net__378_, n_4_net__377_, n_4_net__376_, n_4_net__375_, n_4_net__374_, n_4_net__373_, n_4_net__372_, n_4_net__371_, n_4_net__370_, n_4_net__369_, n_4_net__368_, n_4_net__367_, n_4_net__366_, n_4_net__365_, n_4_net__364_, n_4_net__363_, n_4_net__362_, n_4_net__361_, n_4_net__360_, n_4_net__359_, n_4_net__358_, n_4_net__357_, n_4_net__356_, n_4_net__355_, n_4_net__354_, n_4_net__353_, n_4_net__352_, n_4_net__351_, n_4_net__350_, n_4_net__349_, n_4_net__348_, n_4_net__347_, n_4_net__346_, n_4_net__345_, n_4_net__344_, n_4_net__343_, n_4_net__342_, n_4_net__341_, n_4_net__340_, n_4_net__339_, n_4_net__338_, n_4_net__337_, n_4_net__336_, n_4_net__335_, n_4_net__334_, n_4_net__333_, n_4_net__332_, n_4_net__331_, n_4_net__330_, n_4_net__329_, n_4_net__328_, n_4_net__327_, n_4_net__326_, n_4_net__325_, n_4_net__324_, n_4_net__323_, n_4_net__322_, n_4_net__321_, n_4_net__320_, n_4_net__319_, n_4_net__318_, n_4_net__317_, n_4_net__316_, n_4_net__315_, n_4_net__314_, n_4_net__313_, n_4_net__312_, n_4_net__311_, n_4_net__310_, n_4_net__309_, n_4_net__308_, n_4_net__307_, n_4_net__306_, n_4_net__305_, n_4_net__304_, n_4_net__303_, n_4_net__302_, n_4_net__301_, n_4_net__300_, n_4_net__299_, n_4_net__298_, n_4_net__297_, n_4_net__296_, n_4_net__295_, n_4_net__294_, n_4_net__293_, n_4_net__292_, n_4_net__291_, n_4_net__290_, n_4_net__289_, n_4_net__288_, n_4_net__287_, n_4_net__286_, n_4_net__285_, n_4_net__284_, n_4_net__283_, n_4_net__282_, n_4_net__281_, n_4_net__280_, n_4_net__279_, n_4_net__278_, n_4_net__277_, n_4_net__276_, n_4_net__275_, n_4_net__274_, n_4_net__273_, n_4_net__272_, n_4_net__271_, n_4_net__270_, n_4_net__269_, n_4_net__268_, n_4_net__267_, n_4_net__266_, n_4_net__265_, n_4_net__264_, n_4_net__263_, n_4_net__262_, n_4_net__261_, n_4_net__260_, n_4_net__259_, n_4_net__258_, n_4_net__257_, n_4_net__256_, n_4_net__255_, n_4_net__254_, n_4_net__253_, n_4_net__252_, n_4_net__251_, n_4_net__250_, n_4_net__249_, n_4_net__248_, n_4_net__247_, n_4_net__246_, n_4_net__245_, n_4_net__244_, n_4_net__243_, n_4_net__242_, n_4_net__241_, n_4_net__240_, n_4_net__239_, n_4_net__238_, n_4_net__237_, n_4_net__236_, n_4_net__235_, n_4_net__234_, n_4_net__233_, n_4_net__232_, n_4_net__231_, n_4_net__230_, n_4_net__229_, n_4_net__228_, n_4_net__227_, n_4_net__226_, n_4_net__225_, n_4_net__224_, n_4_net__223_, n_4_net__222_, n_4_net__221_, n_4_net__220_, n_4_net__219_, n_4_net__218_, n_4_net__217_, n_4_net__216_, n_4_net__215_, n_4_net__214_, n_4_net__213_, n_4_net__212_, n_4_net__211_, n_4_net__210_, n_4_net__209_, n_4_net__208_, n_4_net__207_, n_4_net__206_, n_4_net__205_, n_4_net__204_, n_4_net__203_, n_4_net__202_, n_4_net__201_, n_4_net__200_, n_4_net__199_, n_4_net__198_, n_4_net__197_, n_4_net__196_, n_4_net__195_, n_4_net__194_, n_4_net__193_, n_4_net__192_, n_4_net__191_, n_4_net__190_, n_4_net__189_, n_4_net__188_, n_4_net__187_, n_4_net__186_, n_4_net__185_, n_4_net__184_, n_4_net__183_, n_4_net__182_, n_4_net__181_, n_4_net__180_, n_4_net__179_, n_4_net__178_, n_4_net__177_, n_4_net__176_, n_4_net__175_, n_4_net__174_, n_4_net__173_, n_4_net__172_, n_4_net__171_, n_4_net__170_, n_4_net__169_, n_4_net__168_, n_4_net__167_, n_4_net__166_, n_4_net__165_, n_4_net__164_, n_4_net__163_, n_4_net__162_, n_4_net__161_, n_4_net__160_, n_4_net__159_, n_4_net__158_, n_4_net__157_, n_4_net__156_, n_4_net__155_, n_4_net__154_, n_4_net__153_, n_4_net__152_, n_4_net__151_, n_4_net__150_, n_4_net__149_, n_4_net__148_, n_4_net__147_, n_4_net__146_, n_4_net__145_, n_4_net__144_, n_4_net__143_, n_4_net__142_, n_4_net__141_, n_4_net__140_, n_4_net__139_, n_4_net__138_, n_4_net__137_, n_4_net__136_, n_4_net__135_, n_4_net__134_, n_4_net__133_, n_4_net__132_, n_4_net__131_, n_4_net__130_, n_4_net__129_, n_4_net__128_, n_4_net__127_, n_4_net__126_, n_4_net__125_, n_4_net__124_, n_4_net__123_, n_4_net__122_, n_4_net__121_, n_4_net__120_, n_4_net__119_, n_4_net__118_, n_4_net__117_, n_4_net__116_, n_4_net__115_, n_4_net__114_, n_4_net__113_, n_4_net__112_, n_4_net__111_, n_4_net__110_, n_4_net__109_, n_4_net__108_, n_4_net__107_, n_4_net__106_, n_4_net__105_, n_4_net__104_, n_4_net__103_, n_4_net__102_, n_4_net__101_, n_4_net__100_, n_4_net__99_, n_4_net__98_, n_4_net__97_, n_4_net__96_, n_4_net__95_, n_4_net__94_, n_4_net__93_, n_4_net__92_, n_4_net__91_, n_4_net__90_, n_4_net__89_, n_4_net__88_, n_4_net__87_, n_4_net__86_, n_4_net__85_, n_4_net__84_, n_4_net__83_, n_4_net__82_, n_4_net__81_, n_4_net__80_, n_4_net__79_, n_4_net__78_, n_4_net__77_, n_4_net__76_, n_4_net__75_, n_4_net__74_, n_4_net__73_, n_4_net__72_, n_4_net__71_, n_4_net__70_, n_4_net__69_, n_4_net__68_, n_4_net__67_, n_4_net__66_, n_4_net__65_, n_4_net__64_, n_4_net__63_, n_4_net__62_, n_4_net__61_, n_4_net__60_, n_4_net__59_, n_4_net__58_, n_4_net__57_, n_4_net__56_, n_4_net__55_, n_4_net__54_, n_4_net__53_, n_4_net__52_, n_4_net__51_, n_4_net__50_, n_4_net__49_, n_4_net__48_, n_4_net__47_, n_4_net__46_, n_4_net__45_, n_4_net__44_, n_4_net__43_, n_4_net__42_, n_4_net__41_, n_4_net__40_, n_4_net__39_, n_4_net__38_, n_4_net__37_, n_4_net__36_, n_4_net__35_, n_4_net__34_, n_4_net__33_, n_4_net__32_, n_4_net__31_, n_4_net__30_, n_4_net__29_, n_4_net__28_, n_4_net__27_, n_4_net__26_, n_4_net__25_, n_4_net__24_, n_4_net__23_, n_4_net__22_, n_4_net__21_, n_4_net__20_, n_4_net__19_, n_4_net__18_, n_4_net__17_, n_4_net__16_, n_4_net__15_, n_4_net__14_, n_4_net__13_, n_4_net__12_, n_4_net__11_, n_4_net__10_, n_4_net__9_, n_4_net__8_, n_4_net__7_, n_4_net__6_, n_4_net__5_, n_4_net__4_, n_4_net__3_, n_4_net__2_, n_4_net__1_, n_4_net__0_ }),
    .o(oc_7__out_chan_data_head_array)
  );

  assign n_4_net__511_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__511_ : 1'b0;
  assign n_4_net__510_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__510_ : 1'b0;
  assign n_4_net__509_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__509_ : 1'b0;
  assign n_4_net__508_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__508_ : 1'b0;
  assign n_4_net__507_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__507_ : 1'b0;
  assign n_4_net__506_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__506_ : 1'b0;
  assign n_4_net__505_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__505_ : 1'b0;
  assign n_4_net__504_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__504_ : 1'b0;
  assign n_4_net__503_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__503_ : 1'b0;
  assign n_4_net__502_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__502_ : 1'b0;
  assign n_4_net__501_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__501_ : 1'b0;
  assign n_4_net__500_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__500_ : 1'b0;
  assign n_4_net__499_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__499_ : 1'b0;
  assign n_4_net__498_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__498_ : 1'b0;
  assign n_4_net__497_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__497_ : 1'b0;
  assign n_4_net__496_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__496_ : 1'b0;
  assign n_4_net__495_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__495_ : 1'b0;
  assign n_4_net__494_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__494_ : 1'b0;
  assign n_4_net__493_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__493_ : 1'b0;
  assign n_4_net__492_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__492_ : 1'b0;
  assign n_4_net__491_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__491_ : 1'b0;
  assign n_4_net__490_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__490_ : 1'b0;
  assign n_4_net__489_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__489_ : 1'b0;
  assign n_4_net__488_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__488_ : 1'b0;
  assign n_4_net__487_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__487_ : 1'b0;
  assign n_4_net__486_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__486_ : 1'b0;
  assign n_4_net__485_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__485_ : 1'b0;
  assign n_4_net__484_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__484_ : 1'b0;
  assign n_4_net__483_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__483_ : 1'b0;
  assign n_4_net__482_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__482_ : 1'b0;
  assign n_4_net__481_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__481_ : 1'b0;
  assign n_4_net__480_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__480_ : 1'b0;
  assign n_4_net__479_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__479_ : 1'b0;
  assign n_4_net__478_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__478_ : 1'b0;
  assign n_4_net__477_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__477_ : 1'b0;
  assign n_4_net__476_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__476_ : 1'b0;
  assign n_4_net__475_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__475_ : 1'b0;
  assign n_4_net__474_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__474_ : 1'b0;
  assign n_4_net__473_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__473_ : 1'b0;
  assign n_4_net__472_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__472_ : 1'b0;
  assign n_4_net__471_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__471_ : 1'b0;
  assign n_4_net__470_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__470_ : 1'b0;
  assign n_4_net__469_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__469_ : 1'b0;
  assign n_4_net__468_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__468_ : 1'b0;
  assign n_4_net__467_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__467_ : 1'b0;
  assign n_4_net__466_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__466_ : 1'b0;
  assign n_4_net__465_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__465_ : 1'b0;
  assign n_4_net__464_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__464_ : 1'b0;
  assign n_4_net__463_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__463_ : 1'b0;
  assign n_4_net__462_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__462_ : 1'b0;
  assign n_4_net__461_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__461_ : 1'b0;
  assign n_4_net__460_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__460_ : 1'b0;
  assign n_4_net__459_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__459_ : 1'b0;
  assign n_4_net__458_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__458_ : 1'b0;
  assign n_4_net__457_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__457_ : 1'b0;
  assign n_4_net__456_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__456_ : 1'b0;
  assign n_4_net__455_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__455_ : 1'b0;
  assign n_4_net__454_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__454_ : 1'b0;
  assign n_4_net__453_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__453_ : 1'b0;
  assign n_4_net__452_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__452_ : 1'b0;
  assign n_4_net__451_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__451_ : 1'b0;
  assign n_4_net__450_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__450_ : 1'b0;
  assign n_4_net__449_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__449_ : 1'b0;
  assign n_4_net__448_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__448_ : 1'b0;
  assign n_4_net__447_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__447_ : 1'b0;
  assign n_4_net__446_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__446_ : 1'b0;
  assign n_4_net__445_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__445_ : 1'b0;
  assign n_4_net__444_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__444_ : 1'b0;
  assign n_4_net__443_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__443_ : 1'b0;
  assign n_4_net__442_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__442_ : 1'b0;
  assign n_4_net__441_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__441_ : 1'b0;
  assign n_4_net__440_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__440_ : 1'b0;
  assign n_4_net__439_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__439_ : 1'b0;
  assign n_4_net__438_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__438_ : 1'b0;
  assign n_4_net__437_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__437_ : 1'b0;
  assign n_4_net__436_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__436_ : 1'b0;
  assign n_4_net__435_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__435_ : 1'b0;
  assign n_4_net__434_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__434_ : 1'b0;
  assign n_4_net__433_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__433_ : 1'b0;
  assign n_4_net__432_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__432_ : 1'b0;
  assign n_4_net__431_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__431_ : 1'b0;
  assign n_4_net__430_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__430_ : 1'b0;
  assign n_4_net__429_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__429_ : 1'b0;
  assign n_4_net__428_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__428_ : 1'b0;
  assign n_4_net__427_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__427_ : 1'b0;
  assign n_4_net__426_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__426_ : 1'b0;
  assign n_4_net__425_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__425_ : 1'b0;
  assign n_4_net__424_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__424_ : 1'b0;
  assign n_4_net__423_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__423_ : 1'b0;
  assign n_4_net__422_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__422_ : 1'b0;
  assign n_4_net__421_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__421_ : 1'b0;
  assign n_4_net__420_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__420_ : 1'b0;
  assign n_4_net__419_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__419_ : 1'b0;
  assign n_4_net__418_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__418_ : 1'b0;
  assign n_4_net__417_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__417_ : 1'b0;
  assign n_4_net__416_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__416_ : 1'b0;
  assign n_4_net__415_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__415_ : 1'b0;
  assign n_4_net__414_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__414_ : 1'b0;
  assign n_4_net__413_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__413_ : 1'b0;
  assign n_4_net__412_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__412_ : 1'b0;
  assign n_4_net__411_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__411_ : 1'b0;
  assign n_4_net__410_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__410_ : 1'b0;
  assign n_4_net__409_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__409_ : 1'b0;
  assign n_4_net__408_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__408_ : 1'b0;
  assign n_4_net__407_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__407_ : 1'b0;
  assign n_4_net__406_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__406_ : 1'b0;
  assign n_4_net__405_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__405_ : 1'b0;
  assign n_4_net__404_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__404_ : 1'b0;
  assign n_4_net__403_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__403_ : 1'b0;
  assign n_4_net__402_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__402_ : 1'b0;
  assign n_4_net__401_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__401_ : 1'b0;
  assign n_4_net__400_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__400_ : 1'b0;
  assign n_4_net__399_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__399_ : 1'b0;
  assign n_4_net__398_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__398_ : 1'b0;
  assign n_4_net__397_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__397_ : 1'b0;
  assign n_4_net__396_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__396_ : 1'b0;
  assign n_4_net__395_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__395_ : 1'b0;
  assign n_4_net__394_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__394_ : 1'b0;
  assign n_4_net__393_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__393_ : 1'b0;
  assign n_4_net__392_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__392_ : 1'b0;
  assign n_4_net__391_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__391_ : 1'b0;
  assign n_4_net__390_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__390_ : 1'b0;
  assign n_4_net__389_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__389_ : 1'b0;
  assign n_4_net__388_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__388_ : 1'b0;
  assign n_4_net__387_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__387_ : 1'b0;
  assign n_4_net__386_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__386_ : 1'b0;
  assign n_4_net__385_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__385_ : 1'b0;
  assign n_4_net__384_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__384_ : 1'b0;
  assign n_4_net__383_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__383_ : 1'b0;
  assign n_4_net__382_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__382_ : 1'b0;
  assign n_4_net__381_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__381_ : 1'b0;
  assign n_4_net__380_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__380_ : 1'b0;
  assign n_4_net__379_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__379_ : 1'b0;
  assign n_4_net__378_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__378_ : 1'b0;
  assign n_4_net__377_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__377_ : 1'b0;
  assign n_4_net__376_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__376_ : 1'b0;
  assign n_4_net__375_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__375_ : 1'b0;
  assign n_4_net__374_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__374_ : 1'b0;
  assign n_4_net__373_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__373_ : 1'b0;
  assign n_4_net__372_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__372_ : 1'b0;
  assign n_4_net__371_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__371_ : 1'b0;
  assign n_4_net__370_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__370_ : 1'b0;
  assign n_4_net__369_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__369_ : 1'b0;
  assign n_4_net__368_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__368_ : 1'b0;
  assign n_4_net__367_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__367_ : 1'b0;
  assign n_4_net__366_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__366_ : 1'b0;
  assign n_4_net__365_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__365_ : 1'b0;
  assign n_4_net__364_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__364_ : 1'b0;
  assign n_4_net__363_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__363_ : 1'b0;
  assign n_4_net__362_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__362_ : 1'b0;
  assign n_4_net__361_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__361_ : 1'b0;
  assign n_4_net__360_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__360_ : 1'b0;
  assign n_4_net__359_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__359_ : 1'b0;
  assign n_4_net__358_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__358_ : 1'b0;
  assign n_4_net__357_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__357_ : 1'b0;
  assign n_4_net__356_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__356_ : 1'b0;
  assign n_4_net__355_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__355_ : 1'b0;
  assign n_4_net__354_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__354_ : 1'b0;
  assign n_4_net__353_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__353_ : 1'b0;
  assign n_4_net__352_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__352_ : 1'b0;
  assign n_4_net__351_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__351_ : 1'b0;
  assign n_4_net__350_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__350_ : 1'b0;
  assign n_4_net__349_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__349_ : 1'b0;
  assign n_4_net__348_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__348_ : 1'b0;
  assign n_4_net__347_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__347_ : 1'b0;
  assign n_4_net__346_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__346_ : 1'b0;
  assign n_4_net__345_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__345_ : 1'b0;
  assign n_4_net__344_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__344_ : 1'b0;
  assign n_4_net__343_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__343_ : 1'b0;
  assign n_4_net__342_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__342_ : 1'b0;
  assign n_4_net__341_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__341_ : 1'b0;
  assign n_4_net__340_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__340_ : 1'b0;
  assign n_4_net__339_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__339_ : 1'b0;
  assign n_4_net__338_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__338_ : 1'b0;
  assign n_4_net__337_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__337_ : 1'b0;
  assign n_4_net__336_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__336_ : 1'b0;
  assign n_4_net__335_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__335_ : 1'b0;
  assign n_4_net__334_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__334_ : 1'b0;
  assign n_4_net__333_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__333_ : 1'b0;
  assign n_4_net__332_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__332_ : 1'b0;
  assign n_4_net__331_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__331_ : 1'b0;
  assign n_4_net__330_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__330_ : 1'b0;
  assign n_4_net__329_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__329_ : 1'b0;
  assign n_4_net__328_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__328_ : 1'b0;
  assign n_4_net__327_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__327_ : 1'b0;
  assign n_4_net__326_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__326_ : 1'b0;
  assign n_4_net__325_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__325_ : 1'b0;
  assign n_4_net__324_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__324_ : 1'b0;
  assign n_4_net__323_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__323_ : 1'b0;
  assign n_4_net__322_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__322_ : 1'b0;
  assign n_4_net__321_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__321_ : 1'b0;
  assign n_4_net__320_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__320_ : 1'b0;
  assign n_4_net__319_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__319_ : 1'b0;
  assign n_4_net__318_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__318_ : 1'b0;
  assign n_4_net__317_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__317_ : 1'b0;
  assign n_4_net__316_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__316_ : 1'b0;
  assign n_4_net__315_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__315_ : 1'b0;
  assign n_4_net__314_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__314_ : 1'b0;
  assign n_4_net__313_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__313_ : 1'b0;
  assign n_4_net__312_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__312_ : 1'b0;
  assign n_4_net__311_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__311_ : 1'b0;
  assign n_4_net__310_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__310_ : 1'b0;
  assign n_4_net__309_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__309_ : 1'b0;
  assign n_4_net__308_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__308_ : 1'b0;
  assign n_4_net__307_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__307_ : 1'b0;
  assign n_4_net__306_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__306_ : 1'b0;
  assign n_4_net__305_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__305_ : 1'b0;
  assign n_4_net__304_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__304_ : 1'b0;
  assign n_4_net__303_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__303_ : 1'b0;
  assign n_4_net__302_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__302_ : 1'b0;
  assign n_4_net__301_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__301_ : 1'b0;
  assign n_4_net__300_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__300_ : 1'b0;
  assign n_4_net__299_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__299_ : 1'b0;
  assign n_4_net__298_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__298_ : 1'b0;
  assign n_4_net__297_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__297_ : 1'b0;
  assign n_4_net__296_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__296_ : 1'b0;
  assign n_4_net__295_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__295_ : 1'b0;
  assign n_4_net__294_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__294_ : 1'b0;
  assign n_4_net__293_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__293_ : 1'b0;
  assign n_4_net__292_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__292_ : 1'b0;
  assign n_4_net__291_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__291_ : 1'b0;
  assign n_4_net__290_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__290_ : 1'b0;
  assign n_4_net__289_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__289_ : 1'b0;
  assign n_4_net__288_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__288_ : 1'b0;
  assign n_4_net__287_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__287_ : 1'b0;
  assign n_4_net__286_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__286_ : 1'b0;
  assign n_4_net__285_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__285_ : 1'b0;
  assign n_4_net__284_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__284_ : 1'b0;
  assign n_4_net__283_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__283_ : 1'b0;
  assign n_4_net__282_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__282_ : 1'b0;
  assign n_4_net__281_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__281_ : 1'b0;
  assign n_4_net__280_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__280_ : 1'b0;
  assign n_4_net__279_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__279_ : 1'b0;
  assign n_4_net__278_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__278_ : 1'b0;
  assign n_4_net__277_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__277_ : 1'b0;
  assign n_4_net__276_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__276_ : 1'b0;
  assign n_4_net__275_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__275_ : 1'b0;
  assign n_4_net__274_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__274_ : 1'b0;
  assign n_4_net__273_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__273_ : 1'b0;
  assign n_4_net__272_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__272_ : 1'b0;
  assign n_4_net__271_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__271_ : 1'b0;
  assign n_4_net__270_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__270_ : 1'b0;
  assign n_4_net__269_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__269_ : 1'b0;
  assign n_4_net__268_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__268_ : 1'b0;
  assign n_4_net__267_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__267_ : 1'b0;
  assign n_4_net__266_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__266_ : 1'b0;
  assign n_4_net__265_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__265_ : 1'b0;
  assign n_4_net__264_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__264_ : 1'b0;
  assign n_4_net__263_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__263_ : 1'b0;
  assign n_4_net__262_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__262_ : 1'b0;
  assign n_4_net__261_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__261_ : 1'b0;
  assign n_4_net__260_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__260_ : 1'b0;
  assign n_4_net__259_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__259_ : 1'b0;
  assign n_4_net__258_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__258_ : 1'b0;
  assign n_4_net__257_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__257_ : 1'b0;
  assign n_4_net__256_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__256_ : 1'b0;
  assign n_4_net__255_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__255_ : 1'b0;
  assign n_4_net__254_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__254_ : 1'b0;
  assign n_4_net__253_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__253_ : 1'b0;
  assign n_4_net__252_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__252_ : 1'b0;
  assign n_4_net__251_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__251_ : 1'b0;
  assign n_4_net__250_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__250_ : 1'b0;
  assign n_4_net__249_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__249_ : 1'b0;
  assign n_4_net__248_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__248_ : 1'b0;
  assign n_4_net__247_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__247_ : 1'b0;
  assign n_4_net__246_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__246_ : 1'b0;
  assign n_4_net__245_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__245_ : 1'b0;
  assign n_4_net__244_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__244_ : 1'b0;
  assign n_4_net__243_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__243_ : 1'b0;
  assign n_4_net__242_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__242_ : 1'b0;
  assign n_4_net__241_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__241_ : 1'b0;
  assign n_4_net__240_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__240_ : 1'b0;
  assign n_4_net__239_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__239_ : 1'b0;
  assign n_4_net__238_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__238_ : 1'b0;
  assign n_4_net__237_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__237_ : 1'b0;
  assign n_4_net__236_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__236_ : 1'b0;
  assign n_4_net__235_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__235_ : 1'b0;
  assign n_4_net__234_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__234_ : 1'b0;
  assign n_4_net__233_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__233_ : 1'b0;
  assign n_4_net__232_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__232_ : 1'b0;
  assign n_4_net__231_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__231_ : 1'b0;
  assign n_4_net__230_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__230_ : 1'b0;
  assign n_4_net__229_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__229_ : 1'b0;
  assign n_4_net__228_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__228_ : 1'b0;
  assign n_4_net__227_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__227_ : 1'b0;
  assign n_4_net__226_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__226_ : 1'b0;
  assign n_4_net__225_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__225_ : 1'b0;
  assign n_4_net__224_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__224_ : 1'b0;
  assign n_4_net__223_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__223_ : 1'b0;
  assign n_4_net__222_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__222_ : 1'b0;
  assign n_4_net__221_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__221_ : 1'b0;
  assign n_4_net__220_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__220_ : 1'b0;
  assign n_4_net__219_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__219_ : 1'b0;
  assign n_4_net__218_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__218_ : 1'b0;
  assign n_4_net__217_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__217_ : 1'b0;
  assign n_4_net__216_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__216_ : 1'b0;
  assign n_4_net__215_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__215_ : 1'b0;
  assign n_4_net__214_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__214_ : 1'b0;
  assign n_4_net__213_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__213_ : 1'b0;
  assign n_4_net__212_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__212_ : 1'b0;
  assign n_4_net__211_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__211_ : 1'b0;
  assign n_4_net__210_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__210_ : 1'b0;
  assign n_4_net__209_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__209_ : 1'b0;
  assign n_4_net__208_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__208_ : 1'b0;
  assign n_4_net__207_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__207_ : 1'b0;
  assign n_4_net__206_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__206_ : 1'b0;
  assign n_4_net__205_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__205_ : 1'b0;
  assign n_4_net__204_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__204_ : 1'b0;
  assign n_4_net__203_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__203_ : 1'b0;
  assign n_4_net__202_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__202_ : 1'b0;
  assign n_4_net__201_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__201_ : 1'b0;
  assign n_4_net__200_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__200_ : 1'b0;
  assign n_4_net__199_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__199_ : 1'b0;
  assign n_4_net__198_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__198_ : 1'b0;
  assign n_4_net__197_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__197_ : 1'b0;
  assign n_4_net__196_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__196_ : 1'b0;
  assign n_4_net__195_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__195_ : 1'b0;
  assign n_4_net__194_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__194_ : 1'b0;
  assign n_4_net__193_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__193_ : 1'b0;
  assign n_4_net__192_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__192_ : 1'b0;
  assign n_4_net__191_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__191_ : 1'b0;
  assign n_4_net__190_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__190_ : 1'b0;
  assign n_4_net__189_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__189_ : 1'b0;
  assign n_4_net__188_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__188_ : 1'b0;
  assign n_4_net__187_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__187_ : 1'b0;
  assign n_4_net__186_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__186_ : 1'b0;
  assign n_4_net__185_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__185_ : 1'b0;
  assign n_4_net__184_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__184_ : 1'b0;
  assign n_4_net__183_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__183_ : 1'b0;
  assign n_4_net__182_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__182_ : 1'b0;
  assign n_4_net__181_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__181_ : 1'b0;
  assign n_4_net__180_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__180_ : 1'b0;
  assign n_4_net__179_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__179_ : 1'b0;
  assign n_4_net__178_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__178_ : 1'b0;
  assign n_4_net__177_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__177_ : 1'b0;
  assign n_4_net__176_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__176_ : 1'b0;
  assign n_4_net__175_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__175_ : 1'b0;
  assign n_4_net__174_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__174_ : 1'b0;
  assign n_4_net__173_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__173_ : 1'b0;
  assign n_4_net__172_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__172_ : 1'b0;
  assign n_4_net__171_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__171_ : 1'b0;
  assign n_4_net__170_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__170_ : 1'b0;
  assign n_4_net__169_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__169_ : 1'b0;
  assign n_4_net__168_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__168_ : 1'b0;
  assign n_4_net__167_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__167_ : 1'b0;
  assign n_4_net__166_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__166_ : 1'b0;
  assign n_4_net__165_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__165_ : 1'b0;
  assign n_4_net__164_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__164_ : 1'b0;
  assign n_4_net__163_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__163_ : 1'b0;
  assign n_4_net__162_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__162_ : 1'b0;
  assign n_4_net__161_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__161_ : 1'b0;
  assign n_4_net__160_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__160_ : 1'b0;
  assign n_4_net__159_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__159_ : 1'b0;
  assign n_4_net__158_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__158_ : 1'b0;
  assign n_4_net__157_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__157_ : 1'b0;
  assign n_4_net__156_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__156_ : 1'b0;
  assign n_4_net__155_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__155_ : 1'b0;
  assign n_4_net__154_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__154_ : 1'b0;
  assign n_4_net__153_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__153_ : 1'b0;
  assign n_4_net__152_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__152_ : 1'b0;
  assign n_4_net__151_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__151_ : 1'b0;
  assign n_4_net__150_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__150_ : 1'b0;
  assign n_4_net__149_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__149_ : 1'b0;
  assign n_4_net__148_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__148_ : 1'b0;
  assign n_4_net__147_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__147_ : 1'b0;
  assign n_4_net__146_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__146_ : 1'b0;
  assign n_4_net__145_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__145_ : 1'b0;
  assign n_4_net__144_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__144_ : 1'b0;
  assign n_4_net__143_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__143_ : 1'b0;
  assign n_4_net__142_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__142_ : 1'b0;
  assign n_4_net__141_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__141_ : 1'b0;
  assign n_4_net__140_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__140_ : 1'b0;
  assign n_4_net__139_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__139_ : 1'b0;
  assign n_4_net__138_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__138_ : 1'b0;
  assign n_4_net__137_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__137_ : 1'b0;
  assign n_4_net__136_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__136_ : 1'b0;
  assign n_4_net__135_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__135_ : 1'b0;
  assign n_4_net__134_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__134_ : 1'b0;
  assign n_4_net__133_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__133_ : 1'b0;
  assign n_4_net__132_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__132_ : 1'b0;
  assign n_4_net__131_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__131_ : 1'b0;
  assign n_4_net__130_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__130_ : 1'b0;
  assign n_4_net__129_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__129_ : 1'b0;
  assign n_4_net__128_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__128_ : 1'b0;
  assign n_4_net__127_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__127_ : 1'b0;
  assign n_4_net__126_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__126_ : 1'b0;
  assign n_4_net__125_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__125_ : 1'b0;
  assign n_4_net__124_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__124_ : 1'b0;
  assign n_4_net__123_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__123_ : 1'b0;
  assign n_4_net__122_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__122_ : 1'b0;
  assign n_4_net__121_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__121_ : 1'b0;
  assign n_4_net__120_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__120_ : 1'b0;
  assign n_4_net__119_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__119_ : 1'b0;
  assign n_4_net__118_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__118_ : 1'b0;
  assign n_4_net__117_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__117_ : 1'b0;
  assign n_4_net__116_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__116_ : 1'b0;
  assign n_4_net__115_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__115_ : 1'b0;
  assign n_4_net__114_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__114_ : 1'b0;
  assign n_4_net__113_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__113_ : 1'b0;
  assign n_4_net__112_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__112_ : 1'b0;
  assign n_4_net__111_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__111_ : 1'b0;
  assign n_4_net__110_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__110_ : 1'b0;
  assign n_4_net__109_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__109_ : 1'b0;
  assign n_4_net__108_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__108_ : 1'b0;
  assign n_4_net__107_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__107_ : 1'b0;
  assign n_4_net__106_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__106_ : 1'b0;
  assign n_4_net__105_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__105_ : 1'b0;
  assign n_4_net__104_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__104_ : 1'b0;
  assign n_4_net__103_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__103_ : 1'b0;
  assign n_4_net__102_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__102_ : 1'b0;
  assign n_4_net__101_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__101_ : 1'b0;
  assign n_4_net__100_ = (N60)? 1'b0 : 
                         (N62)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N66)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N70)? 1'b0 : 
                         (N72)? 1'b0 : 
                         (N74)? 1'b0 : 
                         (N61)? 1'b0 : 
                         (N63)? 1'b0 : 
                         (N65)? 1'b0 : 
                         (N67)? 1'b0 : 
                         (N69)? 1'b0 : 
                         (N71)? 1'b0 : 
                         (N73)? 1'b0 : 
                         (N75)? data_head_15__100_ : 1'b0;
  assign n_4_net__99_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__99_ : 1'b0;
  assign n_4_net__98_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__98_ : 1'b0;
  assign n_4_net__97_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__97_ : 1'b0;
  assign n_4_net__96_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__96_ : 1'b0;
  assign n_4_net__95_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__95_ : 1'b0;
  assign n_4_net__94_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__94_ : 1'b0;
  assign n_4_net__93_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__93_ : 1'b0;
  assign n_4_net__92_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__92_ : 1'b0;
  assign n_4_net__91_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__91_ : 1'b0;
  assign n_4_net__90_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__90_ : 1'b0;
  assign n_4_net__89_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__89_ : 1'b0;
  assign n_4_net__88_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__88_ : 1'b0;
  assign n_4_net__87_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__87_ : 1'b0;
  assign n_4_net__86_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__86_ : 1'b0;
  assign n_4_net__85_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__85_ : 1'b0;
  assign n_4_net__84_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__84_ : 1'b0;
  assign n_4_net__83_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__83_ : 1'b0;
  assign n_4_net__82_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__82_ : 1'b0;
  assign n_4_net__81_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__81_ : 1'b0;
  assign n_4_net__80_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__80_ : 1'b0;
  assign n_4_net__79_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__79_ : 1'b0;
  assign n_4_net__78_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__78_ : 1'b0;
  assign n_4_net__77_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__77_ : 1'b0;
  assign n_4_net__76_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__76_ : 1'b0;
  assign n_4_net__75_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__75_ : 1'b0;
  assign n_4_net__74_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__74_ : 1'b0;
  assign n_4_net__73_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__73_ : 1'b0;
  assign n_4_net__72_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__72_ : 1'b0;
  assign n_4_net__71_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__71_ : 1'b0;
  assign n_4_net__70_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__70_ : 1'b0;
  assign n_4_net__69_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__69_ : 1'b0;
  assign n_4_net__68_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__68_ : 1'b0;
  assign n_4_net__67_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__67_ : 1'b0;
  assign n_4_net__66_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__66_ : 1'b0;
  assign n_4_net__65_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__65_ : 1'b0;
  assign n_4_net__64_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__64_ : 1'b0;
  assign n_4_net__63_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__63_ : 1'b0;
  assign n_4_net__62_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__62_ : 1'b0;
  assign n_4_net__61_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__61_ : 1'b0;
  assign n_4_net__60_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__60_ : 1'b0;
  assign n_4_net__59_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__59_ : 1'b0;
  assign n_4_net__58_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__58_ : 1'b0;
  assign n_4_net__57_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__57_ : 1'b0;
  assign n_4_net__56_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__56_ : 1'b0;
  assign n_4_net__55_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__55_ : 1'b0;
  assign n_4_net__54_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__54_ : 1'b0;
  assign n_4_net__53_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__53_ : 1'b0;
  assign n_4_net__52_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__52_ : 1'b0;
  assign n_4_net__51_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__51_ : 1'b0;
  assign n_4_net__50_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__50_ : 1'b0;
  assign n_4_net__49_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__49_ : 1'b0;
  assign n_4_net__48_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__48_ : 1'b0;
  assign n_4_net__47_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__47_ : 1'b0;
  assign n_4_net__46_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__46_ : 1'b0;
  assign n_4_net__45_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__45_ : 1'b0;
  assign n_4_net__44_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__44_ : 1'b0;
  assign n_4_net__43_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__43_ : 1'b0;
  assign n_4_net__42_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__42_ : 1'b0;
  assign n_4_net__41_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__41_ : 1'b0;
  assign n_4_net__40_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__40_ : 1'b0;
  assign n_4_net__39_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__39_ : 1'b0;
  assign n_4_net__38_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__38_ : 1'b0;
  assign n_4_net__37_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__37_ : 1'b0;
  assign n_4_net__36_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__36_ : 1'b0;
  assign n_4_net__35_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__35_ : 1'b0;
  assign n_4_net__34_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__34_ : 1'b0;
  assign n_4_net__33_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__33_ : 1'b0;
  assign n_4_net__32_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__32_ : 1'b0;
  assign n_4_net__31_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__31_ : 1'b0;
  assign n_4_net__30_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__30_ : 1'b0;
  assign n_4_net__29_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__29_ : 1'b0;
  assign n_4_net__28_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__28_ : 1'b0;
  assign n_4_net__27_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__27_ : 1'b0;
  assign n_4_net__26_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__26_ : 1'b0;
  assign n_4_net__25_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__25_ : 1'b0;
  assign n_4_net__24_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__24_ : 1'b0;
  assign n_4_net__23_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__23_ : 1'b0;
  assign n_4_net__22_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__22_ : 1'b0;
  assign n_4_net__21_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__21_ : 1'b0;
  assign n_4_net__20_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__20_ : 1'b0;
  assign n_4_net__19_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__19_ : 1'b0;
  assign n_4_net__18_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__18_ : 1'b0;
  assign n_4_net__17_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__17_ : 1'b0;
  assign n_4_net__16_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__16_ : 1'b0;
  assign n_4_net__15_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__15_ : 1'b0;
  assign n_4_net__14_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__14_ : 1'b0;
  assign n_4_net__13_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__13_ : 1'b0;
  assign n_4_net__12_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__12_ : 1'b0;
  assign n_4_net__11_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__11_ : 1'b0;
  assign n_4_net__10_ = (N60)? 1'b0 : 
                        (N62)? 1'b0 : 
                        (N64)? 1'b0 : 
                        (N66)? 1'b0 : 
                        (N68)? 1'b0 : 
                        (N70)? 1'b0 : 
                        (N72)? 1'b0 : 
                        (N74)? 1'b0 : 
                        (N61)? 1'b0 : 
                        (N63)? 1'b0 : 
                        (N65)? 1'b0 : 
                        (N67)? 1'b0 : 
                        (N69)? 1'b0 : 
                        (N71)? 1'b0 : 
                        (N73)? 1'b0 : 
                        (N75)? data_head_15__10_ : 1'b0;
  assign n_4_net__9_ = (N60)? 1'b0 : 
                       (N62)? 1'b0 : 
                       (N64)? 1'b0 : 
                       (N66)? 1'b0 : 
                       (N68)? 1'b0 : 
                       (N70)? 1'b0 : 
                       (N72)? 1'b0 : 
                       (N74)? 1'b0 : 
                       (N61)? 1'b0 : 
                       (N63)? 1'b0 : 
                       (N65)? 1'b0 : 
                       (N67)? 1'b0 : 
                       (N69)? 1'b0 : 
                       (N71)? 1'b0 : 
                       (N73)? 1'b0 : 
                       (N75)? data_head_15__9_ : 1'b0;
  assign n_4_net__8_ = (N60)? 1'b0 : 
                       (N62)? 1'b0 : 
                       (N64)? 1'b0 : 
                       (N66)? 1'b0 : 
                       (N68)? 1'b0 : 
                       (N70)? 1'b0 : 
                       (N72)? 1'b0 : 
                       (N74)? 1'b0 : 
                       (N61)? 1'b0 : 
                       (N63)? 1'b0 : 
                       (N65)? 1'b0 : 
                       (N67)? 1'b0 : 
                       (N69)? 1'b0 : 
                       (N71)? 1'b0 : 
                       (N73)? 1'b0 : 
                       (N75)? data_head_15__8_ : 1'b0;
  assign n_4_net__7_ = (N60)? 1'b0 : 
                       (N62)? 1'b0 : 
                       (N64)? 1'b0 : 
                       (N66)? 1'b0 : 
                       (N68)? 1'b0 : 
                       (N70)? 1'b0 : 
                       (N72)? 1'b0 : 
                       (N74)? 1'b0 : 
                       (N61)? 1'b0 : 
                       (N63)? 1'b0 : 
                       (N65)? 1'b0 : 
                       (N67)? 1'b0 : 
                       (N69)? 1'b0 : 
                       (N71)? 1'b0 : 
                       (N73)? 1'b0 : 
                       (N75)? data_head_15__7_ : 1'b0;
  assign n_4_net__6_ = (N60)? 1'b0 : 
                       (N62)? 1'b0 : 
                       (N64)? 1'b0 : 
                       (N66)? 1'b0 : 
                       (N68)? 1'b0 : 
                       (N70)? 1'b0 : 
                       (N72)? 1'b0 : 
                       (N74)? 1'b0 : 
                       (N61)? 1'b0 : 
                       (N63)? 1'b0 : 
                       (N65)? 1'b0 : 
                       (N67)? 1'b0 : 
                       (N69)? 1'b0 : 
                       (N71)? 1'b0 : 
                       (N73)? 1'b0 : 
                       (N75)? data_head_15__6_ : 1'b0;
  assign n_4_net__5_ = (N60)? 1'b0 : 
                       (N62)? 1'b0 : 
                       (N64)? 1'b0 : 
                       (N66)? 1'b0 : 
                       (N68)? 1'b0 : 
                       (N70)? 1'b0 : 
                       (N72)? 1'b0 : 
                       (N74)? 1'b0 : 
                       (N61)? 1'b0 : 
                       (N63)? 1'b0 : 
                       (N65)? 1'b0 : 
                       (N67)? 1'b0 : 
                       (N69)? 1'b0 : 
                       (N71)? 1'b0 : 
                       (N73)? 1'b0 : 
                       (N75)? data_head_15__5_ : 1'b0;
  assign n_4_net__4_ = (N60)? 1'b0 : 
                       (N62)? 1'b0 : 
                       (N64)? 1'b0 : 
                       (N66)? 1'b0 : 
                       (N68)? 1'b0 : 
                       (N70)? 1'b0 : 
                       (N72)? 1'b0 : 
                       (N74)? 1'b0 : 
                       (N61)? 1'b0 : 
                       (N63)? 1'b0 : 
                       (N65)? 1'b0 : 
                       (N67)? 1'b0 : 
                       (N69)? 1'b0 : 
                       (N71)? 1'b0 : 
                       (N73)? 1'b0 : 
                       (N75)? data_head_15__4_ : 1'b0;
  assign n_4_net__3_ = (N60)? 1'b0 : 
                       (N62)? 1'b0 : 
                       (N64)? 1'b0 : 
                       (N66)? 1'b0 : 
                       (N68)? 1'b0 : 
                       (N70)? 1'b0 : 
                       (N72)? 1'b0 : 
                       (N74)? 1'b0 : 
                       (N61)? 1'b0 : 
                       (N63)? 1'b0 : 
                       (N65)? 1'b0 : 
                       (N67)? 1'b0 : 
                       (N69)? 1'b0 : 
                       (N71)? 1'b0 : 
                       (N73)? 1'b0 : 
                       (N75)? data_head_15__3_ : 1'b0;
  assign n_4_net__2_ = (N60)? 1'b0 : 
                       (N62)? 1'b0 : 
                       (N64)? 1'b0 : 
                       (N66)? 1'b0 : 
                       (N68)? 1'b0 : 
                       (N70)? 1'b0 : 
                       (N72)? 1'b0 : 
                       (N74)? 1'b0 : 
                       (N61)? 1'b0 : 
                       (N63)? 1'b0 : 
                       (N65)? 1'b0 : 
                       (N67)? 1'b0 : 
                       (N69)? 1'b0 : 
                       (N71)? 1'b0 : 
                       (N73)? 1'b0 : 
                       (N75)? data_head_15__2_ : 1'b0;
  assign n_4_net__1_ = (N60)? 1'b0 : 
                       (N62)? 1'b0 : 
                       (N64)? 1'b0 : 
                       (N66)? 1'b0 : 
                       (N68)? 1'b0 : 
                       (N70)? 1'b0 : 
                       (N72)? 1'b0 : 
                       (N74)? 1'b0 : 
                       (N61)? 1'b0 : 
                       (N63)? 1'b0 : 
                       (N65)? 1'b0 : 
                       (N67)? 1'b0 : 
                       (N69)? 1'b0 : 
                       (N71)? 1'b0 : 
                       (N73)? 1'b0 : 
                       (N75)? data_head_15__1_ : 1'b0;
  assign n_4_net__0_ = (N60)? 1'b0 : 
                       (N62)? 1'b0 : 
                       (N64)? 1'b0 : 
                       (N66)? 1'b0 : 
                       (N68)? 1'b0 : 
                       (N70)? 1'b0 : 
                       (N72)? 1'b0 : 
                       (N74)? 1'b0 : 
                       (N61)? 1'b0 : 
                       (N63)? 1'b0 : 
                       (N65)? 1'b0 : 
                       (N67)? 1'b0 : 
                       (N69)? 1'b0 : 
                       (N71)? 1'b0 : 
                       (N73)? 1'b0 : 
                       (N75)? data_head_15__0_ : 1'b0;

  bsg_rr_f2f_output_width_p64_num_out_p8_middle_meet_p8
  oc_7__out_chan_bsg_rr_ff_out
  (
    .clk(clk),
    .reset(n_5_net_),
    .ready_i(ready_i),
    .ready_head_o({ ready_head_7__7_, ready_head_7__6_, ready_head_7__5_, ready_head_7__4_, ready_head_7__3_, ready_head_7__2_, ready_head_7__1_, ready_head_7__0_ }),
    .go_channels_i(go_channels),
    .go_cnt_i(go_cnt),
    .data_head_i(oc_7__out_chan_data_head_array),
    .valid_o({ valid_int_o_7__7_, valid_int_o_7__6_, valid_int_o_7__5_, valid_int_o_7__4_, valid_int_o_7__3_, valid_int_o_7__2_, valid_int_o_7__1_, valid_int_o_7__0_ }),
    .data_o({ data_int_o_7__511_, data_int_o_7__510_, data_int_o_7__509_, data_int_o_7__508_, data_int_o_7__507_, data_int_o_7__506_, data_int_o_7__505_, data_int_o_7__504_, data_int_o_7__503_, data_int_o_7__502_, data_int_o_7__501_, data_int_o_7__500_, data_int_o_7__499_, data_int_o_7__498_, data_int_o_7__497_, data_int_o_7__496_, data_int_o_7__495_, data_int_o_7__494_, data_int_o_7__493_, data_int_o_7__492_, data_int_o_7__491_, data_int_o_7__490_, data_int_o_7__489_, data_int_o_7__488_, data_int_o_7__487_, data_int_o_7__486_, data_int_o_7__485_, data_int_o_7__484_, data_int_o_7__483_, data_int_o_7__482_, data_int_o_7__481_, data_int_o_7__480_, data_int_o_7__479_, data_int_o_7__478_, data_int_o_7__477_, data_int_o_7__476_, data_int_o_7__475_, data_int_o_7__474_, data_int_o_7__473_, data_int_o_7__472_, data_int_o_7__471_, data_int_o_7__470_, data_int_o_7__469_, data_int_o_7__468_, data_int_o_7__467_, data_int_o_7__466_, data_int_o_7__465_, data_int_o_7__464_, data_int_o_7__463_, data_int_o_7__462_, data_int_o_7__461_, data_int_o_7__460_, data_int_o_7__459_, data_int_o_7__458_, data_int_o_7__457_, data_int_o_7__456_, data_int_o_7__455_, data_int_o_7__454_, data_int_o_7__453_, data_int_o_7__452_, data_int_o_7__451_, data_int_o_7__450_, data_int_o_7__449_, data_int_o_7__448_, data_int_o_7__447_, data_int_o_7__446_, data_int_o_7__445_, data_int_o_7__444_, data_int_o_7__443_, data_int_o_7__442_, data_int_o_7__441_, data_int_o_7__440_, data_int_o_7__439_, data_int_o_7__438_, data_int_o_7__437_, data_int_o_7__436_, data_int_o_7__435_, data_int_o_7__434_, data_int_o_7__433_, data_int_o_7__432_, data_int_o_7__431_, data_int_o_7__430_, data_int_o_7__429_, data_int_o_7__428_, data_int_o_7__427_, data_int_o_7__426_, data_int_o_7__425_, data_int_o_7__424_, data_int_o_7__423_, data_int_o_7__422_, data_int_o_7__421_, data_int_o_7__420_, data_int_o_7__419_, data_int_o_7__418_, data_int_o_7__417_, data_int_o_7__416_, data_int_o_7__415_, data_int_o_7__414_, data_int_o_7__413_, data_int_o_7__412_, data_int_o_7__411_, data_int_o_7__410_, data_int_o_7__409_, data_int_o_7__408_, data_int_o_7__407_, data_int_o_7__406_, data_int_o_7__405_, data_int_o_7__404_, data_int_o_7__403_, data_int_o_7__402_, data_int_o_7__401_, data_int_o_7__400_, data_int_o_7__399_, data_int_o_7__398_, data_int_o_7__397_, data_int_o_7__396_, data_int_o_7__395_, data_int_o_7__394_, data_int_o_7__393_, data_int_o_7__392_, data_int_o_7__391_, data_int_o_7__390_, data_int_o_7__389_, data_int_o_7__388_, data_int_o_7__387_, data_int_o_7__386_, data_int_o_7__385_, data_int_o_7__384_, data_int_o_7__383_, data_int_o_7__382_, data_int_o_7__381_, data_int_o_7__380_, data_int_o_7__379_, data_int_o_7__378_, data_int_o_7__377_, data_int_o_7__376_, data_int_o_7__375_, data_int_o_7__374_, data_int_o_7__373_, data_int_o_7__372_, data_int_o_7__371_, data_int_o_7__370_, data_int_o_7__369_, data_int_o_7__368_, data_int_o_7__367_, data_int_o_7__366_, data_int_o_7__365_, data_int_o_7__364_, data_int_o_7__363_, data_int_o_7__362_, data_int_o_7__361_, data_int_o_7__360_, data_int_o_7__359_, data_int_o_7__358_, data_int_o_7__357_, data_int_o_7__356_, data_int_o_7__355_, data_int_o_7__354_, data_int_o_7__353_, data_int_o_7__352_, data_int_o_7__351_, data_int_o_7__350_, data_int_o_7__349_, data_int_o_7__348_, data_int_o_7__347_, data_int_o_7__346_, data_int_o_7__345_, data_int_o_7__344_, data_int_o_7__343_, data_int_o_7__342_, data_int_o_7__341_, data_int_o_7__340_, data_int_o_7__339_, data_int_o_7__338_, data_int_o_7__337_, data_int_o_7__336_, data_int_o_7__335_, data_int_o_7__334_, data_int_o_7__333_, data_int_o_7__332_, data_int_o_7__331_, data_int_o_7__330_, data_int_o_7__329_, data_int_o_7__328_, data_int_o_7__327_, data_int_o_7__326_, data_int_o_7__325_, data_int_o_7__324_, data_int_o_7__323_, data_int_o_7__322_, data_int_o_7__321_, data_int_o_7__320_, data_int_o_7__319_, data_int_o_7__318_, data_int_o_7__317_, data_int_o_7__316_, data_int_o_7__315_, data_int_o_7__314_, data_int_o_7__313_, data_int_o_7__312_, data_int_o_7__311_, data_int_o_7__310_, data_int_o_7__309_, data_int_o_7__308_, data_int_o_7__307_, data_int_o_7__306_, data_int_o_7__305_, data_int_o_7__304_, data_int_o_7__303_, data_int_o_7__302_, data_int_o_7__301_, data_int_o_7__300_, data_int_o_7__299_, data_int_o_7__298_, data_int_o_7__297_, data_int_o_7__296_, data_int_o_7__295_, data_int_o_7__294_, data_int_o_7__293_, data_int_o_7__292_, data_int_o_7__291_, data_int_o_7__290_, data_int_o_7__289_, data_int_o_7__288_, data_int_o_7__287_, data_int_o_7__286_, data_int_o_7__285_, data_int_o_7__284_, data_int_o_7__283_, data_int_o_7__282_, data_int_o_7__281_, data_int_o_7__280_, data_int_o_7__279_, data_int_o_7__278_, data_int_o_7__277_, data_int_o_7__276_, data_int_o_7__275_, data_int_o_7__274_, data_int_o_7__273_, data_int_o_7__272_, data_int_o_7__271_, data_int_o_7__270_, data_int_o_7__269_, data_int_o_7__268_, data_int_o_7__267_, data_int_o_7__266_, data_int_o_7__265_, data_int_o_7__264_, data_int_o_7__263_, data_int_o_7__262_, data_int_o_7__261_, data_int_o_7__260_, data_int_o_7__259_, data_int_o_7__258_, data_int_o_7__257_, data_int_o_7__256_, data_int_o_7__255_, data_int_o_7__254_, data_int_o_7__253_, data_int_o_7__252_, data_int_o_7__251_, data_int_o_7__250_, data_int_o_7__249_, data_int_o_7__248_, data_int_o_7__247_, data_int_o_7__246_, data_int_o_7__245_, data_int_o_7__244_, data_int_o_7__243_, data_int_o_7__242_, data_int_o_7__241_, data_int_o_7__240_, data_int_o_7__239_, data_int_o_7__238_, data_int_o_7__237_, data_int_o_7__236_, data_int_o_7__235_, data_int_o_7__234_, data_int_o_7__233_, data_int_o_7__232_, data_int_o_7__231_, data_int_o_7__230_, data_int_o_7__229_, data_int_o_7__228_, data_int_o_7__227_, data_int_o_7__226_, data_int_o_7__225_, data_int_o_7__224_, data_int_o_7__223_, data_int_o_7__222_, data_int_o_7__221_, data_int_o_7__220_, data_int_o_7__219_, data_int_o_7__218_, data_int_o_7__217_, data_int_o_7__216_, data_int_o_7__215_, data_int_o_7__214_, data_int_o_7__213_, data_int_o_7__212_, data_int_o_7__211_, data_int_o_7__210_, data_int_o_7__209_, data_int_o_7__208_, data_int_o_7__207_, data_int_o_7__206_, data_int_o_7__205_, data_int_o_7__204_, data_int_o_7__203_, data_int_o_7__202_, data_int_o_7__201_, data_int_o_7__200_, data_int_o_7__199_, data_int_o_7__198_, data_int_o_7__197_, data_int_o_7__196_, data_int_o_7__195_, data_int_o_7__194_, data_int_o_7__193_, data_int_o_7__192_, data_int_o_7__191_, data_int_o_7__190_, data_int_o_7__189_, data_int_o_7__188_, data_int_o_7__187_, data_int_o_7__186_, data_int_o_7__185_, data_int_o_7__184_, data_int_o_7__183_, data_int_o_7__182_, data_int_o_7__181_, data_int_o_7__180_, data_int_o_7__179_, data_int_o_7__178_, data_int_o_7__177_, data_int_o_7__176_, data_int_o_7__175_, data_int_o_7__174_, data_int_o_7__173_, data_int_o_7__172_, data_int_o_7__171_, data_int_o_7__170_, data_int_o_7__169_, data_int_o_7__168_, data_int_o_7__167_, data_int_o_7__166_, data_int_o_7__165_, data_int_o_7__164_, data_int_o_7__163_, data_int_o_7__162_, data_int_o_7__161_, data_int_o_7__160_, data_int_o_7__159_, data_int_o_7__158_, data_int_o_7__157_, data_int_o_7__156_, data_int_o_7__155_, data_int_o_7__154_, data_int_o_7__153_, data_int_o_7__152_, data_int_o_7__151_, data_int_o_7__150_, data_int_o_7__149_, data_int_o_7__148_, data_int_o_7__147_, data_int_o_7__146_, data_int_o_7__145_, data_int_o_7__144_, data_int_o_7__143_, data_int_o_7__142_, data_int_o_7__141_, data_int_o_7__140_, data_int_o_7__139_, data_int_o_7__138_, data_int_o_7__137_, data_int_o_7__136_, data_int_o_7__135_, data_int_o_7__134_, data_int_o_7__133_, data_int_o_7__132_, data_int_o_7__131_, data_int_o_7__130_, data_int_o_7__129_, data_int_o_7__128_, data_int_o_7__127_, data_int_o_7__126_, data_int_o_7__125_, data_int_o_7__124_, data_int_o_7__123_, data_int_o_7__122_, data_int_o_7__121_, data_int_o_7__120_, data_int_o_7__119_, data_int_o_7__118_, data_int_o_7__117_, data_int_o_7__116_, data_int_o_7__115_, data_int_o_7__114_, data_int_o_7__113_, data_int_o_7__112_, data_int_o_7__111_, data_int_o_7__110_, data_int_o_7__109_, data_int_o_7__108_, data_int_o_7__107_, data_int_o_7__106_, data_int_o_7__105_, data_int_o_7__104_, data_int_o_7__103_, data_int_o_7__102_, data_int_o_7__101_, data_int_o_7__100_, data_int_o_7__99_, data_int_o_7__98_, data_int_o_7__97_, data_int_o_7__96_, data_int_o_7__95_, data_int_o_7__94_, data_int_o_7__93_, data_int_o_7__92_, data_int_o_7__91_, data_int_o_7__90_, data_int_o_7__89_, data_int_o_7__88_, data_int_o_7__87_, data_int_o_7__86_, data_int_o_7__85_, data_int_o_7__84_, data_int_o_7__83_, data_int_o_7__82_, data_int_o_7__81_, data_int_o_7__80_, data_int_o_7__79_, data_int_o_7__78_, data_int_o_7__77_, data_int_o_7__76_, data_int_o_7__75_, data_int_o_7__74_, data_int_o_7__73_, data_int_o_7__72_, data_int_o_7__71_, data_int_o_7__70_, data_int_o_7__69_, data_int_o_7__68_, data_int_o_7__67_, data_int_o_7__66_, data_int_o_7__65_, data_int_o_7__64_, data_int_o_7__63_, data_int_o_7__62_, data_int_o_7__61_, data_int_o_7__60_, data_int_o_7__59_, data_int_o_7__58_, data_int_o_7__57_, data_int_o_7__56_, data_int_o_7__55_, data_int_o_7__54_, data_int_o_7__53_, data_int_o_7__52_, data_int_o_7__51_, data_int_o_7__50_, data_int_o_7__49_, data_int_o_7__48_, data_int_o_7__47_, data_int_o_7__46_, data_int_o_7__45_, data_int_o_7__44_, data_int_o_7__43_, data_int_o_7__42_, data_int_o_7__41_, data_int_o_7__40_, data_int_o_7__39_, data_int_o_7__38_, data_int_o_7__37_, data_int_o_7__36_, data_int_o_7__35_, data_int_o_7__34_, data_int_o_7__33_, data_int_o_7__32_, data_int_o_7__31_, data_int_o_7__30_, data_int_o_7__29_, data_int_o_7__28_, data_int_o_7__27_, data_int_o_7__26_, data_int_o_7__25_, data_int_o_7__24_, data_int_o_7__23_, data_int_o_7__22_, data_int_o_7__21_, data_int_o_7__20_, data_int_o_7__19_, data_int_o_7__18_, data_int_o_7__17_, data_int_o_7__16_, data_int_o_7__15_, data_int_o_7__14_, data_int_o_7__13_, data_int_o_7__12_, data_int_o_7__11_, data_int_o_7__10_, data_int_o_7__9_, data_int_o_7__8_, data_int_o_7__7_, data_int_o_7__6_, data_int_o_7__5_, data_int_o_7__4_, data_int_o_7__3_, data_int_o_7__2_, data_int_o_7__1_, data_int_o_7__0_ })
  );

  assign N76 = in_top_channel_i[2] & in_top_channel_i[3];
  assign N77 = in_top_channel_i[1] & N76;
  assign N78 = in_top_channel_i[0] & N77;
  assign N79 = ~N78;
  assign N80 = out_top_channel_i[1] & out_top_channel_i[2];
  assign N81 = out_top_channel_i[0] & N80;
  assign N82 = ~N81;
  assign N0 = ~in_top_channel_i[0];
  assign N1 = ~in_top_channel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & in_top_channel_i[1];
  assign N4 = in_top_channel_i[0] & N1;
  assign N5 = in_top_channel_i[0] & in_top_channel_i[1];
  assign N6 = ~in_top_channel_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & in_top_channel_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & in_top_channel_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & in_top_channel_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & in_top_channel_i[2];
  assign N15 = ~in_top_channel_i[3];
  assign N16 = N7 & N15;
  assign N17 = N7 & in_top_channel_i[3];
  assign N18 = N9 & N15;
  assign N19 = N9 & in_top_channel_i[3];
  assign N20 = N11 & N15;
  assign N21 = N11 & in_top_channel_i[3];
  assign N22 = N13 & N15;
  assign N23 = N13 & in_top_channel_i[3];
  assign N24 = N8 & N15;
  assign N25 = N8 & in_top_channel_i[3];
  assign N26 = N10 & N15;
  assign N27 = N10 & in_top_channel_i[3];
  assign N28 = N12 & N15;
  assign N29 = N12 & in_top_channel_i[3];
  assign N30 = N14 & N15;
  assign N31 = N14 & in_top_channel_i[3];
  assign N32 = ~out_top_channel_i[0];
  assign N33 = ~out_top_channel_i[1];
  assign N34 = N32 & N33;
  assign N35 = N32 & out_top_channel_i[1];
  assign N36 = out_top_channel_i[0] & N33;
  assign N37 = out_top_channel_i[0] & out_top_channel_i[1];
  assign N38 = ~out_top_channel_i[2];
  assign N39 = N34 & N38;
  assign N40 = N34 & out_top_channel_i[2];
  assign N41 = N36 & N38;
  assign N42 = N36 & out_top_channel_i[2];
  assign N43 = N35 & N38;
  assign N44 = N35 & out_top_channel_i[2];
  assign N45 = N37 & N38;
  assign N46 = N37 & out_top_channel_i[2];
  assign N47 = N34 & N38;
  assign N48 = N34 & out_top_channel_i[2];
  assign N49 = N36 & N38;
  assign N50 = N36 & out_top_channel_i[2];
  assign N51 = N35 & N38;
  assign N52 = N35 & out_top_channel_i[2];
  assign N53 = N37 & N38;
  assign N54 = N37 & out_top_channel_i[2];
  assign n_0_net_ = reset | N79;
  assign N55 = N37 & N38;
  assign N56 = N37 & out_top_channel_i[2];
  assign N57 = N13 & N15;
  assign N58 = N13 & in_top_channel_i[3];
  assign N59 = N14 & in_top_channel_i[3];
  assign N60 = N7 & N15;
  assign N61 = N7 & in_top_channel_i[3];
  assign N62 = N9 & N15;
  assign N63 = N9 & in_top_channel_i[3];
  assign N64 = N11 & N15;
  assign N65 = N11 & in_top_channel_i[3];
  assign N66 = N13 & N15;
  assign N67 = N13 & in_top_channel_i[3];
  assign N68 = N8 & N15;
  assign N69 = N8 & in_top_channel_i[3];
  assign N70 = N10 & N15;
  assign N71 = N10 & in_top_channel_i[3];
  assign N72 = N12 & N15;
  assign N73 = N12 & in_top_channel_i[3];
  assign N74 = N14 & N15;
  assign N75 = N14 & in_top_channel_i[3];
  assign n_5_net_ = reset | N82;

endmodule

